////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module AES in file /AGEMA/Designs/AES_round-based/AGEMA/AES.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module AES_HPC2_ClockGating_d1 (plaintext_s0, key_s0, clk, reset, key_s1, plaintext_s1, Fresh, ciphertext_s0, done, ciphertext_s1, Synch);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] key_s1 ;
    input [127:0] plaintext_s1 ;
    input [679:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    output Synch ;
    wire n283 ;
    wire n285 ;
    wire n314 ;
    wire n315 ;
    wire n316 ;
    wire n317 ;
    wire n318 ;
    wire n319 ;
    wire n320 ;
    wire n321 ;
    wire n322 ;
    wire n323 ;
    wire n324 ;
    wire n325 ;
    wire n326 ;
    wire n327 ;
    wire n328 ;
    wire n329 ;
    wire n330 ;
    wire n331 ;
    wire n332 ;
    wire n333 ;
    wire n334 ;
    wire n335 ;
    wire n336 ;
    wire n337 ;
    wire n338 ;
    wire n339 ;
    wire RoundReg_Inst_ff_SDE_0_next_state ;
    wire RoundReg_Inst_ff_SDE_1_next_state ;
    wire RoundReg_Inst_ff_SDE_2_next_state ;
    wire RoundReg_Inst_ff_SDE_3_next_state ;
    wire RoundReg_Inst_ff_SDE_4_next_state ;
    wire RoundReg_Inst_ff_SDE_5_next_state ;
    wire RoundReg_Inst_ff_SDE_6_next_state ;
    wire RoundReg_Inst_ff_SDE_7_next_state ;
    wire RoundReg_Inst_ff_SDE_8_next_state ;
    wire RoundReg_Inst_ff_SDE_9_next_state ;
    wire RoundReg_Inst_ff_SDE_10_next_state ;
    wire RoundReg_Inst_ff_SDE_11_next_state ;
    wire RoundReg_Inst_ff_SDE_12_next_state ;
    wire RoundReg_Inst_ff_SDE_13_next_state ;
    wire RoundReg_Inst_ff_SDE_14_next_state ;
    wire RoundReg_Inst_ff_SDE_15_next_state ;
    wire RoundReg_Inst_ff_SDE_16_next_state ;
    wire RoundReg_Inst_ff_SDE_17_next_state ;
    wire RoundReg_Inst_ff_SDE_18_next_state ;
    wire RoundReg_Inst_ff_SDE_19_next_state ;
    wire RoundReg_Inst_ff_SDE_20_next_state ;
    wire RoundReg_Inst_ff_SDE_21_next_state ;
    wire RoundReg_Inst_ff_SDE_22_next_state ;
    wire RoundReg_Inst_ff_SDE_23_next_state ;
    wire RoundReg_Inst_ff_SDE_24_next_state ;
    wire RoundReg_Inst_ff_SDE_25_next_state ;
    wire RoundReg_Inst_ff_SDE_26_next_state ;
    wire RoundReg_Inst_ff_SDE_27_next_state ;
    wire RoundReg_Inst_ff_SDE_28_next_state ;
    wire RoundReg_Inst_ff_SDE_29_next_state ;
    wire RoundReg_Inst_ff_SDE_30_next_state ;
    wire RoundReg_Inst_ff_SDE_31_next_state ;
    wire RoundReg_Inst_ff_SDE_32_next_state ;
    wire RoundReg_Inst_ff_SDE_33_next_state ;
    wire RoundReg_Inst_ff_SDE_34_next_state ;
    wire RoundReg_Inst_ff_SDE_35_next_state ;
    wire RoundReg_Inst_ff_SDE_36_next_state ;
    wire RoundReg_Inst_ff_SDE_37_next_state ;
    wire RoundReg_Inst_ff_SDE_38_next_state ;
    wire RoundReg_Inst_ff_SDE_39_next_state ;
    wire RoundReg_Inst_ff_SDE_40_next_state ;
    wire RoundReg_Inst_ff_SDE_41_next_state ;
    wire RoundReg_Inst_ff_SDE_42_next_state ;
    wire RoundReg_Inst_ff_SDE_43_next_state ;
    wire RoundReg_Inst_ff_SDE_44_next_state ;
    wire RoundReg_Inst_ff_SDE_45_next_state ;
    wire RoundReg_Inst_ff_SDE_46_next_state ;
    wire RoundReg_Inst_ff_SDE_47_next_state ;
    wire RoundReg_Inst_ff_SDE_48_next_state ;
    wire RoundReg_Inst_ff_SDE_49_next_state ;
    wire RoundReg_Inst_ff_SDE_50_next_state ;
    wire RoundReg_Inst_ff_SDE_51_next_state ;
    wire RoundReg_Inst_ff_SDE_52_next_state ;
    wire RoundReg_Inst_ff_SDE_53_next_state ;
    wire RoundReg_Inst_ff_SDE_54_next_state ;
    wire RoundReg_Inst_ff_SDE_55_next_state ;
    wire RoundReg_Inst_ff_SDE_56_next_state ;
    wire RoundReg_Inst_ff_SDE_57_next_state ;
    wire RoundReg_Inst_ff_SDE_58_next_state ;
    wire RoundReg_Inst_ff_SDE_59_next_state ;
    wire RoundReg_Inst_ff_SDE_60_next_state ;
    wire RoundReg_Inst_ff_SDE_61_next_state ;
    wire RoundReg_Inst_ff_SDE_62_next_state ;
    wire RoundReg_Inst_ff_SDE_63_next_state ;
    wire RoundReg_Inst_ff_SDE_64_next_state ;
    wire RoundReg_Inst_ff_SDE_65_next_state ;
    wire RoundReg_Inst_ff_SDE_66_next_state ;
    wire RoundReg_Inst_ff_SDE_67_next_state ;
    wire RoundReg_Inst_ff_SDE_68_next_state ;
    wire RoundReg_Inst_ff_SDE_69_next_state ;
    wire RoundReg_Inst_ff_SDE_70_next_state ;
    wire RoundReg_Inst_ff_SDE_71_next_state ;
    wire RoundReg_Inst_ff_SDE_72_next_state ;
    wire RoundReg_Inst_ff_SDE_73_next_state ;
    wire RoundReg_Inst_ff_SDE_74_next_state ;
    wire RoundReg_Inst_ff_SDE_75_next_state ;
    wire RoundReg_Inst_ff_SDE_76_next_state ;
    wire RoundReg_Inst_ff_SDE_77_next_state ;
    wire RoundReg_Inst_ff_SDE_78_next_state ;
    wire RoundReg_Inst_ff_SDE_79_next_state ;
    wire RoundReg_Inst_ff_SDE_80_next_state ;
    wire RoundReg_Inst_ff_SDE_81_next_state ;
    wire RoundReg_Inst_ff_SDE_82_next_state ;
    wire RoundReg_Inst_ff_SDE_83_next_state ;
    wire RoundReg_Inst_ff_SDE_84_next_state ;
    wire RoundReg_Inst_ff_SDE_85_next_state ;
    wire RoundReg_Inst_ff_SDE_86_next_state ;
    wire RoundReg_Inst_ff_SDE_87_next_state ;
    wire RoundReg_Inst_ff_SDE_88_next_state ;
    wire RoundReg_Inst_ff_SDE_89_next_state ;
    wire RoundReg_Inst_ff_SDE_90_next_state ;
    wire RoundReg_Inst_ff_SDE_91_next_state ;
    wire RoundReg_Inst_ff_SDE_92_next_state ;
    wire RoundReg_Inst_ff_SDE_93_next_state ;
    wire RoundReg_Inst_ff_SDE_94_next_state ;
    wire RoundReg_Inst_ff_SDE_95_next_state ;
    wire RoundReg_Inst_ff_SDE_96_next_state ;
    wire RoundReg_Inst_ff_SDE_97_next_state ;
    wire RoundReg_Inst_ff_SDE_98_next_state ;
    wire RoundReg_Inst_ff_SDE_99_next_state ;
    wire RoundReg_Inst_ff_SDE_100_next_state ;
    wire RoundReg_Inst_ff_SDE_101_next_state ;
    wire RoundReg_Inst_ff_SDE_102_next_state ;
    wire RoundReg_Inst_ff_SDE_103_next_state ;
    wire RoundReg_Inst_ff_SDE_104_next_state ;
    wire RoundReg_Inst_ff_SDE_105_next_state ;
    wire RoundReg_Inst_ff_SDE_106_next_state ;
    wire RoundReg_Inst_ff_SDE_107_next_state ;
    wire RoundReg_Inst_ff_SDE_108_next_state ;
    wire RoundReg_Inst_ff_SDE_109_next_state ;
    wire RoundReg_Inst_ff_SDE_110_next_state ;
    wire RoundReg_Inst_ff_SDE_111_next_state ;
    wire RoundReg_Inst_ff_SDE_112_next_state ;
    wire RoundReg_Inst_ff_SDE_113_next_state ;
    wire RoundReg_Inst_ff_SDE_114_next_state ;
    wire RoundReg_Inst_ff_SDE_115_next_state ;
    wire RoundReg_Inst_ff_SDE_116_next_state ;
    wire RoundReg_Inst_ff_SDE_117_next_state ;
    wire RoundReg_Inst_ff_SDE_118_next_state ;
    wire RoundReg_Inst_ff_SDE_119_next_state ;
    wire RoundReg_Inst_ff_SDE_120_next_state ;
    wire RoundReg_Inst_ff_SDE_121_next_state ;
    wire RoundReg_Inst_ff_SDE_122_next_state ;
    wire RoundReg_Inst_ff_SDE_123_next_state ;
    wire RoundReg_Inst_ff_SDE_124_next_state ;
    wire RoundReg_Inst_ff_SDE_125_next_state ;
    wire RoundReg_Inst_ff_SDE_126_next_state ;
    wire RoundReg_Inst_ff_SDE_127_next_state ;
    wire SubBytesIns_Inst_Sbox_0_L29 ;
    wire SubBytesIns_Inst_Sbox_0_L28 ;
    wire SubBytesIns_Inst_Sbox_0_L27 ;
    wire SubBytesIns_Inst_Sbox_0_L26 ;
    wire SubBytesIns_Inst_Sbox_0_L25 ;
    wire SubBytesIns_Inst_Sbox_0_L24 ;
    wire SubBytesIns_Inst_Sbox_0_L23 ;
    wire SubBytesIns_Inst_Sbox_0_L22 ;
    wire SubBytesIns_Inst_Sbox_0_L21 ;
    wire SubBytesIns_Inst_Sbox_0_L20 ;
    wire SubBytesIns_Inst_Sbox_0_L19 ;
    wire SubBytesIns_Inst_Sbox_0_L18 ;
    wire SubBytesIns_Inst_Sbox_0_L17 ;
    wire SubBytesIns_Inst_Sbox_0_L16 ;
    wire SubBytesIns_Inst_Sbox_0_L15 ;
    wire SubBytesIns_Inst_Sbox_0_L14 ;
    wire SubBytesIns_Inst_Sbox_0_L13 ;
    wire SubBytesIns_Inst_Sbox_0_L12 ;
    wire SubBytesIns_Inst_Sbox_0_L11 ;
    wire SubBytesIns_Inst_Sbox_0_L10 ;
    wire SubBytesIns_Inst_Sbox_0_L9 ;
    wire SubBytesIns_Inst_Sbox_0_L8 ;
    wire SubBytesIns_Inst_Sbox_0_L7 ;
    wire SubBytesIns_Inst_Sbox_0_L6 ;
    wire SubBytesIns_Inst_Sbox_0_L5 ;
    wire SubBytesIns_Inst_Sbox_0_L4 ;
    wire SubBytesIns_Inst_Sbox_0_L3 ;
    wire SubBytesIns_Inst_Sbox_0_L2 ;
    wire SubBytesIns_Inst_Sbox_0_L1 ;
    wire SubBytesIns_Inst_Sbox_0_L0 ;
    wire SubBytesIns_Inst_Sbox_0_M63 ;
    wire SubBytesIns_Inst_Sbox_0_M62 ;
    wire SubBytesIns_Inst_Sbox_0_M61 ;
    wire SubBytesIns_Inst_Sbox_0_M60 ;
    wire SubBytesIns_Inst_Sbox_0_M59 ;
    wire SubBytesIns_Inst_Sbox_0_M58 ;
    wire SubBytesIns_Inst_Sbox_0_M57 ;
    wire SubBytesIns_Inst_Sbox_0_M56 ;
    wire SubBytesIns_Inst_Sbox_0_M55 ;
    wire SubBytesIns_Inst_Sbox_0_M54 ;
    wire SubBytesIns_Inst_Sbox_0_M53 ;
    wire SubBytesIns_Inst_Sbox_0_M52 ;
    wire SubBytesIns_Inst_Sbox_0_M51 ;
    wire SubBytesIns_Inst_Sbox_0_M50 ;
    wire SubBytesIns_Inst_Sbox_0_M49 ;
    wire SubBytesIns_Inst_Sbox_0_M48 ;
    wire SubBytesIns_Inst_Sbox_0_M47 ;
    wire SubBytesIns_Inst_Sbox_0_M46 ;
    wire SubBytesIns_Inst_Sbox_0_M45 ;
    wire SubBytesIns_Inst_Sbox_0_M44 ;
    wire SubBytesIns_Inst_Sbox_0_M43 ;
    wire SubBytesIns_Inst_Sbox_0_M42 ;
    wire SubBytesIns_Inst_Sbox_0_M41 ;
    wire SubBytesIns_Inst_Sbox_0_M40 ;
    wire SubBytesIns_Inst_Sbox_0_M39 ;
    wire SubBytesIns_Inst_Sbox_0_M38 ;
    wire SubBytesIns_Inst_Sbox_0_M37 ;
    wire SubBytesIns_Inst_Sbox_0_M36 ;
    wire SubBytesIns_Inst_Sbox_0_M35 ;
    wire SubBytesIns_Inst_Sbox_0_M34 ;
    wire SubBytesIns_Inst_Sbox_0_M33 ;
    wire SubBytesIns_Inst_Sbox_0_M32 ;
    wire SubBytesIns_Inst_Sbox_0_M31 ;
    wire SubBytesIns_Inst_Sbox_0_M30 ;
    wire SubBytesIns_Inst_Sbox_0_M29 ;
    wire SubBytesIns_Inst_Sbox_0_M28 ;
    wire SubBytesIns_Inst_Sbox_0_M27 ;
    wire SubBytesIns_Inst_Sbox_0_M26 ;
    wire SubBytesIns_Inst_Sbox_0_M25 ;
    wire SubBytesIns_Inst_Sbox_0_M24 ;
    wire SubBytesIns_Inst_Sbox_0_M23 ;
    wire SubBytesIns_Inst_Sbox_0_M22 ;
    wire SubBytesIns_Inst_Sbox_0_M21 ;
    wire SubBytesIns_Inst_Sbox_0_M20 ;
    wire SubBytesIns_Inst_Sbox_0_M19 ;
    wire SubBytesIns_Inst_Sbox_0_M18 ;
    wire SubBytesIns_Inst_Sbox_0_M17 ;
    wire SubBytesIns_Inst_Sbox_0_M16 ;
    wire SubBytesIns_Inst_Sbox_0_M15 ;
    wire SubBytesIns_Inst_Sbox_0_M14 ;
    wire SubBytesIns_Inst_Sbox_0_M13 ;
    wire SubBytesIns_Inst_Sbox_0_M12 ;
    wire SubBytesIns_Inst_Sbox_0_M11 ;
    wire SubBytesIns_Inst_Sbox_0_M10 ;
    wire SubBytesIns_Inst_Sbox_0_M9 ;
    wire SubBytesIns_Inst_Sbox_0_M8 ;
    wire SubBytesIns_Inst_Sbox_0_M7 ;
    wire SubBytesIns_Inst_Sbox_0_M6 ;
    wire SubBytesIns_Inst_Sbox_0_M5 ;
    wire SubBytesIns_Inst_Sbox_0_M4 ;
    wire SubBytesIns_Inst_Sbox_0_M3 ;
    wire SubBytesIns_Inst_Sbox_0_M2 ;
    wire SubBytesIns_Inst_Sbox_0_M1 ;
    wire SubBytesIns_Inst_Sbox_0_T27 ;
    wire SubBytesIns_Inst_Sbox_0_T26 ;
    wire SubBytesIns_Inst_Sbox_0_T25 ;
    wire SubBytesIns_Inst_Sbox_0_T24 ;
    wire SubBytesIns_Inst_Sbox_0_T23 ;
    wire SubBytesIns_Inst_Sbox_0_T22 ;
    wire SubBytesIns_Inst_Sbox_0_T21 ;
    wire SubBytesIns_Inst_Sbox_0_T20 ;
    wire SubBytesIns_Inst_Sbox_0_T19 ;
    wire SubBytesIns_Inst_Sbox_0_T18 ;
    wire SubBytesIns_Inst_Sbox_0_T17 ;
    wire SubBytesIns_Inst_Sbox_0_T16 ;
    wire SubBytesIns_Inst_Sbox_0_T15 ;
    wire SubBytesIns_Inst_Sbox_0_T14 ;
    wire SubBytesIns_Inst_Sbox_0_T13 ;
    wire SubBytesIns_Inst_Sbox_0_T12 ;
    wire SubBytesIns_Inst_Sbox_0_T11 ;
    wire SubBytesIns_Inst_Sbox_0_T10 ;
    wire SubBytesIns_Inst_Sbox_0_T9 ;
    wire SubBytesIns_Inst_Sbox_0_T8 ;
    wire SubBytesIns_Inst_Sbox_0_T7 ;
    wire SubBytesIns_Inst_Sbox_0_T6 ;
    wire SubBytesIns_Inst_Sbox_0_T5 ;
    wire SubBytesIns_Inst_Sbox_0_T4 ;
    wire SubBytesIns_Inst_Sbox_0_T3 ;
    wire SubBytesIns_Inst_Sbox_0_T2 ;
    wire SubBytesIns_Inst_Sbox_0_T1 ;
    wire SubBytesIns_Inst_Sbox_1_L29 ;
    wire SubBytesIns_Inst_Sbox_1_L28 ;
    wire SubBytesIns_Inst_Sbox_1_L27 ;
    wire SubBytesIns_Inst_Sbox_1_L26 ;
    wire SubBytesIns_Inst_Sbox_1_L25 ;
    wire SubBytesIns_Inst_Sbox_1_L24 ;
    wire SubBytesIns_Inst_Sbox_1_L23 ;
    wire SubBytesIns_Inst_Sbox_1_L22 ;
    wire SubBytesIns_Inst_Sbox_1_L21 ;
    wire SubBytesIns_Inst_Sbox_1_L20 ;
    wire SubBytesIns_Inst_Sbox_1_L19 ;
    wire SubBytesIns_Inst_Sbox_1_L18 ;
    wire SubBytesIns_Inst_Sbox_1_L17 ;
    wire SubBytesIns_Inst_Sbox_1_L16 ;
    wire SubBytesIns_Inst_Sbox_1_L15 ;
    wire SubBytesIns_Inst_Sbox_1_L14 ;
    wire SubBytesIns_Inst_Sbox_1_L13 ;
    wire SubBytesIns_Inst_Sbox_1_L12 ;
    wire SubBytesIns_Inst_Sbox_1_L11 ;
    wire SubBytesIns_Inst_Sbox_1_L10 ;
    wire SubBytesIns_Inst_Sbox_1_L9 ;
    wire SubBytesIns_Inst_Sbox_1_L8 ;
    wire SubBytesIns_Inst_Sbox_1_L7 ;
    wire SubBytesIns_Inst_Sbox_1_L6 ;
    wire SubBytesIns_Inst_Sbox_1_L5 ;
    wire SubBytesIns_Inst_Sbox_1_L4 ;
    wire SubBytesIns_Inst_Sbox_1_L3 ;
    wire SubBytesIns_Inst_Sbox_1_L2 ;
    wire SubBytesIns_Inst_Sbox_1_L1 ;
    wire SubBytesIns_Inst_Sbox_1_L0 ;
    wire SubBytesIns_Inst_Sbox_1_M63 ;
    wire SubBytesIns_Inst_Sbox_1_M62 ;
    wire SubBytesIns_Inst_Sbox_1_M61 ;
    wire SubBytesIns_Inst_Sbox_1_M60 ;
    wire SubBytesIns_Inst_Sbox_1_M59 ;
    wire SubBytesIns_Inst_Sbox_1_M58 ;
    wire SubBytesIns_Inst_Sbox_1_M57 ;
    wire SubBytesIns_Inst_Sbox_1_M56 ;
    wire SubBytesIns_Inst_Sbox_1_M55 ;
    wire SubBytesIns_Inst_Sbox_1_M54 ;
    wire SubBytesIns_Inst_Sbox_1_M53 ;
    wire SubBytesIns_Inst_Sbox_1_M52 ;
    wire SubBytesIns_Inst_Sbox_1_M51 ;
    wire SubBytesIns_Inst_Sbox_1_M50 ;
    wire SubBytesIns_Inst_Sbox_1_M49 ;
    wire SubBytesIns_Inst_Sbox_1_M48 ;
    wire SubBytesIns_Inst_Sbox_1_M47 ;
    wire SubBytesIns_Inst_Sbox_1_M46 ;
    wire SubBytesIns_Inst_Sbox_1_M45 ;
    wire SubBytesIns_Inst_Sbox_1_M44 ;
    wire SubBytesIns_Inst_Sbox_1_M43 ;
    wire SubBytesIns_Inst_Sbox_1_M42 ;
    wire SubBytesIns_Inst_Sbox_1_M41 ;
    wire SubBytesIns_Inst_Sbox_1_M40 ;
    wire SubBytesIns_Inst_Sbox_1_M39 ;
    wire SubBytesIns_Inst_Sbox_1_M38 ;
    wire SubBytesIns_Inst_Sbox_1_M37 ;
    wire SubBytesIns_Inst_Sbox_1_M36 ;
    wire SubBytesIns_Inst_Sbox_1_M35 ;
    wire SubBytesIns_Inst_Sbox_1_M34 ;
    wire SubBytesIns_Inst_Sbox_1_M33 ;
    wire SubBytesIns_Inst_Sbox_1_M32 ;
    wire SubBytesIns_Inst_Sbox_1_M31 ;
    wire SubBytesIns_Inst_Sbox_1_M30 ;
    wire SubBytesIns_Inst_Sbox_1_M29 ;
    wire SubBytesIns_Inst_Sbox_1_M28 ;
    wire SubBytesIns_Inst_Sbox_1_M27 ;
    wire SubBytesIns_Inst_Sbox_1_M26 ;
    wire SubBytesIns_Inst_Sbox_1_M25 ;
    wire SubBytesIns_Inst_Sbox_1_M24 ;
    wire SubBytesIns_Inst_Sbox_1_M23 ;
    wire SubBytesIns_Inst_Sbox_1_M22 ;
    wire SubBytesIns_Inst_Sbox_1_M21 ;
    wire SubBytesIns_Inst_Sbox_1_M20 ;
    wire SubBytesIns_Inst_Sbox_1_M19 ;
    wire SubBytesIns_Inst_Sbox_1_M18 ;
    wire SubBytesIns_Inst_Sbox_1_M17 ;
    wire SubBytesIns_Inst_Sbox_1_M16 ;
    wire SubBytesIns_Inst_Sbox_1_M15 ;
    wire SubBytesIns_Inst_Sbox_1_M14 ;
    wire SubBytesIns_Inst_Sbox_1_M13 ;
    wire SubBytesIns_Inst_Sbox_1_M12 ;
    wire SubBytesIns_Inst_Sbox_1_M11 ;
    wire SubBytesIns_Inst_Sbox_1_M10 ;
    wire SubBytesIns_Inst_Sbox_1_M9 ;
    wire SubBytesIns_Inst_Sbox_1_M8 ;
    wire SubBytesIns_Inst_Sbox_1_M7 ;
    wire SubBytesIns_Inst_Sbox_1_M6 ;
    wire SubBytesIns_Inst_Sbox_1_M5 ;
    wire SubBytesIns_Inst_Sbox_1_M4 ;
    wire SubBytesIns_Inst_Sbox_1_M3 ;
    wire SubBytesIns_Inst_Sbox_1_M2 ;
    wire SubBytesIns_Inst_Sbox_1_M1 ;
    wire SubBytesIns_Inst_Sbox_1_T27 ;
    wire SubBytesIns_Inst_Sbox_1_T26 ;
    wire SubBytesIns_Inst_Sbox_1_T25 ;
    wire SubBytesIns_Inst_Sbox_1_T24 ;
    wire SubBytesIns_Inst_Sbox_1_T23 ;
    wire SubBytesIns_Inst_Sbox_1_T22 ;
    wire SubBytesIns_Inst_Sbox_1_T21 ;
    wire SubBytesIns_Inst_Sbox_1_T20 ;
    wire SubBytesIns_Inst_Sbox_1_T19 ;
    wire SubBytesIns_Inst_Sbox_1_T18 ;
    wire SubBytesIns_Inst_Sbox_1_T17 ;
    wire SubBytesIns_Inst_Sbox_1_T16 ;
    wire SubBytesIns_Inst_Sbox_1_T15 ;
    wire SubBytesIns_Inst_Sbox_1_T14 ;
    wire SubBytesIns_Inst_Sbox_1_T13 ;
    wire SubBytesIns_Inst_Sbox_1_T12 ;
    wire SubBytesIns_Inst_Sbox_1_T11 ;
    wire SubBytesIns_Inst_Sbox_1_T10 ;
    wire SubBytesIns_Inst_Sbox_1_T9 ;
    wire SubBytesIns_Inst_Sbox_1_T8 ;
    wire SubBytesIns_Inst_Sbox_1_T7 ;
    wire SubBytesIns_Inst_Sbox_1_T6 ;
    wire SubBytesIns_Inst_Sbox_1_T5 ;
    wire SubBytesIns_Inst_Sbox_1_T4 ;
    wire SubBytesIns_Inst_Sbox_1_T3 ;
    wire SubBytesIns_Inst_Sbox_1_T2 ;
    wire SubBytesIns_Inst_Sbox_1_T1 ;
    wire SubBytesIns_Inst_Sbox_2_L29 ;
    wire SubBytesIns_Inst_Sbox_2_L28 ;
    wire SubBytesIns_Inst_Sbox_2_L27 ;
    wire SubBytesIns_Inst_Sbox_2_L26 ;
    wire SubBytesIns_Inst_Sbox_2_L25 ;
    wire SubBytesIns_Inst_Sbox_2_L24 ;
    wire SubBytesIns_Inst_Sbox_2_L23 ;
    wire SubBytesIns_Inst_Sbox_2_L22 ;
    wire SubBytesIns_Inst_Sbox_2_L21 ;
    wire SubBytesIns_Inst_Sbox_2_L20 ;
    wire SubBytesIns_Inst_Sbox_2_L19 ;
    wire SubBytesIns_Inst_Sbox_2_L18 ;
    wire SubBytesIns_Inst_Sbox_2_L17 ;
    wire SubBytesIns_Inst_Sbox_2_L16 ;
    wire SubBytesIns_Inst_Sbox_2_L15 ;
    wire SubBytesIns_Inst_Sbox_2_L14 ;
    wire SubBytesIns_Inst_Sbox_2_L13 ;
    wire SubBytesIns_Inst_Sbox_2_L12 ;
    wire SubBytesIns_Inst_Sbox_2_L11 ;
    wire SubBytesIns_Inst_Sbox_2_L10 ;
    wire SubBytesIns_Inst_Sbox_2_L9 ;
    wire SubBytesIns_Inst_Sbox_2_L8 ;
    wire SubBytesIns_Inst_Sbox_2_L7 ;
    wire SubBytesIns_Inst_Sbox_2_L6 ;
    wire SubBytesIns_Inst_Sbox_2_L5 ;
    wire SubBytesIns_Inst_Sbox_2_L4 ;
    wire SubBytesIns_Inst_Sbox_2_L3 ;
    wire SubBytesIns_Inst_Sbox_2_L2 ;
    wire SubBytesIns_Inst_Sbox_2_L1 ;
    wire SubBytesIns_Inst_Sbox_2_L0 ;
    wire SubBytesIns_Inst_Sbox_2_M63 ;
    wire SubBytesIns_Inst_Sbox_2_M62 ;
    wire SubBytesIns_Inst_Sbox_2_M61 ;
    wire SubBytesIns_Inst_Sbox_2_M60 ;
    wire SubBytesIns_Inst_Sbox_2_M59 ;
    wire SubBytesIns_Inst_Sbox_2_M58 ;
    wire SubBytesIns_Inst_Sbox_2_M57 ;
    wire SubBytesIns_Inst_Sbox_2_M56 ;
    wire SubBytesIns_Inst_Sbox_2_M55 ;
    wire SubBytesIns_Inst_Sbox_2_M54 ;
    wire SubBytesIns_Inst_Sbox_2_M53 ;
    wire SubBytesIns_Inst_Sbox_2_M52 ;
    wire SubBytesIns_Inst_Sbox_2_M51 ;
    wire SubBytesIns_Inst_Sbox_2_M50 ;
    wire SubBytesIns_Inst_Sbox_2_M49 ;
    wire SubBytesIns_Inst_Sbox_2_M48 ;
    wire SubBytesIns_Inst_Sbox_2_M47 ;
    wire SubBytesIns_Inst_Sbox_2_M46 ;
    wire SubBytesIns_Inst_Sbox_2_M45 ;
    wire SubBytesIns_Inst_Sbox_2_M44 ;
    wire SubBytesIns_Inst_Sbox_2_M43 ;
    wire SubBytesIns_Inst_Sbox_2_M42 ;
    wire SubBytesIns_Inst_Sbox_2_M41 ;
    wire SubBytesIns_Inst_Sbox_2_M40 ;
    wire SubBytesIns_Inst_Sbox_2_M39 ;
    wire SubBytesIns_Inst_Sbox_2_M38 ;
    wire SubBytesIns_Inst_Sbox_2_M37 ;
    wire SubBytesIns_Inst_Sbox_2_M36 ;
    wire SubBytesIns_Inst_Sbox_2_M35 ;
    wire SubBytesIns_Inst_Sbox_2_M34 ;
    wire SubBytesIns_Inst_Sbox_2_M33 ;
    wire SubBytesIns_Inst_Sbox_2_M32 ;
    wire SubBytesIns_Inst_Sbox_2_M31 ;
    wire SubBytesIns_Inst_Sbox_2_M30 ;
    wire SubBytesIns_Inst_Sbox_2_M29 ;
    wire SubBytesIns_Inst_Sbox_2_M28 ;
    wire SubBytesIns_Inst_Sbox_2_M27 ;
    wire SubBytesIns_Inst_Sbox_2_M26 ;
    wire SubBytesIns_Inst_Sbox_2_M25 ;
    wire SubBytesIns_Inst_Sbox_2_M24 ;
    wire SubBytesIns_Inst_Sbox_2_M23 ;
    wire SubBytesIns_Inst_Sbox_2_M22 ;
    wire SubBytesIns_Inst_Sbox_2_M21 ;
    wire SubBytesIns_Inst_Sbox_2_M20 ;
    wire SubBytesIns_Inst_Sbox_2_M19 ;
    wire SubBytesIns_Inst_Sbox_2_M18 ;
    wire SubBytesIns_Inst_Sbox_2_M17 ;
    wire SubBytesIns_Inst_Sbox_2_M16 ;
    wire SubBytesIns_Inst_Sbox_2_M15 ;
    wire SubBytesIns_Inst_Sbox_2_M14 ;
    wire SubBytesIns_Inst_Sbox_2_M13 ;
    wire SubBytesIns_Inst_Sbox_2_M12 ;
    wire SubBytesIns_Inst_Sbox_2_M11 ;
    wire SubBytesIns_Inst_Sbox_2_M10 ;
    wire SubBytesIns_Inst_Sbox_2_M9 ;
    wire SubBytesIns_Inst_Sbox_2_M8 ;
    wire SubBytesIns_Inst_Sbox_2_M7 ;
    wire SubBytesIns_Inst_Sbox_2_M6 ;
    wire SubBytesIns_Inst_Sbox_2_M5 ;
    wire SubBytesIns_Inst_Sbox_2_M4 ;
    wire SubBytesIns_Inst_Sbox_2_M3 ;
    wire SubBytesIns_Inst_Sbox_2_M2 ;
    wire SubBytesIns_Inst_Sbox_2_M1 ;
    wire SubBytesIns_Inst_Sbox_2_T27 ;
    wire SubBytesIns_Inst_Sbox_2_T26 ;
    wire SubBytesIns_Inst_Sbox_2_T25 ;
    wire SubBytesIns_Inst_Sbox_2_T24 ;
    wire SubBytesIns_Inst_Sbox_2_T23 ;
    wire SubBytesIns_Inst_Sbox_2_T22 ;
    wire SubBytesIns_Inst_Sbox_2_T21 ;
    wire SubBytesIns_Inst_Sbox_2_T20 ;
    wire SubBytesIns_Inst_Sbox_2_T19 ;
    wire SubBytesIns_Inst_Sbox_2_T18 ;
    wire SubBytesIns_Inst_Sbox_2_T17 ;
    wire SubBytesIns_Inst_Sbox_2_T16 ;
    wire SubBytesIns_Inst_Sbox_2_T15 ;
    wire SubBytesIns_Inst_Sbox_2_T14 ;
    wire SubBytesIns_Inst_Sbox_2_T13 ;
    wire SubBytesIns_Inst_Sbox_2_T12 ;
    wire SubBytesIns_Inst_Sbox_2_T11 ;
    wire SubBytesIns_Inst_Sbox_2_T10 ;
    wire SubBytesIns_Inst_Sbox_2_T9 ;
    wire SubBytesIns_Inst_Sbox_2_T8 ;
    wire SubBytesIns_Inst_Sbox_2_T7 ;
    wire SubBytesIns_Inst_Sbox_2_T6 ;
    wire SubBytesIns_Inst_Sbox_2_T5 ;
    wire SubBytesIns_Inst_Sbox_2_T4 ;
    wire SubBytesIns_Inst_Sbox_2_T3 ;
    wire SubBytesIns_Inst_Sbox_2_T2 ;
    wire SubBytesIns_Inst_Sbox_2_T1 ;
    wire SubBytesIns_Inst_Sbox_3_L29 ;
    wire SubBytesIns_Inst_Sbox_3_L28 ;
    wire SubBytesIns_Inst_Sbox_3_L27 ;
    wire SubBytesIns_Inst_Sbox_3_L26 ;
    wire SubBytesIns_Inst_Sbox_3_L25 ;
    wire SubBytesIns_Inst_Sbox_3_L24 ;
    wire SubBytesIns_Inst_Sbox_3_L23 ;
    wire SubBytesIns_Inst_Sbox_3_L22 ;
    wire SubBytesIns_Inst_Sbox_3_L21 ;
    wire SubBytesIns_Inst_Sbox_3_L20 ;
    wire SubBytesIns_Inst_Sbox_3_L19 ;
    wire SubBytesIns_Inst_Sbox_3_L18 ;
    wire SubBytesIns_Inst_Sbox_3_L17 ;
    wire SubBytesIns_Inst_Sbox_3_L16 ;
    wire SubBytesIns_Inst_Sbox_3_L15 ;
    wire SubBytesIns_Inst_Sbox_3_L14 ;
    wire SubBytesIns_Inst_Sbox_3_L13 ;
    wire SubBytesIns_Inst_Sbox_3_L12 ;
    wire SubBytesIns_Inst_Sbox_3_L11 ;
    wire SubBytesIns_Inst_Sbox_3_L10 ;
    wire SubBytesIns_Inst_Sbox_3_L9 ;
    wire SubBytesIns_Inst_Sbox_3_L8 ;
    wire SubBytesIns_Inst_Sbox_3_L7 ;
    wire SubBytesIns_Inst_Sbox_3_L6 ;
    wire SubBytesIns_Inst_Sbox_3_L5 ;
    wire SubBytesIns_Inst_Sbox_3_L4 ;
    wire SubBytesIns_Inst_Sbox_3_L3 ;
    wire SubBytesIns_Inst_Sbox_3_L2 ;
    wire SubBytesIns_Inst_Sbox_3_L1 ;
    wire SubBytesIns_Inst_Sbox_3_L0 ;
    wire SubBytesIns_Inst_Sbox_3_M63 ;
    wire SubBytesIns_Inst_Sbox_3_M62 ;
    wire SubBytesIns_Inst_Sbox_3_M61 ;
    wire SubBytesIns_Inst_Sbox_3_M60 ;
    wire SubBytesIns_Inst_Sbox_3_M59 ;
    wire SubBytesIns_Inst_Sbox_3_M58 ;
    wire SubBytesIns_Inst_Sbox_3_M57 ;
    wire SubBytesIns_Inst_Sbox_3_M56 ;
    wire SubBytesIns_Inst_Sbox_3_M55 ;
    wire SubBytesIns_Inst_Sbox_3_M54 ;
    wire SubBytesIns_Inst_Sbox_3_M53 ;
    wire SubBytesIns_Inst_Sbox_3_M52 ;
    wire SubBytesIns_Inst_Sbox_3_M51 ;
    wire SubBytesIns_Inst_Sbox_3_M50 ;
    wire SubBytesIns_Inst_Sbox_3_M49 ;
    wire SubBytesIns_Inst_Sbox_3_M48 ;
    wire SubBytesIns_Inst_Sbox_3_M47 ;
    wire SubBytesIns_Inst_Sbox_3_M46 ;
    wire SubBytesIns_Inst_Sbox_3_M45 ;
    wire SubBytesIns_Inst_Sbox_3_M44 ;
    wire SubBytesIns_Inst_Sbox_3_M43 ;
    wire SubBytesIns_Inst_Sbox_3_M42 ;
    wire SubBytesIns_Inst_Sbox_3_M41 ;
    wire SubBytesIns_Inst_Sbox_3_M40 ;
    wire SubBytesIns_Inst_Sbox_3_M39 ;
    wire SubBytesIns_Inst_Sbox_3_M38 ;
    wire SubBytesIns_Inst_Sbox_3_M37 ;
    wire SubBytesIns_Inst_Sbox_3_M36 ;
    wire SubBytesIns_Inst_Sbox_3_M35 ;
    wire SubBytesIns_Inst_Sbox_3_M34 ;
    wire SubBytesIns_Inst_Sbox_3_M33 ;
    wire SubBytesIns_Inst_Sbox_3_M32 ;
    wire SubBytesIns_Inst_Sbox_3_M31 ;
    wire SubBytesIns_Inst_Sbox_3_M30 ;
    wire SubBytesIns_Inst_Sbox_3_M29 ;
    wire SubBytesIns_Inst_Sbox_3_M28 ;
    wire SubBytesIns_Inst_Sbox_3_M27 ;
    wire SubBytesIns_Inst_Sbox_3_M26 ;
    wire SubBytesIns_Inst_Sbox_3_M25 ;
    wire SubBytesIns_Inst_Sbox_3_M24 ;
    wire SubBytesIns_Inst_Sbox_3_M23 ;
    wire SubBytesIns_Inst_Sbox_3_M22 ;
    wire SubBytesIns_Inst_Sbox_3_M21 ;
    wire SubBytesIns_Inst_Sbox_3_M20 ;
    wire SubBytesIns_Inst_Sbox_3_M19 ;
    wire SubBytesIns_Inst_Sbox_3_M18 ;
    wire SubBytesIns_Inst_Sbox_3_M17 ;
    wire SubBytesIns_Inst_Sbox_3_M16 ;
    wire SubBytesIns_Inst_Sbox_3_M15 ;
    wire SubBytesIns_Inst_Sbox_3_M14 ;
    wire SubBytesIns_Inst_Sbox_3_M13 ;
    wire SubBytesIns_Inst_Sbox_3_M12 ;
    wire SubBytesIns_Inst_Sbox_3_M11 ;
    wire SubBytesIns_Inst_Sbox_3_M10 ;
    wire SubBytesIns_Inst_Sbox_3_M9 ;
    wire SubBytesIns_Inst_Sbox_3_M8 ;
    wire SubBytesIns_Inst_Sbox_3_M7 ;
    wire SubBytesIns_Inst_Sbox_3_M6 ;
    wire SubBytesIns_Inst_Sbox_3_M5 ;
    wire SubBytesIns_Inst_Sbox_3_M4 ;
    wire SubBytesIns_Inst_Sbox_3_M3 ;
    wire SubBytesIns_Inst_Sbox_3_M2 ;
    wire SubBytesIns_Inst_Sbox_3_M1 ;
    wire SubBytesIns_Inst_Sbox_3_T27 ;
    wire SubBytesIns_Inst_Sbox_3_T26 ;
    wire SubBytesIns_Inst_Sbox_3_T25 ;
    wire SubBytesIns_Inst_Sbox_3_T24 ;
    wire SubBytesIns_Inst_Sbox_3_T23 ;
    wire SubBytesIns_Inst_Sbox_3_T22 ;
    wire SubBytesIns_Inst_Sbox_3_T21 ;
    wire SubBytesIns_Inst_Sbox_3_T20 ;
    wire SubBytesIns_Inst_Sbox_3_T19 ;
    wire SubBytesIns_Inst_Sbox_3_T18 ;
    wire SubBytesIns_Inst_Sbox_3_T17 ;
    wire SubBytesIns_Inst_Sbox_3_T16 ;
    wire SubBytesIns_Inst_Sbox_3_T15 ;
    wire SubBytesIns_Inst_Sbox_3_T14 ;
    wire SubBytesIns_Inst_Sbox_3_T13 ;
    wire SubBytesIns_Inst_Sbox_3_T12 ;
    wire SubBytesIns_Inst_Sbox_3_T11 ;
    wire SubBytesIns_Inst_Sbox_3_T10 ;
    wire SubBytesIns_Inst_Sbox_3_T9 ;
    wire SubBytesIns_Inst_Sbox_3_T8 ;
    wire SubBytesIns_Inst_Sbox_3_T7 ;
    wire SubBytesIns_Inst_Sbox_3_T6 ;
    wire SubBytesIns_Inst_Sbox_3_T5 ;
    wire SubBytesIns_Inst_Sbox_3_T4 ;
    wire SubBytesIns_Inst_Sbox_3_T3 ;
    wire SubBytesIns_Inst_Sbox_3_T2 ;
    wire SubBytesIns_Inst_Sbox_3_T1 ;
    wire SubBytesIns_Inst_Sbox_4_L29 ;
    wire SubBytesIns_Inst_Sbox_4_L28 ;
    wire SubBytesIns_Inst_Sbox_4_L27 ;
    wire SubBytesIns_Inst_Sbox_4_L26 ;
    wire SubBytesIns_Inst_Sbox_4_L25 ;
    wire SubBytesIns_Inst_Sbox_4_L24 ;
    wire SubBytesIns_Inst_Sbox_4_L23 ;
    wire SubBytesIns_Inst_Sbox_4_L22 ;
    wire SubBytesIns_Inst_Sbox_4_L21 ;
    wire SubBytesIns_Inst_Sbox_4_L20 ;
    wire SubBytesIns_Inst_Sbox_4_L19 ;
    wire SubBytesIns_Inst_Sbox_4_L18 ;
    wire SubBytesIns_Inst_Sbox_4_L17 ;
    wire SubBytesIns_Inst_Sbox_4_L16 ;
    wire SubBytesIns_Inst_Sbox_4_L15 ;
    wire SubBytesIns_Inst_Sbox_4_L14 ;
    wire SubBytesIns_Inst_Sbox_4_L13 ;
    wire SubBytesIns_Inst_Sbox_4_L12 ;
    wire SubBytesIns_Inst_Sbox_4_L11 ;
    wire SubBytesIns_Inst_Sbox_4_L10 ;
    wire SubBytesIns_Inst_Sbox_4_L9 ;
    wire SubBytesIns_Inst_Sbox_4_L8 ;
    wire SubBytesIns_Inst_Sbox_4_L7 ;
    wire SubBytesIns_Inst_Sbox_4_L6 ;
    wire SubBytesIns_Inst_Sbox_4_L5 ;
    wire SubBytesIns_Inst_Sbox_4_L4 ;
    wire SubBytesIns_Inst_Sbox_4_L3 ;
    wire SubBytesIns_Inst_Sbox_4_L2 ;
    wire SubBytesIns_Inst_Sbox_4_L1 ;
    wire SubBytesIns_Inst_Sbox_4_L0 ;
    wire SubBytesIns_Inst_Sbox_4_M63 ;
    wire SubBytesIns_Inst_Sbox_4_M62 ;
    wire SubBytesIns_Inst_Sbox_4_M61 ;
    wire SubBytesIns_Inst_Sbox_4_M60 ;
    wire SubBytesIns_Inst_Sbox_4_M59 ;
    wire SubBytesIns_Inst_Sbox_4_M58 ;
    wire SubBytesIns_Inst_Sbox_4_M57 ;
    wire SubBytesIns_Inst_Sbox_4_M56 ;
    wire SubBytesIns_Inst_Sbox_4_M55 ;
    wire SubBytesIns_Inst_Sbox_4_M54 ;
    wire SubBytesIns_Inst_Sbox_4_M53 ;
    wire SubBytesIns_Inst_Sbox_4_M52 ;
    wire SubBytesIns_Inst_Sbox_4_M51 ;
    wire SubBytesIns_Inst_Sbox_4_M50 ;
    wire SubBytesIns_Inst_Sbox_4_M49 ;
    wire SubBytesIns_Inst_Sbox_4_M48 ;
    wire SubBytesIns_Inst_Sbox_4_M47 ;
    wire SubBytesIns_Inst_Sbox_4_M46 ;
    wire SubBytesIns_Inst_Sbox_4_M45 ;
    wire SubBytesIns_Inst_Sbox_4_M44 ;
    wire SubBytesIns_Inst_Sbox_4_M43 ;
    wire SubBytesIns_Inst_Sbox_4_M42 ;
    wire SubBytesIns_Inst_Sbox_4_M41 ;
    wire SubBytesIns_Inst_Sbox_4_M40 ;
    wire SubBytesIns_Inst_Sbox_4_M39 ;
    wire SubBytesIns_Inst_Sbox_4_M38 ;
    wire SubBytesIns_Inst_Sbox_4_M37 ;
    wire SubBytesIns_Inst_Sbox_4_M36 ;
    wire SubBytesIns_Inst_Sbox_4_M35 ;
    wire SubBytesIns_Inst_Sbox_4_M34 ;
    wire SubBytesIns_Inst_Sbox_4_M33 ;
    wire SubBytesIns_Inst_Sbox_4_M32 ;
    wire SubBytesIns_Inst_Sbox_4_M31 ;
    wire SubBytesIns_Inst_Sbox_4_M30 ;
    wire SubBytesIns_Inst_Sbox_4_M29 ;
    wire SubBytesIns_Inst_Sbox_4_M28 ;
    wire SubBytesIns_Inst_Sbox_4_M27 ;
    wire SubBytesIns_Inst_Sbox_4_M26 ;
    wire SubBytesIns_Inst_Sbox_4_M25 ;
    wire SubBytesIns_Inst_Sbox_4_M24 ;
    wire SubBytesIns_Inst_Sbox_4_M23 ;
    wire SubBytesIns_Inst_Sbox_4_M22 ;
    wire SubBytesIns_Inst_Sbox_4_M21 ;
    wire SubBytesIns_Inst_Sbox_4_M20 ;
    wire SubBytesIns_Inst_Sbox_4_M19 ;
    wire SubBytesIns_Inst_Sbox_4_M18 ;
    wire SubBytesIns_Inst_Sbox_4_M17 ;
    wire SubBytesIns_Inst_Sbox_4_M16 ;
    wire SubBytesIns_Inst_Sbox_4_M15 ;
    wire SubBytesIns_Inst_Sbox_4_M14 ;
    wire SubBytesIns_Inst_Sbox_4_M13 ;
    wire SubBytesIns_Inst_Sbox_4_M12 ;
    wire SubBytesIns_Inst_Sbox_4_M11 ;
    wire SubBytesIns_Inst_Sbox_4_M10 ;
    wire SubBytesIns_Inst_Sbox_4_M9 ;
    wire SubBytesIns_Inst_Sbox_4_M8 ;
    wire SubBytesIns_Inst_Sbox_4_M7 ;
    wire SubBytesIns_Inst_Sbox_4_M6 ;
    wire SubBytesIns_Inst_Sbox_4_M5 ;
    wire SubBytesIns_Inst_Sbox_4_M4 ;
    wire SubBytesIns_Inst_Sbox_4_M3 ;
    wire SubBytesIns_Inst_Sbox_4_M2 ;
    wire SubBytesIns_Inst_Sbox_4_M1 ;
    wire SubBytesIns_Inst_Sbox_4_T27 ;
    wire SubBytesIns_Inst_Sbox_4_T26 ;
    wire SubBytesIns_Inst_Sbox_4_T25 ;
    wire SubBytesIns_Inst_Sbox_4_T24 ;
    wire SubBytesIns_Inst_Sbox_4_T23 ;
    wire SubBytesIns_Inst_Sbox_4_T22 ;
    wire SubBytesIns_Inst_Sbox_4_T21 ;
    wire SubBytesIns_Inst_Sbox_4_T20 ;
    wire SubBytesIns_Inst_Sbox_4_T19 ;
    wire SubBytesIns_Inst_Sbox_4_T18 ;
    wire SubBytesIns_Inst_Sbox_4_T17 ;
    wire SubBytesIns_Inst_Sbox_4_T16 ;
    wire SubBytesIns_Inst_Sbox_4_T15 ;
    wire SubBytesIns_Inst_Sbox_4_T14 ;
    wire SubBytesIns_Inst_Sbox_4_T13 ;
    wire SubBytesIns_Inst_Sbox_4_T12 ;
    wire SubBytesIns_Inst_Sbox_4_T11 ;
    wire SubBytesIns_Inst_Sbox_4_T10 ;
    wire SubBytesIns_Inst_Sbox_4_T9 ;
    wire SubBytesIns_Inst_Sbox_4_T8 ;
    wire SubBytesIns_Inst_Sbox_4_T7 ;
    wire SubBytesIns_Inst_Sbox_4_T6 ;
    wire SubBytesIns_Inst_Sbox_4_T5 ;
    wire SubBytesIns_Inst_Sbox_4_T4 ;
    wire SubBytesIns_Inst_Sbox_4_T3 ;
    wire SubBytesIns_Inst_Sbox_4_T2 ;
    wire SubBytesIns_Inst_Sbox_4_T1 ;
    wire SubBytesIns_Inst_Sbox_5_L29 ;
    wire SubBytesIns_Inst_Sbox_5_L28 ;
    wire SubBytesIns_Inst_Sbox_5_L27 ;
    wire SubBytesIns_Inst_Sbox_5_L26 ;
    wire SubBytesIns_Inst_Sbox_5_L25 ;
    wire SubBytesIns_Inst_Sbox_5_L24 ;
    wire SubBytesIns_Inst_Sbox_5_L23 ;
    wire SubBytesIns_Inst_Sbox_5_L22 ;
    wire SubBytesIns_Inst_Sbox_5_L21 ;
    wire SubBytesIns_Inst_Sbox_5_L20 ;
    wire SubBytesIns_Inst_Sbox_5_L19 ;
    wire SubBytesIns_Inst_Sbox_5_L18 ;
    wire SubBytesIns_Inst_Sbox_5_L17 ;
    wire SubBytesIns_Inst_Sbox_5_L16 ;
    wire SubBytesIns_Inst_Sbox_5_L15 ;
    wire SubBytesIns_Inst_Sbox_5_L14 ;
    wire SubBytesIns_Inst_Sbox_5_L13 ;
    wire SubBytesIns_Inst_Sbox_5_L12 ;
    wire SubBytesIns_Inst_Sbox_5_L11 ;
    wire SubBytesIns_Inst_Sbox_5_L10 ;
    wire SubBytesIns_Inst_Sbox_5_L9 ;
    wire SubBytesIns_Inst_Sbox_5_L8 ;
    wire SubBytesIns_Inst_Sbox_5_L7 ;
    wire SubBytesIns_Inst_Sbox_5_L6 ;
    wire SubBytesIns_Inst_Sbox_5_L5 ;
    wire SubBytesIns_Inst_Sbox_5_L4 ;
    wire SubBytesIns_Inst_Sbox_5_L3 ;
    wire SubBytesIns_Inst_Sbox_5_L2 ;
    wire SubBytesIns_Inst_Sbox_5_L1 ;
    wire SubBytesIns_Inst_Sbox_5_L0 ;
    wire SubBytesIns_Inst_Sbox_5_M63 ;
    wire SubBytesIns_Inst_Sbox_5_M62 ;
    wire SubBytesIns_Inst_Sbox_5_M61 ;
    wire SubBytesIns_Inst_Sbox_5_M60 ;
    wire SubBytesIns_Inst_Sbox_5_M59 ;
    wire SubBytesIns_Inst_Sbox_5_M58 ;
    wire SubBytesIns_Inst_Sbox_5_M57 ;
    wire SubBytesIns_Inst_Sbox_5_M56 ;
    wire SubBytesIns_Inst_Sbox_5_M55 ;
    wire SubBytesIns_Inst_Sbox_5_M54 ;
    wire SubBytesIns_Inst_Sbox_5_M53 ;
    wire SubBytesIns_Inst_Sbox_5_M52 ;
    wire SubBytesIns_Inst_Sbox_5_M51 ;
    wire SubBytesIns_Inst_Sbox_5_M50 ;
    wire SubBytesIns_Inst_Sbox_5_M49 ;
    wire SubBytesIns_Inst_Sbox_5_M48 ;
    wire SubBytesIns_Inst_Sbox_5_M47 ;
    wire SubBytesIns_Inst_Sbox_5_M46 ;
    wire SubBytesIns_Inst_Sbox_5_M45 ;
    wire SubBytesIns_Inst_Sbox_5_M44 ;
    wire SubBytesIns_Inst_Sbox_5_M43 ;
    wire SubBytesIns_Inst_Sbox_5_M42 ;
    wire SubBytesIns_Inst_Sbox_5_M41 ;
    wire SubBytesIns_Inst_Sbox_5_M40 ;
    wire SubBytesIns_Inst_Sbox_5_M39 ;
    wire SubBytesIns_Inst_Sbox_5_M38 ;
    wire SubBytesIns_Inst_Sbox_5_M37 ;
    wire SubBytesIns_Inst_Sbox_5_M36 ;
    wire SubBytesIns_Inst_Sbox_5_M35 ;
    wire SubBytesIns_Inst_Sbox_5_M34 ;
    wire SubBytesIns_Inst_Sbox_5_M33 ;
    wire SubBytesIns_Inst_Sbox_5_M32 ;
    wire SubBytesIns_Inst_Sbox_5_M31 ;
    wire SubBytesIns_Inst_Sbox_5_M30 ;
    wire SubBytesIns_Inst_Sbox_5_M29 ;
    wire SubBytesIns_Inst_Sbox_5_M28 ;
    wire SubBytesIns_Inst_Sbox_5_M27 ;
    wire SubBytesIns_Inst_Sbox_5_M26 ;
    wire SubBytesIns_Inst_Sbox_5_M25 ;
    wire SubBytesIns_Inst_Sbox_5_M24 ;
    wire SubBytesIns_Inst_Sbox_5_M23 ;
    wire SubBytesIns_Inst_Sbox_5_M22 ;
    wire SubBytesIns_Inst_Sbox_5_M21 ;
    wire SubBytesIns_Inst_Sbox_5_M20 ;
    wire SubBytesIns_Inst_Sbox_5_M19 ;
    wire SubBytesIns_Inst_Sbox_5_M18 ;
    wire SubBytesIns_Inst_Sbox_5_M17 ;
    wire SubBytesIns_Inst_Sbox_5_M16 ;
    wire SubBytesIns_Inst_Sbox_5_M15 ;
    wire SubBytesIns_Inst_Sbox_5_M14 ;
    wire SubBytesIns_Inst_Sbox_5_M13 ;
    wire SubBytesIns_Inst_Sbox_5_M12 ;
    wire SubBytesIns_Inst_Sbox_5_M11 ;
    wire SubBytesIns_Inst_Sbox_5_M10 ;
    wire SubBytesIns_Inst_Sbox_5_M9 ;
    wire SubBytesIns_Inst_Sbox_5_M8 ;
    wire SubBytesIns_Inst_Sbox_5_M7 ;
    wire SubBytesIns_Inst_Sbox_5_M6 ;
    wire SubBytesIns_Inst_Sbox_5_M5 ;
    wire SubBytesIns_Inst_Sbox_5_M4 ;
    wire SubBytesIns_Inst_Sbox_5_M3 ;
    wire SubBytesIns_Inst_Sbox_5_M2 ;
    wire SubBytesIns_Inst_Sbox_5_M1 ;
    wire SubBytesIns_Inst_Sbox_5_T27 ;
    wire SubBytesIns_Inst_Sbox_5_T26 ;
    wire SubBytesIns_Inst_Sbox_5_T25 ;
    wire SubBytesIns_Inst_Sbox_5_T24 ;
    wire SubBytesIns_Inst_Sbox_5_T23 ;
    wire SubBytesIns_Inst_Sbox_5_T22 ;
    wire SubBytesIns_Inst_Sbox_5_T21 ;
    wire SubBytesIns_Inst_Sbox_5_T20 ;
    wire SubBytesIns_Inst_Sbox_5_T19 ;
    wire SubBytesIns_Inst_Sbox_5_T18 ;
    wire SubBytesIns_Inst_Sbox_5_T17 ;
    wire SubBytesIns_Inst_Sbox_5_T16 ;
    wire SubBytesIns_Inst_Sbox_5_T15 ;
    wire SubBytesIns_Inst_Sbox_5_T14 ;
    wire SubBytesIns_Inst_Sbox_5_T13 ;
    wire SubBytesIns_Inst_Sbox_5_T12 ;
    wire SubBytesIns_Inst_Sbox_5_T11 ;
    wire SubBytesIns_Inst_Sbox_5_T10 ;
    wire SubBytesIns_Inst_Sbox_5_T9 ;
    wire SubBytesIns_Inst_Sbox_5_T8 ;
    wire SubBytesIns_Inst_Sbox_5_T7 ;
    wire SubBytesIns_Inst_Sbox_5_T6 ;
    wire SubBytesIns_Inst_Sbox_5_T5 ;
    wire SubBytesIns_Inst_Sbox_5_T4 ;
    wire SubBytesIns_Inst_Sbox_5_T3 ;
    wire SubBytesIns_Inst_Sbox_5_T2 ;
    wire SubBytesIns_Inst_Sbox_5_T1 ;
    wire SubBytesIns_Inst_Sbox_6_L29 ;
    wire SubBytesIns_Inst_Sbox_6_L28 ;
    wire SubBytesIns_Inst_Sbox_6_L27 ;
    wire SubBytesIns_Inst_Sbox_6_L26 ;
    wire SubBytesIns_Inst_Sbox_6_L25 ;
    wire SubBytesIns_Inst_Sbox_6_L24 ;
    wire SubBytesIns_Inst_Sbox_6_L23 ;
    wire SubBytesIns_Inst_Sbox_6_L22 ;
    wire SubBytesIns_Inst_Sbox_6_L21 ;
    wire SubBytesIns_Inst_Sbox_6_L20 ;
    wire SubBytesIns_Inst_Sbox_6_L19 ;
    wire SubBytesIns_Inst_Sbox_6_L18 ;
    wire SubBytesIns_Inst_Sbox_6_L17 ;
    wire SubBytesIns_Inst_Sbox_6_L16 ;
    wire SubBytesIns_Inst_Sbox_6_L15 ;
    wire SubBytesIns_Inst_Sbox_6_L14 ;
    wire SubBytesIns_Inst_Sbox_6_L13 ;
    wire SubBytesIns_Inst_Sbox_6_L12 ;
    wire SubBytesIns_Inst_Sbox_6_L11 ;
    wire SubBytesIns_Inst_Sbox_6_L10 ;
    wire SubBytesIns_Inst_Sbox_6_L9 ;
    wire SubBytesIns_Inst_Sbox_6_L8 ;
    wire SubBytesIns_Inst_Sbox_6_L7 ;
    wire SubBytesIns_Inst_Sbox_6_L6 ;
    wire SubBytesIns_Inst_Sbox_6_L5 ;
    wire SubBytesIns_Inst_Sbox_6_L4 ;
    wire SubBytesIns_Inst_Sbox_6_L3 ;
    wire SubBytesIns_Inst_Sbox_6_L2 ;
    wire SubBytesIns_Inst_Sbox_6_L1 ;
    wire SubBytesIns_Inst_Sbox_6_L0 ;
    wire SubBytesIns_Inst_Sbox_6_M63 ;
    wire SubBytesIns_Inst_Sbox_6_M62 ;
    wire SubBytesIns_Inst_Sbox_6_M61 ;
    wire SubBytesIns_Inst_Sbox_6_M60 ;
    wire SubBytesIns_Inst_Sbox_6_M59 ;
    wire SubBytesIns_Inst_Sbox_6_M58 ;
    wire SubBytesIns_Inst_Sbox_6_M57 ;
    wire SubBytesIns_Inst_Sbox_6_M56 ;
    wire SubBytesIns_Inst_Sbox_6_M55 ;
    wire SubBytesIns_Inst_Sbox_6_M54 ;
    wire SubBytesIns_Inst_Sbox_6_M53 ;
    wire SubBytesIns_Inst_Sbox_6_M52 ;
    wire SubBytesIns_Inst_Sbox_6_M51 ;
    wire SubBytesIns_Inst_Sbox_6_M50 ;
    wire SubBytesIns_Inst_Sbox_6_M49 ;
    wire SubBytesIns_Inst_Sbox_6_M48 ;
    wire SubBytesIns_Inst_Sbox_6_M47 ;
    wire SubBytesIns_Inst_Sbox_6_M46 ;
    wire SubBytesIns_Inst_Sbox_6_M45 ;
    wire SubBytesIns_Inst_Sbox_6_M44 ;
    wire SubBytesIns_Inst_Sbox_6_M43 ;
    wire SubBytesIns_Inst_Sbox_6_M42 ;
    wire SubBytesIns_Inst_Sbox_6_M41 ;
    wire SubBytesIns_Inst_Sbox_6_M40 ;
    wire SubBytesIns_Inst_Sbox_6_M39 ;
    wire SubBytesIns_Inst_Sbox_6_M38 ;
    wire SubBytesIns_Inst_Sbox_6_M37 ;
    wire SubBytesIns_Inst_Sbox_6_M36 ;
    wire SubBytesIns_Inst_Sbox_6_M35 ;
    wire SubBytesIns_Inst_Sbox_6_M34 ;
    wire SubBytesIns_Inst_Sbox_6_M33 ;
    wire SubBytesIns_Inst_Sbox_6_M32 ;
    wire SubBytesIns_Inst_Sbox_6_M31 ;
    wire SubBytesIns_Inst_Sbox_6_M30 ;
    wire SubBytesIns_Inst_Sbox_6_M29 ;
    wire SubBytesIns_Inst_Sbox_6_M28 ;
    wire SubBytesIns_Inst_Sbox_6_M27 ;
    wire SubBytesIns_Inst_Sbox_6_M26 ;
    wire SubBytesIns_Inst_Sbox_6_M25 ;
    wire SubBytesIns_Inst_Sbox_6_M24 ;
    wire SubBytesIns_Inst_Sbox_6_M23 ;
    wire SubBytesIns_Inst_Sbox_6_M22 ;
    wire SubBytesIns_Inst_Sbox_6_M21 ;
    wire SubBytesIns_Inst_Sbox_6_M20 ;
    wire SubBytesIns_Inst_Sbox_6_M19 ;
    wire SubBytesIns_Inst_Sbox_6_M18 ;
    wire SubBytesIns_Inst_Sbox_6_M17 ;
    wire SubBytesIns_Inst_Sbox_6_M16 ;
    wire SubBytesIns_Inst_Sbox_6_M15 ;
    wire SubBytesIns_Inst_Sbox_6_M14 ;
    wire SubBytesIns_Inst_Sbox_6_M13 ;
    wire SubBytesIns_Inst_Sbox_6_M12 ;
    wire SubBytesIns_Inst_Sbox_6_M11 ;
    wire SubBytesIns_Inst_Sbox_6_M10 ;
    wire SubBytesIns_Inst_Sbox_6_M9 ;
    wire SubBytesIns_Inst_Sbox_6_M8 ;
    wire SubBytesIns_Inst_Sbox_6_M7 ;
    wire SubBytesIns_Inst_Sbox_6_M6 ;
    wire SubBytesIns_Inst_Sbox_6_M5 ;
    wire SubBytesIns_Inst_Sbox_6_M4 ;
    wire SubBytesIns_Inst_Sbox_6_M3 ;
    wire SubBytesIns_Inst_Sbox_6_M2 ;
    wire SubBytesIns_Inst_Sbox_6_M1 ;
    wire SubBytesIns_Inst_Sbox_6_T27 ;
    wire SubBytesIns_Inst_Sbox_6_T26 ;
    wire SubBytesIns_Inst_Sbox_6_T25 ;
    wire SubBytesIns_Inst_Sbox_6_T24 ;
    wire SubBytesIns_Inst_Sbox_6_T23 ;
    wire SubBytesIns_Inst_Sbox_6_T22 ;
    wire SubBytesIns_Inst_Sbox_6_T21 ;
    wire SubBytesIns_Inst_Sbox_6_T20 ;
    wire SubBytesIns_Inst_Sbox_6_T19 ;
    wire SubBytesIns_Inst_Sbox_6_T18 ;
    wire SubBytesIns_Inst_Sbox_6_T17 ;
    wire SubBytesIns_Inst_Sbox_6_T16 ;
    wire SubBytesIns_Inst_Sbox_6_T15 ;
    wire SubBytesIns_Inst_Sbox_6_T14 ;
    wire SubBytesIns_Inst_Sbox_6_T13 ;
    wire SubBytesIns_Inst_Sbox_6_T12 ;
    wire SubBytesIns_Inst_Sbox_6_T11 ;
    wire SubBytesIns_Inst_Sbox_6_T10 ;
    wire SubBytesIns_Inst_Sbox_6_T9 ;
    wire SubBytesIns_Inst_Sbox_6_T8 ;
    wire SubBytesIns_Inst_Sbox_6_T7 ;
    wire SubBytesIns_Inst_Sbox_6_T6 ;
    wire SubBytesIns_Inst_Sbox_6_T5 ;
    wire SubBytesIns_Inst_Sbox_6_T4 ;
    wire SubBytesIns_Inst_Sbox_6_T3 ;
    wire SubBytesIns_Inst_Sbox_6_T2 ;
    wire SubBytesIns_Inst_Sbox_6_T1 ;
    wire SubBytesIns_Inst_Sbox_7_L29 ;
    wire SubBytesIns_Inst_Sbox_7_L28 ;
    wire SubBytesIns_Inst_Sbox_7_L27 ;
    wire SubBytesIns_Inst_Sbox_7_L26 ;
    wire SubBytesIns_Inst_Sbox_7_L25 ;
    wire SubBytesIns_Inst_Sbox_7_L24 ;
    wire SubBytesIns_Inst_Sbox_7_L23 ;
    wire SubBytesIns_Inst_Sbox_7_L22 ;
    wire SubBytesIns_Inst_Sbox_7_L21 ;
    wire SubBytesIns_Inst_Sbox_7_L20 ;
    wire SubBytesIns_Inst_Sbox_7_L19 ;
    wire SubBytesIns_Inst_Sbox_7_L18 ;
    wire SubBytesIns_Inst_Sbox_7_L17 ;
    wire SubBytesIns_Inst_Sbox_7_L16 ;
    wire SubBytesIns_Inst_Sbox_7_L15 ;
    wire SubBytesIns_Inst_Sbox_7_L14 ;
    wire SubBytesIns_Inst_Sbox_7_L13 ;
    wire SubBytesIns_Inst_Sbox_7_L12 ;
    wire SubBytesIns_Inst_Sbox_7_L11 ;
    wire SubBytesIns_Inst_Sbox_7_L10 ;
    wire SubBytesIns_Inst_Sbox_7_L9 ;
    wire SubBytesIns_Inst_Sbox_7_L8 ;
    wire SubBytesIns_Inst_Sbox_7_L7 ;
    wire SubBytesIns_Inst_Sbox_7_L6 ;
    wire SubBytesIns_Inst_Sbox_7_L5 ;
    wire SubBytesIns_Inst_Sbox_7_L4 ;
    wire SubBytesIns_Inst_Sbox_7_L3 ;
    wire SubBytesIns_Inst_Sbox_7_L2 ;
    wire SubBytesIns_Inst_Sbox_7_L1 ;
    wire SubBytesIns_Inst_Sbox_7_L0 ;
    wire SubBytesIns_Inst_Sbox_7_M63 ;
    wire SubBytesIns_Inst_Sbox_7_M62 ;
    wire SubBytesIns_Inst_Sbox_7_M61 ;
    wire SubBytesIns_Inst_Sbox_7_M60 ;
    wire SubBytesIns_Inst_Sbox_7_M59 ;
    wire SubBytesIns_Inst_Sbox_7_M58 ;
    wire SubBytesIns_Inst_Sbox_7_M57 ;
    wire SubBytesIns_Inst_Sbox_7_M56 ;
    wire SubBytesIns_Inst_Sbox_7_M55 ;
    wire SubBytesIns_Inst_Sbox_7_M54 ;
    wire SubBytesIns_Inst_Sbox_7_M53 ;
    wire SubBytesIns_Inst_Sbox_7_M52 ;
    wire SubBytesIns_Inst_Sbox_7_M51 ;
    wire SubBytesIns_Inst_Sbox_7_M50 ;
    wire SubBytesIns_Inst_Sbox_7_M49 ;
    wire SubBytesIns_Inst_Sbox_7_M48 ;
    wire SubBytesIns_Inst_Sbox_7_M47 ;
    wire SubBytesIns_Inst_Sbox_7_M46 ;
    wire SubBytesIns_Inst_Sbox_7_M45 ;
    wire SubBytesIns_Inst_Sbox_7_M44 ;
    wire SubBytesIns_Inst_Sbox_7_M43 ;
    wire SubBytesIns_Inst_Sbox_7_M42 ;
    wire SubBytesIns_Inst_Sbox_7_M41 ;
    wire SubBytesIns_Inst_Sbox_7_M40 ;
    wire SubBytesIns_Inst_Sbox_7_M39 ;
    wire SubBytesIns_Inst_Sbox_7_M38 ;
    wire SubBytesIns_Inst_Sbox_7_M37 ;
    wire SubBytesIns_Inst_Sbox_7_M36 ;
    wire SubBytesIns_Inst_Sbox_7_M35 ;
    wire SubBytesIns_Inst_Sbox_7_M34 ;
    wire SubBytesIns_Inst_Sbox_7_M33 ;
    wire SubBytesIns_Inst_Sbox_7_M32 ;
    wire SubBytesIns_Inst_Sbox_7_M31 ;
    wire SubBytesIns_Inst_Sbox_7_M30 ;
    wire SubBytesIns_Inst_Sbox_7_M29 ;
    wire SubBytesIns_Inst_Sbox_7_M28 ;
    wire SubBytesIns_Inst_Sbox_7_M27 ;
    wire SubBytesIns_Inst_Sbox_7_M26 ;
    wire SubBytesIns_Inst_Sbox_7_M25 ;
    wire SubBytesIns_Inst_Sbox_7_M24 ;
    wire SubBytesIns_Inst_Sbox_7_M23 ;
    wire SubBytesIns_Inst_Sbox_7_M22 ;
    wire SubBytesIns_Inst_Sbox_7_M21 ;
    wire SubBytesIns_Inst_Sbox_7_M20 ;
    wire SubBytesIns_Inst_Sbox_7_M19 ;
    wire SubBytesIns_Inst_Sbox_7_M18 ;
    wire SubBytesIns_Inst_Sbox_7_M17 ;
    wire SubBytesIns_Inst_Sbox_7_M16 ;
    wire SubBytesIns_Inst_Sbox_7_M15 ;
    wire SubBytesIns_Inst_Sbox_7_M14 ;
    wire SubBytesIns_Inst_Sbox_7_M13 ;
    wire SubBytesIns_Inst_Sbox_7_M12 ;
    wire SubBytesIns_Inst_Sbox_7_M11 ;
    wire SubBytesIns_Inst_Sbox_7_M10 ;
    wire SubBytesIns_Inst_Sbox_7_M9 ;
    wire SubBytesIns_Inst_Sbox_7_M8 ;
    wire SubBytesIns_Inst_Sbox_7_M7 ;
    wire SubBytesIns_Inst_Sbox_7_M6 ;
    wire SubBytesIns_Inst_Sbox_7_M5 ;
    wire SubBytesIns_Inst_Sbox_7_M4 ;
    wire SubBytesIns_Inst_Sbox_7_M3 ;
    wire SubBytesIns_Inst_Sbox_7_M2 ;
    wire SubBytesIns_Inst_Sbox_7_M1 ;
    wire SubBytesIns_Inst_Sbox_7_T27 ;
    wire SubBytesIns_Inst_Sbox_7_T26 ;
    wire SubBytesIns_Inst_Sbox_7_T25 ;
    wire SubBytesIns_Inst_Sbox_7_T24 ;
    wire SubBytesIns_Inst_Sbox_7_T23 ;
    wire SubBytesIns_Inst_Sbox_7_T22 ;
    wire SubBytesIns_Inst_Sbox_7_T21 ;
    wire SubBytesIns_Inst_Sbox_7_T20 ;
    wire SubBytesIns_Inst_Sbox_7_T19 ;
    wire SubBytesIns_Inst_Sbox_7_T18 ;
    wire SubBytesIns_Inst_Sbox_7_T17 ;
    wire SubBytesIns_Inst_Sbox_7_T16 ;
    wire SubBytesIns_Inst_Sbox_7_T15 ;
    wire SubBytesIns_Inst_Sbox_7_T14 ;
    wire SubBytesIns_Inst_Sbox_7_T13 ;
    wire SubBytesIns_Inst_Sbox_7_T12 ;
    wire SubBytesIns_Inst_Sbox_7_T11 ;
    wire SubBytesIns_Inst_Sbox_7_T10 ;
    wire SubBytesIns_Inst_Sbox_7_T9 ;
    wire SubBytesIns_Inst_Sbox_7_T8 ;
    wire SubBytesIns_Inst_Sbox_7_T7 ;
    wire SubBytesIns_Inst_Sbox_7_T6 ;
    wire SubBytesIns_Inst_Sbox_7_T5 ;
    wire SubBytesIns_Inst_Sbox_7_T4 ;
    wire SubBytesIns_Inst_Sbox_7_T3 ;
    wire SubBytesIns_Inst_Sbox_7_T2 ;
    wire SubBytesIns_Inst_Sbox_7_T1 ;
    wire SubBytesIns_Inst_Sbox_8_L29 ;
    wire SubBytesIns_Inst_Sbox_8_L28 ;
    wire SubBytesIns_Inst_Sbox_8_L27 ;
    wire SubBytesIns_Inst_Sbox_8_L26 ;
    wire SubBytesIns_Inst_Sbox_8_L25 ;
    wire SubBytesIns_Inst_Sbox_8_L24 ;
    wire SubBytesIns_Inst_Sbox_8_L23 ;
    wire SubBytesIns_Inst_Sbox_8_L22 ;
    wire SubBytesIns_Inst_Sbox_8_L21 ;
    wire SubBytesIns_Inst_Sbox_8_L20 ;
    wire SubBytesIns_Inst_Sbox_8_L19 ;
    wire SubBytesIns_Inst_Sbox_8_L18 ;
    wire SubBytesIns_Inst_Sbox_8_L17 ;
    wire SubBytesIns_Inst_Sbox_8_L16 ;
    wire SubBytesIns_Inst_Sbox_8_L15 ;
    wire SubBytesIns_Inst_Sbox_8_L14 ;
    wire SubBytesIns_Inst_Sbox_8_L13 ;
    wire SubBytesIns_Inst_Sbox_8_L12 ;
    wire SubBytesIns_Inst_Sbox_8_L11 ;
    wire SubBytesIns_Inst_Sbox_8_L10 ;
    wire SubBytesIns_Inst_Sbox_8_L9 ;
    wire SubBytesIns_Inst_Sbox_8_L8 ;
    wire SubBytesIns_Inst_Sbox_8_L7 ;
    wire SubBytesIns_Inst_Sbox_8_L6 ;
    wire SubBytesIns_Inst_Sbox_8_L5 ;
    wire SubBytesIns_Inst_Sbox_8_L4 ;
    wire SubBytesIns_Inst_Sbox_8_L3 ;
    wire SubBytesIns_Inst_Sbox_8_L2 ;
    wire SubBytesIns_Inst_Sbox_8_L1 ;
    wire SubBytesIns_Inst_Sbox_8_L0 ;
    wire SubBytesIns_Inst_Sbox_8_M63 ;
    wire SubBytesIns_Inst_Sbox_8_M62 ;
    wire SubBytesIns_Inst_Sbox_8_M61 ;
    wire SubBytesIns_Inst_Sbox_8_M60 ;
    wire SubBytesIns_Inst_Sbox_8_M59 ;
    wire SubBytesIns_Inst_Sbox_8_M58 ;
    wire SubBytesIns_Inst_Sbox_8_M57 ;
    wire SubBytesIns_Inst_Sbox_8_M56 ;
    wire SubBytesIns_Inst_Sbox_8_M55 ;
    wire SubBytesIns_Inst_Sbox_8_M54 ;
    wire SubBytesIns_Inst_Sbox_8_M53 ;
    wire SubBytesIns_Inst_Sbox_8_M52 ;
    wire SubBytesIns_Inst_Sbox_8_M51 ;
    wire SubBytesIns_Inst_Sbox_8_M50 ;
    wire SubBytesIns_Inst_Sbox_8_M49 ;
    wire SubBytesIns_Inst_Sbox_8_M48 ;
    wire SubBytesIns_Inst_Sbox_8_M47 ;
    wire SubBytesIns_Inst_Sbox_8_M46 ;
    wire SubBytesIns_Inst_Sbox_8_M45 ;
    wire SubBytesIns_Inst_Sbox_8_M44 ;
    wire SubBytesIns_Inst_Sbox_8_M43 ;
    wire SubBytesIns_Inst_Sbox_8_M42 ;
    wire SubBytesIns_Inst_Sbox_8_M41 ;
    wire SubBytesIns_Inst_Sbox_8_M40 ;
    wire SubBytesIns_Inst_Sbox_8_M39 ;
    wire SubBytesIns_Inst_Sbox_8_M38 ;
    wire SubBytesIns_Inst_Sbox_8_M37 ;
    wire SubBytesIns_Inst_Sbox_8_M36 ;
    wire SubBytesIns_Inst_Sbox_8_M35 ;
    wire SubBytesIns_Inst_Sbox_8_M34 ;
    wire SubBytesIns_Inst_Sbox_8_M33 ;
    wire SubBytesIns_Inst_Sbox_8_M32 ;
    wire SubBytesIns_Inst_Sbox_8_M31 ;
    wire SubBytesIns_Inst_Sbox_8_M30 ;
    wire SubBytesIns_Inst_Sbox_8_M29 ;
    wire SubBytesIns_Inst_Sbox_8_M28 ;
    wire SubBytesIns_Inst_Sbox_8_M27 ;
    wire SubBytesIns_Inst_Sbox_8_M26 ;
    wire SubBytesIns_Inst_Sbox_8_M25 ;
    wire SubBytesIns_Inst_Sbox_8_M24 ;
    wire SubBytesIns_Inst_Sbox_8_M23 ;
    wire SubBytesIns_Inst_Sbox_8_M22 ;
    wire SubBytesIns_Inst_Sbox_8_M21 ;
    wire SubBytesIns_Inst_Sbox_8_M20 ;
    wire SubBytesIns_Inst_Sbox_8_M19 ;
    wire SubBytesIns_Inst_Sbox_8_M18 ;
    wire SubBytesIns_Inst_Sbox_8_M17 ;
    wire SubBytesIns_Inst_Sbox_8_M16 ;
    wire SubBytesIns_Inst_Sbox_8_M15 ;
    wire SubBytesIns_Inst_Sbox_8_M14 ;
    wire SubBytesIns_Inst_Sbox_8_M13 ;
    wire SubBytesIns_Inst_Sbox_8_M12 ;
    wire SubBytesIns_Inst_Sbox_8_M11 ;
    wire SubBytesIns_Inst_Sbox_8_M10 ;
    wire SubBytesIns_Inst_Sbox_8_M9 ;
    wire SubBytesIns_Inst_Sbox_8_M8 ;
    wire SubBytesIns_Inst_Sbox_8_M7 ;
    wire SubBytesIns_Inst_Sbox_8_M6 ;
    wire SubBytesIns_Inst_Sbox_8_M5 ;
    wire SubBytesIns_Inst_Sbox_8_M4 ;
    wire SubBytesIns_Inst_Sbox_8_M3 ;
    wire SubBytesIns_Inst_Sbox_8_M2 ;
    wire SubBytesIns_Inst_Sbox_8_M1 ;
    wire SubBytesIns_Inst_Sbox_8_T27 ;
    wire SubBytesIns_Inst_Sbox_8_T26 ;
    wire SubBytesIns_Inst_Sbox_8_T25 ;
    wire SubBytesIns_Inst_Sbox_8_T24 ;
    wire SubBytesIns_Inst_Sbox_8_T23 ;
    wire SubBytesIns_Inst_Sbox_8_T22 ;
    wire SubBytesIns_Inst_Sbox_8_T21 ;
    wire SubBytesIns_Inst_Sbox_8_T20 ;
    wire SubBytesIns_Inst_Sbox_8_T19 ;
    wire SubBytesIns_Inst_Sbox_8_T18 ;
    wire SubBytesIns_Inst_Sbox_8_T17 ;
    wire SubBytesIns_Inst_Sbox_8_T16 ;
    wire SubBytesIns_Inst_Sbox_8_T15 ;
    wire SubBytesIns_Inst_Sbox_8_T14 ;
    wire SubBytesIns_Inst_Sbox_8_T13 ;
    wire SubBytesIns_Inst_Sbox_8_T12 ;
    wire SubBytesIns_Inst_Sbox_8_T11 ;
    wire SubBytesIns_Inst_Sbox_8_T10 ;
    wire SubBytesIns_Inst_Sbox_8_T9 ;
    wire SubBytesIns_Inst_Sbox_8_T8 ;
    wire SubBytesIns_Inst_Sbox_8_T7 ;
    wire SubBytesIns_Inst_Sbox_8_T6 ;
    wire SubBytesIns_Inst_Sbox_8_T5 ;
    wire SubBytesIns_Inst_Sbox_8_T4 ;
    wire SubBytesIns_Inst_Sbox_8_T3 ;
    wire SubBytesIns_Inst_Sbox_8_T2 ;
    wire SubBytesIns_Inst_Sbox_8_T1 ;
    wire SubBytesIns_Inst_Sbox_9_L29 ;
    wire SubBytesIns_Inst_Sbox_9_L28 ;
    wire SubBytesIns_Inst_Sbox_9_L27 ;
    wire SubBytesIns_Inst_Sbox_9_L26 ;
    wire SubBytesIns_Inst_Sbox_9_L25 ;
    wire SubBytesIns_Inst_Sbox_9_L24 ;
    wire SubBytesIns_Inst_Sbox_9_L23 ;
    wire SubBytesIns_Inst_Sbox_9_L22 ;
    wire SubBytesIns_Inst_Sbox_9_L21 ;
    wire SubBytesIns_Inst_Sbox_9_L20 ;
    wire SubBytesIns_Inst_Sbox_9_L19 ;
    wire SubBytesIns_Inst_Sbox_9_L18 ;
    wire SubBytesIns_Inst_Sbox_9_L17 ;
    wire SubBytesIns_Inst_Sbox_9_L16 ;
    wire SubBytesIns_Inst_Sbox_9_L15 ;
    wire SubBytesIns_Inst_Sbox_9_L14 ;
    wire SubBytesIns_Inst_Sbox_9_L13 ;
    wire SubBytesIns_Inst_Sbox_9_L12 ;
    wire SubBytesIns_Inst_Sbox_9_L11 ;
    wire SubBytesIns_Inst_Sbox_9_L10 ;
    wire SubBytesIns_Inst_Sbox_9_L9 ;
    wire SubBytesIns_Inst_Sbox_9_L8 ;
    wire SubBytesIns_Inst_Sbox_9_L7 ;
    wire SubBytesIns_Inst_Sbox_9_L6 ;
    wire SubBytesIns_Inst_Sbox_9_L5 ;
    wire SubBytesIns_Inst_Sbox_9_L4 ;
    wire SubBytesIns_Inst_Sbox_9_L3 ;
    wire SubBytesIns_Inst_Sbox_9_L2 ;
    wire SubBytesIns_Inst_Sbox_9_L1 ;
    wire SubBytesIns_Inst_Sbox_9_L0 ;
    wire SubBytesIns_Inst_Sbox_9_M63 ;
    wire SubBytesIns_Inst_Sbox_9_M62 ;
    wire SubBytesIns_Inst_Sbox_9_M61 ;
    wire SubBytesIns_Inst_Sbox_9_M60 ;
    wire SubBytesIns_Inst_Sbox_9_M59 ;
    wire SubBytesIns_Inst_Sbox_9_M58 ;
    wire SubBytesIns_Inst_Sbox_9_M57 ;
    wire SubBytesIns_Inst_Sbox_9_M56 ;
    wire SubBytesIns_Inst_Sbox_9_M55 ;
    wire SubBytesIns_Inst_Sbox_9_M54 ;
    wire SubBytesIns_Inst_Sbox_9_M53 ;
    wire SubBytesIns_Inst_Sbox_9_M52 ;
    wire SubBytesIns_Inst_Sbox_9_M51 ;
    wire SubBytesIns_Inst_Sbox_9_M50 ;
    wire SubBytesIns_Inst_Sbox_9_M49 ;
    wire SubBytesIns_Inst_Sbox_9_M48 ;
    wire SubBytesIns_Inst_Sbox_9_M47 ;
    wire SubBytesIns_Inst_Sbox_9_M46 ;
    wire SubBytesIns_Inst_Sbox_9_M45 ;
    wire SubBytesIns_Inst_Sbox_9_M44 ;
    wire SubBytesIns_Inst_Sbox_9_M43 ;
    wire SubBytesIns_Inst_Sbox_9_M42 ;
    wire SubBytesIns_Inst_Sbox_9_M41 ;
    wire SubBytesIns_Inst_Sbox_9_M40 ;
    wire SubBytesIns_Inst_Sbox_9_M39 ;
    wire SubBytesIns_Inst_Sbox_9_M38 ;
    wire SubBytesIns_Inst_Sbox_9_M37 ;
    wire SubBytesIns_Inst_Sbox_9_M36 ;
    wire SubBytesIns_Inst_Sbox_9_M35 ;
    wire SubBytesIns_Inst_Sbox_9_M34 ;
    wire SubBytesIns_Inst_Sbox_9_M33 ;
    wire SubBytesIns_Inst_Sbox_9_M32 ;
    wire SubBytesIns_Inst_Sbox_9_M31 ;
    wire SubBytesIns_Inst_Sbox_9_M30 ;
    wire SubBytesIns_Inst_Sbox_9_M29 ;
    wire SubBytesIns_Inst_Sbox_9_M28 ;
    wire SubBytesIns_Inst_Sbox_9_M27 ;
    wire SubBytesIns_Inst_Sbox_9_M26 ;
    wire SubBytesIns_Inst_Sbox_9_M25 ;
    wire SubBytesIns_Inst_Sbox_9_M24 ;
    wire SubBytesIns_Inst_Sbox_9_M23 ;
    wire SubBytesIns_Inst_Sbox_9_M22 ;
    wire SubBytesIns_Inst_Sbox_9_M21 ;
    wire SubBytesIns_Inst_Sbox_9_M20 ;
    wire SubBytesIns_Inst_Sbox_9_M19 ;
    wire SubBytesIns_Inst_Sbox_9_M18 ;
    wire SubBytesIns_Inst_Sbox_9_M17 ;
    wire SubBytesIns_Inst_Sbox_9_M16 ;
    wire SubBytesIns_Inst_Sbox_9_M15 ;
    wire SubBytesIns_Inst_Sbox_9_M14 ;
    wire SubBytesIns_Inst_Sbox_9_M13 ;
    wire SubBytesIns_Inst_Sbox_9_M12 ;
    wire SubBytesIns_Inst_Sbox_9_M11 ;
    wire SubBytesIns_Inst_Sbox_9_M10 ;
    wire SubBytesIns_Inst_Sbox_9_M9 ;
    wire SubBytesIns_Inst_Sbox_9_M8 ;
    wire SubBytesIns_Inst_Sbox_9_M7 ;
    wire SubBytesIns_Inst_Sbox_9_M6 ;
    wire SubBytesIns_Inst_Sbox_9_M5 ;
    wire SubBytesIns_Inst_Sbox_9_M4 ;
    wire SubBytesIns_Inst_Sbox_9_M3 ;
    wire SubBytesIns_Inst_Sbox_9_M2 ;
    wire SubBytesIns_Inst_Sbox_9_M1 ;
    wire SubBytesIns_Inst_Sbox_9_T27 ;
    wire SubBytesIns_Inst_Sbox_9_T26 ;
    wire SubBytesIns_Inst_Sbox_9_T25 ;
    wire SubBytesIns_Inst_Sbox_9_T24 ;
    wire SubBytesIns_Inst_Sbox_9_T23 ;
    wire SubBytesIns_Inst_Sbox_9_T22 ;
    wire SubBytesIns_Inst_Sbox_9_T21 ;
    wire SubBytesIns_Inst_Sbox_9_T20 ;
    wire SubBytesIns_Inst_Sbox_9_T19 ;
    wire SubBytesIns_Inst_Sbox_9_T18 ;
    wire SubBytesIns_Inst_Sbox_9_T17 ;
    wire SubBytesIns_Inst_Sbox_9_T16 ;
    wire SubBytesIns_Inst_Sbox_9_T15 ;
    wire SubBytesIns_Inst_Sbox_9_T14 ;
    wire SubBytesIns_Inst_Sbox_9_T13 ;
    wire SubBytesIns_Inst_Sbox_9_T12 ;
    wire SubBytesIns_Inst_Sbox_9_T11 ;
    wire SubBytesIns_Inst_Sbox_9_T10 ;
    wire SubBytesIns_Inst_Sbox_9_T9 ;
    wire SubBytesIns_Inst_Sbox_9_T8 ;
    wire SubBytesIns_Inst_Sbox_9_T7 ;
    wire SubBytesIns_Inst_Sbox_9_T6 ;
    wire SubBytesIns_Inst_Sbox_9_T5 ;
    wire SubBytesIns_Inst_Sbox_9_T4 ;
    wire SubBytesIns_Inst_Sbox_9_T3 ;
    wire SubBytesIns_Inst_Sbox_9_T2 ;
    wire SubBytesIns_Inst_Sbox_9_T1 ;
    wire SubBytesIns_Inst_Sbox_10_L29 ;
    wire SubBytesIns_Inst_Sbox_10_L28 ;
    wire SubBytesIns_Inst_Sbox_10_L27 ;
    wire SubBytesIns_Inst_Sbox_10_L26 ;
    wire SubBytesIns_Inst_Sbox_10_L25 ;
    wire SubBytesIns_Inst_Sbox_10_L24 ;
    wire SubBytesIns_Inst_Sbox_10_L23 ;
    wire SubBytesIns_Inst_Sbox_10_L22 ;
    wire SubBytesIns_Inst_Sbox_10_L21 ;
    wire SubBytesIns_Inst_Sbox_10_L20 ;
    wire SubBytesIns_Inst_Sbox_10_L19 ;
    wire SubBytesIns_Inst_Sbox_10_L18 ;
    wire SubBytesIns_Inst_Sbox_10_L17 ;
    wire SubBytesIns_Inst_Sbox_10_L16 ;
    wire SubBytesIns_Inst_Sbox_10_L15 ;
    wire SubBytesIns_Inst_Sbox_10_L14 ;
    wire SubBytesIns_Inst_Sbox_10_L13 ;
    wire SubBytesIns_Inst_Sbox_10_L12 ;
    wire SubBytesIns_Inst_Sbox_10_L11 ;
    wire SubBytesIns_Inst_Sbox_10_L10 ;
    wire SubBytesIns_Inst_Sbox_10_L9 ;
    wire SubBytesIns_Inst_Sbox_10_L8 ;
    wire SubBytesIns_Inst_Sbox_10_L7 ;
    wire SubBytesIns_Inst_Sbox_10_L6 ;
    wire SubBytesIns_Inst_Sbox_10_L5 ;
    wire SubBytesIns_Inst_Sbox_10_L4 ;
    wire SubBytesIns_Inst_Sbox_10_L3 ;
    wire SubBytesIns_Inst_Sbox_10_L2 ;
    wire SubBytesIns_Inst_Sbox_10_L1 ;
    wire SubBytesIns_Inst_Sbox_10_L0 ;
    wire SubBytesIns_Inst_Sbox_10_M63 ;
    wire SubBytesIns_Inst_Sbox_10_M62 ;
    wire SubBytesIns_Inst_Sbox_10_M61 ;
    wire SubBytesIns_Inst_Sbox_10_M60 ;
    wire SubBytesIns_Inst_Sbox_10_M59 ;
    wire SubBytesIns_Inst_Sbox_10_M58 ;
    wire SubBytesIns_Inst_Sbox_10_M57 ;
    wire SubBytesIns_Inst_Sbox_10_M56 ;
    wire SubBytesIns_Inst_Sbox_10_M55 ;
    wire SubBytesIns_Inst_Sbox_10_M54 ;
    wire SubBytesIns_Inst_Sbox_10_M53 ;
    wire SubBytesIns_Inst_Sbox_10_M52 ;
    wire SubBytesIns_Inst_Sbox_10_M51 ;
    wire SubBytesIns_Inst_Sbox_10_M50 ;
    wire SubBytesIns_Inst_Sbox_10_M49 ;
    wire SubBytesIns_Inst_Sbox_10_M48 ;
    wire SubBytesIns_Inst_Sbox_10_M47 ;
    wire SubBytesIns_Inst_Sbox_10_M46 ;
    wire SubBytesIns_Inst_Sbox_10_M45 ;
    wire SubBytesIns_Inst_Sbox_10_M44 ;
    wire SubBytesIns_Inst_Sbox_10_M43 ;
    wire SubBytesIns_Inst_Sbox_10_M42 ;
    wire SubBytesIns_Inst_Sbox_10_M41 ;
    wire SubBytesIns_Inst_Sbox_10_M40 ;
    wire SubBytesIns_Inst_Sbox_10_M39 ;
    wire SubBytesIns_Inst_Sbox_10_M38 ;
    wire SubBytesIns_Inst_Sbox_10_M37 ;
    wire SubBytesIns_Inst_Sbox_10_M36 ;
    wire SubBytesIns_Inst_Sbox_10_M35 ;
    wire SubBytesIns_Inst_Sbox_10_M34 ;
    wire SubBytesIns_Inst_Sbox_10_M33 ;
    wire SubBytesIns_Inst_Sbox_10_M32 ;
    wire SubBytesIns_Inst_Sbox_10_M31 ;
    wire SubBytesIns_Inst_Sbox_10_M30 ;
    wire SubBytesIns_Inst_Sbox_10_M29 ;
    wire SubBytesIns_Inst_Sbox_10_M28 ;
    wire SubBytesIns_Inst_Sbox_10_M27 ;
    wire SubBytesIns_Inst_Sbox_10_M26 ;
    wire SubBytesIns_Inst_Sbox_10_M25 ;
    wire SubBytesIns_Inst_Sbox_10_M24 ;
    wire SubBytesIns_Inst_Sbox_10_M23 ;
    wire SubBytesIns_Inst_Sbox_10_M22 ;
    wire SubBytesIns_Inst_Sbox_10_M21 ;
    wire SubBytesIns_Inst_Sbox_10_M20 ;
    wire SubBytesIns_Inst_Sbox_10_M19 ;
    wire SubBytesIns_Inst_Sbox_10_M18 ;
    wire SubBytesIns_Inst_Sbox_10_M17 ;
    wire SubBytesIns_Inst_Sbox_10_M16 ;
    wire SubBytesIns_Inst_Sbox_10_M15 ;
    wire SubBytesIns_Inst_Sbox_10_M14 ;
    wire SubBytesIns_Inst_Sbox_10_M13 ;
    wire SubBytesIns_Inst_Sbox_10_M12 ;
    wire SubBytesIns_Inst_Sbox_10_M11 ;
    wire SubBytesIns_Inst_Sbox_10_M10 ;
    wire SubBytesIns_Inst_Sbox_10_M9 ;
    wire SubBytesIns_Inst_Sbox_10_M8 ;
    wire SubBytesIns_Inst_Sbox_10_M7 ;
    wire SubBytesIns_Inst_Sbox_10_M6 ;
    wire SubBytesIns_Inst_Sbox_10_M5 ;
    wire SubBytesIns_Inst_Sbox_10_M4 ;
    wire SubBytesIns_Inst_Sbox_10_M3 ;
    wire SubBytesIns_Inst_Sbox_10_M2 ;
    wire SubBytesIns_Inst_Sbox_10_M1 ;
    wire SubBytesIns_Inst_Sbox_10_T27 ;
    wire SubBytesIns_Inst_Sbox_10_T26 ;
    wire SubBytesIns_Inst_Sbox_10_T25 ;
    wire SubBytesIns_Inst_Sbox_10_T24 ;
    wire SubBytesIns_Inst_Sbox_10_T23 ;
    wire SubBytesIns_Inst_Sbox_10_T22 ;
    wire SubBytesIns_Inst_Sbox_10_T21 ;
    wire SubBytesIns_Inst_Sbox_10_T20 ;
    wire SubBytesIns_Inst_Sbox_10_T19 ;
    wire SubBytesIns_Inst_Sbox_10_T18 ;
    wire SubBytesIns_Inst_Sbox_10_T17 ;
    wire SubBytesIns_Inst_Sbox_10_T16 ;
    wire SubBytesIns_Inst_Sbox_10_T15 ;
    wire SubBytesIns_Inst_Sbox_10_T14 ;
    wire SubBytesIns_Inst_Sbox_10_T13 ;
    wire SubBytesIns_Inst_Sbox_10_T12 ;
    wire SubBytesIns_Inst_Sbox_10_T11 ;
    wire SubBytesIns_Inst_Sbox_10_T10 ;
    wire SubBytesIns_Inst_Sbox_10_T9 ;
    wire SubBytesIns_Inst_Sbox_10_T8 ;
    wire SubBytesIns_Inst_Sbox_10_T7 ;
    wire SubBytesIns_Inst_Sbox_10_T6 ;
    wire SubBytesIns_Inst_Sbox_10_T5 ;
    wire SubBytesIns_Inst_Sbox_10_T4 ;
    wire SubBytesIns_Inst_Sbox_10_T3 ;
    wire SubBytesIns_Inst_Sbox_10_T2 ;
    wire SubBytesIns_Inst_Sbox_10_T1 ;
    wire SubBytesIns_Inst_Sbox_11_L29 ;
    wire SubBytesIns_Inst_Sbox_11_L28 ;
    wire SubBytesIns_Inst_Sbox_11_L27 ;
    wire SubBytesIns_Inst_Sbox_11_L26 ;
    wire SubBytesIns_Inst_Sbox_11_L25 ;
    wire SubBytesIns_Inst_Sbox_11_L24 ;
    wire SubBytesIns_Inst_Sbox_11_L23 ;
    wire SubBytesIns_Inst_Sbox_11_L22 ;
    wire SubBytesIns_Inst_Sbox_11_L21 ;
    wire SubBytesIns_Inst_Sbox_11_L20 ;
    wire SubBytesIns_Inst_Sbox_11_L19 ;
    wire SubBytesIns_Inst_Sbox_11_L18 ;
    wire SubBytesIns_Inst_Sbox_11_L17 ;
    wire SubBytesIns_Inst_Sbox_11_L16 ;
    wire SubBytesIns_Inst_Sbox_11_L15 ;
    wire SubBytesIns_Inst_Sbox_11_L14 ;
    wire SubBytesIns_Inst_Sbox_11_L13 ;
    wire SubBytesIns_Inst_Sbox_11_L12 ;
    wire SubBytesIns_Inst_Sbox_11_L11 ;
    wire SubBytesIns_Inst_Sbox_11_L10 ;
    wire SubBytesIns_Inst_Sbox_11_L9 ;
    wire SubBytesIns_Inst_Sbox_11_L8 ;
    wire SubBytesIns_Inst_Sbox_11_L7 ;
    wire SubBytesIns_Inst_Sbox_11_L6 ;
    wire SubBytesIns_Inst_Sbox_11_L5 ;
    wire SubBytesIns_Inst_Sbox_11_L4 ;
    wire SubBytesIns_Inst_Sbox_11_L3 ;
    wire SubBytesIns_Inst_Sbox_11_L2 ;
    wire SubBytesIns_Inst_Sbox_11_L1 ;
    wire SubBytesIns_Inst_Sbox_11_L0 ;
    wire SubBytesIns_Inst_Sbox_11_M63 ;
    wire SubBytesIns_Inst_Sbox_11_M62 ;
    wire SubBytesIns_Inst_Sbox_11_M61 ;
    wire SubBytesIns_Inst_Sbox_11_M60 ;
    wire SubBytesIns_Inst_Sbox_11_M59 ;
    wire SubBytesIns_Inst_Sbox_11_M58 ;
    wire SubBytesIns_Inst_Sbox_11_M57 ;
    wire SubBytesIns_Inst_Sbox_11_M56 ;
    wire SubBytesIns_Inst_Sbox_11_M55 ;
    wire SubBytesIns_Inst_Sbox_11_M54 ;
    wire SubBytesIns_Inst_Sbox_11_M53 ;
    wire SubBytesIns_Inst_Sbox_11_M52 ;
    wire SubBytesIns_Inst_Sbox_11_M51 ;
    wire SubBytesIns_Inst_Sbox_11_M50 ;
    wire SubBytesIns_Inst_Sbox_11_M49 ;
    wire SubBytesIns_Inst_Sbox_11_M48 ;
    wire SubBytesIns_Inst_Sbox_11_M47 ;
    wire SubBytesIns_Inst_Sbox_11_M46 ;
    wire SubBytesIns_Inst_Sbox_11_M45 ;
    wire SubBytesIns_Inst_Sbox_11_M44 ;
    wire SubBytesIns_Inst_Sbox_11_M43 ;
    wire SubBytesIns_Inst_Sbox_11_M42 ;
    wire SubBytesIns_Inst_Sbox_11_M41 ;
    wire SubBytesIns_Inst_Sbox_11_M40 ;
    wire SubBytesIns_Inst_Sbox_11_M39 ;
    wire SubBytesIns_Inst_Sbox_11_M38 ;
    wire SubBytesIns_Inst_Sbox_11_M37 ;
    wire SubBytesIns_Inst_Sbox_11_M36 ;
    wire SubBytesIns_Inst_Sbox_11_M35 ;
    wire SubBytesIns_Inst_Sbox_11_M34 ;
    wire SubBytesIns_Inst_Sbox_11_M33 ;
    wire SubBytesIns_Inst_Sbox_11_M32 ;
    wire SubBytesIns_Inst_Sbox_11_M31 ;
    wire SubBytesIns_Inst_Sbox_11_M30 ;
    wire SubBytesIns_Inst_Sbox_11_M29 ;
    wire SubBytesIns_Inst_Sbox_11_M28 ;
    wire SubBytesIns_Inst_Sbox_11_M27 ;
    wire SubBytesIns_Inst_Sbox_11_M26 ;
    wire SubBytesIns_Inst_Sbox_11_M25 ;
    wire SubBytesIns_Inst_Sbox_11_M24 ;
    wire SubBytesIns_Inst_Sbox_11_M23 ;
    wire SubBytesIns_Inst_Sbox_11_M22 ;
    wire SubBytesIns_Inst_Sbox_11_M21 ;
    wire SubBytesIns_Inst_Sbox_11_M20 ;
    wire SubBytesIns_Inst_Sbox_11_M19 ;
    wire SubBytesIns_Inst_Sbox_11_M18 ;
    wire SubBytesIns_Inst_Sbox_11_M17 ;
    wire SubBytesIns_Inst_Sbox_11_M16 ;
    wire SubBytesIns_Inst_Sbox_11_M15 ;
    wire SubBytesIns_Inst_Sbox_11_M14 ;
    wire SubBytesIns_Inst_Sbox_11_M13 ;
    wire SubBytesIns_Inst_Sbox_11_M12 ;
    wire SubBytesIns_Inst_Sbox_11_M11 ;
    wire SubBytesIns_Inst_Sbox_11_M10 ;
    wire SubBytesIns_Inst_Sbox_11_M9 ;
    wire SubBytesIns_Inst_Sbox_11_M8 ;
    wire SubBytesIns_Inst_Sbox_11_M7 ;
    wire SubBytesIns_Inst_Sbox_11_M6 ;
    wire SubBytesIns_Inst_Sbox_11_M5 ;
    wire SubBytesIns_Inst_Sbox_11_M4 ;
    wire SubBytesIns_Inst_Sbox_11_M3 ;
    wire SubBytesIns_Inst_Sbox_11_M2 ;
    wire SubBytesIns_Inst_Sbox_11_M1 ;
    wire SubBytesIns_Inst_Sbox_11_T27 ;
    wire SubBytesIns_Inst_Sbox_11_T26 ;
    wire SubBytesIns_Inst_Sbox_11_T25 ;
    wire SubBytesIns_Inst_Sbox_11_T24 ;
    wire SubBytesIns_Inst_Sbox_11_T23 ;
    wire SubBytesIns_Inst_Sbox_11_T22 ;
    wire SubBytesIns_Inst_Sbox_11_T21 ;
    wire SubBytesIns_Inst_Sbox_11_T20 ;
    wire SubBytesIns_Inst_Sbox_11_T19 ;
    wire SubBytesIns_Inst_Sbox_11_T18 ;
    wire SubBytesIns_Inst_Sbox_11_T17 ;
    wire SubBytesIns_Inst_Sbox_11_T16 ;
    wire SubBytesIns_Inst_Sbox_11_T15 ;
    wire SubBytesIns_Inst_Sbox_11_T14 ;
    wire SubBytesIns_Inst_Sbox_11_T13 ;
    wire SubBytesIns_Inst_Sbox_11_T12 ;
    wire SubBytesIns_Inst_Sbox_11_T11 ;
    wire SubBytesIns_Inst_Sbox_11_T10 ;
    wire SubBytesIns_Inst_Sbox_11_T9 ;
    wire SubBytesIns_Inst_Sbox_11_T8 ;
    wire SubBytesIns_Inst_Sbox_11_T7 ;
    wire SubBytesIns_Inst_Sbox_11_T6 ;
    wire SubBytesIns_Inst_Sbox_11_T5 ;
    wire SubBytesIns_Inst_Sbox_11_T4 ;
    wire SubBytesIns_Inst_Sbox_11_T3 ;
    wire SubBytesIns_Inst_Sbox_11_T2 ;
    wire SubBytesIns_Inst_Sbox_11_T1 ;
    wire SubBytesIns_Inst_Sbox_12_L29 ;
    wire SubBytesIns_Inst_Sbox_12_L28 ;
    wire SubBytesIns_Inst_Sbox_12_L27 ;
    wire SubBytesIns_Inst_Sbox_12_L26 ;
    wire SubBytesIns_Inst_Sbox_12_L25 ;
    wire SubBytesIns_Inst_Sbox_12_L24 ;
    wire SubBytesIns_Inst_Sbox_12_L23 ;
    wire SubBytesIns_Inst_Sbox_12_L22 ;
    wire SubBytesIns_Inst_Sbox_12_L21 ;
    wire SubBytesIns_Inst_Sbox_12_L20 ;
    wire SubBytesIns_Inst_Sbox_12_L19 ;
    wire SubBytesIns_Inst_Sbox_12_L18 ;
    wire SubBytesIns_Inst_Sbox_12_L17 ;
    wire SubBytesIns_Inst_Sbox_12_L16 ;
    wire SubBytesIns_Inst_Sbox_12_L15 ;
    wire SubBytesIns_Inst_Sbox_12_L14 ;
    wire SubBytesIns_Inst_Sbox_12_L13 ;
    wire SubBytesIns_Inst_Sbox_12_L12 ;
    wire SubBytesIns_Inst_Sbox_12_L11 ;
    wire SubBytesIns_Inst_Sbox_12_L10 ;
    wire SubBytesIns_Inst_Sbox_12_L9 ;
    wire SubBytesIns_Inst_Sbox_12_L8 ;
    wire SubBytesIns_Inst_Sbox_12_L7 ;
    wire SubBytesIns_Inst_Sbox_12_L6 ;
    wire SubBytesIns_Inst_Sbox_12_L5 ;
    wire SubBytesIns_Inst_Sbox_12_L4 ;
    wire SubBytesIns_Inst_Sbox_12_L3 ;
    wire SubBytesIns_Inst_Sbox_12_L2 ;
    wire SubBytesIns_Inst_Sbox_12_L1 ;
    wire SubBytesIns_Inst_Sbox_12_L0 ;
    wire SubBytesIns_Inst_Sbox_12_M63 ;
    wire SubBytesIns_Inst_Sbox_12_M62 ;
    wire SubBytesIns_Inst_Sbox_12_M61 ;
    wire SubBytesIns_Inst_Sbox_12_M60 ;
    wire SubBytesIns_Inst_Sbox_12_M59 ;
    wire SubBytesIns_Inst_Sbox_12_M58 ;
    wire SubBytesIns_Inst_Sbox_12_M57 ;
    wire SubBytesIns_Inst_Sbox_12_M56 ;
    wire SubBytesIns_Inst_Sbox_12_M55 ;
    wire SubBytesIns_Inst_Sbox_12_M54 ;
    wire SubBytesIns_Inst_Sbox_12_M53 ;
    wire SubBytesIns_Inst_Sbox_12_M52 ;
    wire SubBytesIns_Inst_Sbox_12_M51 ;
    wire SubBytesIns_Inst_Sbox_12_M50 ;
    wire SubBytesIns_Inst_Sbox_12_M49 ;
    wire SubBytesIns_Inst_Sbox_12_M48 ;
    wire SubBytesIns_Inst_Sbox_12_M47 ;
    wire SubBytesIns_Inst_Sbox_12_M46 ;
    wire SubBytesIns_Inst_Sbox_12_M45 ;
    wire SubBytesIns_Inst_Sbox_12_M44 ;
    wire SubBytesIns_Inst_Sbox_12_M43 ;
    wire SubBytesIns_Inst_Sbox_12_M42 ;
    wire SubBytesIns_Inst_Sbox_12_M41 ;
    wire SubBytesIns_Inst_Sbox_12_M40 ;
    wire SubBytesIns_Inst_Sbox_12_M39 ;
    wire SubBytesIns_Inst_Sbox_12_M38 ;
    wire SubBytesIns_Inst_Sbox_12_M37 ;
    wire SubBytesIns_Inst_Sbox_12_M36 ;
    wire SubBytesIns_Inst_Sbox_12_M35 ;
    wire SubBytesIns_Inst_Sbox_12_M34 ;
    wire SubBytesIns_Inst_Sbox_12_M33 ;
    wire SubBytesIns_Inst_Sbox_12_M32 ;
    wire SubBytesIns_Inst_Sbox_12_M31 ;
    wire SubBytesIns_Inst_Sbox_12_M30 ;
    wire SubBytesIns_Inst_Sbox_12_M29 ;
    wire SubBytesIns_Inst_Sbox_12_M28 ;
    wire SubBytesIns_Inst_Sbox_12_M27 ;
    wire SubBytesIns_Inst_Sbox_12_M26 ;
    wire SubBytesIns_Inst_Sbox_12_M25 ;
    wire SubBytesIns_Inst_Sbox_12_M24 ;
    wire SubBytesIns_Inst_Sbox_12_M23 ;
    wire SubBytesIns_Inst_Sbox_12_M22 ;
    wire SubBytesIns_Inst_Sbox_12_M21 ;
    wire SubBytesIns_Inst_Sbox_12_M20 ;
    wire SubBytesIns_Inst_Sbox_12_M19 ;
    wire SubBytesIns_Inst_Sbox_12_M18 ;
    wire SubBytesIns_Inst_Sbox_12_M17 ;
    wire SubBytesIns_Inst_Sbox_12_M16 ;
    wire SubBytesIns_Inst_Sbox_12_M15 ;
    wire SubBytesIns_Inst_Sbox_12_M14 ;
    wire SubBytesIns_Inst_Sbox_12_M13 ;
    wire SubBytesIns_Inst_Sbox_12_M12 ;
    wire SubBytesIns_Inst_Sbox_12_M11 ;
    wire SubBytesIns_Inst_Sbox_12_M10 ;
    wire SubBytesIns_Inst_Sbox_12_M9 ;
    wire SubBytesIns_Inst_Sbox_12_M8 ;
    wire SubBytesIns_Inst_Sbox_12_M7 ;
    wire SubBytesIns_Inst_Sbox_12_M6 ;
    wire SubBytesIns_Inst_Sbox_12_M5 ;
    wire SubBytesIns_Inst_Sbox_12_M4 ;
    wire SubBytesIns_Inst_Sbox_12_M3 ;
    wire SubBytesIns_Inst_Sbox_12_M2 ;
    wire SubBytesIns_Inst_Sbox_12_M1 ;
    wire SubBytesIns_Inst_Sbox_12_T27 ;
    wire SubBytesIns_Inst_Sbox_12_T26 ;
    wire SubBytesIns_Inst_Sbox_12_T25 ;
    wire SubBytesIns_Inst_Sbox_12_T24 ;
    wire SubBytesIns_Inst_Sbox_12_T23 ;
    wire SubBytesIns_Inst_Sbox_12_T22 ;
    wire SubBytesIns_Inst_Sbox_12_T21 ;
    wire SubBytesIns_Inst_Sbox_12_T20 ;
    wire SubBytesIns_Inst_Sbox_12_T19 ;
    wire SubBytesIns_Inst_Sbox_12_T18 ;
    wire SubBytesIns_Inst_Sbox_12_T17 ;
    wire SubBytesIns_Inst_Sbox_12_T16 ;
    wire SubBytesIns_Inst_Sbox_12_T15 ;
    wire SubBytesIns_Inst_Sbox_12_T14 ;
    wire SubBytesIns_Inst_Sbox_12_T13 ;
    wire SubBytesIns_Inst_Sbox_12_T12 ;
    wire SubBytesIns_Inst_Sbox_12_T11 ;
    wire SubBytesIns_Inst_Sbox_12_T10 ;
    wire SubBytesIns_Inst_Sbox_12_T9 ;
    wire SubBytesIns_Inst_Sbox_12_T8 ;
    wire SubBytesIns_Inst_Sbox_12_T7 ;
    wire SubBytesIns_Inst_Sbox_12_T6 ;
    wire SubBytesIns_Inst_Sbox_12_T5 ;
    wire SubBytesIns_Inst_Sbox_12_T4 ;
    wire SubBytesIns_Inst_Sbox_12_T3 ;
    wire SubBytesIns_Inst_Sbox_12_T2 ;
    wire SubBytesIns_Inst_Sbox_12_T1 ;
    wire SubBytesIns_Inst_Sbox_13_L29 ;
    wire SubBytesIns_Inst_Sbox_13_L28 ;
    wire SubBytesIns_Inst_Sbox_13_L27 ;
    wire SubBytesIns_Inst_Sbox_13_L26 ;
    wire SubBytesIns_Inst_Sbox_13_L25 ;
    wire SubBytesIns_Inst_Sbox_13_L24 ;
    wire SubBytesIns_Inst_Sbox_13_L23 ;
    wire SubBytesIns_Inst_Sbox_13_L22 ;
    wire SubBytesIns_Inst_Sbox_13_L21 ;
    wire SubBytesIns_Inst_Sbox_13_L20 ;
    wire SubBytesIns_Inst_Sbox_13_L19 ;
    wire SubBytesIns_Inst_Sbox_13_L18 ;
    wire SubBytesIns_Inst_Sbox_13_L17 ;
    wire SubBytesIns_Inst_Sbox_13_L16 ;
    wire SubBytesIns_Inst_Sbox_13_L15 ;
    wire SubBytesIns_Inst_Sbox_13_L14 ;
    wire SubBytesIns_Inst_Sbox_13_L13 ;
    wire SubBytesIns_Inst_Sbox_13_L12 ;
    wire SubBytesIns_Inst_Sbox_13_L11 ;
    wire SubBytesIns_Inst_Sbox_13_L10 ;
    wire SubBytesIns_Inst_Sbox_13_L9 ;
    wire SubBytesIns_Inst_Sbox_13_L8 ;
    wire SubBytesIns_Inst_Sbox_13_L7 ;
    wire SubBytesIns_Inst_Sbox_13_L6 ;
    wire SubBytesIns_Inst_Sbox_13_L5 ;
    wire SubBytesIns_Inst_Sbox_13_L4 ;
    wire SubBytesIns_Inst_Sbox_13_L3 ;
    wire SubBytesIns_Inst_Sbox_13_L2 ;
    wire SubBytesIns_Inst_Sbox_13_L1 ;
    wire SubBytesIns_Inst_Sbox_13_L0 ;
    wire SubBytesIns_Inst_Sbox_13_M63 ;
    wire SubBytesIns_Inst_Sbox_13_M62 ;
    wire SubBytesIns_Inst_Sbox_13_M61 ;
    wire SubBytesIns_Inst_Sbox_13_M60 ;
    wire SubBytesIns_Inst_Sbox_13_M59 ;
    wire SubBytesIns_Inst_Sbox_13_M58 ;
    wire SubBytesIns_Inst_Sbox_13_M57 ;
    wire SubBytesIns_Inst_Sbox_13_M56 ;
    wire SubBytesIns_Inst_Sbox_13_M55 ;
    wire SubBytesIns_Inst_Sbox_13_M54 ;
    wire SubBytesIns_Inst_Sbox_13_M53 ;
    wire SubBytesIns_Inst_Sbox_13_M52 ;
    wire SubBytesIns_Inst_Sbox_13_M51 ;
    wire SubBytesIns_Inst_Sbox_13_M50 ;
    wire SubBytesIns_Inst_Sbox_13_M49 ;
    wire SubBytesIns_Inst_Sbox_13_M48 ;
    wire SubBytesIns_Inst_Sbox_13_M47 ;
    wire SubBytesIns_Inst_Sbox_13_M46 ;
    wire SubBytesIns_Inst_Sbox_13_M45 ;
    wire SubBytesIns_Inst_Sbox_13_M44 ;
    wire SubBytesIns_Inst_Sbox_13_M43 ;
    wire SubBytesIns_Inst_Sbox_13_M42 ;
    wire SubBytesIns_Inst_Sbox_13_M41 ;
    wire SubBytesIns_Inst_Sbox_13_M40 ;
    wire SubBytesIns_Inst_Sbox_13_M39 ;
    wire SubBytesIns_Inst_Sbox_13_M38 ;
    wire SubBytesIns_Inst_Sbox_13_M37 ;
    wire SubBytesIns_Inst_Sbox_13_M36 ;
    wire SubBytesIns_Inst_Sbox_13_M35 ;
    wire SubBytesIns_Inst_Sbox_13_M34 ;
    wire SubBytesIns_Inst_Sbox_13_M33 ;
    wire SubBytesIns_Inst_Sbox_13_M32 ;
    wire SubBytesIns_Inst_Sbox_13_M31 ;
    wire SubBytesIns_Inst_Sbox_13_M30 ;
    wire SubBytesIns_Inst_Sbox_13_M29 ;
    wire SubBytesIns_Inst_Sbox_13_M28 ;
    wire SubBytesIns_Inst_Sbox_13_M27 ;
    wire SubBytesIns_Inst_Sbox_13_M26 ;
    wire SubBytesIns_Inst_Sbox_13_M25 ;
    wire SubBytesIns_Inst_Sbox_13_M24 ;
    wire SubBytesIns_Inst_Sbox_13_M23 ;
    wire SubBytesIns_Inst_Sbox_13_M22 ;
    wire SubBytesIns_Inst_Sbox_13_M21 ;
    wire SubBytesIns_Inst_Sbox_13_M20 ;
    wire SubBytesIns_Inst_Sbox_13_M19 ;
    wire SubBytesIns_Inst_Sbox_13_M18 ;
    wire SubBytesIns_Inst_Sbox_13_M17 ;
    wire SubBytesIns_Inst_Sbox_13_M16 ;
    wire SubBytesIns_Inst_Sbox_13_M15 ;
    wire SubBytesIns_Inst_Sbox_13_M14 ;
    wire SubBytesIns_Inst_Sbox_13_M13 ;
    wire SubBytesIns_Inst_Sbox_13_M12 ;
    wire SubBytesIns_Inst_Sbox_13_M11 ;
    wire SubBytesIns_Inst_Sbox_13_M10 ;
    wire SubBytesIns_Inst_Sbox_13_M9 ;
    wire SubBytesIns_Inst_Sbox_13_M8 ;
    wire SubBytesIns_Inst_Sbox_13_M7 ;
    wire SubBytesIns_Inst_Sbox_13_M6 ;
    wire SubBytesIns_Inst_Sbox_13_M5 ;
    wire SubBytesIns_Inst_Sbox_13_M4 ;
    wire SubBytesIns_Inst_Sbox_13_M3 ;
    wire SubBytesIns_Inst_Sbox_13_M2 ;
    wire SubBytesIns_Inst_Sbox_13_M1 ;
    wire SubBytesIns_Inst_Sbox_13_T27 ;
    wire SubBytesIns_Inst_Sbox_13_T26 ;
    wire SubBytesIns_Inst_Sbox_13_T25 ;
    wire SubBytesIns_Inst_Sbox_13_T24 ;
    wire SubBytesIns_Inst_Sbox_13_T23 ;
    wire SubBytesIns_Inst_Sbox_13_T22 ;
    wire SubBytesIns_Inst_Sbox_13_T21 ;
    wire SubBytesIns_Inst_Sbox_13_T20 ;
    wire SubBytesIns_Inst_Sbox_13_T19 ;
    wire SubBytesIns_Inst_Sbox_13_T18 ;
    wire SubBytesIns_Inst_Sbox_13_T17 ;
    wire SubBytesIns_Inst_Sbox_13_T16 ;
    wire SubBytesIns_Inst_Sbox_13_T15 ;
    wire SubBytesIns_Inst_Sbox_13_T14 ;
    wire SubBytesIns_Inst_Sbox_13_T13 ;
    wire SubBytesIns_Inst_Sbox_13_T12 ;
    wire SubBytesIns_Inst_Sbox_13_T11 ;
    wire SubBytesIns_Inst_Sbox_13_T10 ;
    wire SubBytesIns_Inst_Sbox_13_T9 ;
    wire SubBytesIns_Inst_Sbox_13_T8 ;
    wire SubBytesIns_Inst_Sbox_13_T7 ;
    wire SubBytesIns_Inst_Sbox_13_T6 ;
    wire SubBytesIns_Inst_Sbox_13_T5 ;
    wire SubBytesIns_Inst_Sbox_13_T4 ;
    wire SubBytesIns_Inst_Sbox_13_T3 ;
    wire SubBytesIns_Inst_Sbox_13_T2 ;
    wire SubBytesIns_Inst_Sbox_13_T1 ;
    wire SubBytesIns_Inst_Sbox_14_L29 ;
    wire SubBytesIns_Inst_Sbox_14_L28 ;
    wire SubBytesIns_Inst_Sbox_14_L27 ;
    wire SubBytesIns_Inst_Sbox_14_L26 ;
    wire SubBytesIns_Inst_Sbox_14_L25 ;
    wire SubBytesIns_Inst_Sbox_14_L24 ;
    wire SubBytesIns_Inst_Sbox_14_L23 ;
    wire SubBytesIns_Inst_Sbox_14_L22 ;
    wire SubBytesIns_Inst_Sbox_14_L21 ;
    wire SubBytesIns_Inst_Sbox_14_L20 ;
    wire SubBytesIns_Inst_Sbox_14_L19 ;
    wire SubBytesIns_Inst_Sbox_14_L18 ;
    wire SubBytesIns_Inst_Sbox_14_L17 ;
    wire SubBytesIns_Inst_Sbox_14_L16 ;
    wire SubBytesIns_Inst_Sbox_14_L15 ;
    wire SubBytesIns_Inst_Sbox_14_L14 ;
    wire SubBytesIns_Inst_Sbox_14_L13 ;
    wire SubBytesIns_Inst_Sbox_14_L12 ;
    wire SubBytesIns_Inst_Sbox_14_L11 ;
    wire SubBytesIns_Inst_Sbox_14_L10 ;
    wire SubBytesIns_Inst_Sbox_14_L9 ;
    wire SubBytesIns_Inst_Sbox_14_L8 ;
    wire SubBytesIns_Inst_Sbox_14_L7 ;
    wire SubBytesIns_Inst_Sbox_14_L6 ;
    wire SubBytesIns_Inst_Sbox_14_L5 ;
    wire SubBytesIns_Inst_Sbox_14_L4 ;
    wire SubBytesIns_Inst_Sbox_14_L3 ;
    wire SubBytesIns_Inst_Sbox_14_L2 ;
    wire SubBytesIns_Inst_Sbox_14_L1 ;
    wire SubBytesIns_Inst_Sbox_14_L0 ;
    wire SubBytesIns_Inst_Sbox_14_M63 ;
    wire SubBytesIns_Inst_Sbox_14_M62 ;
    wire SubBytesIns_Inst_Sbox_14_M61 ;
    wire SubBytesIns_Inst_Sbox_14_M60 ;
    wire SubBytesIns_Inst_Sbox_14_M59 ;
    wire SubBytesIns_Inst_Sbox_14_M58 ;
    wire SubBytesIns_Inst_Sbox_14_M57 ;
    wire SubBytesIns_Inst_Sbox_14_M56 ;
    wire SubBytesIns_Inst_Sbox_14_M55 ;
    wire SubBytesIns_Inst_Sbox_14_M54 ;
    wire SubBytesIns_Inst_Sbox_14_M53 ;
    wire SubBytesIns_Inst_Sbox_14_M52 ;
    wire SubBytesIns_Inst_Sbox_14_M51 ;
    wire SubBytesIns_Inst_Sbox_14_M50 ;
    wire SubBytesIns_Inst_Sbox_14_M49 ;
    wire SubBytesIns_Inst_Sbox_14_M48 ;
    wire SubBytesIns_Inst_Sbox_14_M47 ;
    wire SubBytesIns_Inst_Sbox_14_M46 ;
    wire SubBytesIns_Inst_Sbox_14_M45 ;
    wire SubBytesIns_Inst_Sbox_14_M44 ;
    wire SubBytesIns_Inst_Sbox_14_M43 ;
    wire SubBytesIns_Inst_Sbox_14_M42 ;
    wire SubBytesIns_Inst_Sbox_14_M41 ;
    wire SubBytesIns_Inst_Sbox_14_M40 ;
    wire SubBytesIns_Inst_Sbox_14_M39 ;
    wire SubBytesIns_Inst_Sbox_14_M38 ;
    wire SubBytesIns_Inst_Sbox_14_M37 ;
    wire SubBytesIns_Inst_Sbox_14_M36 ;
    wire SubBytesIns_Inst_Sbox_14_M35 ;
    wire SubBytesIns_Inst_Sbox_14_M34 ;
    wire SubBytesIns_Inst_Sbox_14_M33 ;
    wire SubBytesIns_Inst_Sbox_14_M32 ;
    wire SubBytesIns_Inst_Sbox_14_M31 ;
    wire SubBytesIns_Inst_Sbox_14_M30 ;
    wire SubBytesIns_Inst_Sbox_14_M29 ;
    wire SubBytesIns_Inst_Sbox_14_M28 ;
    wire SubBytesIns_Inst_Sbox_14_M27 ;
    wire SubBytesIns_Inst_Sbox_14_M26 ;
    wire SubBytesIns_Inst_Sbox_14_M25 ;
    wire SubBytesIns_Inst_Sbox_14_M24 ;
    wire SubBytesIns_Inst_Sbox_14_M23 ;
    wire SubBytesIns_Inst_Sbox_14_M22 ;
    wire SubBytesIns_Inst_Sbox_14_M21 ;
    wire SubBytesIns_Inst_Sbox_14_M20 ;
    wire SubBytesIns_Inst_Sbox_14_M19 ;
    wire SubBytesIns_Inst_Sbox_14_M18 ;
    wire SubBytesIns_Inst_Sbox_14_M17 ;
    wire SubBytesIns_Inst_Sbox_14_M16 ;
    wire SubBytesIns_Inst_Sbox_14_M15 ;
    wire SubBytesIns_Inst_Sbox_14_M14 ;
    wire SubBytesIns_Inst_Sbox_14_M13 ;
    wire SubBytesIns_Inst_Sbox_14_M12 ;
    wire SubBytesIns_Inst_Sbox_14_M11 ;
    wire SubBytesIns_Inst_Sbox_14_M10 ;
    wire SubBytesIns_Inst_Sbox_14_M9 ;
    wire SubBytesIns_Inst_Sbox_14_M8 ;
    wire SubBytesIns_Inst_Sbox_14_M7 ;
    wire SubBytesIns_Inst_Sbox_14_M6 ;
    wire SubBytesIns_Inst_Sbox_14_M5 ;
    wire SubBytesIns_Inst_Sbox_14_M4 ;
    wire SubBytesIns_Inst_Sbox_14_M3 ;
    wire SubBytesIns_Inst_Sbox_14_M2 ;
    wire SubBytesIns_Inst_Sbox_14_M1 ;
    wire SubBytesIns_Inst_Sbox_14_T27 ;
    wire SubBytesIns_Inst_Sbox_14_T26 ;
    wire SubBytesIns_Inst_Sbox_14_T25 ;
    wire SubBytesIns_Inst_Sbox_14_T24 ;
    wire SubBytesIns_Inst_Sbox_14_T23 ;
    wire SubBytesIns_Inst_Sbox_14_T22 ;
    wire SubBytesIns_Inst_Sbox_14_T21 ;
    wire SubBytesIns_Inst_Sbox_14_T20 ;
    wire SubBytesIns_Inst_Sbox_14_T19 ;
    wire SubBytesIns_Inst_Sbox_14_T18 ;
    wire SubBytesIns_Inst_Sbox_14_T17 ;
    wire SubBytesIns_Inst_Sbox_14_T16 ;
    wire SubBytesIns_Inst_Sbox_14_T15 ;
    wire SubBytesIns_Inst_Sbox_14_T14 ;
    wire SubBytesIns_Inst_Sbox_14_T13 ;
    wire SubBytesIns_Inst_Sbox_14_T12 ;
    wire SubBytesIns_Inst_Sbox_14_T11 ;
    wire SubBytesIns_Inst_Sbox_14_T10 ;
    wire SubBytesIns_Inst_Sbox_14_T9 ;
    wire SubBytesIns_Inst_Sbox_14_T8 ;
    wire SubBytesIns_Inst_Sbox_14_T7 ;
    wire SubBytesIns_Inst_Sbox_14_T6 ;
    wire SubBytesIns_Inst_Sbox_14_T5 ;
    wire SubBytesIns_Inst_Sbox_14_T4 ;
    wire SubBytesIns_Inst_Sbox_14_T3 ;
    wire SubBytesIns_Inst_Sbox_14_T2 ;
    wire SubBytesIns_Inst_Sbox_14_T1 ;
    wire SubBytesIns_Inst_Sbox_15_L29 ;
    wire SubBytesIns_Inst_Sbox_15_L28 ;
    wire SubBytesIns_Inst_Sbox_15_L27 ;
    wire SubBytesIns_Inst_Sbox_15_L26 ;
    wire SubBytesIns_Inst_Sbox_15_L25 ;
    wire SubBytesIns_Inst_Sbox_15_L24 ;
    wire SubBytesIns_Inst_Sbox_15_L23 ;
    wire SubBytesIns_Inst_Sbox_15_L22 ;
    wire SubBytesIns_Inst_Sbox_15_L21 ;
    wire SubBytesIns_Inst_Sbox_15_L20 ;
    wire SubBytesIns_Inst_Sbox_15_L19 ;
    wire SubBytesIns_Inst_Sbox_15_L18 ;
    wire SubBytesIns_Inst_Sbox_15_L17 ;
    wire SubBytesIns_Inst_Sbox_15_L16 ;
    wire SubBytesIns_Inst_Sbox_15_L15 ;
    wire SubBytesIns_Inst_Sbox_15_L14 ;
    wire SubBytesIns_Inst_Sbox_15_L13 ;
    wire SubBytesIns_Inst_Sbox_15_L12 ;
    wire SubBytesIns_Inst_Sbox_15_L11 ;
    wire SubBytesIns_Inst_Sbox_15_L10 ;
    wire SubBytesIns_Inst_Sbox_15_L9 ;
    wire SubBytesIns_Inst_Sbox_15_L8 ;
    wire SubBytesIns_Inst_Sbox_15_L7 ;
    wire SubBytesIns_Inst_Sbox_15_L6 ;
    wire SubBytesIns_Inst_Sbox_15_L5 ;
    wire SubBytesIns_Inst_Sbox_15_L4 ;
    wire SubBytesIns_Inst_Sbox_15_L3 ;
    wire SubBytesIns_Inst_Sbox_15_L2 ;
    wire SubBytesIns_Inst_Sbox_15_L1 ;
    wire SubBytesIns_Inst_Sbox_15_L0 ;
    wire SubBytesIns_Inst_Sbox_15_M63 ;
    wire SubBytesIns_Inst_Sbox_15_M62 ;
    wire SubBytesIns_Inst_Sbox_15_M61 ;
    wire SubBytesIns_Inst_Sbox_15_M60 ;
    wire SubBytesIns_Inst_Sbox_15_M59 ;
    wire SubBytesIns_Inst_Sbox_15_M58 ;
    wire SubBytesIns_Inst_Sbox_15_M57 ;
    wire SubBytesIns_Inst_Sbox_15_M56 ;
    wire SubBytesIns_Inst_Sbox_15_M55 ;
    wire SubBytesIns_Inst_Sbox_15_M54 ;
    wire SubBytesIns_Inst_Sbox_15_M53 ;
    wire SubBytesIns_Inst_Sbox_15_M52 ;
    wire SubBytesIns_Inst_Sbox_15_M51 ;
    wire SubBytesIns_Inst_Sbox_15_M50 ;
    wire SubBytesIns_Inst_Sbox_15_M49 ;
    wire SubBytesIns_Inst_Sbox_15_M48 ;
    wire SubBytesIns_Inst_Sbox_15_M47 ;
    wire SubBytesIns_Inst_Sbox_15_M46 ;
    wire SubBytesIns_Inst_Sbox_15_M45 ;
    wire SubBytesIns_Inst_Sbox_15_M44 ;
    wire SubBytesIns_Inst_Sbox_15_M43 ;
    wire SubBytesIns_Inst_Sbox_15_M42 ;
    wire SubBytesIns_Inst_Sbox_15_M41 ;
    wire SubBytesIns_Inst_Sbox_15_M40 ;
    wire SubBytesIns_Inst_Sbox_15_M39 ;
    wire SubBytesIns_Inst_Sbox_15_M38 ;
    wire SubBytesIns_Inst_Sbox_15_M37 ;
    wire SubBytesIns_Inst_Sbox_15_M36 ;
    wire SubBytesIns_Inst_Sbox_15_M35 ;
    wire SubBytesIns_Inst_Sbox_15_M34 ;
    wire SubBytesIns_Inst_Sbox_15_M33 ;
    wire SubBytesIns_Inst_Sbox_15_M32 ;
    wire SubBytesIns_Inst_Sbox_15_M31 ;
    wire SubBytesIns_Inst_Sbox_15_M30 ;
    wire SubBytesIns_Inst_Sbox_15_M29 ;
    wire SubBytesIns_Inst_Sbox_15_M28 ;
    wire SubBytesIns_Inst_Sbox_15_M27 ;
    wire SubBytesIns_Inst_Sbox_15_M26 ;
    wire SubBytesIns_Inst_Sbox_15_M25 ;
    wire SubBytesIns_Inst_Sbox_15_M24 ;
    wire SubBytesIns_Inst_Sbox_15_M23 ;
    wire SubBytesIns_Inst_Sbox_15_M22 ;
    wire SubBytesIns_Inst_Sbox_15_M21 ;
    wire SubBytesIns_Inst_Sbox_15_M20 ;
    wire SubBytesIns_Inst_Sbox_15_M19 ;
    wire SubBytesIns_Inst_Sbox_15_M18 ;
    wire SubBytesIns_Inst_Sbox_15_M17 ;
    wire SubBytesIns_Inst_Sbox_15_M16 ;
    wire SubBytesIns_Inst_Sbox_15_M15 ;
    wire SubBytesIns_Inst_Sbox_15_M14 ;
    wire SubBytesIns_Inst_Sbox_15_M13 ;
    wire SubBytesIns_Inst_Sbox_15_M12 ;
    wire SubBytesIns_Inst_Sbox_15_M11 ;
    wire SubBytesIns_Inst_Sbox_15_M10 ;
    wire SubBytesIns_Inst_Sbox_15_M9 ;
    wire SubBytesIns_Inst_Sbox_15_M8 ;
    wire SubBytesIns_Inst_Sbox_15_M7 ;
    wire SubBytesIns_Inst_Sbox_15_M6 ;
    wire SubBytesIns_Inst_Sbox_15_M5 ;
    wire SubBytesIns_Inst_Sbox_15_M4 ;
    wire SubBytesIns_Inst_Sbox_15_M3 ;
    wire SubBytesIns_Inst_Sbox_15_M2 ;
    wire SubBytesIns_Inst_Sbox_15_M1 ;
    wire SubBytesIns_Inst_Sbox_15_T27 ;
    wire SubBytesIns_Inst_Sbox_15_T26 ;
    wire SubBytesIns_Inst_Sbox_15_T25 ;
    wire SubBytesIns_Inst_Sbox_15_T24 ;
    wire SubBytesIns_Inst_Sbox_15_T23 ;
    wire SubBytesIns_Inst_Sbox_15_T22 ;
    wire SubBytesIns_Inst_Sbox_15_T21 ;
    wire SubBytesIns_Inst_Sbox_15_T20 ;
    wire SubBytesIns_Inst_Sbox_15_T19 ;
    wire SubBytesIns_Inst_Sbox_15_T18 ;
    wire SubBytesIns_Inst_Sbox_15_T17 ;
    wire SubBytesIns_Inst_Sbox_15_T16 ;
    wire SubBytesIns_Inst_Sbox_15_T15 ;
    wire SubBytesIns_Inst_Sbox_15_T14 ;
    wire SubBytesIns_Inst_Sbox_15_T13 ;
    wire SubBytesIns_Inst_Sbox_15_T12 ;
    wire SubBytesIns_Inst_Sbox_15_T11 ;
    wire SubBytesIns_Inst_Sbox_15_T10 ;
    wire SubBytesIns_Inst_Sbox_15_T9 ;
    wire SubBytesIns_Inst_Sbox_15_T8 ;
    wire SubBytesIns_Inst_Sbox_15_T7 ;
    wire SubBytesIns_Inst_Sbox_15_T6 ;
    wire SubBytesIns_Inst_Sbox_15_T5 ;
    wire SubBytesIns_Inst_Sbox_15_T4 ;
    wire SubBytesIns_Inst_Sbox_15_T3 ;
    wire SubBytesIns_Inst_Sbox_15_T2 ;
    wire SubBytesIns_Inst_Sbox_15_T1 ;
    wire MixColumnsIns_MixOneColumnInst_0_n64 ;
    wire MixColumnsIns_MixOneColumnInst_0_n63 ;
    wire MixColumnsIns_MixOneColumnInst_0_n62 ;
    wire MixColumnsIns_MixOneColumnInst_0_n61 ;
    wire MixColumnsIns_MixOneColumnInst_0_n60 ;
    wire MixColumnsIns_MixOneColumnInst_0_n59 ;
    wire MixColumnsIns_MixOneColumnInst_0_n58 ;
    wire MixColumnsIns_MixOneColumnInst_0_n57 ;
    wire MixColumnsIns_MixOneColumnInst_0_n56 ;
    wire MixColumnsIns_MixOneColumnInst_0_n55 ;
    wire MixColumnsIns_MixOneColumnInst_0_n54 ;
    wire MixColumnsIns_MixOneColumnInst_0_n53 ;
    wire MixColumnsIns_MixOneColumnInst_0_n52 ;
    wire MixColumnsIns_MixOneColumnInst_0_n51 ;
    wire MixColumnsIns_MixOneColumnInst_0_n50 ;
    wire MixColumnsIns_MixOneColumnInst_0_n49 ;
    wire MixColumnsIns_MixOneColumnInst_0_n48 ;
    wire MixColumnsIns_MixOneColumnInst_0_n47 ;
    wire MixColumnsIns_MixOneColumnInst_0_n46 ;
    wire MixColumnsIns_MixOneColumnInst_0_n45 ;
    wire MixColumnsIns_MixOneColumnInst_0_n44 ;
    wire MixColumnsIns_MixOneColumnInst_0_n43 ;
    wire MixColumnsIns_MixOneColumnInst_0_n42 ;
    wire MixColumnsIns_MixOneColumnInst_0_n41 ;
    wire MixColumnsIns_MixOneColumnInst_0_n40 ;
    wire MixColumnsIns_MixOneColumnInst_0_n39 ;
    wire MixColumnsIns_MixOneColumnInst_0_n38 ;
    wire MixColumnsIns_MixOneColumnInst_0_n37 ;
    wire MixColumnsIns_MixOneColumnInst_0_n36 ;
    wire MixColumnsIns_MixOneColumnInst_0_n35 ;
    wire MixColumnsIns_MixOneColumnInst_0_n34 ;
    wire MixColumnsIns_MixOneColumnInst_0_n33 ;
    wire MixColumnsIns_MixOneColumnInst_0_n32 ;
    wire MixColumnsIns_MixOneColumnInst_0_n31 ;
    wire MixColumnsIns_MixOneColumnInst_0_n30 ;
    wire MixColumnsIns_MixOneColumnInst_0_n29 ;
    wire MixColumnsIns_MixOneColumnInst_0_n28 ;
    wire MixColumnsIns_MixOneColumnInst_0_n27 ;
    wire MixColumnsIns_MixOneColumnInst_0_n26 ;
    wire MixColumnsIns_MixOneColumnInst_0_n25 ;
    wire MixColumnsIns_MixOneColumnInst_0_n24 ;
    wire MixColumnsIns_MixOneColumnInst_0_n23 ;
    wire MixColumnsIns_MixOneColumnInst_0_n22 ;
    wire MixColumnsIns_MixOneColumnInst_0_n21 ;
    wire MixColumnsIns_MixOneColumnInst_0_n20 ;
    wire MixColumnsIns_MixOneColumnInst_0_n19 ;
    wire MixColumnsIns_MixOneColumnInst_0_n18 ;
    wire MixColumnsIns_MixOneColumnInst_0_n17 ;
    wire MixColumnsIns_MixOneColumnInst_0_n16 ;
    wire MixColumnsIns_MixOneColumnInst_0_n15 ;
    wire MixColumnsIns_MixOneColumnInst_0_n14 ;
    wire MixColumnsIns_MixOneColumnInst_0_n13 ;
    wire MixColumnsIns_MixOneColumnInst_0_n12 ;
    wire MixColumnsIns_MixOneColumnInst_0_n11 ;
    wire MixColumnsIns_MixOneColumnInst_0_n10 ;
    wire MixColumnsIns_MixOneColumnInst_0_n9 ;
    wire MixColumnsIns_MixOneColumnInst_0_n8 ;
    wire MixColumnsIns_MixOneColumnInst_0_n7 ;
    wire MixColumnsIns_MixOneColumnInst_0_n6 ;
    wire MixColumnsIns_MixOneColumnInst_0_n5 ;
    wire MixColumnsIns_MixOneColumnInst_0_n4 ;
    wire MixColumnsIns_MixOneColumnInst_0_n3 ;
    wire MixColumnsIns_MixOneColumnInst_0_n2 ;
    wire MixColumnsIns_MixOneColumnInst_0_n1 ;
    wire MixColumnsIns_MixOneColumnInst_1_n64 ;
    wire MixColumnsIns_MixOneColumnInst_1_n63 ;
    wire MixColumnsIns_MixOneColumnInst_1_n62 ;
    wire MixColumnsIns_MixOneColumnInst_1_n61 ;
    wire MixColumnsIns_MixOneColumnInst_1_n60 ;
    wire MixColumnsIns_MixOneColumnInst_1_n59 ;
    wire MixColumnsIns_MixOneColumnInst_1_n58 ;
    wire MixColumnsIns_MixOneColumnInst_1_n57 ;
    wire MixColumnsIns_MixOneColumnInst_1_n56 ;
    wire MixColumnsIns_MixOneColumnInst_1_n55 ;
    wire MixColumnsIns_MixOneColumnInst_1_n54 ;
    wire MixColumnsIns_MixOneColumnInst_1_n53 ;
    wire MixColumnsIns_MixOneColumnInst_1_n52 ;
    wire MixColumnsIns_MixOneColumnInst_1_n51 ;
    wire MixColumnsIns_MixOneColumnInst_1_n50 ;
    wire MixColumnsIns_MixOneColumnInst_1_n49 ;
    wire MixColumnsIns_MixOneColumnInst_1_n48 ;
    wire MixColumnsIns_MixOneColumnInst_1_n47 ;
    wire MixColumnsIns_MixOneColumnInst_1_n46 ;
    wire MixColumnsIns_MixOneColumnInst_1_n45 ;
    wire MixColumnsIns_MixOneColumnInst_1_n44 ;
    wire MixColumnsIns_MixOneColumnInst_1_n43 ;
    wire MixColumnsIns_MixOneColumnInst_1_n42 ;
    wire MixColumnsIns_MixOneColumnInst_1_n41 ;
    wire MixColumnsIns_MixOneColumnInst_1_n40 ;
    wire MixColumnsIns_MixOneColumnInst_1_n39 ;
    wire MixColumnsIns_MixOneColumnInst_1_n38 ;
    wire MixColumnsIns_MixOneColumnInst_1_n37 ;
    wire MixColumnsIns_MixOneColumnInst_1_n36 ;
    wire MixColumnsIns_MixOneColumnInst_1_n35 ;
    wire MixColumnsIns_MixOneColumnInst_1_n34 ;
    wire MixColumnsIns_MixOneColumnInst_1_n33 ;
    wire MixColumnsIns_MixOneColumnInst_1_n32 ;
    wire MixColumnsIns_MixOneColumnInst_1_n31 ;
    wire MixColumnsIns_MixOneColumnInst_1_n30 ;
    wire MixColumnsIns_MixOneColumnInst_1_n29 ;
    wire MixColumnsIns_MixOneColumnInst_1_n28 ;
    wire MixColumnsIns_MixOneColumnInst_1_n27 ;
    wire MixColumnsIns_MixOneColumnInst_1_n26 ;
    wire MixColumnsIns_MixOneColumnInst_1_n25 ;
    wire MixColumnsIns_MixOneColumnInst_1_n24 ;
    wire MixColumnsIns_MixOneColumnInst_1_n23 ;
    wire MixColumnsIns_MixOneColumnInst_1_n22 ;
    wire MixColumnsIns_MixOneColumnInst_1_n21 ;
    wire MixColumnsIns_MixOneColumnInst_1_n20 ;
    wire MixColumnsIns_MixOneColumnInst_1_n19 ;
    wire MixColumnsIns_MixOneColumnInst_1_n18 ;
    wire MixColumnsIns_MixOneColumnInst_1_n17 ;
    wire MixColumnsIns_MixOneColumnInst_1_n16 ;
    wire MixColumnsIns_MixOneColumnInst_1_n15 ;
    wire MixColumnsIns_MixOneColumnInst_1_n14 ;
    wire MixColumnsIns_MixOneColumnInst_1_n13 ;
    wire MixColumnsIns_MixOneColumnInst_1_n12 ;
    wire MixColumnsIns_MixOneColumnInst_1_n11 ;
    wire MixColumnsIns_MixOneColumnInst_1_n10 ;
    wire MixColumnsIns_MixOneColumnInst_1_n9 ;
    wire MixColumnsIns_MixOneColumnInst_1_n8 ;
    wire MixColumnsIns_MixOneColumnInst_1_n7 ;
    wire MixColumnsIns_MixOneColumnInst_1_n6 ;
    wire MixColumnsIns_MixOneColumnInst_1_n5 ;
    wire MixColumnsIns_MixOneColumnInst_1_n4 ;
    wire MixColumnsIns_MixOneColumnInst_1_n3 ;
    wire MixColumnsIns_MixOneColumnInst_1_n2 ;
    wire MixColumnsIns_MixOneColumnInst_1_n1 ;
    wire MixColumnsIns_MixOneColumnInst_2_n64 ;
    wire MixColumnsIns_MixOneColumnInst_2_n63 ;
    wire MixColumnsIns_MixOneColumnInst_2_n62 ;
    wire MixColumnsIns_MixOneColumnInst_2_n61 ;
    wire MixColumnsIns_MixOneColumnInst_2_n60 ;
    wire MixColumnsIns_MixOneColumnInst_2_n59 ;
    wire MixColumnsIns_MixOneColumnInst_2_n58 ;
    wire MixColumnsIns_MixOneColumnInst_2_n57 ;
    wire MixColumnsIns_MixOneColumnInst_2_n56 ;
    wire MixColumnsIns_MixOneColumnInst_2_n55 ;
    wire MixColumnsIns_MixOneColumnInst_2_n54 ;
    wire MixColumnsIns_MixOneColumnInst_2_n53 ;
    wire MixColumnsIns_MixOneColumnInst_2_n52 ;
    wire MixColumnsIns_MixOneColumnInst_2_n51 ;
    wire MixColumnsIns_MixOneColumnInst_2_n50 ;
    wire MixColumnsIns_MixOneColumnInst_2_n49 ;
    wire MixColumnsIns_MixOneColumnInst_2_n48 ;
    wire MixColumnsIns_MixOneColumnInst_2_n47 ;
    wire MixColumnsIns_MixOneColumnInst_2_n46 ;
    wire MixColumnsIns_MixOneColumnInst_2_n45 ;
    wire MixColumnsIns_MixOneColumnInst_2_n44 ;
    wire MixColumnsIns_MixOneColumnInst_2_n43 ;
    wire MixColumnsIns_MixOneColumnInst_2_n42 ;
    wire MixColumnsIns_MixOneColumnInst_2_n41 ;
    wire MixColumnsIns_MixOneColumnInst_2_n40 ;
    wire MixColumnsIns_MixOneColumnInst_2_n39 ;
    wire MixColumnsIns_MixOneColumnInst_2_n38 ;
    wire MixColumnsIns_MixOneColumnInst_2_n37 ;
    wire MixColumnsIns_MixOneColumnInst_2_n36 ;
    wire MixColumnsIns_MixOneColumnInst_2_n35 ;
    wire MixColumnsIns_MixOneColumnInst_2_n34 ;
    wire MixColumnsIns_MixOneColumnInst_2_n33 ;
    wire MixColumnsIns_MixOneColumnInst_2_n32 ;
    wire MixColumnsIns_MixOneColumnInst_2_n31 ;
    wire MixColumnsIns_MixOneColumnInst_2_n30 ;
    wire MixColumnsIns_MixOneColumnInst_2_n29 ;
    wire MixColumnsIns_MixOneColumnInst_2_n28 ;
    wire MixColumnsIns_MixOneColumnInst_2_n27 ;
    wire MixColumnsIns_MixOneColumnInst_2_n26 ;
    wire MixColumnsIns_MixOneColumnInst_2_n25 ;
    wire MixColumnsIns_MixOneColumnInst_2_n24 ;
    wire MixColumnsIns_MixOneColumnInst_2_n23 ;
    wire MixColumnsIns_MixOneColumnInst_2_n22 ;
    wire MixColumnsIns_MixOneColumnInst_2_n21 ;
    wire MixColumnsIns_MixOneColumnInst_2_n20 ;
    wire MixColumnsIns_MixOneColumnInst_2_n19 ;
    wire MixColumnsIns_MixOneColumnInst_2_n18 ;
    wire MixColumnsIns_MixOneColumnInst_2_n17 ;
    wire MixColumnsIns_MixOneColumnInst_2_n16 ;
    wire MixColumnsIns_MixOneColumnInst_2_n15 ;
    wire MixColumnsIns_MixOneColumnInst_2_n14 ;
    wire MixColumnsIns_MixOneColumnInst_2_n13 ;
    wire MixColumnsIns_MixOneColumnInst_2_n12 ;
    wire MixColumnsIns_MixOneColumnInst_2_n11 ;
    wire MixColumnsIns_MixOneColumnInst_2_n10 ;
    wire MixColumnsIns_MixOneColumnInst_2_n9 ;
    wire MixColumnsIns_MixOneColumnInst_2_n8 ;
    wire MixColumnsIns_MixOneColumnInst_2_n7 ;
    wire MixColumnsIns_MixOneColumnInst_2_n6 ;
    wire MixColumnsIns_MixOneColumnInst_2_n5 ;
    wire MixColumnsIns_MixOneColumnInst_2_n4 ;
    wire MixColumnsIns_MixOneColumnInst_2_n3 ;
    wire MixColumnsIns_MixOneColumnInst_2_n2 ;
    wire MixColumnsIns_MixOneColumnInst_2_n1 ;
    wire MixColumnsIns_MixOneColumnInst_3_n64 ;
    wire MixColumnsIns_MixOneColumnInst_3_n63 ;
    wire MixColumnsIns_MixOneColumnInst_3_n62 ;
    wire MixColumnsIns_MixOneColumnInst_3_n61 ;
    wire MixColumnsIns_MixOneColumnInst_3_n60 ;
    wire MixColumnsIns_MixOneColumnInst_3_n59 ;
    wire MixColumnsIns_MixOneColumnInst_3_n58 ;
    wire MixColumnsIns_MixOneColumnInst_3_n57 ;
    wire MixColumnsIns_MixOneColumnInst_3_n56 ;
    wire MixColumnsIns_MixOneColumnInst_3_n55 ;
    wire MixColumnsIns_MixOneColumnInst_3_n54 ;
    wire MixColumnsIns_MixOneColumnInst_3_n53 ;
    wire MixColumnsIns_MixOneColumnInst_3_n52 ;
    wire MixColumnsIns_MixOneColumnInst_3_n51 ;
    wire MixColumnsIns_MixOneColumnInst_3_n50 ;
    wire MixColumnsIns_MixOneColumnInst_3_n49 ;
    wire MixColumnsIns_MixOneColumnInst_3_n48 ;
    wire MixColumnsIns_MixOneColumnInst_3_n47 ;
    wire MixColumnsIns_MixOneColumnInst_3_n46 ;
    wire MixColumnsIns_MixOneColumnInst_3_n45 ;
    wire MixColumnsIns_MixOneColumnInst_3_n44 ;
    wire MixColumnsIns_MixOneColumnInst_3_n43 ;
    wire MixColumnsIns_MixOneColumnInst_3_n42 ;
    wire MixColumnsIns_MixOneColumnInst_3_n41 ;
    wire MixColumnsIns_MixOneColumnInst_3_n40 ;
    wire MixColumnsIns_MixOneColumnInst_3_n39 ;
    wire MixColumnsIns_MixOneColumnInst_3_n38 ;
    wire MixColumnsIns_MixOneColumnInst_3_n37 ;
    wire MixColumnsIns_MixOneColumnInst_3_n36 ;
    wire MixColumnsIns_MixOneColumnInst_3_n35 ;
    wire MixColumnsIns_MixOneColumnInst_3_n34 ;
    wire MixColumnsIns_MixOneColumnInst_3_n33 ;
    wire MixColumnsIns_MixOneColumnInst_3_n32 ;
    wire MixColumnsIns_MixOneColumnInst_3_n31 ;
    wire MixColumnsIns_MixOneColumnInst_3_n30 ;
    wire MixColumnsIns_MixOneColumnInst_3_n29 ;
    wire MixColumnsIns_MixOneColumnInst_3_n28 ;
    wire MixColumnsIns_MixOneColumnInst_3_n27 ;
    wire MixColumnsIns_MixOneColumnInst_3_n26 ;
    wire MixColumnsIns_MixOneColumnInst_3_n25 ;
    wire MixColumnsIns_MixOneColumnInst_3_n24 ;
    wire MixColumnsIns_MixOneColumnInst_3_n23 ;
    wire MixColumnsIns_MixOneColumnInst_3_n22 ;
    wire MixColumnsIns_MixOneColumnInst_3_n21 ;
    wire MixColumnsIns_MixOneColumnInst_3_n20 ;
    wire MixColumnsIns_MixOneColumnInst_3_n19 ;
    wire MixColumnsIns_MixOneColumnInst_3_n18 ;
    wire MixColumnsIns_MixOneColumnInst_3_n17 ;
    wire MixColumnsIns_MixOneColumnInst_3_n16 ;
    wire MixColumnsIns_MixOneColumnInst_3_n15 ;
    wire MixColumnsIns_MixOneColumnInst_3_n14 ;
    wire MixColumnsIns_MixOneColumnInst_3_n13 ;
    wire MixColumnsIns_MixOneColumnInst_3_n12 ;
    wire MixColumnsIns_MixOneColumnInst_3_n11 ;
    wire MixColumnsIns_MixOneColumnInst_3_n10 ;
    wire MixColumnsIns_MixOneColumnInst_3_n9 ;
    wire MixColumnsIns_MixOneColumnInst_3_n8 ;
    wire MixColumnsIns_MixOneColumnInst_3_n7 ;
    wire MixColumnsIns_MixOneColumnInst_3_n6 ;
    wire MixColumnsIns_MixOneColumnInst_3_n5 ;
    wire MixColumnsIns_MixOneColumnInst_3_n4 ;
    wire MixColumnsIns_MixOneColumnInst_3_n3 ;
    wire MixColumnsIns_MixOneColumnInst_3_n2 ;
    wire MixColumnsIns_MixOneColumnInst_3_n1 ;
    wire KeyReg_Inst_ff_SDE_0_next_state ;
    wire KeyReg_Inst_ff_SDE_1_next_state ;
    wire KeyReg_Inst_ff_SDE_2_next_state ;
    wire KeyReg_Inst_ff_SDE_3_next_state ;
    wire KeyReg_Inst_ff_SDE_4_next_state ;
    wire KeyReg_Inst_ff_SDE_5_next_state ;
    wire KeyReg_Inst_ff_SDE_6_next_state ;
    wire KeyReg_Inst_ff_SDE_7_next_state ;
    wire KeyReg_Inst_ff_SDE_8_next_state ;
    wire KeyReg_Inst_ff_SDE_9_next_state ;
    wire KeyReg_Inst_ff_SDE_10_next_state ;
    wire KeyReg_Inst_ff_SDE_11_next_state ;
    wire KeyReg_Inst_ff_SDE_12_next_state ;
    wire KeyReg_Inst_ff_SDE_13_next_state ;
    wire KeyReg_Inst_ff_SDE_14_next_state ;
    wire KeyReg_Inst_ff_SDE_15_next_state ;
    wire KeyReg_Inst_ff_SDE_16_next_state ;
    wire KeyReg_Inst_ff_SDE_17_next_state ;
    wire KeyReg_Inst_ff_SDE_18_next_state ;
    wire KeyReg_Inst_ff_SDE_19_next_state ;
    wire KeyReg_Inst_ff_SDE_20_next_state ;
    wire KeyReg_Inst_ff_SDE_21_next_state ;
    wire KeyReg_Inst_ff_SDE_22_next_state ;
    wire KeyReg_Inst_ff_SDE_23_next_state ;
    wire KeyReg_Inst_ff_SDE_24_next_state ;
    wire KeyReg_Inst_ff_SDE_25_next_state ;
    wire KeyReg_Inst_ff_SDE_26_next_state ;
    wire KeyReg_Inst_ff_SDE_27_next_state ;
    wire KeyReg_Inst_ff_SDE_28_next_state ;
    wire KeyReg_Inst_ff_SDE_29_next_state ;
    wire KeyReg_Inst_ff_SDE_30_next_state ;
    wire KeyReg_Inst_ff_SDE_31_next_state ;
    wire KeyReg_Inst_ff_SDE_32_next_state ;
    wire KeyReg_Inst_ff_SDE_33_next_state ;
    wire KeyReg_Inst_ff_SDE_34_next_state ;
    wire KeyReg_Inst_ff_SDE_35_next_state ;
    wire KeyReg_Inst_ff_SDE_36_next_state ;
    wire KeyReg_Inst_ff_SDE_37_next_state ;
    wire KeyReg_Inst_ff_SDE_38_next_state ;
    wire KeyReg_Inst_ff_SDE_39_next_state ;
    wire KeyReg_Inst_ff_SDE_40_next_state ;
    wire KeyReg_Inst_ff_SDE_41_next_state ;
    wire KeyReg_Inst_ff_SDE_42_next_state ;
    wire KeyReg_Inst_ff_SDE_43_next_state ;
    wire KeyReg_Inst_ff_SDE_44_next_state ;
    wire KeyReg_Inst_ff_SDE_45_next_state ;
    wire KeyReg_Inst_ff_SDE_46_next_state ;
    wire KeyReg_Inst_ff_SDE_47_next_state ;
    wire KeyReg_Inst_ff_SDE_48_next_state ;
    wire KeyReg_Inst_ff_SDE_49_next_state ;
    wire KeyReg_Inst_ff_SDE_50_next_state ;
    wire KeyReg_Inst_ff_SDE_51_next_state ;
    wire KeyReg_Inst_ff_SDE_52_next_state ;
    wire KeyReg_Inst_ff_SDE_53_next_state ;
    wire KeyReg_Inst_ff_SDE_54_next_state ;
    wire KeyReg_Inst_ff_SDE_55_next_state ;
    wire KeyReg_Inst_ff_SDE_56_next_state ;
    wire KeyReg_Inst_ff_SDE_57_next_state ;
    wire KeyReg_Inst_ff_SDE_58_next_state ;
    wire KeyReg_Inst_ff_SDE_59_next_state ;
    wire KeyReg_Inst_ff_SDE_60_next_state ;
    wire KeyReg_Inst_ff_SDE_61_next_state ;
    wire KeyReg_Inst_ff_SDE_62_next_state ;
    wire KeyReg_Inst_ff_SDE_63_next_state ;
    wire KeyReg_Inst_ff_SDE_64_next_state ;
    wire KeyReg_Inst_ff_SDE_65_next_state ;
    wire KeyReg_Inst_ff_SDE_66_next_state ;
    wire KeyReg_Inst_ff_SDE_67_next_state ;
    wire KeyReg_Inst_ff_SDE_68_next_state ;
    wire KeyReg_Inst_ff_SDE_69_next_state ;
    wire KeyReg_Inst_ff_SDE_70_next_state ;
    wire KeyReg_Inst_ff_SDE_71_next_state ;
    wire KeyReg_Inst_ff_SDE_72_next_state ;
    wire KeyReg_Inst_ff_SDE_73_next_state ;
    wire KeyReg_Inst_ff_SDE_74_next_state ;
    wire KeyReg_Inst_ff_SDE_75_next_state ;
    wire KeyReg_Inst_ff_SDE_76_next_state ;
    wire KeyReg_Inst_ff_SDE_77_next_state ;
    wire KeyReg_Inst_ff_SDE_78_next_state ;
    wire KeyReg_Inst_ff_SDE_79_next_state ;
    wire KeyReg_Inst_ff_SDE_80_next_state ;
    wire KeyReg_Inst_ff_SDE_81_next_state ;
    wire KeyReg_Inst_ff_SDE_82_next_state ;
    wire KeyReg_Inst_ff_SDE_83_next_state ;
    wire KeyReg_Inst_ff_SDE_84_next_state ;
    wire KeyReg_Inst_ff_SDE_85_next_state ;
    wire KeyReg_Inst_ff_SDE_86_next_state ;
    wire KeyReg_Inst_ff_SDE_87_next_state ;
    wire KeyReg_Inst_ff_SDE_88_next_state ;
    wire KeyReg_Inst_ff_SDE_89_next_state ;
    wire KeyReg_Inst_ff_SDE_90_next_state ;
    wire KeyReg_Inst_ff_SDE_91_next_state ;
    wire KeyReg_Inst_ff_SDE_92_next_state ;
    wire KeyReg_Inst_ff_SDE_93_next_state ;
    wire KeyReg_Inst_ff_SDE_94_next_state ;
    wire KeyReg_Inst_ff_SDE_95_next_state ;
    wire KeyReg_Inst_ff_SDE_96_next_state ;
    wire KeyReg_Inst_ff_SDE_97_next_state ;
    wire KeyReg_Inst_ff_SDE_98_next_state ;
    wire KeyReg_Inst_ff_SDE_99_next_state ;
    wire KeyReg_Inst_ff_SDE_100_next_state ;
    wire KeyReg_Inst_ff_SDE_101_next_state ;
    wire KeyReg_Inst_ff_SDE_102_next_state ;
    wire KeyReg_Inst_ff_SDE_103_next_state ;
    wire KeyReg_Inst_ff_SDE_104_next_state ;
    wire KeyReg_Inst_ff_SDE_105_next_state ;
    wire KeyReg_Inst_ff_SDE_106_next_state ;
    wire KeyReg_Inst_ff_SDE_107_next_state ;
    wire KeyReg_Inst_ff_SDE_108_next_state ;
    wire KeyReg_Inst_ff_SDE_109_next_state ;
    wire KeyReg_Inst_ff_SDE_110_next_state ;
    wire KeyReg_Inst_ff_SDE_111_next_state ;
    wire KeyReg_Inst_ff_SDE_112_next_state ;
    wire KeyReg_Inst_ff_SDE_113_next_state ;
    wire KeyReg_Inst_ff_SDE_114_next_state ;
    wire KeyReg_Inst_ff_SDE_115_next_state ;
    wire KeyReg_Inst_ff_SDE_116_next_state ;
    wire KeyReg_Inst_ff_SDE_117_next_state ;
    wire KeyReg_Inst_ff_SDE_118_next_state ;
    wire KeyReg_Inst_ff_SDE_119_next_state ;
    wire KeyReg_Inst_ff_SDE_120_next_state ;
    wire KeyReg_Inst_ff_SDE_121_next_state ;
    wire KeyReg_Inst_ff_SDE_122_next_state ;
    wire KeyReg_Inst_ff_SDE_123_next_state ;
    wire KeyReg_Inst_ff_SDE_124_next_state ;
    wire KeyReg_Inst_ff_SDE_125_next_state ;
    wire KeyReg_Inst_ff_SDE_126_next_state ;
    wire KeyReg_Inst_ff_SDE_127_next_state ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_ ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1 ;
    wire RoundCounterIns_n13 ;
    wire RoundCounterIns_n12 ;
    wire RoundCounterIns_n11 ;
    wire RoundCounterIns_n10 ;
    wire RoundCounterIns_n9 ;
    wire RoundCounterIns_n8 ;
    wire RoundCounterIns_n7 ;
    wire RoundCounterIns_n4 ;
    wire RoundCounterIns_n3 ;
    wire RoundCounterIns_n2 ;
    wire RoundCounterIns_n1 ;
    wire RoundCounterIns_N10 ;
    wire RoundCounterIns_n5 ;
    wire RoundCounterIns_N8 ;
    wire RoundCounterIns_n6 ;
    wire RoundCounterIns_N7 ;
    wire [127:0] RoundOutput ;
    wire [127:0] RoundInput ;
    wire [123:0] MixColumnsInput ;
    wire [127:0] MixColumnsOutput ;
    wire [127:0] KeyExpansionOutput ;
    wire [127:0] RoundKey ;
    wire [5:0] Rcon ;
    wire [3:0] RoundCounter ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_0_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_1_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_2_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_3_DoubleBytes ;
    wire [31:0] KeyExpansionIns_tmp ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5195 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5202 ;
    wire new_AGEMA_signal_5203 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5207 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5213 ;
    wire new_AGEMA_signal_5214 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5219 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5226 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5231 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5238 ;
    wire new_AGEMA_signal_5239 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5249 ;
    wire new_AGEMA_signal_5250 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5255 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5262 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5273 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5291 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5303 ;
    wire new_AGEMA_signal_5304 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5309 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6654 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;
    wire new_AGEMA_signal_6672 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6677 ;
    wire new_AGEMA_signal_6678 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6682 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6688 ;
    wire new_AGEMA_signal_6689 ;
    wire new_AGEMA_signal_6690 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6695 ;
    wire new_AGEMA_signal_6696 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6700 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6706 ;
    wire new_AGEMA_signal_6707 ;
    wire new_AGEMA_signal_6708 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6713 ;
    wire new_AGEMA_signal_6714 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6718 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6724 ;
    wire new_AGEMA_signal_6725 ;
    wire new_AGEMA_signal_6726 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7036 ;
    wire new_AGEMA_signal_7037 ;
    wire new_AGEMA_signal_7038 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7042 ;
    wire new_AGEMA_signal_7043 ;
    wire new_AGEMA_signal_7044 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7048 ;
    wire new_AGEMA_signal_7049 ;
    wire new_AGEMA_signal_7050 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7054 ;
    wire new_AGEMA_signal_7055 ;
    wire new_AGEMA_signal_7056 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7060 ;
    wire new_AGEMA_signal_7061 ;
    wire new_AGEMA_signal_7062 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7066 ;
    wire new_AGEMA_signal_7067 ;
    wire new_AGEMA_signal_7068 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7072 ;
    wire new_AGEMA_signal_7073 ;
    wire new_AGEMA_signal_7074 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7078 ;
    wire new_AGEMA_signal_7079 ;
    wire new_AGEMA_signal_7080 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7084 ;
    wire new_AGEMA_signal_7085 ;
    wire new_AGEMA_signal_7086 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7090 ;
    wire new_AGEMA_signal_7091 ;
    wire new_AGEMA_signal_7092 ;
    wire new_AGEMA_signal_7093 ;
    wire new_AGEMA_signal_7094 ;
    wire new_AGEMA_signal_7095 ;
    wire new_AGEMA_signal_7096 ;
    wire new_AGEMA_signal_7097 ;
    wire new_AGEMA_signal_7098 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7102 ;
    wire new_AGEMA_signal_7103 ;
    wire new_AGEMA_signal_7104 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7108 ;
    wire new_AGEMA_signal_7109 ;
    wire new_AGEMA_signal_7110 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7114 ;
    wire new_AGEMA_signal_7115 ;
    wire new_AGEMA_signal_7116 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7120 ;
    wire new_AGEMA_signal_7121 ;
    wire new_AGEMA_signal_7122 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7126 ;
    wire new_AGEMA_signal_7127 ;
    wire new_AGEMA_signal_7128 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7132 ;
    wire new_AGEMA_signal_7133 ;
    wire new_AGEMA_signal_7134 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7138 ;
    wire new_AGEMA_signal_7139 ;
    wire new_AGEMA_signal_7140 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7144 ;
    wire new_AGEMA_signal_7145 ;
    wire new_AGEMA_signal_7146 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7150 ;
    wire new_AGEMA_signal_7151 ;
    wire new_AGEMA_signal_7152 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7156 ;
    wire new_AGEMA_signal_7157 ;
    wire new_AGEMA_signal_7158 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7162 ;
    wire new_AGEMA_signal_7163 ;
    wire new_AGEMA_signal_7164 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7168 ;
    wire new_AGEMA_signal_7169 ;
    wire new_AGEMA_signal_7170 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7174 ;
    wire new_AGEMA_signal_7175 ;
    wire new_AGEMA_signal_7176 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7180 ;
    wire new_AGEMA_signal_7181 ;
    wire new_AGEMA_signal_7182 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7186 ;
    wire new_AGEMA_signal_7187 ;
    wire new_AGEMA_signal_7188 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7192 ;
    wire new_AGEMA_signal_7193 ;
    wire new_AGEMA_signal_7194 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7198 ;
    wire new_AGEMA_signal_7199 ;
    wire new_AGEMA_signal_7200 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7204 ;
    wire new_AGEMA_signal_7205 ;
    wire new_AGEMA_signal_7206 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7489 ;
    wire new_AGEMA_signal_7490 ;
    wire new_AGEMA_signal_7491 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7495 ;
    wire new_AGEMA_signal_7496 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7502 ;
    wire new_AGEMA_signal_7503 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7507 ;
    wire new_AGEMA_signal_7508 ;
    wire new_AGEMA_signal_7509 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7513 ;
    wire new_AGEMA_signal_7514 ;
    wire new_AGEMA_signal_7515 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7519 ;
    wire new_AGEMA_signal_7520 ;
    wire new_AGEMA_signal_7521 ;
    wire new_AGEMA_signal_7522 ;
    wire new_AGEMA_signal_7523 ;
    wire new_AGEMA_signal_7524 ;
    wire new_AGEMA_signal_7525 ;
    wire new_AGEMA_signal_7526 ;
    wire new_AGEMA_signal_7527 ;
    wire new_AGEMA_signal_7528 ;
    wire new_AGEMA_signal_7529 ;
    wire new_AGEMA_signal_7530 ;
    wire new_AGEMA_signal_7531 ;
    wire new_AGEMA_signal_7532 ;
    wire new_AGEMA_signal_7533 ;
    wire new_AGEMA_signal_7534 ;
    wire new_AGEMA_signal_7535 ;
    wire new_AGEMA_signal_7536 ;
    wire new_AGEMA_signal_7537 ;
    wire new_AGEMA_signal_7538 ;
    wire new_AGEMA_signal_7539 ;
    wire new_AGEMA_signal_7540 ;
    wire new_AGEMA_signal_7541 ;
    wire new_AGEMA_signal_7542 ;
    wire new_AGEMA_signal_7543 ;
    wire new_AGEMA_signal_7544 ;
    wire new_AGEMA_signal_7545 ;
    wire new_AGEMA_signal_7546 ;
    wire new_AGEMA_signal_7547 ;
    wire new_AGEMA_signal_7548 ;
    wire new_AGEMA_signal_7549 ;
    wire new_AGEMA_signal_7550 ;
    wire new_AGEMA_signal_7551 ;
    wire new_AGEMA_signal_7552 ;
    wire new_AGEMA_signal_7553 ;
    wire new_AGEMA_signal_7554 ;
    wire new_AGEMA_signal_7555 ;
    wire new_AGEMA_signal_7556 ;
    wire new_AGEMA_signal_7557 ;
    wire new_AGEMA_signal_7558 ;
    wire new_AGEMA_signal_7559 ;
    wire new_AGEMA_signal_7560 ;
    wire new_AGEMA_signal_7561 ;
    wire new_AGEMA_signal_7562 ;
    wire new_AGEMA_signal_7563 ;
    wire new_AGEMA_signal_7564 ;
    wire new_AGEMA_signal_7565 ;
    wire new_AGEMA_signal_7566 ;
    wire new_AGEMA_signal_7567 ;
    wire new_AGEMA_signal_7568 ;
    wire new_AGEMA_signal_7569 ;
    wire new_AGEMA_signal_7570 ;
    wire new_AGEMA_signal_7571 ;
    wire new_AGEMA_signal_7572 ;
    wire new_AGEMA_signal_7573 ;
    wire new_AGEMA_signal_7574 ;
    wire new_AGEMA_signal_7575 ;
    wire new_AGEMA_signal_7576 ;
    wire new_AGEMA_signal_7577 ;
    wire new_AGEMA_signal_7578 ;
    wire new_AGEMA_signal_7579 ;
    wire new_AGEMA_signal_7580 ;
    wire new_AGEMA_signal_7581 ;
    wire new_AGEMA_signal_7582 ;
    wire new_AGEMA_signal_7583 ;
    wire new_AGEMA_signal_7584 ;
    wire new_AGEMA_signal_7585 ;
    wire new_AGEMA_signal_7586 ;
    wire new_AGEMA_signal_7587 ;
    wire new_AGEMA_signal_7588 ;
    wire new_AGEMA_signal_7589 ;
    wire new_AGEMA_signal_7590 ;
    wire new_AGEMA_signal_7591 ;
    wire new_AGEMA_signal_7592 ;
    wire new_AGEMA_signal_7593 ;
    wire new_AGEMA_signal_7594 ;
    wire new_AGEMA_signal_7595 ;
    wire new_AGEMA_signal_7596 ;
    wire new_AGEMA_signal_7597 ;
    wire new_AGEMA_signal_7598 ;
    wire new_AGEMA_signal_7599 ;
    wire new_AGEMA_signal_7600 ;
    wire new_AGEMA_signal_7601 ;
    wire new_AGEMA_signal_7602 ;
    wire new_AGEMA_signal_7603 ;
    wire new_AGEMA_signal_7604 ;
    wire new_AGEMA_signal_7605 ;
    wire new_AGEMA_signal_7606 ;
    wire new_AGEMA_signal_7607 ;
    wire new_AGEMA_signal_7608 ;
    wire new_AGEMA_signal_7609 ;
    wire new_AGEMA_signal_7610 ;
    wire new_AGEMA_signal_7611 ;
    wire new_AGEMA_signal_7612 ;
    wire new_AGEMA_signal_7613 ;
    wire new_AGEMA_signal_7614 ;
    wire new_AGEMA_signal_7615 ;
    wire new_AGEMA_signal_7616 ;
    wire new_AGEMA_signal_7617 ;
    wire new_AGEMA_signal_7618 ;
    wire new_AGEMA_signal_7619 ;
    wire new_AGEMA_signal_7620 ;
    wire new_AGEMA_signal_7621 ;
    wire new_AGEMA_signal_7622 ;
    wire new_AGEMA_signal_7623 ;
    wire new_AGEMA_signal_7624 ;
    wire new_AGEMA_signal_7625 ;
    wire new_AGEMA_signal_7626 ;
    wire new_AGEMA_signal_7627 ;
    wire new_AGEMA_signal_7628 ;
    wire new_AGEMA_signal_7629 ;
    wire new_AGEMA_signal_7630 ;
    wire new_AGEMA_signal_7631 ;
    wire new_AGEMA_signal_7632 ;
    wire new_AGEMA_signal_7633 ;
    wire new_AGEMA_signal_7634 ;
    wire new_AGEMA_signal_7635 ;
    wire new_AGEMA_signal_7636 ;
    wire new_AGEMA_signal_7637 ;
    wire new_AGEMA_signal_7638 ;
    wire new_AGEMA_signal_7639 ;
    wire new_AGEMA_signal_7640 ;
    wire new_AGEMA_signal_7641 ;
    wire new_AGEMA_signal_7642 ;
    wire new_AGEMA_signal_7643 ;
    wire new_AGEMA_signal_7644 ;
    wire new_AGEMA_signal_7645 ;
    wire new_AGEMA_signal_7646 ;
    wire new_AGEMA_signal_7647 ;
    wire new_AGEMA_signal_7648 ;
    wire new_AGEMA_signal_7649 ;
    wire new_AGEMA_signal_7650 ;
    wire new_AGEMA_signal_7651 ;
    wire new_AGEMA_signal_7652 ;
    wire new_AGEMA_signal_7653 ;
    wire new_AGEMA_signal_7654 ;
    wire new_AGEMA_signal_7655 ;
    wire new_AGEMA_signal_7656 ;
    wire new_AGEMA_signal_7657 ;
    wire new_AGEMA_signal_7658 ;
    wire new_AGEMA_signal_7659 ;
    wire new_AGEMA_signal_7660 ;
    wire new_AGEMA_signal_7661 ;
    wire new_AGEMA_signal_7662 ;
    wire new_AGEMA_signal_7664 ;
    wire new_AGEMA_signal_7666 ;
    wire new_AGEMA_signal_7668 ;
    wire new_AGEMA_signal_7670 ;
    wire new_AGEMA_signal_7672 ;
    wire new_AGEMA_signal_7674 ;
    wire new_AGEMA_signal_7676 ;
    wire new_AGEMA_signal_7678 ;
    wire new_AGEMA_signal_7680 ;
    wire new_AGEMA_signal_7682 ;
    wire new_AGEMA_signal_7684 ;
    wire new_AGEMA_signal_7686 ;
    wire new_AGEMA_signal_7688 ;
    wire new_AGEMA_signal_7690 ;
    wire new_AGEMA_signal_7692 ;
    wire new_AGEMA_signal_7694 ;
    wire new_AGEMA_signal_7696 ;
    wire new_AGEMA_signal_7698 ;
    wire new_AGEMA_signal_7700 ;
    wire new_AGEMA_signal_7702 ;
    wire new_AGEMA_signal_7704 ;
    wire new_AGEMA_signal_7706 ;
    wire new_AGEMA_signal_7708 ;
    wire new_AGEMA_signal_7710 ;
    wire new_AGEMA_signal_7712 ;
    wire new_AGEMA_signal_7713 ;
    wire new_AGEMA_signal_7714 ;
    wire new_AGEMA_signal_7715 ;
    wire new_AGEMA_signal_7716 ;
    wire new_AGEMA_signal_7717 ;
    wire new_AGEMA_signal_7718 ;
    wire new_AGEMA_signal_7719 ;
    wire new_AGEMA_signal_7720 ;
    wire new_AGEMA_signal_7721 ;
    wire new_AGEMA_signal_7722 ;
    wire new_AGEMA_signal_7723 ;
    wire new_AGEMA_signal_7724 ;
    wire new_AGEMA_signal_7725 ;
    wire new_AGEMA_signal_7726 ;
    wire new_AGEMA_signal_7727 ;
    wire new_AGEMA_signal_7728 ;
    wire new_AGEMA_signal_7729 ;
    wire new_AGEMA_signal_7730 ;
    wire new_AGEMA_signal_7731 ;
    wire new_AGEMA_signal_7732 ;
    wire new_AGEMA_signal_7733 ;
    wire new_AGEMA_signal_7734 ;
    wire new_AGEMA_signal_7735 ;
    wire new_AGEMA_signal_7736 ;
    wire new_AGEMA_signal_7737 ;
    wire new_AGEMA_signal_7738 ;
    wire new_AGEMA_signal_7739 ;
    wire new_AGEMA_signal_7740 ;
    wire new_AGEMA_signal_7741 ;
    wire new_AGEMA_signal_7742 ;
    wire new_AGEMA_signal_7743 ;
    wire new_AGEMA_signal_7744 ;
    wire new_AGEMA_signal_7745 ;
    wire new_AGEMA_signal_7746 ;
    wire new_AGEMA_signal_7747 ;
    wire new_AGEMA_signal_7748 ;
    wire new_AGEMA_signal_7749 ;
    wire new_AGEMA_signal_7750 ;
    wire new_AGEMA_signal_7751 ;
    wire new_AGEMA_signal_7752 ;
    wire new_AGEMA_signal_7753 ;
    wire new_AGEMA_signal_7754 ;
    wire new_AGEMA_signal_7755 ;
    wire new_AGEMA_signal_7756 ;
    wire new_AGEMA_signal_7757 ;
    wire new_AGEMA_signal_7758 ;
    wire new_AGEMA_signal_7759 ;
    wire new_AGEMA_signal_7760 ;
    wire new_AGEMA_signal_7761 ;
    wire new_AGEMA_signal_7762 ;
    wire new_AGEMA_signal_7763 ;
    wire new_AGEMA_signal_7764 ;
    wire new_AGEMA_signal_7765 ;
    wire new_AGEMA_signal_7766 ;
    wire new_AGEMA_signal_7767 ;
    wire new_AGEMA_signal_7768 ;
    wire new_AGEMA_signal_7769 ;
    wire new_AGEMA_signal_7770 ;
    wire new_AGEMA_signal_7771 ;
    wire new_AGEMA_signal_7772 ;
    wire new_AGEMA_signal_7773 ;
    wire new_AGEMA_signal_7774 ;
    wire new_AGEMA_signal_7775 ;
    wire new_AGEMA_signal_7776 ;
    wire new_AGEMA_signal_7777 ;
    wire new_AGEMA_signal_7778 ;
    wire new_AGEMA_signal_7779 ;
    wire new_AGEMA_signal_7780 ;
    wire new_AGEMA_signal_7781 ;
    wire new_AGEMA_signal_7782 ;
    wire new_AGEMA_signal_7783 ;
    wire new_AGEMA_signal_7784 ;
    wire new_AGEMA_signal_7785 ;
    wire new_AGEMA_signal_7786 ;
    wire new_AGEMA_signal_7787 ;
    wire new_AGEMA_signal_7788 ;
    wire new_AGEMA_signal_7789 ;
    wire new_AGEMA_signal_7790 ;
    wire new_AGEMA_signal_7791 ;
    wire new_AGEMA_signal_7792 ;
    wire new_AGEMA_signal_7793 ;
    wire new_AGEMA_signal_7794 ;
    wire new_AGEMA_signal_7795 ;
    wire new_AGEMA_signal_7796 ;
    wire new_AGEMA_signal_7797 ;
    wire new_AGEMA_signal_7798 ;
    wire new_AGEMA_signal_7799 ;
    wire new_AGEMA_signal_7800 ;
    wire new_AGEMA_signal_7801 ;
    wire new_AGEMA_signal_7802 ;
    wire new_AGEMA_signal_7803 ;
    wire new_AGEMA_signal_7804 ;
    wire new_AGEMA_signal_7805 ;
    wire new_AGEMA_signal_7806 ;
    wire new_AGEMA_signal_7807 ;
    wire new_AGEMA_signal_7808 ;
    wire new_AGEMA_signal_7809 ;
    wire new_AGEMA_signal_7810 ;
    wire new_AGEMA_signal_7811 ;
    wire new_AGEMA_signal_7812 ;
    wire new_AGEMA_signal_7813 ;
    wire new_AGEMA_signal_7814 ;
    wire new_AGEMA_signal_7815 ;
    wire new_AGEMA_signal_7816 ;
    wire new_AGEMA_signal_7817 ;
    wire new_AGEMA_signal_7818 ;
    wire new_AGEMA_signal_7819 ;
    wire new_AGEMA_signal_7820 ;
    wire new_AGEMA_signal_7821 ;
    wire new_AGEMA_signal_7822 ;
    wire new_AGEMA_signal_7823 ;
    wire new_AGEMA_signal_7824 ;
    wire new_AGEMA_signal_7825 ;
    wire new_AGEMA_signal_7826 ;
    wire new_AGEMA_signal_7827 ;
    wire new_AGEMA_signal_7828 ;
    wire new_AGEMA_signal_7829 ;
    wire new_AGEMA_signal_7830 ;
    wire new_AGEMA_signal_7831 ;
    wire new_AGEMA_signal_7832 ;
    wire new_AGEMA_signal_7833 ;
    wire new_AGEMA_signal_7834 ;
    wire new_AGEMA_signal_7835 ;
    wire new_AGEMA_signal_7836 ;
    wire new_AGEMA_signal_7837 ;
    wire new_AGEMA_signal_7838 ;
    wire new_AGEMA_signal_7839 ;
    wire new_AGEMA_signal_7840 ;
    wire new_AGEMA_signal_7841 ;
    wire new_AGEMA_signal_7842 ;
    wire new_AGEMA_signal_7843 ;
    wire new_AGEMA_signal_7844 ;
    wire new_AGEMA_signal_7845 ;
    wire new_AGEMA_signal_7846 ;
    wire new_AGEMA_signal_7847 ;
    wire new_AGEMA_signal_7848 ;
    wire new_AGEMA_signal_7849 ;
    wire new_AGEMA_signal_7850 ;
    wire new_AGEMA_signal_7851 ;
    wire new_AGEMA_signal_7852 ;
    wire new_AGEMA_signal_7853 ;
    wire new_AGEMA_signal_7854 ;
    wire new_AGEMA_signal_7855 ;
    wire new_AGEMA_signal_7856 ;
    wire new_AGEMA_signal_7857 ;
    wire new_AGEMA_signal_7858 ;
    wire new_AGEMA_signal_7859 ;
    wire new_AGEMA_signal_7860 ;
    wire new_AGEMA_signal_7861 ;
    wire new_AGEMA_signal_7862 ;
    wire new_AGEMA_signal_7863 ;
    wire new_AGEMA_signal_7864 ;
    wire new_AGEMA_signal_7865 ;
    wire new_AGEMA_signal_7866 ;
    wire new_AGEMA_signal_7867 ;
    wire new_AGEMA_signal_7868 ;
    wire new_AGEMA_signal_7869 ;
    wire new_AGEMA_signal_7870 ;
    wire new_AGEMA_signal_7871 ;
    wire new_AGEMA_signal_7872 ;
    wire new_AGEMA_signal_7874 ;
    wire new_AGEMA_signal_7876 ;
    wire new_AGEMA_signal_7878 ;
    wire new_AGEMA_signal_7880 ;
    wire new_AGEMA_signal_7882 ;
    wire new_AGEMA_signal_7884 ;
    wire new_AGEMA_signal_7886 ;
    wire new_AGEMA_signal_7888 ;
    wire new_AGEMA_signal_7890 ;
    wire new_AGEMA_signal_7892 ;
    wire new_AGEMA_signal_7894 ;
    wire new_AGEMA_signal_7896 ;
    wire new_AGEMA_signal_7898 ;
    wire new_AGEMA_signal_7900 ;
    wire new_AGEMA_signal_7902 ;
    wire new_AGEMA_signal_7904 ;
    wire new_AGEMA_signal_7906 ;
    wire new_AGEMA_signal_7908 ;
    wire new_AGEMA_signal_7910 ;
    wire new_AGEMA_signal_7912 ;
    wire new_AGEMA_signal_7914 ;
    wire new_AGEMA_signal_7916 ;
    wire new_AGEMA_signal_7918 ;
    wire new_AGEMA_signal_7920 ;
    wire new_AGEMA_signal_7922 ;
    wire new_AGEMA_signal_7924 ;
    wire new_AGEMA_signal_7926 ;
    wire new_AGEMA_signal_7928 ;
    wire new_AGEMA_signal_7930 ;
    wire new_AGEMA_signal_7932 ;
    wire new_AGEMA_signal_7934 ;
    wire new_AGEMA_signal_7936 ;
    wire new_AGEMA_signal_7937 ;
    wire new_AGEMA_signal_7938 ;
    wire new_AGEMA_signal_7939 ;
    wire new_AGEMA_signal_7940 ;
    wire new_AGEMA_signal_7941 ;
    wire new_AGEMA_signal_7942 ;
    wire new_AGEMA_signal_7943 ;
    wire new_AGEMA_signal_7944 ;
    wire new_AGEMA_signal_7945 ;
    wire new_AGEMA_signal_7946 ;
    wire new_AGEMA_signal_7947 ;
    wire new_AGEMA_signal_7948 ;
    wire new_AGEMA_signal_7949 ;
    wire new_AGEMA_signal_7950 ;
    wire new_AGEMA_signal_7951 ;
    wire new_AGEMA_signal_7952 ;
    wire new_AGEMA_signal_7953 ;
    wire new_AGEMA_signal_7954 ;
    wire new_AGEMA_signal_7955 ;
    wire new_AGEMA_signal_7956 ;
    wire new_AGEMA_signal_7957 ;
    wire new_AGEMA_signal_7958 ;
    wire new_AGEMA_signal_7959 ;
    wire new_AGEMA_signal_7960 ;
    wire new_AGEMA_signal_7961 ;
    wire new_AGEMA_signal_7962 ;
    wire new_AGEMA_signal_7963 ;
    wire new_AGEMA_signal_7964 ;
    wire new_AGEMA_signal_7965 ;
    wire new_AGEMA_signal_7966 ;
    wire new_AGEMA_signal_7967 ;
    wire new_AGEMA_signal_7968 ;
    wire new_AGEMA_signal_7969 ;
    wire new_AGEMA_signal_7970 ;
    wire new_AGEMA_signal_7971 ;
    wire new_AGEMA_signal_7972 ;
    wire new_AGEMA_signal_7973 ;
    wire new_AGEMA_signal_7974 ;
    wire new_AGEMA_signal_7975 ;
    wire new_AGEMA_signal_7976 ;
    wire new_AGEMA_signal_7977 ;
    wire new_AGEMA_signal_7978 ;
    wire new_AGEMA_signal_7979 ;
    wire new_AGEMA_signal_7980 ;
    wire new_AGEMA_signal_7981 ;
    wire new_AGEMA_signal_7982 ;
    wire new_AGEMA_signal_7983 ;
    wire new_AGEMA_signal_7984 ;
    wire new_AGEMA_signal_7985 ;
    wire new_AGEMA_signal_7986 ;
    wire new_AGEMA_signal_7987 ;
    wire new_AGEMA_signal_7988 ;
    wire new_AGEMA_signal_7989 ;
    wire new_AGEMA_signal_7990 ;
    wire new_AGEMA_signal_7991 ;
    wire new_AGEMA_signal_7992 ;
    wire new_AGEMA_signal_7993 ;
    wire new_AGEMA_signal_7994 ;
    wire new_AGEMA_signal_7995 ;
    wire new_AGEMA_signal_7996 ;
    wire new_AGEMA_signal_7997 ;
    wire new_AGEMA_signal_7998 ;
    wire new_AGEMA_signal_7999 ;
    wire new_AGEMA_signal_8000 ;
    wire new_AGEMA_signal_8001 ;
    wire new_AGEMA_signal_8002 ;
    wire new_AGEMA_signal_8003 ;
    wire new_AGEMA_signal_8004 ;
    wire new_AGEMA_signal_8005 ;
    wire new_AGEMA_signal_8006 ;
    wire new_AGEMA_signal_8007 ;
    wire new_AGEMA_signal_8008 ;
    wire new_AGEMA_signal_8009 ;
    wire new_AGEMA_signal_8010 ;
    wire new_AGEMA_signal_8011 ;
    wire new_AGEMA_signal_8012 ;
    wire new_AGEMA_signal_8013 ;
    wire new_AGEMA_signal_8014 ;
    wire new_AGEMA_signal_8015 ;
    wire new_AGEMA_signal_8016 ;
    wire new_AGEMA_signal_8017 ;
    wire new_AGEMA_signal_8018 ;
    wire new_AGEMA_signal_8019 ;
    wire new_AGEMA_signal_8020 ;
    wire new_AGEMA_signal_8021 ;
    wire new_AGEMA_signal_8022 ;
    wire new_AGEMA_signal_8023 ;
    wire new_AGEMA_signal_8024 ;
    wire new_AGEMA_signal_8025 ;
    wire new_AGEMA_signal_8026 ;
    wire new_AGEMA_signal_8027 ;
    wire new_AGEMA_signal_8028 ;
    wire new_AGEMA_signal_8029 ;
    wire new_AGEMA_signal_8030 ;
    wire new_AGEMA_signal_8031 ;
    wire new_AGEMA_signal_8032 ;
    wire new_AGEMA_signal_8033 ;
    wire new_AGEMA_signal_8034 ;
    wire new_AGEMA_signal_8035 ;
    wire new_AGEMA_signal_8036 ;
    wire new_AGEMA_signal_8037 ;
    wire new_AGEMA_signal_8038 ;
    wire new_AGEMA_signal_8039 ;
    wire new_AGEMA_signal_8040 ;
    wire new_AGEMA_signal_8041 ;
    wire new_AGEMA_signal_8042 ;
    wire new_AGEMA_signal_8043 ;
    wire new_AGEMA_signal_8044 ;
    wire new_AGEMA_signal_8045 ;
    wire new_AGEMA_signal_8046 ;
    wire new_AGEMA_signal_8047 ;
    wire new_AGEMA_signal_8048 ;
    wire new_AGEMA_signal_8049 ;
    wire new_AGEMA_signal_8050 ;
    wire new_AGEMA_signal_8051 ;
    wire new_AGEMA_signal_8052 ;
    wire new_AGEMA_signal_8053 ;
    wire new_AGEMA_signal_8054 ;
    wire new_AGEMA_signal_8055 ;
    wire new_AGEMA_signal_8056 ;
    wire new_AGEMA_signal_8057 ;
    wire new_AGEMA_signal_8058 ;
    wire new_AGEMA_signal_8059 ;
    wire new_AGEMA_signal_8060 ;
    wire new_AGEMA_signal_8061 ;
    wire new_AGEMA_signal_8062 ;
    wire new_AGEMA_signal_8063 ;
    wire new_AGEMA_signal_8064 ;
    wire new_AGEMA_signal_8065 ;
    wire new_AGEMA_signal_8066 ;
    wire new_AGEMA_signal_8067 ;
    wire new_AGEMA_signal_8068 ;
    wire new_AGEMA_signal_8069 ;
    wire new_AGEMA_signal_8070 ;
    wire new_AGEMA_signal_8071 ;
    wire new_AGEMA_signal_8072 ;
    wire new_AGEMA_signal_8073 ;
    wire new_AGEMA_signal_8074 ;
    wire new_AGEMA_signal_8075 ;
    wire new_AGEMA_signal_8076 ;
    wire new_AGEMA_signal_8077 ;
    wire new_AGEMA_signal_8078 ;
    wire new_AGEMA_signal_8079 ;
    wire new_AGEMA_signal_8080 ;
    wire new_AGEMA_signal_8081 ;
    wire new_AGEMA_signal_8082 ;
    wire new_AGEMA_signal_8083 ;
    wire new_AGEMA_signal_8084 ;
    wire new_AGEMA_signal_8085 ;
    wire new_AGEMA_signal_8086 ;
    wire new_AGEMA_signal_8087 ;
    wire new_AGEMA_signal_8088 ;
    wire new_AGEMA_signal_8089 ;
    wire new_AGEMA_signal_8090 ;
    wire new_AGEMA_signal_8091 ;
    wire new_AGEMA_signal_8092 ;
    wire new_AGEMA_signal_8093 ;
    wire new_AGEMA_signal_8094 ;
    wire new_AGEMA_signal_8095 ;
    wire new_AGEMA_signal_8096 ;
    wire new_AGEMA_signal_8098 ;
    wire new_AGEMA_signal_8100 ;
    wire new_AGEMA_signal_8102 ;
    wire new_AGEMA_signal_8104 ;
    wire new_AGEMA_signal_8106 ;
    wire new_AGEMA_signal_8108 ;
    wire new_AGEMA_signal_8110 ;
    wire new_AGEMA_signal_8112 ;
    wire new_AGEMA_signal_8114 ;
    wire new_AGEMA_signal_8116 ;
    wire new_AGEMA_signal_8118 ;
    wire new_AGEMA_signal_8120 ;
    wire new_AGEMA_signal_8122 ;
    wire new_AGEMA_signal_8124 ;
    wire new_AGEMA_signal_8126 ;
    wire new_AGEMA_signal_8128 ;
    wire new_AGEMA_signal_8130 ;
    wire new_AGEMA_signal_8132 ;
    wire new_AGEMA_signal_8134 ;
    wire new_AGEMA_signal_8136 ;
    wire new_AGEMA_signal_8138 ;
    wire new_AGEMA_signal_8140 ;
    wire new_AGEMA_signal_8142 ;
    wire new_AGEMA_signal_8144 ;
    wire new_AGEMA_signal_8146 ;
    wire new_AGEMA_signal_8148 ;
    wire new_AGEMA_signal_8150 ;
    wire new_AGEMA_signal_8152 ;
    wire new_AGEMA_signal_8154 ;
    wire new_AGEMA_signal_8156 ;
    wire new_AGEMA_signal_8158 ;
    wire new_AGEMA_signal_8160 ;
    wire new_AGEMA_signal_8161 ;
    wire new_AGEMA_signal_8162 ;
    wire new_AGEMA_signal_8163 ;
    wire new_AGEMA_signal_8164 ;
    wire new_AGEMA_signal_8165 ;
    wire new_AGEMA_signal_8166 ;
    wire new_AGEMA_signal_8167 ;
    wire new_AGEMA_signal_8168 ;
    wire new_AGEMA_signal_8169 ;
    wire new_AGEMA_signal_8170 ;
    wire new_AGEMA_signal_8171 ;
    wire new_AGEMA_signal_8172 ;
    wire new_AGEMA_signal_8173 ;
    wire new_AGEMA_signal_8174 ;
    wire new_AGEMA_signal_8175 ;
    wire new_AGEMA_signal_8176 ;
    wire new_AGEMA_signal_8177 ;
    wire new_AGEMA_signal_8178 ;
    wire new_AGEMA_signal_8179 ;
    wire new_AGEMA_signal_8180 ;
    wire new_AGEMA_signal_8181 ;
    wire new_AGEMA_signal_8182 ;
    wire new_AGEMA_signal_8183 ;
    wire new_AGEMA_signal_8184 ;
    wire new_AGEMA_signal_8185 ;
    wire new_AGEMA_signal_8186 ;
    wire new_AGEMA_signal_8187 ;
    wire new_AGEMA_signal_8188 ;
    wire new_AGEMA_signal_8189 ;
    wire new_AGEMA_signal_8190 ;
    wire new_AGEMA_signal_8191 ;
    wire new_AGEMA_signal_8192 ;
    wire new_AGEMA_signal_8193 ;
    wire new_AGEMA_signal_8194 ;
    wire new_AGEMA_signal_8195 ;
    wire new_AGEMA_signal_8196 ;
    wire new_AGEMA_signal_8197 ;
    wire new_AGEMA_signal_8198 ;
    wire new_AGEMA_signal_8199 ;
    wire new_AGEMA_signal_8200 ;
    wire new_AGEMA_signal_8201 ;
    wire new_AGEMA_signal_8202 ;
    wire new_AGEMA_signal_8203 ;
    wire new_AGEMA_signal_8204 ;
    wire new_AGEMA_signal_8205 ;
    wire new_AGEMA_signal_8206 ;
    wire new_AGEMA_signal_8207 ;
    wire new_AGEMA_signal_8208 ;
    wire new_AGEMA_signal_8209 ;
    wire new_AGEMA_signal_8210 ;
    wire new_AGEMA_signal_8211 ;
    wire new_AGEMA_signal_8212 ;
    wire new_AGEMA_signal_8213 ;
    wire new_AGEMA_signal_8214 ;
    wire new_AGEMA_signal_8215 ;
    wire new_AGEMA_signal_8216 ;
    wire new_AGEMA_signal_8217 ;
    wire new_AGEMA_signal_8218 ;
    wire new_AGEMA_signal_8219 ;
    wire new_AGEMA_signal_8220 ;
    wire new_AGEMA_signal_8221 ;
    wire new_AGEMA_signal_8222 ;
    wire new_AGEMA_signal_8223 ;
    wire new_AGEMA_signal_8224 ;
    wire new_AGEMA_signal_8225 ;
    wire new_AGEMA_signal_8226 ;
    wire new_AGEMA_signal_8227 ;
    wire new_AGEMA_signal_8228 ;
    wire new_AGEMA_signal_8229 ;
    wire new_AGEMA_signal_8230 ;
    wire new_AGEMA_signal_8231 ;
    wire new_AGEMA_signal_8232 ;
    wire new_AGEMA_signal_8233 ;
    wire new_AGEMA_signal_8234 ;
    wire new_AGEMA_signal_8235 ;
    wire new_AGEMA_signal_8236 ;
    wire new_AGEMA_signal_8237 ;
    wire new_AGEMA_signal_8238 ;
    wire new_AGEMA_signal_8239 ;
    wire new_AGEMA_signal_8240 ;
    wire new_AGEMA_signal_8241 ;
    wire new_AGEMA_signal_8242 ;
    wire new_AGEMA_signal_8243 ;
    wire new_AGEMA_signal_8244 ;
    wire new_AGEMA_signal_8245 ;
    wire new_AGEMA_signal_8246 ;
    wire new_AGEMA_signal_8247 ;
    wire new_AGEMA_signal_8248 ;
    wire new_AGEMA_signal_8249 ;
    wire new_AGEMA_signal_8250 ;
    wire new_AGEMA_signal_8251 ;
    wire new_AGEMA_signal_8252 ;
    wire new_AGEMA_signal_8253 ;
    wire new_AGEMA_signal_8254 ;
    wire new_AGEMA_signal_8255 ;
    wire new_AGEMA_signal_8256 ;
    wire new_AGEMA_signal_8257 ;
    wire new_AGEMA_signal_8258 ;
    wire new_AGEMA_signal_8259 ;
    wire new_AGEMA_signal_8260 ;
    wire new_AGEMA_signal_8261 ;
    wire new_AGEMA_signal_8262 ;
    wire new_AGEMA_signal_8263 ;
    wire new_AGEMA_signal_8264 ;
    wire new_AGEMA_signal_8265 ;
    wire new_AGEMA_signal_8266 ;
    wire new_AGEMA_signal_8267 ;
    wire new_AGEMA_signal_8268 ;
    wire new_AGEMA_signal_8269 ;
    wire new_AGEMA_signal_8270 ;
    wire new_AGEMA_signal_8271 ;
    wire new_AGEMA_signal_8272 ;
    wire new_AGEMA_signal_8273 ;
    wire new_AGEMA_signal_8274 ;
    wire new_AGEMA_signal_8275 ;
    wire new_AGEMA_signal_8276 ;
    wire new_AGEMA_signal_8277 ;
    wire new_AGEMA_signal_8278 ;
    wire new_AGEMA_signal_8279 ;
    wire new_AGEMA_signal_8280 ;
    wire new_AGEMA_signal_8281 ;
    wire new_AGEMA_signal_8282 ;
    wire new_AGEMA_signal_8283 ;
    wire new_AGEMA_signal_8284 ;
    wire new_AGEMA_signal_8285 ;
    wire new_AGEMA_signal_8286 ;
    wire new_AGEMA_signal_8287 ;
    wire new_AGEMA_signal_8288 ;
    wire new_AGEMA_signal_8289 ;
    wire new_AGEMA_signal_8290 ;
    wire new_AGEMA_signal_8291 ;
    wire new_AGEMA_signal_8292 ;
    wire new_AGEMA_signal_8293 ;
    wire new_AGEMA_signal_8294 ;
    wire new_AGEMA_signal_8295 ;
    wire new_AGEMA_signal_8296 ;
    wire new_AGEMA_signal_8297 ;
    wire new_AGEMA_signal_8298 ;
    wire new_AGEMA_signal_8299 ;
    wire new_AGEMA_signal_8300 ;
    wire new_AGEMA_signal_8301 ;
    wire new_AGEMA_signal_8302 ;
    wire new_AGEMA_signal_8303 ;
    wire new_AGEMA_signal_8304 ;
    wire new_AGEMA_signal_8305 ;
    wire new_AGEMA_signal_8306 ;
    wire new_AGEMA_signal_8307 ;
    wire new_AGEMA_signal_8308 ;
    wire new_AGEMA_signal_8309 ;
    wire new_AGEMA_signal_8310 ;
    wire new_AGEMA_signal_8311 ;
    wire new_AGEMA_signal_8312 ;
    wire new_AGEMA_signal_8313 ;
    wire new_AGEMA_signal_8314 ;
    wire new_AGEMA_signal_8315 ;
    wire new_AGEMA_signal_8316 ;
    wire new_AGEMA_signal_8317 ;
    wire new_AGEMA_signal_8319 ;
    wire new_AGEMA_signal_8321 ;
    wire new_AGEMA_signal_8323 ;
    wire new_AGEMA_signal_8325 ;
    wire new_AGEMA_signal_8327 ;
    wire new_AGEMA_signal_8329 ;
    wire new_AGEMA_signal_8331 ;
    wire new_AGEMA_signal_8333 ;
    wire new_AGEMA_signal_8335 ;
    wire new_AGEMA_signal_8337 ;
    wire new_AGEMA_signal_8339 ;
    wire new_AGEMA_signal_8341 ;
    wire new_AGEMA_signal_8343 ;
    wire new_AGEMA_signal_8345 ;
    wire new_AGEMA_signal_8347 ;
    wire new_AGEMA_signal_8349 ;
    wire new_AGEMA_signal_8351 ;
    wire new_AGEMA_signal_8353 ;
    wire new_AGEMA_signal_8355 ;
    wire new_AGEMA_signal_8357 ;
    wire new_AGEMA_signal_8359 ;
    wire new_AGEMA_signal_8361 ;
    wire new_AGEMA_signal_8363 ;
    wire new_AGEMA_signal_8365 ;
    wire new_AGEMA_signal_8367 ;
    wire new_AGEMA_signal_8369 ;
    wire new_AGEMA_signal_8371 ;
    wire new_AGEMA_signal_8373 ;
    wire new_AGEMA_signal_8375 ;
    wire new_AGEMA_signal_8376 ;
    wire new_AGEMA_signal_8377 ;
    wire new_AGEMA_signal_8378 ;
    wire new_AGEMA_signal_8379 ;
    wire new_AGEMA_signal_8380 ;
    wire new_AGEMA_signal_8381 ;
    wire new_AGEMA_signal_8382 ;
    wire new_AGEMA_signal_8383 ;
    wire new_AGEMA_signal_8384 ;
    wire new_AGEMA_signal_8385 ;
    wire new_AGEMA_signal_8386 ;
    wire new_AGEMA_signal_8387 ;
    wire new_AGEMA_signal_8388 ;
    wire new_AGEMA_signal_8389 ;
    wire new_AGEMA_signal_8390 ;
    wire new_AGEMA_signal_8391 ;
    wire new_AGEMA_signal_8392 ;
    wire new_AGEMA_signal_8393 ;
    wire new_AGEMA_signal_8394 ;
    wire new_AGEMA_signal_8395 ;
    wire new_AGEMA_signal_8396 ;
    wire new_AGEMA_signal_8397 ;
    wire new_AGEMA_signal_8398 ;
    wire new_AGEMA_signal_8399 ;
    wire new_AGEMA_signal_8400 ;
    wire new_AGEMA_signal_8401 ;
    wire new_AGEMA_signal_8402 ;
    wire new_AGEMA_signal_8403 ;
    wire new_AGEMA_signal_8404 ;
    wire new_AGEMA_signal_8405 ;
    wire new_AGEMA_signal_8406 ;
    wire new_AGEMA_signal_8407 ;
    wire new_AGEMA_signal_8408 ;
    wire new_AGEMA_signal_8409 ;
    wire new_AGEMA_signal_8410 ;
    wire new_AGEMA_signal_8411 ;
    wire new_AGEMA_signal_8412 ;
    wire new_AGEMA_signal_8413 ;
    wire new_AGEMA_signal_8414 ;
    wire new_AGEMA_signal_8415 ;
    wire new_AGEMA_signal_8416 ;
    wire new_AGEMA_signal_8417 ;
    wire new_AGEMA_signal_8418 ;
    wire new_AGEMA_signal_8419 ;
    wire new_AGEMA_signal_8420 ;
    wire new_AGEMA_signal_8421 ;
    wire new_AGEMA_signal_8422 ;
    wire new_AGEMA_signal_8423 ;
    wire new_AGEMA_signal_8424 ;
    wire new_AGEMA_signal_8425 ;
    wire new_AGEMA_signal_8426 ;
    wire new_AGEMA_signal_8427 ;
    wire new_AGEMA_signal_8428 ;
    wire new_AGEMA_signal_8429 ;
    wire new_AGEMA_signal_8430 ;
    wire new_AGEMA_signal_8432 ;
    wire new_AGEMA_signal_8434 ;
    wire new_AGEMA_signal_8436 ;
    wire new_AGEMA_signal_8438 ;
    wire new_AGEMA_signal_8440 ;
    wire new_AGEMA_signal_8442 ;
    wire new_AGEMA_signal_8444 ;
    wire new_AGEMA_signal_8446 ;
    wire new_AGEMA_signal_8448 ;
    wire new_AGEMA_signal_8450 ;
    wire new_AGEMA_signal_8452 ;
    wire new_AGEMA_signal_8454 ;
    wire new_AGEMA_signal_8456 ;
    wire new_AGEMA_signal_8458 ;
    wire new_AGEMA_signal_8460 ;
    wire new_AGEMA_signal_8462 ;
    wire new_AGEMA_signal_8464 ;
    wire new_AGEMA_signal_8466 ;
    wire new_AGEMA_signal_8468 ;
    wire new_AGEMA_signal_8470 ;
    wire new_AGEMA_signal_8472 ;
    wire new_AGEMA_signal_8474 ;
    wire new_AGEMA_signal_8476 ;
    wire new_AGEMA_signal_8478 ;
    wire new_AGEMA_signal_8480 ;
    wire new_AGEMA_signal_8482 ;
    wire new_AGEMA_signal_8484 ;
    wire new_AGEMA_signal_8486 ;
    wire new_AGEMA_signal_8488 ;
    wire new_AGEMA_signal_8490 ;
    wire new_AGEMA_signal_8492 ;
    wire new_AGEMA_signal_8494 ;
    wire new_AGEMA_signal_8496 ;
    wire new_AGEMA_signal_8498 ;
    wire new_AGEMA_signal_8500 ;
    wire new_AGEMA_signal_8502 ;
    wire new_AGEMA_signal_8504 ;
    wire new_AGEMA_signal_8506 ;
    wire new_AGEMA_signal_8508 ;
    wire new_AGEMA_signal_8510 ;
    wire new_AGEMA_signal_8512 ;
    wire new_AGEMA_signal_8514 ;
    wire new_AGEMA_signal_8516 ;
    wire new_AGEMA_signal_8518 ;
    wire new_AGEMA_signal_8520 ;
    wire new_AGEMA_signal_8522 ;
    wire new_AGEMA_signal_8524 ;
    wire new_AGEMA_signal_8526 ;
    wire new_AGEMA_signal_8528 ;
    wire new_AGEMA_signal_8530 ;
    wire new_AGEMA_signal_8532 ;
    wire new_AGEMA_signal_8534 ;
    wire new_AGEMA_signal_8536 ;
    wire new_AGEMA_signal_8538 ;
    wire new_AGEMA_signal_8540 ;
    wire new_AGEMA_signal_8542 ;
    wire new_AGEMA_signal_8544 ;
    wire new_AGEMA_signal_8546 ;
    wire new_AGEMA_signal_8548 ;
    wire new_AGEMA_signal_8550 ;
    wire new_AGEMA_signal_8552 ;
    wire new_AGEMA_signal_8554 ;
    wire new_AGEMA_signal_8556 ;
    wire new_AGEMA_signal_8558 ;
    wire new_AGEMA_signal_8560 ;
    wire new_AGEMA_signal_8562 ;
    wire new_AGEMA_signal_8564 ;
    wire new_AGEMA_signal_8566 ;
    wire new_AGEMA_signal_8568 ;
    wire new_AGEMA_signal_8570 ;
    wire new_AGEMA_signal_8572 ;
    wire new_AGEMA_signal_8574 ;
    wire new_AGEMA_signal_8576 ;
    wire new_AGEMA_signal_8578 ;
    wire new_AGEMA_signal_8580 ;
    wire new_AGEMA_signal_8582 ;
    wire new_AGEMA_signal_8584 ;
    wire new_AGEMA_signal_8586 ;
    wire new_AGEMA_signal_8588 ;
    wire new_AGEMA_signal_8590 ;
    wire new_AGEMA_signal_8592 ;
    wire new_AGEMA_signal_8594 ;
    wire new_AGEMA_signal_8596 ;
    wire new_AGEMA_signal_8598 ;
    wire new_AGEMA_signal_8600 ;
    wire new_AGEMA_signal_8602 ;
    wire new_AGEMA_signal_8604 ;
    wire new_AGEMA_signal_8606 ;
    wire new_AGEMA_signal_8608 ;
    wire new_AGEMA_signal_8610 ;
    wire new_AGEMA_signal_8612 ;
    wire new_AGEMA_signal_8614 ;
    wire new_AGEMA_signal_8616 ;
    wire new_AGEMA_signal_8618 ;
    wire new_AGEMA_signal_8620 ;
    wire new_AGEMA_signal_8622 ;
    wire new_AGEMA_signal_8624 ;
    wire new_AGEMA_signal_8626 ;
    wire new_AGEMA_signal_8628 ;
    wire new_AGEMA_signal_8630 ;
    wire new_AGEMA_signal_8632 ;
    wire new_AGEMA_signal_8634 ;
    wire new_AGEMA_signal_8636 ;
    wire new_AGEMA_signal_8638 ;
    wire new_AGEMA_signal_8640 ;
    wire new_AGEMA_signal_8642 ;
    wire new_AGEMA_signal_8644 ;
    wire new_AGEMA_signal_8646 ;
    wire new_AGEMA_signal_8648 ;
    wire new_AGEMA_signal_8650 ;
    wire new_AGEMA_signal_8652 ;
    wire new_AGEMA_signal_8654 ;
    wire new_AGEMA_signal_8656 ;
    wire new_AGEMA_signal_8658 ;
    wire new_AGEMA_signal_8660 ;
    wire new_AGEMA_signal_8662 ;
    wire new_AGEMA_signal_8664 ;
    wire new_AGEMA_signal_8666 ;
    wire new_AGEMA_signal_8668 ;
    wire new_AGEMA_signal_8670 ;
    wire new_AGEMA_signal_8672 ;
    wire new_AGEMA_signal_8674 ;
    wire new_AGEMA_signal_8676 ;
    wire new_AGEMA_signal_8678 ;
    wire new_AGEMA_signal_8680 ;
    wire new_AGEMA_signal_8682 ;
    wire new_AGEMA_signal_8684 ;
    wire new_AGEMA_signal_8686 ;
    wire new_AGEMA_signal_8688 ;
    wire new_AGEMA_signal_8690 ;
    wire new_AGEMA_signal_8692 ;
    wire new_AGEMA_signal_8694 ;
    wire new_AGEMA_signal_8696 ;
    wire new_AGEMA_signal_8698 ;
    wire new_AGEMA_signal_8700 ;
    wire clk_gated ;

    /* cells in depth 0 */
    INV_X1 U830 ( .A (n314), .ZN (n319) ) ;
    INV_X1 U831 ( .A (n314), .ZN (n320) ) ;
    INV_X1 U832 ( .A (n314), .ZN (n317) ) ;
    INV_X1 U833 ( .A (n314), .ZN (n315) ) ;
    INV_X1 U834 ( .A (n314), .ZN (n316) ) ;
    INV_X1 U835 ( .A (n314), .ZN (n318) ) ;
    NOR2_X1 U836 ( .A1 (n325), .A2 (n330), .ZN (n314) ) ;
    INV_X1 U837 ( .A (RoundCounter[0]), .ZN (n325) ) ;
    INV_X1 U838 ( .A (n314), .ZN (n321) ) ;
    NOR2_X1 U839 ( .A1 (RoundCounter[2]), .A2 (RoundCounter[1]), .ZN (n323) ) ;
    INV_X1 U840 ( .A (n323), .ZN (n322) ) ;
    NOR2_X1 U841 ( .A1 (RoundCounter[0]), .A2 (n322), .ZN (Rcon[0]) ) ;
    NOR2_X1 U842 ( .A1 (RoundCounter[0]), .A2 (RoundCounter[3]), .ZN (n337) ) ;
    NOR2_X1 U843 ( .A1 (n337), .A2 (n322), .ZN (Rcon[1]) ) ;
    NAND2_X1 U844 ( .A1 (RoundCounter[3]), .A2 (n323), .ZN (n330) ) ;
    INV_X1 U845 ( .A (RoundCounter[2]), .ZN (n328) ) ;
    AND2_X1 U846 ( .A1 (n328), .A2 (RoundCounter[1]), .ZN (n333) ) ;
    NAND2_X1 U847 ( .A1 (n337), .A2 (n333), .ZN (n324) ) ;
    NAND2_X1 U848 ( .A1 (n321), .A2 (n324), .ZN (Rcon[2]) ) ;
    NOR2_X1 U849 ( .A1 (RoundCounter[3]), .A2 (n325), .ZN (n335) ) ;
    NAND2_X1 U850 ( .A1 (n333), .A2 (n335), .ZN (n327) ) ;
    NAND2_X1 U851 ( .A1 (RoundCounter[3]), .A2 (Rcon[0]), .ZN (n326) ) ;
    NAND2_X1 U852 ( .A1 (n327), .A2 (n326), .ZN (Rcon[3]) ) ;
    NOR2_X1 U853 ( .A1 (RoundCounter[1]), .A2 (n328), .ZN (n331) ) ;
    NAND2_X1 U854 ( .A1 (n337), .A2 (n331), .ZN (n329) ) ;
    NAND2_X1 U855 ( .A1 (n330), .A2 (n329), .ZN (Rcon[4]) ) ;
    NAND2_X1 U856 ( .A1 (n335), .A2 (n331), .ZN (n332) ) ;
    NAND2_X1 U857 ( .A1 (n321), .A2 (n332), .ZN (Rcon[5]) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U986 ( .a ({new_AGEMA_signal_4549, RoundInput[0]}), .b ({new_AGEMA_signal_4550, RoundKey[0]}), .c ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U987 ( .a ({new_AGEMA_signal_4552, RoundInput[100]}), .b ({new_AGEMA_signal_4553, RoundKey[100]}), .c ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U988 ( .a ({new_AGEMA_signal_4555, RoundInput[101]}), .b ({new_AGEMA_signal_4556, RoundKey[101]}), .c ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U989 ( .a ({new_AGEMA_signal_4558, RoundInput[102]}), .b ({new_AGEMA_signal_4559, RoundKey[102]}), .c ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U990 ( .a ({new_AGEMA_signal_4561, RoundInput[103]}), .b ({new_AGEMA_signal_4562, RoundKey[103]}), .c ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U991 ( .a ({new_AGEMA_signal_4564, RoundInput[104]}), .b ({new_AGEMA_signal_4565, RoundKey[104]}), .c ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U992 ( .a ({new_AGEMA_signal_4567, RoundInput[105]}), .b ({new_AGEMA_signal_4568, RoundKey[105]}), .c ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U993 ( .a ({new_AGEMA_signal_4570, RoundInput[106]}), .b ({new_AGEMA_signal_4571, RoundKey[106]}), .c ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U994 ( .a ({new_AGEMA_signal_4573, RoundInput[107]}), .b ({new_AGEMA_signal_4574, RoundKey[107]}), .c ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U995 ( .a ({new_AGEMA_signal_4576, RoundInput[108]}), .b ({new_AGEMA_signal_4577, RoundKey[108]}), .c ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U996 ( .a ({new_AGEMA_signal_4579, RoundInput[109]}), .b ({new_AGEMA_signal_4580, RoundKey[109]}), .c ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U997 ( .a ({new_AGEMA_signal_4582, RoundInput[10]}), .b ({new_AGEMA_signal_4583, RoundKey[10]}), .c ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U998 ( .a ({new_AGEMA_signal_4585, RoundInput[110]}), .b ({new_AGEMA_signal_4586, RoundKey[110]}), .c ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U999 ( .a ({new_AGEMA_signal_4588, RoundInput[111]}), .b ({new_AGEMA_signal_4589, RoundKey[111]}), .c ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1000 ( .a ({new_AGEMA_signal_4591, RoundInput[112]}), .b ({new_AGEMA_signal_4592, RoundKey[112]}), .c ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1001 ( .a ({new_AGEMA_signal_4594, RoundInput[113]}), .b ({new_AGEMA_signal_4595, RoundKey[113]}), .c ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1002 ( .a ({new_AGEMA_signal_4597, RoundInput[114]}), .b ({new_AGEMA_signal_4598, RoundKey[114]}), .c ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1003 ( .a ({new_AGEMA_signal_4600, RoundInput[115]}), .b ({new_AGEMA_signal_4601, RoundKey[115]}), .c ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1004 ( .a ({new_AGEMA_signal_4603, RoundInput[116]}), .b ({new_AGEMA_signal_4604, RoundKey[116]}), .c ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1005 ( .a ({new_AGEMA_signal_4606, RoundInput[117]}), .b ({new_AGEMA_signal_4607, RoundKey[117]}), .c ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1006 ( .a ({new_AGEMA_signal_4609, RoundInput[118]}), .b ({new_AGEMA_signal_4610, RoundKey[118]}), .c ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1007 ( .a ({new_AGEMA_signal_4612, RoundInput[119]}), .b ({new_AGEMA_signal_4613, RoundKey[119]}), .c ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1008 ( .a ({new_AGEMA_signal_4615, RoundInput[11]}), .b ({new_AGEMA_signal_4616, RoundKey[11]}), .c ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1009 ( .a ({new_AGEMA_signal_4618, RoundInput[120]}), .b ({new_AGEMA_signal_4619, RoundKey[120]}), .c ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1010 ( .a ({new_AGEMA_signal_4621, RoundInput[121]}), .b ({new_AGEMA_signal_4622, RoundKey[121]}), .c ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1011 ( .a ({new_AGEMA_signal_4624, RoundInput[122]}), .b ({new_AGEMA_signal_4625, RoundKey[122]}), .c ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1012 ( .a ({new_AGEMA_signal_4627, RoundInput[123]}), .b ({new_AGEMA_signal_4628, RoundKey[123]}), .c ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1013 ( .a ({new_AGEMA_signal_4630, RoundInput[124]}), .b ({new_AGEMA_signal_4631, RoundKey[124]}), .c ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1014 ( .a ({new_AGEMA_signal_4633, RoundInput[125]}), .b ({new_AGEMA_signal_4634, RoundKey[125]}), .c ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1015 ( .a ({new_AGEMA_signal_4636, RoundInput[126]}), .b ({new_AGEMA_signal_4637, RoundKey[126]}), .c ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1016 ( .a ({new_AGEMA_signal_4639, RoundInput[127]}), .b ({new_AGEMA_signal_4640, RoundKey[127]}), .c ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1017 ( .a ({new_AGEMA_signal_4642, RoundInput[12]}), .b ({new_AGEMA_signal_4643, RoundKey[12]}), .c ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1018 ( .a ({new_AGEMA_signal_4645, RoundInput[13]}), .b ({new_AGEMA_signal_4646, RoundKey[13]}), .c ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1019 ( .a ({new_AGEMA_signal_4648, RoundInput[14]}), .b ({new_AGEMA_signal_4649, RoundKey[14]}), .c ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1020 ( .a ({new_AGEMA_signal_4651, RoundInput[15]}), .b ({new_AGEMA_signal_4652, RoundKey[15]}), .c ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1021 ( .a ({new_AGEMA_signal_4654, RoundInput[16]}), .b ({new_AGEMA_signal_4655, RoundKey[16]}), .c ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1022 ( .a ({new_AGEMA_signal_4657, RoundInput[17]}), .b ({new_AGEMA_signal_4658, RoundKey[17]}), .c ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1023 ( .a ({new_AGEMA_signal_4660, RoundInput[18]}), .b ({new_AGEMA_signal_4661, RoundKey[18]}), .c ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1024 ( .a ({new_AGEMA_signal_4663, RoundInput[19]}), .b ({new_AGEMA_signal_4664, RoundKey[19]}), .c ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1025 ( .a ({new_AGEMA_signal_4666, RoundInput[1]}), .b ({new_AGEMA_signal_4667, RoundKey[1]}), .c ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1026 ( .a ({new_AGEMA_signal_4669, RoundInput[20]}), .b ({new_AGEMA_signal_4670, RoundKey[20]}), .c ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1027 ( .a ({new_AGEMA_signal_4672, RoundInput[21]}), .b ({new_AGEMA_signal_4673, RoundKey[21]}), .c ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1028 ( .a ({new_AGEMA_signal_4675, RoundInput[22]}), .b ({new_AGEMA_signal_4676, RoundKey[22]}), .c ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1029 ( .a ({new_AGEMA_signal_4678, RoundInput[23]}), .b ({new_AGEMA_signal_4679, RoundKey[23]}), .c ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1030 ( .a ({new_AGEMA_signal_4681, RoundInput[24]}), .b ({new_AGEMA_signal_4682, RoundKey[24]}), .c ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1031 ( .a ({new_AGEMA_signal_4684, RoundInput[25]}), .b ({new_AGEMA_signal_4685, RoundKey[25]}), .c ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1032 ( .a ({new_AGEMA_signal_4687, RoundInput[26]}), .b ({new_AGEMA_signal_4688, RoundKey[26]}), .c ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1033 ( .a ({new_AGEMA_signal_4690, RoundInput[27]}), .b ({new_AGEMA_signal_4691, RoundKey[27]}), .c ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1034 ( .a ({new_AGEMA_signal_4693, RoundInput[28]}), .b ({new_AGEMA_signal_4694, RoundKey[28]}), .c ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1035 ( .a ({new_AGEMA_signal_4696, RoundInput[29]}), .b ({new_AGEMA_signal_4697, RoundKey[29]}), .c ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1036 ( .a ({new_AGEMA_signal_4699, RoundInput[2]}), .b ({new_AGEMA_signal_4700, RoundKey[2]}), .c ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1037 ( .a ({new_AGEMA_signal_4702, RoundInput[30]}), .b ({new_AGEMA_signal_4703, RoundKey[30]}), .c ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1038 ( .a ({new_AGEMA_signal_4705, RoundInput[31]}), .b ({new_AGEMA_signal_4706, RoundKey[31]}), .c ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1039 ( .a ({new_AGEMA_signal_4708, RoundInput[32]}), .b ({new_AGEMA_signal_4709, RoundKey[32]}), .c ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1040 ( .a ({new_AGEMA_signal_4711, RoundInput[33]}), .b ({new_AGEMA_signal_4712, RoundKey[33]}), .c ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1041 ( .a ({new_AGEMA_signal_4714, RoundInput[34]}), .b ({new_AGEMA_signal_4715, RoundKey[34]}), .c ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1042 ( .a ({new_AGEMA_signal_4717, RoundInput[35]}), .b ({new_AGEMA_signal_4718, RoundKey[35]}), .c ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1043 ( .a ({new_AGEMA_signal_4720, RoundInput[36]}), .b ({new_AGEMA_signal_4721, RoundKey[36]}), .c ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1044 ( .a ({new_AGEMA_signal_4723, RoundInput[37]}), .b ({new_AGEMA_signal_4724, RoundKey[37]}), .c ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1045 ( .a ({new_AGEMA_signal_4726, RoundInput[38]}), .b ({new_AGEMA_signal_4727, RoundKey[38]}), .c ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1046 ( .a ({new_AGEMA_signal_4729, RoundInput[39]}), .b ({new_AGEMA_signal_4730, RoundKey[39]}), .c ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1047 ( .a ({new_AGEMA_signal_4732, RoundInput[3]}), .b ({new_AGEMA_signal_4733, RoundKey[3]}), .c ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1048 ( .a ({new_AGEMA_signal_4735, RoundInput[40]}), .b ({new_AGEMA_signal_4736, RoundKey[40]}), .c ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1049 ( .a ({new_AGEMA_signal_4738, RoundInput[41]}), .b ({new_AGEMA_signal_4739, RoundKey[41]}), .c ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1050 ( .a ({new_AGEMA_signal_4741, RoundInput[42]}), .b ({new_AGEMA_signal_4742, RoundKey[42]}), .c ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1051 ( .a ({new_AGEMA_signal_4744, RoundInput[43]}), .b ({new_AGEMA_signal_4745, RoundKey[43]}), .c ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1052 ( .a ({new_AGEMA_signal_4747, RoundInput[44]}), .b ({new_AGEMA_signal_4748, RoundKey[44]}), .c ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1053 ( .a ({new_AGEMA_signal_4750, RoundInput[45]}), .b ({new_AGEMA_signal_4751, RoundKey[45]}), .c ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1054 ( .a ({new_AGEMA_signal_4753, RoundInput[46]}), .b ({new_AGEMA_signal_4754, RoundKey[46]}), .c ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1055 ( .a ({new_AGEMA_signal_4756, RoundInput[47]}), .b ({new_AGEMA_signal_4757, RoundKey[47]}), .c ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1056 ( .a ({new_AGEMA_signal_4759, RoundInput[48]}), .b ({new_AGEMA_signal_4760, RoundKey[48]}), .c ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1057 ( .a ({new_AGEMA_signal_4762, RoundInput[49]}), .b ({new_AGEMA_signal_4763, RoundKey[49]}), .c ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1058 ( .a ({new_AGEMA_signal_4765, RoundInput[4]}), .b ({new_AGEMA_signal_4766, RoundKey[4]}), .c ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1059 ( .a ({new_AGEMA_signal_4768, RoundInput[50]}), .b ({new_AGEMA_signal_4769, RoundKey[50]}), .c ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1060 ( .a ({new_AGEMA_signal_4771, RoundInput[51]}), .b ({new_AGEMA_signal_4772, RoundKey[51]}), .c ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1061 ( .a ({new_AGEMA_signal_4774, RoundInput[52]}), .b ({new_AGEMA_signal_4775, RoundKey[52]}), .c ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1062 ( .a ({new_AGEMA_signal_4777, RoundInput[53]}), .b ({new_AGEMA_signal_4778, RoundKey[53]}), .c ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1063 ( .a ({new_AGEMA_signal_4780, RoundInput[54]}), .b ({new_AGEMA_signal_4781, RoundKey[54]}), .c ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1064 ( .a ({new_AGEMA_signal_4783, RoundInput[55]}), .b ({new_AGEMA_signal_4784, RoundKey[55]}), .c ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1065 ( .a ({new_AGEMA_signal_4786, RoundInput[56]}), .b ({new_AGEMA_signal_4787, RoundKey[56]}), .c ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1066 ( .a ({new_AGEMA_signal_4789, RoundInput[57]}), .b ({new_AGEMA_signal_4790, RoundKey[57]}), .c ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1067 ( .a ({new_AGEMA_signal_4792, RoundInput[58]}), .b ({new_AGEMA_signal_4793, RoundKey[58]}), .c ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1068 ( .a ({new_AGEMA_signal_4795, RoundInput[59]}), .b ({new_AGEMA_signal_4796, RoundKey[59]}), .c ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1069 ( .a ({new_AGEMA_signal_4798, RoundInput[5]}), .b ({new_AGEMA_signal_4799, RoundKey[5]}), .c ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1070 ( .a ({new_AGEMA_signal_4801, RoundInput[60]}), .b ({new_AGEMA_signal_4802, RoundKey[60]}), .c ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1071 ( .a ({new_AGEMA_signal_4804, RoundInput[61]}), .b ({new_AGEMA_signal_4805, RoundKey[61]}), .c ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1072 ( .a ({new_AGEMA_signal_4807, RoundInput[62]}), .b ({new_AGEMA_signal_4808, RoundKey[62]}), .c ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1073 ( .a ({new_AGEMA_signal_4810, RoundInput[63]}), .b ({new_AGEMA_signal_4811, RoundKey[63]}), .c ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1074 ( .a ({new_AGEMA_signal_4813, RoundInput[64]}), .b ({new_AGEMA_signal_4814, RoundKey[64]}), .c ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1075 ( .a ({new_AGEMA_signal_4816, RoundInput[65]}), .b ({new_AGEMA_signal_4817, RoundKey[65]}), .c ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1076 ( .a ({new_AGEMA_signal_4819, RoundInput[66]}), .b ({new_AGEMA_signal_4820, RoundKey[66]}), .c ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1077 ( .a ({new_AGEMA_signal_4822, RoundInput[67]}), .b ({new_AGEMA_signal_4823, RoundKey[67]}), .c ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1078 ( .a ({new_AGEMA_signal_4825, RoundInput[68]}), .b ({new_AGEMA_signal_4826, RoundKey[68]}), .c ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1079 ( .a ({new_AGEMA_signal_4828, RoundInput[69]}), .b ({new_AGEMA_signal_4829, RoundKey[69]}), .c ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1080 ( .a ({new_AGEMA_signal_4831, RoundInput[6]}), .b ({new_AGEMA_signal_4832, RoundKey[6]}), .c ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1081 ( .a ({new_AGEMA_signal_4834, RoundInput[70]}), .b ({new_AGEMA_signal_4835, RoundKey[70]}), .c ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1082 ( .a ({new_AGEMA_signal_4837, RoundInput[71]}), .b ({new_AGEMA_signal_4838, RoundKey[71]}), .c ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1083 ( .a ({new_AGEMA_signal_4840, RoundInput[72]}), .b ({new_AGEMA_signal_4841, RoundKey[72]}), .c ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1084 ( .a ({new_AGEMA_signal_4843, RoundInput[73]}), .b ({new_AGEMA_signal_4844, RoundKey[73]}), .c ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1085 ( .a ({new_AGEMA_signal_4846, RoundInput[74]}), .b ({new_AGEMA_signal_4847, RoundKey[74]}), .c ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1086 ( .a ({new_AGEMA_signal_4849, RoundInput[75]}), .b ({new_AGEMA_signal_4850, RoundKey[75]}), .c ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1087 ( .a ({new_AGEMA_signal_4852, RoundInput[76]}), .b ({new_AGEMA_signal_4853, RoundKey[76]}), .c ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1088 ( .a ({new_AGEMA_signal_4855, RoundInput[77]}), .b ({new_AGEMA_signal_4856, RoundKey[77]}), .c ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1089 ( .a ({new_AGEMA_signal_4858, RoundInput[78]}), .b ({new_AGEMA_signal_4859, RoundKey[78]}), .c ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1090 ( .a ({new_AGEMA_signal_4861, RoundInput[79]}), .b ({new_AGEMA_signal_4862, RoundKey[79]}), .c ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1091 ( .a ({new_AGEMA_signal_4864, RoundInput[7]}), .b ({new_AGEMA_signal_4865, RoundKey[7]}), .c ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1092 ( .a ({new_AGEMA_signal_4867, RoundInput[80]}), .b ({new_AGEMA_signal_4868, RoundKey[80]}), .c ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1093 ( .a ({new_AGEMA_signal_4870, RoundInput[81]}), .b ({new_AGEMA_signal_4871, RoundKey[81]}), .c ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1094 ( .a ({new_AGEMA_signal_4873, RoundInput[82]}), .b ({new_AGEMA_signal_4874, RoundKey[82]}), .c ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1095 ( .a ({new_AGEMA_signal_4876, RoundInput[83]}), .b ({new_AGEMA_signal_4877, RoundKey[83]}), .c ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1096 ( .a ({new_AGEMA_signal_4879, RoundInput[84]}), .b ({new_AGEMA_signal_4880, RoundKey[84]}), .c ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1097 ( .a ({new_AGEMA_signal_4882, RoundInput[85]}), .b ({new_AGEMA_signal_4883, RoundKey[85]}), .c ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1098 ( .a ({new_AGEMA_signal_4885, RoundInput[86]}), .b ({new_AGEMA_signal_4886, RoundKey[86]}), .c ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1099 ( .a ({new_AGEMA_signal_4888, RoundInput[87]}), .b ({new_AGEMA_signal_4889, RoundKey[87]}), .c ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1100 ( .a ({new_AGEMA_signal_4891, RoundInput[88]}), .b ({new_AGEMA_signal_4892, RoundKey[88]}), .c ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1101 ( .a ({new_AGEMA_signal_4894, RoundInput[89]}), .b ({new_AGEMA_signal_4895, RoundKey[89]}), .c ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1102 ( .a ({new_AGEMA_signal_4897, RoundInput[8]}), .b ({new_AGEMA_signal_4898, RoundKey[8]}), .c ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1103 ( .a ({new_AGEMA_signal_4900, RoundInput[90]}), .b ({new_AGEMA_signal_4901, RoundKey[90]}), .c ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1104 ( .a ({new_AGEMA_signal_4903, RoundInput[91]}), .b ({new_AGEMA_signal_4904, RoundKey[91]}), .c ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1105 ( .a ({new_AGEMA_signal_4906, RoundInput[92]}), .b ({new_AGEMA_signal_4907, RoundKey[92]}), .c ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1106 ( .a ({new_AGEMA_signal_4909, RoundInput[93]}), .b ({new_AGEMA_signal_4910, RoundKey[93]}), .c ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1107 ( .a ({new_AGEMA_signal_4912, RoundInput[94]}), .b ({new_AGEMA_signal_4913, RoundKey[94]}), .c ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1108 ( .a ({new_AGEMA_signal_4915, RoundInput[95]}), .b ({new_AGEMA_signal_4916, RoundKey[95]}), .c ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1109 ( .a ({new_AGEMA_signal_4918, RoundInput[96]}), .b ({new_AGEMA_signal_4919, RoundKey[96]}), .c ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1110 ( .a ({new_AGEMA_signal_4921, RoundInput[97]}), .b ({new_AGEMA_signal_4922, RoundKey[97]}), .c ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1111 ( .a ({new_AGEMA_signal_4924, RoundInput[98]}), .b ({new_AGEMA_signal_4925, RoundKey[98]}), .c ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1112 ( .a ({new_AGEMA_signal_4927, RoundInput[99]}), .b ({new_AGEMA_signal_4928, RoundKey[99]}), .c ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U1113 ( .a ({new_AGEMA_signal_4930, RoundInput[9]}), .b ({new_AGEMA_signal_4931, RoundKey[9]}), .c ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    NAND2_X1 U1114 ( .A1 (RoundCounter[3]), .A2 (n333), .ZN (n334) ) ;
    NOR2_X1 U1115 ( .A1 (RoundCounter[0]), .A2 (n334), .ZN (done) ) ;
    INV_X1 U1116 ( .A (n335), .ZN (n336) ) ;
    NAND2_X1 U1117 ( .A1 (RoundCounter[2]), .A2 (RoundCounter[1]), .ZN (n338) ) ;
    NOR2_X1 U1118 ( .A1 (n336), .A2 (n338), .ZN (n283) ) ;
    INV_X1 U1119 ( .A (n337), .ZN (n339) ) ;
    NOR2_X1 U1120 ( .A1 (n339), .A2 (n338), .ZN (n285) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T1_U1 ( .a ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({ciphertext_s1[4], ciphertext_s0[4]}), .c ({new_AGEMA_signal_4973, SubBytesIns_Inst_Sbox_0_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T2_U1 ( .a ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_4974, SubBytesIns_Inst_Sbox_0_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T3_U1 ( .a ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_4975, SubBytesIns_Inst_Sbox_0_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T4_U1 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_4976, SubBytesIns_Inst_Sbox_0_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T5_U1 ( .a ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_4977, SubBytesIns_Inst_Sbox_0_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T6_U1 ( .a ({new_AGEMA_signal_4973, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_4977, SubBytesIns_Inst_Sbox_0_T5}), .c ({new_AGEMA_signal_5165, SubBytesIns_Inst_Sbox_0_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T7_U1 ( .a ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({ciphertext_s1[5], ciphertext_s0[5]}), .c ({new_AGEMA_signal_4978, SubBytesIns_Inst_Sbox_0_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T8_U1 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_5165, SubBytesIns_Inst_Sbox_0_T6}), .c ({new_AGEMA_signal_5345, SubBytesIns_Inst_Sbox_0_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T9_U1 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_4978, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_5166, SubBytesIns_Inst_Sbox_0_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T10_U1 ( .a ({new_AGEMA_signal_5165, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_4978, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_5346, SubBytesIns_Inst_Sbox_0_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T11_U1 ( .a ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_4979, SubBytesIns_Inst_Sbox_0_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T12_U1 ( .a ({ciphertext_s1[5], ciphertext_s0[5]}), .b ({ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_4980, SubBytesIns_Inst_Sbox_0_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T13_U1 ( .a ({new_AGEMA_signal_4975, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_4976, SubBytesIns_Inst_Sbox_0_T4}), .c ({new_AGEMA_signal_5167, SubBytesIns_Inst_Sbox_0_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T14_U1 ( .a ({new_AGEMA_signal_5165, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_4979, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_5347, SubBytesIns_Inst_Sbox_0_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T15_U1 ( .a ({new_AGEMA_signal_4977, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_4979, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_5168, SubBytesIns_Inst_Sbox_0_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T16_U1 ( .a ({new_AGEMA_signal_4977, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_4980, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_5169, SubBytesIns_Inst_Sbox_0_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T17_U1 ( .a ({new_AGEMA_signal_5166, SubBytesIns_Inst_Sbox_0_T9}), .b ({new_AGEMA_signal_5169, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_5348, SubBytesIns_Inst_Sbox_0_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T18_U1 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_4981, SubBytesIns_Inst_Sbox_0_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T19_U1 ( .a ({new_AGEMA_signal_4978, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_4981, SubBytesIns_Inst_Sbox_0_T18}), .c ({new_AGEMA_signal_5170, SubBytesIns_Inst_Sbox_0_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T20_U1 ( .a ({new_AGEMA_signal_4973, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5170, SubBytesIns_Inst_Sbox_0_T19}), .c ({new_AGEMA_signal_5349, SubBytesIns_Inst_Sbox_0_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T21_U1 ( .a ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_4982, SubBytesIns_Inst_Sbox_0_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T22_U1 ( .a ({new_AGEMA_signal_4978, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_4982, SubBytesIns_Inst_Sbox_0_T21}), .c ({new_AGEMA_signal_5171, SubBytesIns_Inst_Sbox_0_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T23_U1 ( .a ({new_AGEMA_signal_4974, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_5171, SubBytesIns_Inst_Sbox_0_T22}), .c ({new_AGEMA_signal_5350, SubBytesIns_Inst_Sbox_0_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T24_U1 ( .a ({new_AGEMA_signal_4974, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_5346, SubBytesIns_Inst_Sbox_0_T10}), .c ({new_AGEMA_signal_5589, SubBytesIns_Inst_Sbox_0_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T25_U1 ( .a ({new_AGEMA_signal_5349, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_5348, SubBytesIns_Inst_Sbox_0_T17}), .c ({new_AGEMA_signal_5590, SubBytesIns_Inst_Sbox_0_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T26_U1 ( .a ({new_AGEMA_signal_4975, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5169, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_5351, SubBytesIns_Inst_Sbox_0_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T27_U1 ( .a ({new_AGEMA_signal_4973, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_4980, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_5172, SubBytesIns_Inst_Sbox_0_T27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T1_U1 ( .a ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s1[12], ciphertext_s0[12]}), .c ({new_AGEMA_signal_4983, SubBytesIns_Inst_Sbox_1_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T2_U1 ( .a ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_4984, SubBytesIns_Inst_Sbox_1_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T3_U1 ( .a ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({new_AGEMA_signal_4985, SubBytesIns_Inst_Sbox_1_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T4_U1 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_4986, SubBytesIns_Inst_Sbox_1_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T5_U1 ( .a ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({new_AGEMA_signal_4987, SubBytesIns_Inst_Sbox_1_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T6_U1 ( .a ({new_AGEMA_signal_4983, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_4987, SubBytesIns_Inst_Sbox_1_T5}), .c ({new_AGEMA_signal_5173, SubBytesIns_Inst_Sbox_1_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T7_U1 ( .a ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({ciphertext_s1[13], ciphertext_s0[13]}), .c ({new_AGEMA_signal_4988, SubBytesIns_Inst_Sbox_1_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T8_U1 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_5173, SubBytesIns_Inst_Sbox_1_T6}), .c ({new_AGEMA_signal_5358, SubBytesIns_Inst_Sbox_1_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T9_U1 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_4988, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_5174, SubBytesIns_Inst_Sbox_1_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T10_U1 ( .a ({new_AGEMA_signal_5173, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_4988, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_5359, SubBytesIns_Inst_Sbox_1_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T11_U1 ( .a ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_4989, SubBytesIns_Inst_Sbox_1_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T12_U1 ( .a ({ciphertext_s1[13], ciphertext_s0[13]}), .b ({ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_4990, SubBytesIns_Inst_Sbox_1_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T13_U1 ( .a ({new_AGEMA_signal_4985, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_4986, SubBytesIns_Inst_Sbox_1_T4}), .c ({new_AGEMA_signal_5175, SubBytesIns_Inst_Sbox_1_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T14_U1 ( .a ({new_AGEMA_signal_5173, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_4989, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_5360, SubBytesIns_Inst_Sbox_1_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T15_U1 ( .a ({new_AGEMA_signal_4987, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_4989, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_5176, SubBytesIns_Inst_Sbox_1_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T16_U1 ( .a ({new_AGEMA_signal_4987, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_4990, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_5177, SubBytesIns_Inst_Sbox_1_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T17_U1 ( .a ({new_AGEMA_signal_5174, SubBytesIns_Inst_Sbox_1_T9}), .b ({new_AGEMA_signal_5177, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_5361, SubBytesIns_Inst_Sbox_1_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T18_U1 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s1[8], ciphertext_s0[8]}), .c ({new_AGEMA_signal_4991, SubBytesIns_Inst_Sbox_1_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T19_U1 ( .a ({new_AGEMA_signal_4988, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_4991, SubBytesIns_Inst_Sbox_1_T18}), .c ({new_AGEMA_signal_5178, SubBytesIns_Inst_Sbox_1_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T20_U1 ( .a ({new_AGEMA_signal_4983, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5178, SubBytesIns_Inst_Sbox_1_T19}), .c ({new_AGEMA_signal_5362, SubBytesIns_Inst_Sbox_1_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T21_U1 ( .a ({ciphertext_s1[9], ciphertext_s0[9]}), .b ({ciphertext_s1[8], ciphertext_s0[8]}), .c ({new_AGEMA_signal_4992, SubBytesIns_Inst_Sbox_1_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T22_U1 ( .a ({new_AGEMA_signal_4988, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_4992, SubBytesIns_Inst_Sbox_1_T21}), .c ({new_AGEMA_signal_5179, SubBytesIns_Inst_Sbox_1_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T23_U1 ( .a ({new_AGEMA_signal_4984, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_5179, SubBytesIns_Inst_Sbox_1_T22}), .c ({new_AGEMA_signal_5363, SubBytesIns_Inst_Sbox_1_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T24_U1 ( .a ({new_AGEMA_signal_4984, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_5359, SubBytesIns_Inst_Sbox_1_T10}), .c ({new_AGEMA_signal_5598, SubBytesIns_Inst_Sbox_1_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T25_U1 ( .a ({new_AGEMA_signal_5362, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_5361, SubBytesIns_Inst_Sbox_1_T17}), .c ({new_AGEMA_signal_5599, SubBytesIns_Inst_Sbox_1_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T26_U1 ( .a ({new_AGEMA_signal_4985, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5177, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_5364, SubBytesIns_Inst_Sbox_1_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T27_U1 ( .a ({new_AGEMA_signal_4983, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_4990, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_5180, SubBytesIns_Inst_Sbox_1_T27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T1_U1 ( .a ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({ciphertext_s1[20], ciphertext_s0[20]}), .c ({new_AGEMA_signal_4993, SubBytesIns_Inst_Sbox_2_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T2_U1 ( .a ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_4994, SubBytesIns_Inst_Sbox_2_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T3_U1 ( .a ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_4995, SubBytesIns_Inst_Sbox_2_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T4_U1 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_4996, SubBytesIns_Inst_Sbox_2_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T5_U1 ( .a ({ciphertext_s1[19], ciphertext_s0[19]}), .b ({ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_4997, SubBytesIns_Inst_Sbox_2_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T6_U1 ( .a ({new_AGEMA_signal_4993, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_4997, SubBytesIns_Inst_Sbox_2_T5}), .c ({new_AGEMA_signal_5181, SubBytesIns_Inst_Sbox_2_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T7_U1 ( .a ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({ciphertext_s1[21], ciphertext_s0[21]}), .c ({new_AGEMA_signal_4998, SubBytesIns_Inst_Sbox_2_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T8_U1 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_5181, SubBytesIns_Inst_Sbox_2_T6}), .c ({new_AGEMA_signal_5371, SubBytesIns_Inst_Sbox_2_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T9_U1 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_4998, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_5182, SubBytesIns_Inst_Sbox_2_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T10_U1 ( .a ({new_AGEMA_signal_5181, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_4998, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_5372, SubBytesIns_Inst_Sbox_2_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T11_U1 ( .a ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_4999, SubBytesIns_Inst_Sbox_2_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T12_U1 ( .a ({ciphertext_s1[21], ciphertext_s0[21]}), .b ({ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_5000, SubBytesIns_Inst_Sbox_2_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T13_U1 ( .a ({new_AGEMA_signal_4995, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_4996, SubBytesIns_Inst_Sbox_2_T4}), .c ({new_AGEMA_signal_5183, SubBytesIns_Inst_Sbox_2_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T14_U1 ( .a ({new_AGEMA_signal_5181, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_4999, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_5373, SubBytesIns_Inst_Sbox_2_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T15_U1 ( .a ({new_AGEMA_signal_4997, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_4999, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_5184, SubBytesIns_Inst_Sbox_2_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T16_U1 ( .a ({new_AGEMA_signal_4997, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_5000, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_5185, SubBytesIns_Inst_Sbox_2_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T17_U1 ( .a ({new_AGEMA_signal_5182, SubBytesIns_Inst_Sbox_2_T9}), .b ({new_AGEMA_signal_5185, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_5374, SubBytesIns_Inst_Sbox_2_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T18_U1 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_5001, SubBytesIns_Inst_Sbox_2_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T19_U1 ( .a ({new_AGEMA_signal_4998, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5001, SubBytesIns_Inst_Sbox_2_T18}), .c ({new_AGEMA_signal_5186, SubBytesIns_Inst_Sbox_2_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T20_U1 ( .a ({new_AGEMA_signal_4993, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5186, SubBytesIns_Inst_Sbox_2_T19}), .c ({new_AGEMA_signal_5375, SubBytesIns_Inst_Sbox_2_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T21_U1 ( .a ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_5002, SubBytesIns_Inst_Sbox_2_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T22_U1 ( .a ({new_AGEMA_signal_4998, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5002, SubBytesIns_Inst_Sbox_2_T21}), .c ({new_AGEMA_signal_5187, SubBytesIns_Inst_Sbox_2_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T23_U1 ( .a ({new_AGEMA_signal_4994, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_5187, SubBytesIns_Inst_Sbox_2_T22}), .c ({new_AGEMA_signal_5376, SubBytesIns_Inst_Sbox_2_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T24_U1 ( .a ({new_AGEMA_signal_4994, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_5372, SubBytesIns_Inst_Sbox_2_T10}), .c ({new_AGEMA_signal_5607, SubBytesIns_Inst_Sbox_2_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T25_U1 ( .a ({new_AGEMA_signal_5375, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_5374, SubBytesIns_Inst_Sbox_2_T17}), .c ({new_AGEMA_signal_5608, SubBytesIns_Inst_Sbox_2_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T26_U1 ( .a ({new_AGEMA_signal_4995, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5185, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_5377, SubBytesIns_Inst_Sbox_2_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T27_U1 ( .a ({new_AGEMA_signal_4993, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5000, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_5188, SubBytesIns_Inst_Sbox_2_T27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T1_U1 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_5003, SubBytesIns_Inst_Sbox_3_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T2_U1 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5004, SubBytesIns_Inst_Sbox_3_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T3_U1 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_5005, SubBytesIns_Inst_Sbox_3_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T4_U1 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5006, SubBytesIns_Inst_Sbox_3_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T5_U1 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_5007, SubBytesIns_Inst_Sbox_3_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T6_U1 ( .a ({new_AGEMA_signal_5003, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5007, SubBytesIns_Inst_Sbox_3_T5}), .c ({new_AGEMA_signal_5189, SubBytesIns_Inst_Sbox_3_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T7_U1 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_5008, SubBytesIns_Inst_Sbox_3_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T8_U1 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_5189, SubBytesIns_Inst_Sbox_3_T6}), .c ({new_AGEMA_signal_5384, SubBytesIns_Inst_Sbox_3_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T9_U1 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_5008, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_5190, SubBytesIns_Inst_Sbox_3_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T10_U1 ( .a ({new_AGEMA_signal_5189, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5008, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_5385, SubBytesIns_Inst_Sbox_3_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T11_U1 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5009, SubBytesIns_Inst_Sbox_3_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T12_U1 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5010, SubBytesIns_Inst_Sbox_3_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T13_U1 ( .a ({new_AGEMA_signal_5005, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5006, SubBytesIns_Inst_Sbox_3_T4}), .c ({new_AGEMA_signal_5191, SubBytesIns_Inst_Sbox_3_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T14_U1 ( .a ({new_AGEMA_signal_5189, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5009, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_5386, SubBytesIns_Inst_Sbox_3_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T15_U1 ( .a ({new_AGEMA_signal_5007, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5009, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_5192, SubBytesIns_Inst_Sbox_3_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T16_U1 ( .a ({new_AGEMA_signal_5007, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5010, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_5193, SubBytesIns_Inst_Sbox_3_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T17_U1 ( .a ({new_AGEMA_signal_5190, SubBytesIns_Inst_Sbox_3_T9}), .b ({new_AGEMA_signal_5193, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_5387, SubBytesIns_Inst_Sbox_3_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T18_U1 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_5011, SubBytesIns_Inst_Sbox_3_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T19_U1 ( .a ({new_AGEMA_signal_5008, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5011, SubBytesIns_Inst_Sbox_3_T18}), .c ({new_AGEMA_signal_5194, SubBytesIns_Inst_Sbox_3_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T20_U1 ( .a ({new_AGEMA_signal_5003, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5194, SubBytesIns_Inst_Sbox_3_T19}), .c ({new_AGEMA_signal_5388, SubBytesIns_Inst_Sbox_3_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T21_U1 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_5012, SubBytesIns_Inst_Sbox_3_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T22_U1 ( .a ({new_AGEMA_signal_5008, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5012, SubBytesIns_Inst_Sbox_3_T21}), .c ({new_AGEMA_signal_5195, SubBytesIns_Inst_Sbox_3_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T23_U1 ( .a ({new_AGEMA_signal_5004, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_5195, SubBytesIns_Inst_Sbox_3_T22}), .c ({new_AGEMA_signal_5389, SubBytesIns_Inst_Sbox_3_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T24_U1 ( .a ({new_AGEMA_signal_5004, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_5385, SubBytesIns_Inst_Sbox_3_T10}), .c ({new_AGEMA_signal_5616, SubBytesIns_Inst_Sbox_3_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T25_U1 ( .a ({new_AGEMA_signal_5388, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_5387, SubBytesIns_Inst_Sbox_3_T17}), .c ({new_AGEMA_signal_5617, SubBytesIns_Inst_Sbox_3_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T26_U1 ( .a ({new_AGEMA_signal_5005, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5193, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_5390, SubBytesIns_Inst_Sbox_3_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T27_U1 ( .a ({new_AGEMA_signal_5003, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5010, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_5196, SubBytesIns_Inst_Sbox_3_T27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T1_U1 ( .a ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({ciphertext_s1[36], ciphertext_s0[36]}), .c ({new_AGEMA_signal_5013, SubBytesIns_Inst_Sbox_4_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T2_U1 ( .a ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5014, SubBytesIns_Inst_Sbox_4_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T3_U1 ( .a ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_5015, SubBytesIns_Inst_Sbox_4_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T4_U1 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5016, SubBytesIns_Inst_Sbox_4_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T5_U1 ( .a ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_5017, SubBytesIns_Inst_Sbox_4_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T6_U1 ( .a ({new_AGEMA_signal_5013, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5017, SubBytesIns_Inst_Sbox_4_T5}), .c ({new_AGEMA_signal_5197, SubBytesIns_Inst_Sbox_4_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T7_U1 ( .a ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({ciphertext_s1[37], ciphertext_s0[37]}), .c ({new_AGEMA_signal_5018, SubBytesIns_Inst_Sbox_4_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T8_U1 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_5197, SubBytesIns_Inst_Sbox_4_T6}), .c ({new_AGEMA_signal_5397, SubBytesIns_Inst_Sbox_4_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T9_U1 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_5018, SubBytesIns_Inst_Sbox_4_T7}), .c ({new_AGEMA_signal_5198, SubBytesIns_Inst_Sbox_4_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T10_U1 ( .a ({new_AGEMA_signal_5197, SubBytesIns_Inst_Sbox_4_T6}), .b ({new_AGEMA_signal_5018, SubBytesIns_Inst_Sbox_4_T7}), .c ({new_AGEMA_signal_5398, SubBytesIns_Inst_Sbox_4_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T11_U1 ( .a ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5019, SubBytesIns_Inst_Sbox_4_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T12_U1 ( .a ({ciphertext_s1[37], ciphertext_s0[37]}), .b ({ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5020, SubBytesIns_Inst_Sbox_4_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T13_U1 ( .a ({new_AGEMA_signal_5015, SubBytesIns_Inst_Sbox_4_T3}), .b ({new_AGEMA_signal_5016, SubBytesIns_Inst_Sbox_4_T4}), .c ({new_AGEMA_signal_5199, SubBytesIns_Inst_Sbox_4_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T14_U1 ( .a ({new_AGEMA_signal_5197, SubBytesIns_Inst_Sbox_4_T6}), .b ({new_AGEMA_signal_5019, SubBytesIns_Inst_Sbox_4_T11}), .c ({new_AGEMA_signal_5399, SubBytesIns_Inst_Sbox_4_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T15_U1 ( .a ({new_AGEMA_signal_5017, SubBytesIns_Inst_Sbox_4_T5}), .b ({new_AGEMA_signal_5019, SubBytesIns_Inst_Sbox_4_T11}), .c ({new_AGEMA_signal_5200, SubBytesIns_Inst_Sbox_4_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T16_U1 ( .a ({new_AGEMA_signal_5017, SubBytesIns_Inst_Sbox_4_T5}), .b ({new_AGEMA_signal_5020, SubBytesIns_Inst_Sbox_4_T12}), .c ({new_AGEMA_signal_5201, SubBytesIns_Inst_Sbox_4_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T17_U1 ( .a ({new_AGEMA_signal_5198, SubBytesIns_Inst_Sbox_4_T9}), .b ({new_AGEMA_signal_5201, SubBytesIns_Inst_Sbox_4_T16}), .c ({new_AGEMA_signal_5400, SubBytesIns_Inst_Sbox_4_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T18_U1 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_5021, SubBytesIns_Inst_Sbox_4_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T19_U1 ( .a ({new_AGEMA_signal_5018, SubBytesIns_Inst_Sbox_4_T7}), .b ({new_AGEMA_signal_5021, SubBytesIns_Inst_Sbox_4_T18}), .c ({new_AGEMA_signal_5202, SubBytesIns_Inst_Sbox_4_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T20_U1 ( .a ({new_AGEMA_signal_5013, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5202, SubBytesIns_Inst_Sbox_4_T19}), .c ({new_AGEMA_signal_5401, SubBytesIns_Inst_Sbox_4_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T21_U1 ( .a ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_5022, SubBytesIns_Inst_Sbox_4_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T22_U1 ( .a ({new_AGEMA_signal_5018, SubBytesIns_Inst_Sbox_4_T7}), .b ({new_AGEMA_signal_5022, SubBytesIns_Inst_Sbox_4_T21}), .c ({new_AGEMA_signal_5203, SubBytesIns_Inst_Sbox_4_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T23_U1 ( .a ({new_AGEMA_signal_5014, SubBytesIns_Inst_Sbox_4_T2}), .b ({new_AGEMA_signal_5203, SubBytesIns_Inst_Sbox_4_T22}), .c ({new_AGEMA_signal_5402, SubBytesIns_Inst_Sbox_4_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T24_U1 ( .a ({new_AGEMA_signal_5014, SubBytesIns_Inst_Sbox_4_T2}), .b ({new_AGEMA_signal_5398, SubBytesIns_Inst_Sbox_4_T10}), .c ({new_AGEMA_signal_5625, SubBytesIns_Inst_Sbox_4_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T25_U1 ( .a ({new_AGEMA_signal_5401, SubBytesIns_Inst_Sbox_4_T20}), .b ({new_AGEMA_signal_5400, SubBytesIns_Inst_Sbox_4_T17}), .c ({new_AGEMA_signal_5626, SubBytesIns_Inst_Sbox_4_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T26_U1 ( .a ({new_AGEMA_signal_5015, SubBytesIns_Inst_Sbox_4_T3}), .b ({new_AGEMA_signal_5201, SubBytesIns_Inst_Sbox_4_T16}), .c ({new_AGEMA_signal_5403, SubBytesIns_Inst_Sbox_4_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T27_U1 ( .a ({new_AGEMA_signal_5013, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5020, SubBytesIns_Inst_Sbox_4_T12}), .c ({new_AGEMA_signal_5204, SubBytesIns_Inst_Sbox_4_T27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T1_U1 ( .a ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({ciphertext_s1[44], ciphertext_s0[44]}), .c ({new_AGEMA_signal_5023, SubBytesIns_Inst_Sbox_5_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T2_U1 ( .a ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5024, SubBytesIns_Inst_Sbox_5_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T3_U1 ( .a ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_5025, SubBytesIns_Inst_Sbox_5_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T4_U1 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5026, SubBytesIns_Inst_Sbox_5_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T5_U1 ( .a ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_5027, SubBytesIns_Inst_Sbox_5_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T6_U1 ( .a ({new_AGEMA_signal_5023, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5027, SubBytesIns_Inst_Sbox_5_T5}), .c ({new_AGEMA_signal_5205, SubBytesIns_Inst_Sbox_5_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T7_U1 ( .a ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({ciphertext_s1[45], ciphertext_s0[45]}), .c ({new_AGEMA_signal_5028, SubBytesIns_Inst_Sbox_5_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T8_U1 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_5205, SubBytesIns_Inst_Sbox_5_T6}), .c ({new_AGEMA_signal_5410, SubBytesIns_Inst_Sbox_5_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T9_U1 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_5028, SubBytesIns_Inst_Sbox_5_T7}), .c ({new_AGEMA_signal_5206, SubBytesIns_Inst_Sbox_5_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T10_U1 ( .a ({new_AGEMA_signal_5205, SubBytesIns_Inst_Sbox_5_T6}), .b ({new_AGEMA_signal_5028, SubBytesIns_Inst_Sbox_5_T7}), .c ({new_AGEMA_signal_5411, SubBytesIns_Inst_Sbox_5_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T11_U1 ( .a ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5029, SubBytesIns_Inst_Sbox_5_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T12_U1 ( .a ({ciphertext_s1[45], ciphertext_s0[45]}), .b ({ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5030, SubBytesIns_Inst_Sbox_5_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T13_U1 ( .a ({new_AGEMA_signal_5025, SubBytesIns_Inst_Sbox_5_T3}), .b ({new_AGEMA_signal_5026, SubBytesIns_Inst_Sbox_5_T4}), .c ({new_AGEMA_signal_5207, SubBytesIns_Inst_Sbox_5_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T14_U1 ( .a ({new_AGEMA_signal_5205, SubBytesIns_Inst_Sbox_5_T6}), .b ({new_AGEMA_signal_5029, SubBytesIns_Inst_Sbox_5_T11}), .c ({new_AGEMA_signal_5412, SubBytesIns_Inst_Sbox_5_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T15_U1 ( .a ({new_AGEMA_signal_5027, SubBytesIns_Inst_Sbox_5_T5}), .b ({new_AGEMA_signal_5029, SubBytesIns_Inst_Sbox_5_T11}), .c ({new_AGEMA_signal_5208, SubBytesIns_Inst_Sbox_5_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T16_U1 ( .a ({new_AGEMA_signal_5027, SubBytesIns_Inst_Sbox_5_T5}), .b ({new_AGEMA_signal_5030, SubBytesIns_Inst_Sbox_5_T12}), .c ({new_AGEMA_signal_5209, SubBytesIns_Inst_Sbox_5_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T17_U1 ( .a ({new_AGEMA_signal_5206, SubBytesIns_Inst_Sbox_5_T9}), .b ({new_AGEMA_signal_5209, SubBytesIns_Inst_Sbox_5_T16}), .c ({new_AGEMA_signal_5413, SubBytesIns_Inst_Sbox_5_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T18_U1 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_5031, SubBytesIns_Inst_Sbox_5_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T19_U1 ( .a ({new_AGEMA_signal_5028, SubBytesIns_Inst_Sbox_5_T7}), .b ({new_AGEMA_signal_5031, SubBytesIns_Inst_Sbox_5_T18}), .c ({new_AGEMA_signal_5210, SubBytesIns_Inst_Sbox_5_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T20_U1 ( .a ({new_AGEMA_signal_5023, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5210, SubBytesIns_Inst_Sbox_5_T19}), .c ({new_AGEMA_signal_5414, SubBytesIns_Inst_Sbox_5_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T21_U1 ( .a ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_5032, SubBytesIns_Inst_Sbox_5_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T22_U1 ( .a ({new_AGEMA_signal_5028, SubBytesIns_Inst_Sbox_5_T7}), .b ({new_AGEMA_signal_5032, SubBytesIns_Inst_Sbox_5_T21}), .c ({new_AGEMA_signal_5211, SubBytesIns_Inst_Sbox_5_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T23_U1 ( .a ({new_AGEMA_signal_5024, SubBytesIns_Inst_Sbox_5_T2}), .b ({new_AGEMA_signal_5211, SubBytesIns_Inst_Sbox_5_T22}), .c ({new_AGEMA_signal_5415, SubBytesIns_Inst_Sbox_5_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T24_U1 ( .a ({new_AGEMA_signal_5024, SubBytesIns_Inst_Sbox_5_T2}), .b ({new_AGEMA_signal_5411, SubBytesIns_Inst_Sbox_5_T10}), .c ({new_AGEMA_signal_5634, SubBytesIns_Inst_Sbox_5_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T25_U1 ( .a ({new_AGEMA_signal_5414, SubBytesIns_Inst_Sbox_5_T20}), .b ({new_AGEMA_signal_5413, SubBytesIns_Inst_Sbox_5_T17}), .c ({new_AGEMA_signal_5635, SubBytesIns_Inst_Sbox_5_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T26_U1 ( .a ({new_AGEMA_signal_5025, SubBytesIns_Inst_Sbox_5_T3}), .b ({new_AGEMA_signal_5209, SubBytesIns_Inst_Sbox_5_T16}), .c ({new_AGEMA_signal_5416, SubBytesIns_Inst_Sbox_5_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T27_U1 ( .a ({new_AGEMA_signal_5023, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5030, SubBytesIns_Inst_Sbox_5_T12}), .c ({new_AGEMA_signal_5212, SubBytesIns_Inst_Sbox_5_T27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T1_U1 ( .a ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({ciphertext_s1[52], ciphertext_s0[52]}), .c ({new_AGEMA_signal_5033, SubBytesIns_Inst_Sbox_6_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T2_U1 ( .a ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_5034, SubBytesIns_Inst_Sbox_6_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T3_U1 ( .a ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_5035, SubBytesIns_Inst_Sbox_6_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T4_U1 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_5036, SubBytesIns_Inst_Sbox_6_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T5_U1 ( .a ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_5037, SubBytesIns_Inst_Sbox_6_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T6_U1 ( .a ({new_AGEMA_signal_5033, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_5037, SubBytesIns_Inst_Sbox_6_T5}), .c ({new_AGEMA_signal_5213, SubBytesIns_Inst_Sbox_6_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T7_U1 ( .a ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({ciphertext_s1[53], ciphertext_s0[53]}), .c ({new_AGEMA_signal_5038, SubBytesIns_Inst_Sbox_6_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T8_U1 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_5213, SubBytesIns_Inst_Sbox_6_T6}), .c ({new_AGEMA_signal_5423, SubBytesIns_Inst_Sbox_6_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T9_U1 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_5038, SubBytesIns_Inst_Sbox_6_T7}), .c ({new_AGEMA_signal_5214, SubBytesIns_Inst_Sbox_6_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T10_U1 ( .a ({new_AGEMA_signal_5213, SubBytesIns_Inst_Sbox_6_T6}), .b ({new_AGEMA_signal_5038, SubBytesIns_Inst_Sbox_6_T7}), .c ({new_AGEMA_signal_5424, SubBytesIns_Inst_Sbox_6_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T11_U1 ( .a ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_5039, SubBytesIns_Inst_Sbox_6_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T12_U1 ( .a ({ciphertext_s1[53], ciphertext_s0[53]}), .b ({ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_5040, SubBytesIns_Inst_Sbox_6_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T13_U1 ( .a ({new_AGEMA_signal_5035, SubBytesIns_Inst_Sbox_6_T3}), .b ({new_AGEMA_signal_5036, SubBytesIns_Inst_Sbox_6_T4}), .c ({new_AGEMA_signal_5215, SubBytesIns_Inst_Sbox_6_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T14_U1 ( .a ({new_AGEMA_signal_5213, SubBytesIns_Inst_Sbox_6_T6}), .b ({new_AGEMA_signal_5039, SubBytesIns_Inst_Sbox_6_T11}), .c ({new_AGEMA_signal_5425, SubBytesIns_Inst_Sbox_6_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T15_U1 ( .a ({new_AGEMA_signal_5037, SubBytesIns_Inst_Sbox_6_T5}), .b ({new_AGEMA_signal_5039, SubBytesIns_Inst_Sbox_6_T11}), .c ({new_AGEMA_signal_5216, SubBytesIns_Inst_Sbox_6_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T16_U1 ( .a ({new_AGEMA_signal_5037, SubBytesIns_Inst_Sbox_6_T5}), .b ({new_AGEMA_signal_5040, SubBytesIns_Inst_Sbox_6_T12}), .c ({new_AGEMA_signal_5217, SubBytesIns_Inst_Sbox_6_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T17_U1 ( .a ({new_AGEMA_signal_5214, SubBytesIns_Inst_Sbox_6_T9}), .b ({new_AGEMA_signal_5217, SubBytesIns_Inst_Sbox_6_T16}), .c ({new_AGEMA_signal_5426, SubBytesIns_Inst_Sbox_6_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T18_U1 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_5041, SubBytesIns_Inst_Sbox_6_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T19_U1 ( .a ({new_AGEMA_signal_5038, SubBytesIns_Inst_Sbox_6_T7}), .b ({new_AGEMA_signal_5041, SubBytesIns_Inst_Sbox_6_T18}), .c ({new_AGEMA_signal_5218, SubBytesIns_Inst_Sbox_6_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T20_U1 ( .a ({new_AGEMA_signal_5033, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_5218, SubBytesIns_Inst_Sbox_6_T19}), .c ({new_AGEMA_signal_5427, SubBytesIns_Inst_Sbox_6_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T21_U1 ( .a ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_5042, SubBytesIns_Inst_Sbox_6_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T22_U1 ( .a ({new_AGEMA_signal_5038, SubBytesIns_Inst_Sbox_6_T7}), .b ({new_AGEMA_signal_5042, SubBytesIns_Inst_Sbox_6_T21}), .c ({new_AGEMA_signal_5219, SubBytesIns_Inst_Sbox_6_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T23_U1 ( .a ({new_AGEMA_signal_5034, SubBytesIns_Inst_Sbox_6_T2}), .b ({new_AGEMA_signal_5219, SubBytesIns_Inst_Sbox_6_T22}), .c ({new_AGEMA_signal_5428, SubBytesIns_Inst_Sbox_6_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T24_U1 ( .a ({new_AGEMA_signal_5034, SubBytesIns_Inst_Sbox_6_T2}), .b ({new_AGEMA_signal_5424, SubBytesIns_Inst_Sbox_6_T10}), .c ({new_AGEMA_signal_5643, SubBytesIns_Inst_Sbox_6_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T25_U1 ( .a ({new_AGEMA_signal_5427, SubBytesIns_Inst_Sbox_6_T20}), .b ({new_AGEMA_signal_5426, SubBytesIns_Inst_Sbox_6_T17}), .c ({new_AGEMA_signal_5644, SubBytesIns_Inst_Sbox_6_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T26_U1 ( .a ({new_AGEMA_signal_5035, SubBytesIns_Inst_Sbox_6_T3}), .b ({new_AGEMA_signal_5217, SubBytesIns_Inst_Sbox_6_T16}), .c ({new_AGEMA_signal_5429, SubBytesIns_Inst_Sbox_6_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T27_U1 ( .a ({new_AGEMA_signal_5033, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_5040, SubBytesIns_Inst_Sbox_6_T12}), .c ({new_AGEMA_signal_5220, SubBytesIns_Inst_Sbox_6_T27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T1_U1 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_5043, SubBytesIns_Inst_Sbox_7_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T2_U1 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_5044, SubBytesIns_Inst_Sbox_7_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T3_U1 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_5045, SubBytesIns_Inst_Sbox_7_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T4_U1 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_5046, SubBytesIns_Inst_Sbox_7_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T5_U1 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_5047, SubBytesIns_Inst_Sbox_7_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T6_U1 ( .a ({new_AGEMA_signal_5043, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_5047, SubBytesIns_Inst_Sbox_7_T5}), .c ({new_AGEMA_signal_5221, SubBytesIns_Inst_Sbox_7_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T7_U1 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_5048, SubBytesIns_Inst_Sbox_7_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T8_U1 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_5221, SubBytesIns_Inst_Sbox_7_T6}), .c ({new_AGEMA_signal_5436, SubBytesIns_Inst_Sbox_7_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T9_U1 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_5048, SubBytesIns_Inst_Sbox_7_T7}), .c ({new_AGEMA_signal_5222, SubBytesIns_Inst_Sbox_7_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T10_U1 ( .a ({new_AGEMA_signal_5221, SubBytesIns_Inst_Sbox_7_T6}), .b ({new_AGEMA_signal_5048, SubBytesIns_Inst_Sbox_7_T7}), .c ({new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_7_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T11_U1 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_5049, SubBytesIns_Inst_Sbox_7_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T12_U1 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_5050, SubBytesIns_Inst_Sbox_7_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T13_U1 ( .a ({new_AGEMA_signal_5045, SubBytesIns_Inst_Sbox_7_T3}), .b ({new_AGEMA_signal_5046, SubBytesIns_Inst_Sbox_7_T4}), .c ({new_AGEMA_signal_5223, SubBytesIns_Inst_Sbox_7_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T14_U1 ( .a ({new_AGEMA_signal_5221, SubBytesIns_Inst_Sbox_7_T6}), .b ({new_AGEMA_signal_5049, SubBytesIns_Inst_Sbox_7_T11}), .c ({new_AGEMA_signal_5438, SubBytesIns_Inst_Sbox_7_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T15_U1 ( .a ({new_AGEMA_signal_5047, SubBytesIns_Inst_Sbox_7_T5}), .b ({new_AGEMA_signal_5049, SubBytesIns_Inst_Sbox_7_T11}), .c ({new_AGEMA_signal_5224, SubBytesIns_Inst_Sbox_7_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T16_U1 ( .a ({new_AGEMA_signal_5047, SubBytesIns_Inst_Sbox_7_T5}), .b ({new_AGEMA_signal_5050, SubBytesIns_Inst_Sbox_7_T12}), .c ({new_AGEMA_signal_5225, SubBytesIns_Inst_Sbox_7_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T17_U1 ( .a ({new_AGEMA_signal_5222, SubBytesIns_Inst_Sbox_7_T9}), .b ({new_AGEMA_signal_5225, SubBytesIns_Inst_Sbox_7_T16}), .c ({new_AGEMA_signal_5439, SubBytesIns_Inst_Sbox_7_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T18_U1 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_5051, SubBytesIns_Inst_Sbox_7_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T19_U1 ( .a ({new_AGEMA_signal_5048, SubBytesIns_Inst_Sbox_7_T7}), .b ({new_AGEMA_signal_5051, SubBytesIns_Inst_Sbox_7_T18}), .c ({new_AGEMA_signal_5226, SubBytesIns_Inst_Sbox_7_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T20_U1 ( .a ({new_AGEMA_signal_5043, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_5226, SubBytesIns_Inst_Sbox_7_T19}), .c ({new_AGEMA_signal_5440, SubBytesIns_Inst_Sbox_7_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T21_U1 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_5052, SubBytesIns_Inst_Sbox_7_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T22_U1 ( .a ({new_AGEMA_signal_5048, SubBytesIns_Inst_Sbox_7_T7}), .b ({new_AGEMA_signal_5052, SubBytesIns_Inst_Sbox_7_T21}), .c ({new_AGEMA_signal_5227, SubBytesIns_Inst_Sbox_7_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T23_U1 ( .a ({new_AGEMA_signal_5044, SubBytesIns_Inst_Sbox_7_T2}), .b ({new_AGEMA_signal_5227, SubBytesIns_Inst_Sbox_7_T22}), .c ({new_AGEMA_signal_5441, SubBytesIns_Inst_Sbox_7_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T24_U1 ( .a ({new_AGEMA_signal_5044, SubBytesIns_Inst_Sbox_7_T2}), .b ({new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_7_T10}), .c ({new_AGEMA_signal_5652, SubBytesIns_Inst_Sbox_7_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T25_U1 ( .a ({new_AGEMA_signal_5440, SubBytesIns_Inst_Sbox_7_T20}), .b ({new_AGEMA_signal_5439, SubBytesIns_Inst_Sbox_7_T17}), .c ({new_AGEMA_signal_5653, SubBytesIns_Inst_Sbox_7_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T26_U1 ( .a ({new_AGEMA_signal_5045, SubBytesIns_Inst_Sbox_7_T3}), .b ({new_AGEMA_signal_5225, SubBytesIns_Inst_Sbox_7_T16}), .c ({new_AGEMA_signal_5442, SubBytesIns_Inst_Sbox_7_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T27_U1 ( .a ({new_AGEMA_signal_5043, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_5050, SubBytesIns_Inst_Sbox_7_T12}), .c ({new_AGEMA_signal_5228, SubBytesIns_Inst_Sbox_7_T27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T1_U1 ( .a ({ciphertext_s1[71], ciphertext_s0[71]}), .b ({ciphertext_s1[68], ciphertext_s0[68]}), .c ({new_AGEMA_signal_5053, SubBytesIns_Inst_Sbox_8_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T2_U1 ( .a ({ciphertext_s1[71], ciphertext_s0[71]}), .b ({ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_5054, SubBytesIns_Inst_Sbox_8_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T3_U1 ( .a ({ciphertext_s1[71], ciphertext_s0[71]}), .b ({ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_5055, SubBytesIns_Inst_Sbox_8_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T4_U1 ( .a ({ciphertext_s1[68], ciphertext_s0[68]}), .b ({ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_5056, SubBytesIns_Inst_Sbox_8_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T5_U1 ( .a ({ciphertext_s1[67], ciphertext_s0[67]}), .b ({ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_5057, SubBytesIns_Inst_Sbox_8_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T6_U1 ( .a ({new_AGEMA_signal_5053, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_5057, SubBytesIns_Inst_Sbox_8_T5}), .c ({new_AGEMA_signal_5229, SubBytesIns_Inst_Sbox_8_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T7_U1 ( .a ({ciphertext_s1[70], ciphertext_s0[70]}), .b ({ciphertext_s1[69], ciphertext_s0[69]}), .c ({new_AGEMA_signal_5058, SubBytesIns_Inst_Sbox_8_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T8_U1 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({new_AGEMA_signal_5229, SubBytesIns_Inst_Sbox_8_T6}), .c ({new_AGEMA_signal_5449, SubBytesIns_Inst_Sbox_8_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T9_U1 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({new_AGEMA_signal_5058, SubBytesIns_Inst_Sbox_8_T7}), .c ({new_AGEMA_signal_5230, SubBytesIns_Inst_Sbox_8_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T10_U1 ( .a ({new_AGEMA_signal_5229, SubBytesIns_Inst_Sbox_8_T6}), .b ({new_AGEMA_signal_5058, SubBytesIns_Inst_Sbox_8_T7}), .c ({new_AGEMA_signal_5450, SubBytesIns_Inst_Sbox_8_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T11_U1 ( .a ({ciphertext_s1[70], ciphertext_s0[70]}), .b ({ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_5059, SubBytesIns_Inst_Sbox_8_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T12_U1 ( .a ({ciphertext_s1[69], ciphertext_s0[69]}), .b ({ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_5060, SubBytesIns_Inst_Sbox_8_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T13_U1 ( .a ({new_AGEMA_signal_5055, SubBytesIns_Inst_Sbox_8_T3}), .b ({new_AGEMA_signal_5056, SubBytesIns_Inst_Sbox_8_T4}), .c ({new_AGEMA_signal_5231, SubBytesIns_Inst_Sbox_8_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T14_U1 ( .a ({new_AGEMA_signal_5229, SubBytesIns_Inst_Sbox_8_T6}), .b ({new_AGEMA_signal_5059, SubBytesIns_Inst_Sbox_8_T11}), .c ({new_AGEMA_signal_5451, SubBytesIns_Inst_Sbox_8_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T15_U1 ( .a ({new_AGEMA_signal_5057, SubBytesIns_Inst_Sbox_8_T5}), .b ({new_AGEMA_signal_5059, SubBytesIns_Inst_Sbox_8_T11}), .c ({new_AGEMA_signal_5232, SubBytesIns_Inst_Sbox_8_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T16_U1 ( .a ({new_AGEMA_signal_5057, SubBytesIns_Inst_Sbox_8_T5}), .b ({new_AGEMA_signal_5060, SubBytesIns_Inst_Sbox_8_T12}), .c ({new_AGEMA_signal_5233, SubBytesIns_Inst_Sbox_8_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T17_U1 ( .a ({new_AGEMA_signal_5230, SubBytesIns_Inst_Sbox_8_T9}), .b ({new_AGEMA_signal_5233, SubBytesIns_Inst_Sbox_8_T16}), .c ({new_AGEMA_signal_5452, SubBytesIns_Inst_Sbox_8_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T18_U1 ( .a ({ciphertext_s1[68], ciphertext_s0[68]}), .b ({ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_5061, SubBytesIns_Inst_Sbox_8_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T19_U1 ( .a ({new_AGEMA_signal_5058, SubBytesIns_Inst_Sbox_8_T7}), .b ({new_AGEMA_signal_5061, SubBytesIns_Inst_Sbox_8_T18}), .c ({new_AGEMA_signal_5234, SubBytesIns_Inst_Sbox_8_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T20_U1 ( .a ({new_AGEMA_signal_5053, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_5234, SubBytesIns_Inst_Sbox_8_T19}), .c ({new_AGEMA_signal_5453, SubBytesIns_Inst_Sbox_8_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T21_U1 ( .a ({ciphertext_s1[65], ciphertext_s0[65]}), .b ({ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_5062, SubBytesIns_Inst_Sbox_8_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T22_U1 ( .a ({new_AGEMA_signal_5058, SubBytesIns_Inst_Sbox_8_T7}), .b ({new_AGEMA_signal_5062, SubBytesIns_Inst_Sbox_8_T21}), .c ({new_AGEMA_signal_5235, SubBytesIns_Inst_Sbox_8_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T23_U1 ( .a ({new_AGEMA_signal_5054, SubBytesIns_Inst_Sbox_8_T2}), .b ({new_AGEMA_signal_5235, SubBytesIns_Inst_Sbox_8_T22}), .c ({new_AGEMA_signal_5454, SubBytesIns_Inst_Sbox_8_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T24_U1 ( .a ({new_AGEMA_signal_5054, SubBytesIns_Inst_Sbox_8_T2}), .b ({new_AGEMA_signal_5450, SubBytesIns_Inst_Sbox_8_T10}), .c ({new_AGEMA_signal_5661, SubBytesIns_Inst_Sbox_8_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T25_U1 ( .a ({new_AGEMA_signal_5453, SubBytesIns_Inst_Sbox_8_T20}), .b ({new_AGEMA_signal_5452, SubBytesIns_Inst_Sbox_8_T17}), .c ({new_AGEMA_signal_5662, SubBytesIns_Inst_Sbox_8_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T26_U1 ( .a ({new_AGEMA_signal_5055, SubBytesIns_Inst_Sbox_8_T3}), .b ({new_AGEMA_signal_5233, SubBytesIns_Inst_Sbox_8_T16}), .c ({new_AGEMA_signal_5455, SubBytesIns_Inst_Sbox_8_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T27_U1 ( .a ({new_AGEMA_signal_5053, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_5060, SubBytesIns_Inst_Sbox_8_T12}), .c ({new_AGEMA_signal_5236, SubBytesIns_Inst_Sbox_8_T27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T1_U1 ( .a ({ciphertext_s1[79], ciphertext_s0[79]}), .b ({ciphertext_s1[76], ciphertext_s0[76]}), .c ({new_AGEMA_signal_5063, SubBytesIns_Inst_Sbox_9_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T2_U1 ( .a ({ciphertext_s1[79], ciphertext_s0[79]}), .b ({ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_5064, SubBytesIns_Inst_Sbox_9_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T3_U1 ( .a ({ciphertext_s1[79], ciphertext_s0[79]}), .b ({ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_5065, SubBytesIns_Inst_Sbox_9_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T4_U1 ( .a ({ciphertext_s1[76], ciphertext_s0[76]}), .b ({ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_5066, SubBytesIns_Inst_Sbox_9_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T5_U1 ( .a ({ciphertext_s1[75], ciphertext_s0[75]}), .b ({ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_5067, SubBytesIns_Inst_Sbox_9_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T6_U1 ( .a ({new_AGEMA_signal_5063, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_5067, SubBytesIns_Inst_Sbox_9_T5}), .c ({new_AGEMA_signal_5237, SubBytesIns_Inst_Sbox_9_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T7_U1 ( .a ({ciphertext_s1[78], ciphertext_s0[78]}), .b ({ciphertext_s1[77], ciphertext_s0[77]}), .c ({new_AGEMA_signal_5068, SubBytesIns_Inst_Sbox_9_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T8_U1 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({new_AGEMA_signal_5237, SubBytesIns_Inst_Sbox_9_T6}), .c ({new_AGEMA_signal_5462, SubBytesIns_Inst_Sbox_9_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T9_U1 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({new_AGEMA_signal_5068, SubBytesIns_Inst_Sbox_9_T7}), .c ({new_AGEMA_signal_5238, SubBytesIns_Inst_Sbox_9_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T10_U1 ( .a ({new_AGEMA_signal_5237, SubBytesIns_Inst_Sbox_9_T6}), .b ({new_AGEMA_signal_5068, SubBytesIns_Inst_Sbox_9_T7}), .c ({new_AGEMA_signal_5463, SubBytesIns_Inst_Sbox_9_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T11_U1 ( .a ({ciphertext_s1[78], ciphertext_s0[78]}), .b ({ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_5069, SubBytesIns_Inst_Sbox_9_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T12_U1 ( .a ({ciphertext_s1[77], ciphertext_s0[77]}), .b ({ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_5070, SubBytesIns_Inst_Sbox_9_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T13_U1 ( .a ({new_AGEMA_signal_5065, SubBytesIns_Inst_Sbox_9_T3}), .b ({new_AGEMA_signal_5066, SubBytesIns_Inst_Sbox_9_T4}), .c ({new_AGEMA_signal_5239, SubBytesIns_Inst_Sbox_9_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T14_U1 ( .a ({new_AGEMA_signal_5237, SubBytesIns_Inst_Sbox_9_T6}), .b ({new_AGEMA_signal_5069, SubBytesIns_Inst_Sbox_9_T11}), .c ({new_AGEMA_signal_5464, SubBytesIns_Inst_Sbox_9_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T15_U1 ( .a ({new_AGEMA_signal_5067, SubBytesIns_Inst_Sbox_9_T5}), .b ({new_AGEMA_signal_5069, SubBytesIns_Inst_Sbox_9_T11}), .c ({new_AGEMA_signal_5240, SubBytesIns_Inst_Sbox_9_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T16_U1 ( .a ({new_AGEMA_signal_5067, SubBytesIns_Inst_Sbox_9_T5}), .b ({new_AGEMA_signal_5070, SubBytesIns_Inst_Sbox_9_T12}), .c ({new_AGEMA_signal_5241, SubBytesIns_Inst_Sbox_9_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T17_U1 ( .a ({new_AGEMA_signal_5238, SubBytesIns_Inst_Sbox_9_T9}), .b ({new_AGEMA_signal_5241, SubBytesIns_Inst_Sbox_9_T16}), .c ({new_AGEMA_signal_5465, SubBytesIns_Inst_Sbox_9_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T18_U1 ( .a ({ciphertext_s1[76], ciphertext_s0[76]}), .b ({ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_5071, SubBytesIns_Inst_Sbox_9_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T19_U1 ( .a ({new_AGEMA_signal_5068, SubBytesIns_Inst_Sbox_9_T7}), .b ({new_AGEMA_signal_5071, SubBytesIns_Inst_Sbox_9_T18}), .c ({new_AGEMA_signal_5242, SubBytesIns_Inst_Sbox_9_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T20_U1 ( .a ({new_AGEMA_signal_5063, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_5242, SubBytesIns_Inst_Sbox_9_T19}), .c ({new_AGEMA_signal_5466, SubBytesIns_Inst_Sbox_9_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T21_U1 ( .a ({ciphertext_s1[73], ciphertext_s0[73]}), .b ({ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_5072, SubBytesIns_Inst_Sbox_9_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T22_U1 ( .a ({new_AGEMA_signal_5068, SubBytesIns_Inst_Sbox_9_T7}), .b ({new_AGEMA_signal_5072, SubBytesIns_Inst_Sbox_9_T21}), .c ({new_AGEMA_signal_5243, SubBytesIns_Inst_Sbox_9_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T23_U1 ( .a ({new_AGEMA_signal_5064, SubBytesIns_Inst_Sbox_9_T2}), .b ({new_AGEMA_signal_5243, SubBytesIns_Inst_Sbox_9_T22}), .c ({new_AGEMA_signal_5467, SubBytesIns_Inst_Sbox_9_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T24_U1 ( .a ({new_AGEMA_signal_5064, SubBytesIns_Inst_Sbox_9_T2}), .b ({new_AGEMA_signal_5463, SubBytesIns_Inst_Sbox_9_T10}), .c ({new_AGEMA_signal_5670, SubBytesIns_Inst_Sbox_9_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T25_U1 ( .a ({new_AGEMA_signal_5466, SubBytesIns_Inst_Sbox_9_T20}), .b ({new_AGEMA_signal_5465, SubBytesIns_Inst_Sbox_9_T17}), .c ({new_AGEMA_signal_5671, SubBytesIns_Inst_Sbox_9_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T26_U1 ( .a ({new_AGEMA_signal_5065, SubBytesIns_Inst_Sbox_9_T3}), .b ({new_AGEMA_signal_5241, SubBytesIns_Inst_Sbox_9_T16}), .c ({new_AGEMA_signal_5468, SubBytesIns_Inst_Sbox_9_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T27_U1 ( .a ({new_AGEMA_signal_5063, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_5070, SubBytesIns_Inst_Sbox_9_T12}), .c ({new_AGEMA_signal_5244, SubBytesIns_Inst_Sbox_9_T27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T1_U1 ( .a ({ciphertext_s1[87], ciphertext_s0[87]}), .b ({ciphertext_s1[84], ciphertext_s0[84]}), .c ({new_AGEMA_signal_5073, SubBytesIns_Inst_Sbox_10_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T2_U1 ( .a ({ciphertext_s1[87], ciphertext_s0[87]}), .b ({ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_5074, SubBytesIns_Inst_Sbox_10_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T3_U1 ( .a ({ciphertext_s1[87], ciphertext_s0[87]}), .b ({ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_5075, SubBytesIns_Inst_Sbox_10_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T4_U1 ( .a ({ciphertext_s1[84], ciphertext_s0[84]}), .b ({ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_5076, SubBytesIns_Inst_Sbox_10_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T5_U1 ( .a ({ciphertext_s1[83], ciphertext_s0[83]}), .b ({ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_5077, SubBytesIns_Inst_Sbox_10_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T6_U1 ( .a ({new_AGEMA_signal_5073, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_5077, SubBytesIns_Inst_Sbox_10_T5}), .c ({new_AGEMA_signal_5245, SubBytesIns_Inst_Sbox_10_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T7_U1 ( .a ({ciphertext_s1[86], ciphertext_s0[86]}), .b ({ciphertext_s1[85], ciphertext_s0[85]}), .c ({new_AGEMA_signal_5078, SubBytesIns_Inst_Sbox_10_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T8_U1 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({new_AGEMA_signal_5245, SubBytesIns_Inst_Sbox_10_T6}), .c ({new_AGEMA_signal_5475, SubBytesIns_Inst_Sbox_10_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T9_U1 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({new_AGEMA_signal_5078, SubBytesIns_Inst_Sbox_10_T7}), .c ({new_AGEMA_signal_5246, SubBytesIns_Inst_Sbox_10_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T10_U1 ( .a ({new_AGEMA_signal_5245, SubBytesIns_Inst_Sbox_10_T6}), .b ({new_AGEMA_signal_5078, SubBytesIns_Inst_Sbox_10_T7}), .c ({new_AGEMA_signal_5476, SubBytesIns_Inst_Sbox_10_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T11_U1 ( .a ({ciphertext_s1[86], ciphertext_s0[86]}), .b ({ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_5079, SubBytesIns_Inst_Sbox_10_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T12_U1 ( .a ({ciphertext_s1[85], ciphertext_s0[85]}), .b ({ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_5080, SubBytesIns_Inst_Sbox_10_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T13_U1 ( .a ({new_AGEMA_signal_5075, SubBytesIns_Inst_Sbox_10_T3}), .b ({new_AGEMA_signal_5076, SubBytesIns_Inst_Sbox_10_T4}), .c ({new_AGEMA_signal_5247, SubBytesIns_Inst_Sbox_10_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T14_U1 ( .a ({new_AGEMA_signal_5245, SubBytesIns_Inst_Sbox_10_T6}), .b ({new_AGEMA_signal_5079, SubBytesIns_Inst_Sbox_10_T11}), .c ({new_AGEMA_signal_5477, SubBytesIns_Inst_Sbox_10_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T15_U1 ( .a ({new_AGEMA_signal_5077, SubBytesIns_Inst_Sbox_10_T5}), .b ({new_AGEMA_signal_5079, SubBytesIns_Inst_Sbox_10_T11}), .c ({new_AGEMA_signal_5248, SubBytesIns_Inst_Sbox_10_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T16_U1 ( .a ({new_AGEMA_signal_5077, SubBytesIns_Inst_Sbox_10_T5}), .b ({new_AGEMA_signal_5080, SubBytesIns_Inst_Sbox_10_T12}), .c ({new_AGEMA_signal_5249, SubBytesIns_Inst_Sbox_10_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T17_U1 ( .a ({new_AGEMA_signal_5246, SubBytesIns_Inst_Sbox_10_T9}), .b ({new_AGEMA_signal_5249, SubBytesIns_Inst_Sbox_10_T16}), .c ({new_AGEMA_signal_5478, SubBytesIns_Inst_Sbox_10_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T18_U1 ( .a ({ciphertext_s1[84], ciphertext_s0[84]}), .b ({ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_5081, SubBytesIns_Inst_Sbox_10_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T19_U1 ( .a ({new_AGEMA_signal_5078, SubBytesIns_Inst_Sbox_10_T7}), .b ({new_AGEMA_signal_5081, SubBytesIns_Inst_Sbox_10_T18}), .c ({new_AGEMA_signal_5250, SubBytesIns_Inst_Sbox_10_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T20_U1 ( .a ({new_AGEMA_signal_5073, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_5250, SubBytesIns_Inst_Sbox_10_T19}), .c ({new_AGEMA_signal_5479, SubBytesIns_Inst_Sbox_10_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T21_U1 ( .a ({ciphertext_s1[81], ciphertext_s0[81]}), .b ({ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_5082, SubBytesIns_Inst_Sbox_10_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T22_U1 ( .a ({new_AGEMA_signal_5078, SubBytesIns_Inst_Sbox_10_T7}), .b ({new_AGEMA_signal_5082, SubBytesIns_Inst_Sbox_10_T21}), .c ({new_AGEMA_signal_5251, SubBytesIns_Inst_Sbox_10_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T23_U1 ( .a ({new_AGEMA_signal_5074, SubBytesIns_Inst_Sbox_10_T2}), .b ({new_AGEMA_signal_5251, SubBytesIns_Inst_Sbox_10_T22}), .c ({new_AGEMA_signal_5480, SubBytesIns_Inst_Sbox_10_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T24_U1 ( .a ({new_AGEMA_signal_5074, SubBytesIns_Inst_Sbox_10_T2}), .b ({new_AGEMA_signal_5476, SubBytesIns_Inst_Sbox_10_T10}), .c ({new_AGEMA_signal_5679, SubBytesIns_Inst_Sbox_10_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T25_U1 ( .a ({new_AGEMA_signal_5479, SubBytesIns_Inst_Sbox_10_T20}), .b ({new_AGEMA_signal_5478, SubBytesIns_Inst_Sbox_10_T17}), .c ({new_AGEMA_signal_5680, SubBytesIns_Inst_Sbox_10_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T26_U1 ( .a ({new_AGEMA_signal_5075, SubBytesIns_Inst_Sbox_10_T3}), .b ({new_AGEMA_signal_5249, SubBytesIns_Inst_Sbox_10_T16}), .c ({new_AGEMA_signal_5481, SubBytesIns_Inst_Sbox_10_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T27_U1 ( .a ({new_AGEMA_signal_5073, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_5080, SubBytesIns_Inst_Sbox_10_T12}), .c ({new_AGEMA_signal_5252, SubBytesIns_Inst_Sbox_10_T27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T1_U1 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_5083, SubBytesIns_Inst_Sbox_11_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T2_U1 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_5084, SubBytesIns_Inst_Sbox_11_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T3_U1 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_5085, SubBytesIns_Inst_Sbox_11_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T4_U1 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_5086, SubBytesIns_Inst_Sbox_11_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T5_U1 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_5087, SubBytesIns_Inst_Sbox_11_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T6_U1 ( .a ({new_AGEMA_signal_5083, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_5087, SubBytesIns_Inst_Sbox_11_T5}), .c ({new_AGEMA_signal_5253, SubBytesIns_Inst_Sbox_11_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T7_U1 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_5088, SubBytesIns_Inst_Sbox_11_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T8_U1 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({new_AGEMA_signal_5253, SubBytesIns_Inst_Sbox_11_T6}), .c ({new_AGEMA_signal_5488, SubBytesIns_Inst_Sbox_11_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T9_U1 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({new_AGEMA_signal_5088, SubBytesIns_Inst_Sbox_11_T7}), .c ({new_AGEMA_signal_5254, SubBytesIns_Inst_Sbox_11_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T10_U1 ( .a ({new_AGEMA_signal_5253, SubBytesIns_Inst_Sbox_11_T6}), .b ({new_AGEMA_signal_5088, SubBytesIns_Inst_Sbox_11_T7}), .c ({new_AGEMA_signal_5489, SubBytesIns_Inst_Sbox_11_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T11_U1 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_5089, SubBytesIns_Inst_Sbox_11_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T12_U1 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_5090, SubBytesIns_Inst_Sbox_11_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T13_U1 ( .a ({new_AGEMA_signal_5085, SubBytesIns_Inst_Sbox_11_T3}), .b ({new_AGEMA_signal_5086, SubBytesIns_Inst_Sbox_11_T4}), .c ({new_AGEMA_signal_5255, SubBytesIns_Inst_Sbox_11_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T14_U1 ( .a ({new_AGEMA_signal_5253, SubBytesIns_Inst_Sbox_11_T6}), .b ({new_AGEMA_signal_5089, SubBytesIns_Inst_Sbox_11_T11}), .c ({new_AGEMA_signal_5490, SubBytesIns_Inst_Sbox_11_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T15_U1 ( .a ({new_AGEMA_signal_5087, SubBytesIns_Inst_Sbox_11_T5}), .b ({new_AGEMA_signal_5089, SubBytesIns_Inst_Sbox_11_T11}), .c ({new_AGEMA_signal_5256, SubBytesIns_Inst_Sbox_11_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T16_U1 ( .a ({new_AGEMA_signal_5087, SubBytesIns_Inst_Sbox_11_T5}), .b ({new_AGEMA_signal_5090, SubBytesIns_Inst_Sbox_11_T12}), .c ({new_AGEMA_signal_5257, SubBytesIns_Inst_Sbox_11_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T17_U1 ( .a ({new_AGEMA_signal_5254, SubBytesIns_Inst_Sbox_11_T9}), .b ({new_AGEMA_signal_5257, SubBytesIns_Inst_Sbox_11_T16}), .c ({new_AGEMA_signal_5491, SubBytesIns_Inst_Sbox_11_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T18_U1 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_5091, SubBytesIns_Inst_Sbox_11_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T19_U1 ( .a ({new_AGEMA_signal_5088, SubBytesIns_Inst_Sbox_11_T7}), .b ({new_AGEMA_signal_5091, SubBytesIns_Inst_Sbox_11_T18}), .c ({new_AGEMA_signal_5258, SubBytesIns_Inst_Sbox_11_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T20_U1 ( .a ({new_AGEMA_signal_5083, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_5258, SubBytesIns_Inst_Sbox_11_T19}), .c ({new_AGEMA_signal_5492, SubBytesIns_Inst_Sbox_11_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T21_U1 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_5092, SubBytesIns_Inst_Sbox_11_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T22_U1 ( .a ({new_AGEMA_signal_5088, SubBytesIns_Inst_Sbox_11_T7}), .b ({new_AGEMA_signal_5092, SubBytesIns_Inst_Sbox_11_T21}), .c ({new_AGEMA_signal_5259, SubBytesIns_Inst_Sbox_11_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T23_U1 ( .a ({new_AGEMA_signal_5084, SubBytesIns_Inst_Sbox_11_T2}), .b ({new_AGEMA_signal_5259, SubBytesIns_Inst_Sbox_11_T22}), .c ({new_AGEMA_signal_5493, SubBytesIns_Inst_Sbox_11_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T24_U1 ( .a ({new_AGEMA_signal_5084, SubBytesIns_Inst_Sbox_11_T2}), .b ({new_AGEMA_signal_5489, SubBytesIns_Inst_Sbox_11_T10}), .c ({new_AGEMA_signal_5688, SubBytesIns_Inst_Sbox_11_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T25_U1 ( .a ({new_AGEMA_signal_5492, SubBytesIns_Inst_Sbox_11_T20}), .b ({new_AGEMA_signal_5491, SubBytesIns_Inst_Sbox_11_T17}), .c ({new_AGEMA_signal_5689, SubBytesIns_Inst_Sbox_11_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T26_U1 ( .a ({new_AGEMA_signal_5085, SubBytesIns_Inst_Sbox_11_T3}), .b ({new_AGEMA_signal_5257, SubBytesIns_Inst_Sbox_11_T16}), .c ({new_AGEMA_signal_5494, SubBytesIns_Inst_Sbox_11_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T27_U1 ( .a ({new_AGEMA_signal_5083, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_5090, SubBytesIns_Inst_Sbox_11_T12}), .c ({new_AGEMA_signal_5260, SubBytesIns_Inst_Sbox_11_T27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T1_U1 ( .a ({ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s1[100], ciphertext_s0[100]}), .c ({new_AGEMA_signal_5093, SubBytesIns_Inst_Sbox_12_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T2_U1 ( .a ({ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_5094, SubBytesIns_Inst_Sbox_12_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T3_U1 ( .a ({ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_5095, SubBytesIns_Inst_Sbox_12_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T4_U1 ( .a ({ciphertext_s1[100], ciphertext_s0[100]}), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_5096, SubBytesIns_Inst_Sbox_12_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T5_U1 ( .a ({ciphertext_s1[99], ciphertext_s0[99]}), .b ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_5097, SubBytesIns_Inst_Sbox_12_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T6_U1 ( .a ({new_AGEMA_signal_5093, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_5097, SubBytesIns_Inst_Sbox_12_T5}), .c ({new_AGEMA_signal_5261, SubBytesIns_Inst_Sbox_12_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T7_U1 ( .a ({ciphertext_s1[102], ciphertext_s0[102]}), .b ({ciphertext_s1[101], ciphertext_s0[101]}), .c ({new_AGEMA_signal_5098, SubBytesIns_Inst_Sbox_12_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T8_U1 ( .a ({ciphertext_s1[96], ciphertext_s0[96]}), .b ({new_AGEMA_signal_5261, SubBytesIns_Inst_Sbox_12_T6}), .c ({new_AGEMA_signal_5501, SubBytesIns_Inst_Sbox_12_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T9_U1 ( .a ({ciphertext_s1[96], ciphertext_s0[96]}), .b ({new_AGEMA_signal_5098, SubBytesIns_Inst_Sbox_12_T7}), .c ({new_AGEMA_signal_5262, SubBytesIns_Inst_Sbox_12_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T10_U1 ( .a ({new_AGEMA_signal_5261, SubBytesIns_Inst_Sbox_12_T6}), .b ({new_AGEMA_signal_5098, SubBytesIns_Inst_Sbox_12_T7}), .c ({new_AGEMA_signal_5502, SubBytesIns_Inst_Sbox_12_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T11_U1 ( .a ({ciphertext_s1[102], ciphertext_s0[102]}), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_5099, SubBytesIns_Inst_Sbox_12_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T12_U1 ( .a ({ciphertext_s1[101], ciphertext_s0[101]}), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_5100, SubBytesIns_Inst_Sbox_12_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T13_U1 ( .a ({new_AGEMA_signal_5095, SubBytesIns_Inst_Sbox_12_T3}), .b ({new_AGEMA_signal_5096, SubBytesIns_Inst_Sbox_12_T4}), .c ({new_AGEMA_signal_5263, SubBytesIns_Inst_Sbox_12_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T14_U1 ( .a ({new_AGEMA_signal_5261, SubBytesIns_Inst_Sbox_12_T6}), .b ({new_AGEMA_signal_5099, SubBytesIns_Inst_Sbox_12_T11}), .c ({new_AGEMA_signal_5503, SubBytesIns_Inst_Sbox_12_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T15_U1 ( .a ({new_AGEMA_signal_5097, SubBytesIns_Inst_Sbox_12_T5}), .b ({new_AGEMA_signal_5099, SubBytesIns_Inst_Sbox_12_T11}), .c ({new_AGEMA_signal_5264, SubBytesIns_Inst_Sbox_12_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T16_U1 ( .a ({new_AGEMA_signal_5097, SubBytesIns_Inst_Sbox_12_T5}), .b ({new_AGEMA_signal_5100, SubBytesIns_Inst_Sbox_12_T12}), .c ({new_AGEMA_signal_5265, SubBytesIns_Inst_Sbox_12_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T17_U1 ( .a ({new_AGEMA_signal_5262, SubBytesIns_Inst_Sbox_12_T9}), .b ({new_AGEMA_signal_5265, SubBytesIns_Inst_Sbox_12_T16}), .c ({new_AGEMA_signal_5504, SubBytesIns_Inst_Sbox_12_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T18_U1 ( .a ({ciphertext_s1[100], ciphertext_s0[100]}), .b ({ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_5101, SubBytesIns_Inst_Sbox_12_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T19_U1 ( .a ({new_AGEMA_signal_5098, SubBytesIns_Inst_Sbox_12_T7}), .b ({new_AGEMA_signal_5101, SubBytesIns_Inst_Sbox_12_T18}), .c ({new_AGEMA_signal_5266, SubBytesIns_Inst_Sbox_12_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T20_U1 ( .a ({new_AGEMA_signal_5093, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_5266, SubBytesIns_Inst_Sbox_12_T19}), .c ({new_AGEMA_signal_5505, SubBytesIns_Inst_Sbox_12_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T21_U1 ( .a ({ciphertext_s1[97], ciphertext_s0[97]}), .b ({ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_5102, SubBytesIns_Inst_Sbox_12_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T22_U1 ( .a ({new_AGEMA_signal_5098, SubBytesIns_Inst_Sbox_12_T7}), .b ({new_AGEMA_signal_5102, SubBytesIns_Inst_Sbox_12_T21}), .c ({new_AGEMA_signal_5267, SubBytesIns_Inst_Sbox_12_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T23_U1 ( .a ({new_AGEMA_signal_5094, SubBytesIns_Inst_Sbox_12_T2}), .b ({new_AGEMA_signal_5267, SubBytesIns_Inst_Sbox_12_T22}), .c ({new_AGEMA_signal_5506, SubBytesIns_Inst_Sbox_12_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T24_U1 ( .a ({new_AGEMA_signal_5094, SubBytesIns_Inst_Sbox_12_T2}), .b ({new_AGEMA_signal_5502, SubBytesIns_Inst_Sbox_12_T10}), .c ({new_AGEMA_signal_5697, SubBytesIns_Inst_Sbox_12_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T25_U1 ( .a ({new_AGEMA_signal_5505, SubBytesIns_Inst_Sbox_12_T20}), .b ({new_AGEMA_signal_5504, SubBytesIns_Inst_Sbox_12_T17}), .c ({new_AGEMA_signal_5698, SubBytesIns_Inst_Sbox_12_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T26_U1 ( .a ({new_AGEMA_signal_5095, SubBytesIns_Inst_Sbox_12_T3}), .b ({new_AGEMA_signal_5265, SubBytesIns_Inst_Sbox_12_T16}), .c ({new_AGEMA_signal_5507, SubBytesIns_Inst_Sbox_12_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T27_U1 ( .a ({new_AGEMA_signal_5093, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_5100, SubBytesIns_Inst_Sbox_12_T12}), .c ({new_AGEMA_signal_5268, SubBytesIns_Inst_Sbox_12_T27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T1_U1 ( .a ({ciphertext_s1[111], ciphertext_s0[111]}), .b ({ciphertext_s1[108], ciphertext_s0[108]}), .c ({new_AGEMA_signal_5103, SubBytesIns_Inst_Sbox_13_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T2_U1 ( .a ({ciphertext_s1[111], ciphertext_s0[111]}), .b ({ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_5104, SubBytesIns_Inst_Sbox_13_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T3_U1 ( .a ({ciphertext_s1[111], ciphertext_s0[111]}), .b ({ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_5105, SubBytesIns_Inst_Sbox_13_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T4_U1 ( .a ({ciphertext_s1[108], ciphertext_s0[108]}), .b ({ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_5106, SubBytesIns_Inst_Sbox_13_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T5_U1 ( .a ({ciphertext_s1[107], ciphertext_s0[107]}), .b ({ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_5107, SubBytesIns_Inst_Sbox_13_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T6_U1 ( .a ({new_AGEMA_signal_5103, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_5107, SubBytesIns_Inst_Sbox_13_T5}), .c ({new_AGEMA_signal_5269, SubBytesIns_Inst_Sbox_13_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T7_U1 ( .a ({ciphertext_s1[110], ciphertext_s0[110]}), .b ({ciphertext_s1[109], ciphertext_s0[109]}), .c ({new_AGEMA_signal_5108, SubBytesIns_Inst_Sbox_13_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T8_U1 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({new_AGEMA_signal_5269, SubBytesIns_Inst_Sbox_13_T6}), .c ({new_AGEMA_signal_5514, SubBytesIns_Inst_Sbox_13_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T9_U1 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({new_AGEMA_signal_5108, SubBytesIns_Inst_Sbox_13_T7}), .c ({new_AGEMA_signal_5270, SubBytesIns_Inst_Sbox_13_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T10_U1 ( .a ({new_AGEMA_signal_5269, SubBytesIns_Inst_Sbox_13_T6}), .b ({new_AGEMA_signal_5108, SubBytesIns_Inst_Sbox_13_T7}), .c ({new_AGEMA_signal_5515, SubBytesIns_Inst_Sbox_13_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T11_U1 ( .a ({ciphertext_s1[110], ciphertext_s0[110]}), .b ({ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_5109, SubBytesIns_Inst_Sbox_13_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T12_U1 ( .a ({ciphertext_s1[109], ciphertext_s0[109]}), .b ({ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_5110, SubBytesIns_Inst_Sbox_13_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T13_U1 ( .a ({new_AGEMA_signal_5105, SubBytesIns_Inst_Sbox_13_T3}), .b ({new_AGEMA_signal_5106, SubBytesIns_Inst_Sbox_13_T4}), .c ({new_AGEMA_signal_5271, SubBytesIns_Inst_Sbox_13_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T14_U1 ( .a ({new_AGEMA_signal_5269, SubBytesIns_Inst_Sbox_13_T6}), .b ({new_AGEMA_signal_5109, SubBytesIns_Inst_Sbox_13_T11}), .c ({new_AGEMA_signal_5516, SubBytesIns_Inst_Sbox_13_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T15_U1 ( .a ({new_AGEMA_signal_5107, SubBytesIns_Inst_Sbox_13_T5}), .b ({new_AGEMA_signal_5109, SubBytesIns_Inst_Sbox_13_T11}), .c ({new_AGEMA_signal_5272, SubBytesIns_Inst_Sbox_13_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T16_U1 ( .a ({new_AGEMA_signal_5107, SubBytesIns_Inst_Sbox_13_T5}), .b ({new_AGEMA_signal_5110, SubBytesIns_Inst_Sbox_13_T12}), .c ({new_AGEMA_signal_5273, SubBytesIns_Inst_Sbox_13_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T17_U1 ( .a ({new_AGEMA_signal_5270, SubBytesIns_Inst_Sbox_13_T9}), .b ({new_AGEMA_signal_5273, SubBytesIns_Inst_Sbox_13_T16}), .c ({new_AGEMA_signal_5517, SubBytesIns_Inst_Sbox_13_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T18_U1 ( .a ({ciphertext_s1[108], ciphertext_s0[108]}), .b ({ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_5111, SubBytesIns_Inst_Sbox_13_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T19_U1 ( .a ({new_AGEMA_signal_5108, SubBytesIns_Inst_Sbox_13_T7}), .b ({new_AGEMA_signal_5111, SubBytesIns_Inst_Sbox_13_T18}), .c ({new_AGEMA_signal_5274, SubBytesIns_Inst_Sbox_13_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T20_U1 ( .a ({new_AGEMA_signal_5103, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_5274, SubBytesIns_Inst_Sbox_13_T19}), .c ({new_AGEMA_signal_5518, SubBytesIns_Inst_Sbox_13_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T21_U1 ( .a ({ciphertext_s1[105], ciphertext_s0[105]}), .b ({ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_5112, SubBytesIns_Inst_Sbox_13_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T22_U1 ( .a ({new_AGEMA_signal_5108, SubBytesIns_Inst_Sbox_13_T7}), .b ({new_AGEMA_signal_5112, SubBytesIns_Inst_Sbox_13_T21}), .c ({new_AGEMA_signal_5275, SubBytesIns_Inst_Sbox_13_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T23_U1 ( .a ({new_AGEMA_signal_5104, SubBytesIns_Inst_Sbox_13_T2}), .b ({new_AGEMA_signal_5275, SubBytesIns_Inst_Sbox_13_T22}), .c ({new_AGEMA_signal_5519, SubBytesIns_Inst_Sbox_13_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T24_U1 ( .a ({new_AGEMA_signal_5104, SubBytesIns_Inst_Sbox_13_T2}), .b ({new_AGEMA_signal_5515, SubBytesIns_Inst_Sbox_13_T10}), .c ({new_AGEMA_signal_5706, SubBytesIns_Inst_Sbox_13_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T25_U1 ( .a ({new_AGEMA_signal_5518, SubBytesIns_Inst_Sbox_13_T20}), .b ({new_AGEMA_signal_5517, SubBytesIns_Inst_Sbox_13_T17}), .c ({new_AGEMA_signal_5707, SubBytesIns_Inst_Sbox_13_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T26_U1 ( .a ({new_AGEMA_signal_5105, SubBytesIns_Inst_Sbox_13_T3}), .b ({new_AGEMA_signal_5273, SubBytesIns_Inst_Sbox_13_T16}), .c ({new_AGEMA_signal_5520, SubBytesIns_Inst_Sbox_13_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T27_U1 ( .a ({new_AGEMA_signal_5103, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_5110, SubBytesIns_Inst_Sbox_13_T12}), .c ({new_AGEMA_signal_5276, SubBytesIns_Inst_Sbox_13_T27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T1_U1 ( .a ({ciphertext_s1[119], ciphertext_s0[119]}), .b ({ciphertext_s1[116], ciphertext_s0[116]}), .c ({new_AGEMA_signal_5113, SubBytesIns_Inst_Sbox_14_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T2_U1 ( .a ({ciphertext_s1[119], ciphertext_s0[119]}), .b ({ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_5114, SubBytesIns_Inst_Sbox_14_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T3_U1 ( .a ({ciphertext_s1[119], ciphertext_s0[119]}), .b ({ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_5115, SubBytesIns_Inst_Sbox_14_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T4_U1 ( .a ({ciphertext_s1[116], ciphertext_s0[116]}), .b ({ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_5116, SubBytesIns_Inst_Sbox_14_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T5_U1 ( .a ({ciphertext_s1[115], ciphertext_s0[115]}), .b ({ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_5117, SubBytesIns_Inst_Sbox_14_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T6_U1 ( .a ({new_AGEMA_signal_5113, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_5117, SubBytesIns_Inst_Sbox_14_T5}), .c ({new_AGEMA_signal_5277, SubBytesIns_Inst_Sbox_14_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T7_U1 ( .a ({ciphertext_s1[118], ciphertext_s0[118]}), .b ({ciphertext_s1[117], ciphertext_s0[117]}), .c ({new_AGEMA_signal_5118, SubBytesIns_Inst_Sbox_14_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T8_U1 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({new_AGEMA_signal_5277, SubBytesIns_Inst_Sbox_14_T6}), .c ({new_AGEMA_signal_5527, SubBytesIns_Inst_Sbox_14_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T9_U1 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({new_AGEMA_signal_5118, SubBytesIns_Inst_Sbox_14_T7}), .c ({new_AGEMA_signal_5278, SubBytesIns_Inst_Sbox_14_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T10_U1 ( .a ({new_AGEMA_signal_5277, SubBytesIns_Inst_Sbox_14_T6}), .b ({new_AGEMA_signal_5118, SubBytesIns_Inst_Sbox_14_T7}), .c ({new_AGEMA_signal_5528, SubBytesIns_Inst_Sbox_14_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T11_U1 ( .a ({ciphertext_s1[118], ciphertext_s0[118]}), .b ({ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_5119, SubBytesIns_Inst_Sbox_14_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T12_U1 ( .a ({ciphertext_s1[117], ciphertext_s0[117]}), .b ({ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_5120, SubBytesIns_Inst_Sbox_14_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T13_U1 ( .a ({new_AGEMA_signal_5115, SubBytesIns_Inst_Sbox_14_T3}), .b ({new_AGEMA_signal_5116, SubBytesIns_Inst_Sbox_14_T4}), .c ({new_AGEMA_signal_5279, SubBytesIns_Inst_Sbox_14_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T14_U1 ( .a ({new_AGEMA_signal_5277, SubBytesIns_Inst_Sbox_14_T6}), .b ({new_AGEMA_signal_5119, SubBytesIns_Inst_Sbox_14_T11}), .c ({new_AGEMA_signal_5529, SubBytesIns_Inst_Sbox_14_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T15_U1 ( .a ({new_AGEMA_signal_5117, SubBytesIns_Inst_Sbox_14_T5}), .b ({new_AGEMA_signal_5119, SubBytesIns_Inst_Sbox_14_T11}), .c ({new_AGEMA_signal_5280, SubBytesIns_Inst_Sbox_14_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T16_U1 ( .a ({new_AGEMA_signal_5117, SubBytesIns_Inst_Sbox_14_T5}), .b ({new_AGEMA_signal_5120, SubBytesIns_Inst_Sbox_14_T12}), .c ({new_AGEMA_signal_5281, SubBytesIns_Inst_Sbox_14_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T17_U1 ( .a ({new_AGEMA_signal_5278, SubBytesIns_Inst_Sbox_14_T9}), .b ({new_AGEMA_signal_5281, SubBytesIns_Inst_Sbox_14_T16}), .c ({new_AGEMA_signal_5530, SubBytesIns_Inst_Sbox_14_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T18_U1 ( .a ({ciphertext_s1[116], ciphertext_s0[116]}), .b ({ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_5121, SubBytesIns_Inst_Sbox_14_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T19_U1 ( .a ({new_AGEMA_signal_5118, SubBytesIns_Inst_Sbox_14_T7}), .b ({new_AGEMA_signal_5121, SubBytesIns_Inst_Sbox_14_T18}), .c ({new_AGEMA_signal_5282, SubBytesIns_Inst_Sbox_14_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T20_U1 ( .a ({new_AGEMA_signal_5113, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_5282, SubBytesIns_Inst_Sbox_14_T19}), .c ({new_AGEMA_signal_5531, SubBytesIns_Inst_Sbox_14_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T21_U1 ( .a ({ciphertext_s1[113], ciphertext_s0[113]}), .b ({ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_5122, SubBytesIns_Inst_Sbox_14_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T22_U1 ( .a ({new_AGEMA_signal_5118, SubBytesIns_Inst_Sbox_14_T7}), .b ({new_AGEMA_signal_5122, SubBytesIns_Inst_Sbox_14_T21}), .c ({new_AGEMA_signal_5283, SubBytesIns_Inst_Sbox_14_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T23_U1 ( .a ({new_AGEMA_signal_5114, SubBytesIns_Inst_Sbox_14_T2}), .b ({new_AGEMA_signal_5283, SubBytesIns_Inst_Sbox_14_T22}), .c ({new_AGEMA_signal_5532, SubBytesIns_Inst_Sbox_14_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T24_U1 ( .a ({new_AGEMA_signal_5114, SubBytesIns_Inst_Sbox_14_T2}), .b ({new_AGEMA_signal_5528, SubBytesIns_Inst_Sbox_14_T10}), .c ({new_AGEMA_signal_5715, SubBytesIns_Inst_Sbox_14_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T25_U1 ( .a ({new_AGEMA_signal_5531, SubBytesIns_Inst_Sbox_14_T20}), .b ({new_AGEMA_signal_5530, SubBytesIns_Inst_Sbox_14_T17}), .c ({new_AGEMA_signal_5716, SubBytesIns_Inst_Sbox_14_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T26_U1 ( .a ({new_AGEMA_signal_5115, SubBytesIns_Inst_Sbox_14_T3}), .b ({new_AGEMA_signal_5281, SubBytesIns_Inst_Sbox_14_T16}), .c ({new_AGEMA_signal_5533, SubBytesIns_Inst_Sbox_14_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T27_U1 ( .a ({new_AGEMA_signal_5113, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_5120, SubBytesIns_Inst_Sbox_14_T12}), .c ({new_AGEMA_signal_5284, SubBytesIns_Inst_Sbox_14_T27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T1_U1 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_5123, SubBytesIns_Inst_Sbox_15_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T2_U1 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_5124, SubBytesIns_Inst_Sbox_15_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T3_U1 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_5125, SubBytesIns_Inst_Sbox_15_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T4_U1 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_5126, SubBytesIns_Inst_Sbox_15_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T5_U1 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_5127, SubBytesIns_Inst_Sbox_15_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T6_U1 ( .a ({new_AGEMA_signal_5123, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_5127, SubBytesIns_Inst_Sbox_15_T5}), .c ({new_AGEMA_signal_5285, SubBytesIns_Inst_Sbox_15_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T7_U1 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_5128, SubBytesIns_Inst_Sbox_15_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T8_U1 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_5285, SubBytesIns_Inst_Sbox_15_T6}), .c ({new_AGEMA_signal_5540, SubBytesIns_Inst_Sbox_15_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T9_U1 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_5128, SubBytesIns_Inst_Sbox_15_T7}), .c ({new_AGEMA_signal_5286, SubBytesIns_Inst_Sbox_15_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T10_U1 ( .a ({new_AGEMA_signal_5285, SubBytesIns_Inst_Sbox_15_T6}), .b ({new_AGEMA_signal_5128, SubBytesIns_Inst_Sbox_15_T7}), .c ({new_AGEMA_signal_5541, SubBytesIns_Inst_Sbox_15_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T11_U1 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_5129, SubBytesIns_Inst_Sbox_15_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T12_U1 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_5130, SubBytesIns_Inst_Sbox_15_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T13_U1 ( .a ({new_AGEMA_signal_5125, SubBytesIns_Inst_Sbox_15_T3}), .b ({new_AGEMA_signal_5126, SubBytesIns_Inst_Sbox_15_T4}), .c ({new_AGEMA_signal_5287, SubBytesIns_Inst_Sbox_15_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T14_U1 ( .a ({new_AGEMA_signal_5285, SubBytesIns_Inst_Sbox_15_T6}), .b ({new_AGEMA_signal_5129, SubBytesIns_Inst_Sbox_15_T11}), .c ({new_AGEMA_signal_5542, SubBytesIns_Inst_Sbox_15_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T15_U1 ( .a ({new_AGEMA_signal_5127, SubBytesIns_Inst_Sbox_15_T5}), .b ({new_AGEMA_signal_5129, SubBytesIns_Inst_Sbox_15_T11}), .c ({new_AGEMA_signal_5288, SubBytesIns_Inst_Sbox_15_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T16_U1 ( .a ({new_AGEMA_signal_5127, SubBytesIns_Inst_Sbox_15_T5}), .b ({new_AGEMA_signal_5130, SubBytesIns_Inst_Sbox_15_T12}), .c ({new_AGEMA_signal_5289, SubBytesIns_Inst_Sbox_15_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T17_U1 ( .a ({new_AGEMA_signal_5286, SubBytesIns_Inst_Sbox_15_T9}), .b ({new_AGEMA_signal_5289, SubBytesIns_Inst_Sbox_15_T16}), .c ({new_AGEMA_signal_5543, SubBytesIns_Inst_Sbox_15_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T18_U1 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_5131, SubBytesIns_Inst_Sbox_15_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T19_U1 ( .a ({new_AGEMA_signal_5128, SubBytesIns_Inst_Sbox_15_T7}), .b ({new_AGEMA_signal_5131, SubBytesIns_Inst_Sbox_15_T18}), .c ({new_AGEMA_signal_5290, SubBytesIns_Inst_Sbox_15_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T20_U1 ( .a ({new_AGEMA_signal_5123, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_5290, SubBytesIns_Inst_Sbox_15_T19}), .c ({new_AGEMA_signal_5544, SubBytesIns_Inst_Sbox_15_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T21_U1 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_5132, SubBytesIns_Inst_Sbox_15_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T22_U1 ( .a ({new_AGEMA_signal_5128, SubBytesIns_Inst_Sbox_15_T7}), .b ({new_AGEMA_signal_5132, SubBytesIns_Inst_Sbox_15_T21}), .c ({new_AGEMA_signal_5291, SubBytesIns_Inst_Sbox_15_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T23_U1 ( .a ({new_AGEMA_signal_5124, SubBytesIns_Inst_Sbox_15_T2}), .b ({new_AGEMA_signal_5291, SubBytesIns_Inst_Sbox_15_T22}), .c ({new_AGEMA_signal_5545, SubBytesIns_Inst_Sbox_15_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T24_U1 ( .a ({new_AGEMA_signal_5124, SubBytesIns_Inst_Sbox_15_T2}), .b ({new_AGEMA_signal_5541, SubBytesIns_Inst_Sbox_15_T10}), .c ({new_AGEMA_signal_5724, SubBytesIns_Inst_Sbox_15_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T25_U1 ( .a ({new_AGEMA_signal_5544, SubBytesIns_Inst_Sbox_15_T20}), .b ({new_AGEMA_signal_5543, SubBytesIns_Inst_Sbox_15_T17}), .c ({new_AGEMA_signal_5725, SubBytesIns_Inst_Sbox_15_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T26_U1 ( .a ({new_AGEMA_signal_5125, SubBytesIns_Inst_Sbox_15_T3}), .b ({new_AGEMA_signal_5289, SubBytesIns_Inst_Sbox_15_T16}), .c ({new_AGEMA_signal_5546, SubBytesIns_Inst_Sbox_15_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T27_U1 ( .a ({new_AGEMA_signal_5123, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_5130, SubBytesIns_Inst_Sbox_15_T12}), .c ({new_AGEMA_signal_5292, SubBytesIns_Inst_Sbox_15_T27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T1_U1 ( .a ({new_AGEMA_signal_4679, RoundKey[23]}), .b ({new_AGEMA_signal_4670, RoundKey[20]}), .c ({new_AGEMA_signal_4933, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T2_U1 ( .a ({new_AGEMA_signal_4679, RoundKey[23]}), .b ({new_AGEMA_signal_4661, RoundKey[18]}), .c ({new_AGEMA_signal_4934, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T3_U1 ( .a ({new_AGEMA_signal_4679, RoundKey[23]}), .b ({new_AGEMA_signal_4658, RoundKey[17]}), .c ({new_AGEMA_signal_4935, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T4_U1 ( .a ({new_AGEMA_signal_4670, RoundKey[20]}), .b ({new_AGEMA_signal_4661, RoundKey[18]}), .c ({new_AGEMA_signal_4936, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T5_U1 ( .a ({new_AGEMA_signal_4664, RoundKey[19]}), .b ({new_AGEMA_signal_4658, RoundKey[17]}), .c ({new_AGEMA_signal_4937, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T6_U1 ( .a ({new_AGEMA_signal_4933, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_4937, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}), .c ({new_AGEMA_signal_5133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T7_U1 ( .a ({new_AGEMA_signal_4676, RoundKey[22]}), .b ({new_AGEMA_signal_4673, RoundKey[21]}), .c ({new_AGEMA_signal_4938, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T8_U1 ( .a ({new_AGEMA_signal_4655, RoundKey[16]}), .b ({new_AGEMA_signal_5133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .c ({new_AGEMA_signal_5293, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T9_U1 ( .a ({new_AGEMA_signal_4655, RoundKey[16]}), .b ({new_AGEMA_signal_4938, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_5134, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T10_U1 ( .a ({new_AGEMA_signal_5133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_4938, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_5294, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T11_U1 ( .a ({new_AGEMA_signal_4676, RoundKey[22]}), .b ({new_AGEMA_signal_4661, RoundKey[18]}), .c ({new_AGEMA_signal_4939, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T12_U1 ( .a ({new_AGEMA_signal_4673, RoundKey[21]}), .b ({new_AGEMA_signal_4661, RoundKey[18]}), .c ({new_AGEMA_signal_4940, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T13_U1 ( .a ({new_AGEMA_signal_4935, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_4936, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}), .c ({new_AGEMA_signal_5135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T14_U1 ( .a ({new_AGEMA_signal_5133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_4939, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_5295, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T15_U1 ( .a ({new_AGEMA_signal_4937, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_4939, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_5136, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T16_U1 ( .a ({new_AGEMA_signal_4937, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_4940, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_5137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T17_U1 ( .a ({new_AGEMA_signal_5134, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}), .b ({new_AGEMA_signal_5137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_5296, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T18_U1 ( .a ({new_AGEMA_signal_4670, RoundKey[20]}), .b ({new_AGEMA_signal_4655, RoundKey[16]}), .c ({new_AGEMA_signal_4941, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T19_U1 ( .a ({new_AGEMA_signal_4938, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_4941, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18}), .c ({new_AGEMA_signal_5138, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T20_U1 ( .a ({new_AGEMA_signal_4933, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5138, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}), .c ({new_AGEMA_signal_5297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T21_U1 ( .a ({new_AGEMA_signal_4658, RoundKey[17]}), .b ({new_AGEMA_signal_4655, RoundKey[16]}), .c ({new_AGEMA_signal_4942, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T22_U1 ( .a ({new_AGEMA_signal_4938, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_4942, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21}), .c ({new_AGEMA_signal_5139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T23_U1 ( .a ({new_AGEMA_signal_4934, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_5139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}), .c ({new_AGEMA_signal_5298, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T24_U1 ( .a ({new_AGEMA_signal_4934, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_5294, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}), .c ({new_AGEMA_signal_5553, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T25_U1 ( .a ({new_AGEMA_signal_5297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_5296, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}), .c ({new_AGEMA_signal_5554, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T26_U1 ( .a ({new_AGEMA_signal_4935, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_5299, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T27_U1 ( .a ({new_AGEMA_signal_4933, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_4940, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_5140, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T1_U1 ( .a ({new_AGEMA_signal_4652, RoundKey[15]}), .b ({new_AGEMA_signal_4643, RoundKey[12]}), .c ({new_AGEMA_signal_4943, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T2_U1 ( .a ({new_AGEMA_signal_4652, RoundKey[15]}), .b ({new_AGEMA_signal_4583, RoundKey[10]}), .c ({new_AGEMA_signal_4944, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T3_U1 ( .a ({new_AGEMA_signal_4652, RoundKey[15]}), .b ({new_AGEMA_signal_4931, RoundKey[9]}), .c ({new_AGEMA_signal_4945, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T4_U1 ( .a ({new_AGEMA_signal_4643, RoundKey[12]}), .b ({new_AGEMA_signal_4583, RoundKey[10]}), .c ({new_AGEMA_signal_4946, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T5_U1 ( .a ({new_AGEMA_signal_4616, RoundKey[11]}), .b ({new_AGEMA_signal_4931, RoundKey[9]}), .c ({new_AGEMA_signal_4947, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T6_U1 ( .a ({new_AGEMA_signal_4943, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_4947, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}), .c ({new_AGEMA_signal_5141, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T7_U1 ( .a ({new_AGEMA_signal_4649, RoundKey[14]}), .b ({new_AGEMA_signal_4646, RoundKey[13]}), .c ({new_AGEMA_signal_4948, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T8_U1 ( .a ({new_AGEMA_signal_4898, RoundKey[8]}), .b ({new_AGEMA_signal_5141, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .c ({new_AGEMA_signal_5306, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T9_U1 ( .a ({new_AGEMA_signal_4898, RoundKey[8]}), .b ({new_AGEMA_signal_4948, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_5142, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T10_U1 ( .a ({new_AGEMA_signal_5141, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_4948, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_5307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T11_U1 ( .a ({new_AGEMA_signal_4649, RoundKey[14]}), .b ({new_AGEMA_signal_4583, RoundKey[10]}), .c ({new_AGEMA_signal_4949, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T12_U1 ( .a ({new_AGEMA_signal_4646, RoundKey[13]}), .b ({new_AGEMA_signal_4583, RoundKey[10]}), .c ({new_AGEMA_signal_4950, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T13_U1 ( .a ({new_AGEMA_signal_4945, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_4946, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}), .c ({new_AGEMA_signal_5143, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T14_U1 ( .a ({new_AGEMA_signal_5141, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_4949, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_5308, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T15_U1 ( .a ({new_AGEMA_signal_4947, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_4949, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_5144, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T16_U1 ( .a ({new_AGEMA_signal_4947, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_4950, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_5145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T17_U1 ( .a ({new_AGEMA_signal_5142, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}), .b ({new_AGEMA_signal_5145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_5309, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T18_U1 ( .a ({new_AGEMA_signal_4643, RoundKey[12]}), .b ({new_AGEMA_signal_4898, RoundKey[8]}), .c ({new_AGEMA_signal_4951, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T19_U1 ( .a ({new_AGEMA_signal_4948, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_4951, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18}), .c ({new_AGEMA_signal_5146, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T20_U1 ( .a ({new_AGEMA_signal_4943, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5146, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}), .c ({new_AGEMA_signal_5310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T21_U1 ( .a ({new_AGEMA_signal_4931, RoundKey[9]}), .b ({new_AGEMA_signal_4898, RoundKey[8]}), .c ({new_AGEMA_signal_4952, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T22_U1 ( .a ({new_AGEMA_signal_4948, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_4952, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21}), .c ({new_AGEMA_signal_5147, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T23_U1 ( .a ({new_AGEMA_signal_4944, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_5147, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}), .c ({new_AGEMA_signal_5311, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T24_U1 ( .a ({new_AGEMA_signal_4944, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_5307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}), .c ({new_AGEMA_signal_5562, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T25_U1 ( .a ({new_AGEMA_signal_5310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_5309, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}), .c ({new_AGEMA_signal_5563, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T26_U1 ( .a ({new_AGEMA_signal_4945, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_5312, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T27_U1 ( .a ({new_AGEMA_signal_4943, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_4950, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_5148, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T1_U1 ( .a ({new_AGEMA_signal_4865, RoundKey[7]}), .b ({new_AGEMA_signal_4766, RoundKey[4]}), .c ({new_AGEMA_signal_4953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T2_U1 ( .a ({new_AGEMA_signal_4865, RoundKey[7]}), .b ({new_AGEMA_signal_4700, RoundKey[2]}), .c ({new_AGEMA_signal_4954, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T3_U1 ( .a ({new_AGEMA_signal_4865, RoundKey[7]}), .b ({new_AGEMA_signal_4667, RoundKey[1]}), .c ({new_AGEMA_signal_4955, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T4_U1 ( .a ({new_AGEMA_signal_4766, RoundKey[4]}), .b ({new_AGEMA_signal_4700, RoundKey[2]}), .c ({new_AGEMA_signal_4956, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T5_U1 ( .a ({new_AGEMA_signal_4733, RoundKey[3]}), .b ({new_AGEMA_signal_4667, RoundKey[1]}), .c ({new_AGEMA_signal_4957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T6_U1 ( .a ({new_AGEMA_signal_4953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_4957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}), .c ({new_AGEMA_signal_5149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T7_U1 ( .a ({new_AGEMA_signal_4832, RoundKey[6]}), .b ({new_AGEMA_signal_4799, RoundKey[5]}), .c ({new_AGEMA_signal_4958, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T8_U1 ( .a ({new_AGEMA_signal_4550, RoundKey[0]}), .b ({new_AGEMA_signal_5149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .c ({new_AGEMA_signal_5319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T9_U1 ( .a ({new_AGEMA_signal_4550, RoundKey[0]}), .b ({new_AGEMA_signal_4958, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_5150, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T10_U1 ( .a ({new_AGEMA_signal_5149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_4958, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_5320, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T11_U1 ( .a ({new_AGEMA_signal_4832, RoundKey[6]}), .b ({new_AGEMA_signal_4700, RoundKey[2]}), .c ({new_AGEMA_signal_4959, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T12_U1 ( .a ({new_AGEMA_signal_4799, RoundKey[5]}), .b ({new_AGEMA_signal_4700, RoundKey[2]}), .c ({new_AGEMA_signal_4960, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T13_U1 ( .a ({new_AGEMA_signal_4955, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_4956, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}), .c ({new_AGEMA_signal_5151, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T14_U1 ( .a ({new_AGEMA_signal_5149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_4959, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_5321, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T15_U1 ( .a ({new_AGEMA_signal_4957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_4959, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_5152, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T16_U1 ( .a ({new_AGEMA_signal_4957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_4960, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_5153, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T17_U1 ( .a ({new_AGEMA_signal_5150, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}), .b ({new_AGEMA_signal_5153, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_5322, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T18_U1 ( .a ({new_AGEMA_signal_4766, RoundKey[4]}), .b ({new_AGEMA_signal_4550, RoundKey[0]}), .c ({new_AGEMA_signal_4961, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T19_U1 ( .a ({new_AGEMA_signal_4958, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_4961, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18}), .c ({new_AGEMA_signal_5154, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T20_U1 ( .a ({new_AGEMA_signal_4953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5154, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}), .c ({new_AGEMA_signal_5323, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T21_U1 ( .a ({new_AGEMA_signal_4667, RoundKey[1]}), .b ({new_AGEMA_signal_4550, RoundKey[0]}), .c ({new_AGEMA_signal_4962, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T22_U1 ( .a ({new_AGEMA_signal_4958, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_4962, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21}), .c ({new_AGEMA_signal_5155, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T23_U1 ( .a ({new_AGEMA_signal_4954, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_5155, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}), .c ({new_AGEMA_signal_5324, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T24_U1 ( .a ({new_AGEMA_signal_4954, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_5320, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}), .c ({new_AGEMA_signal_5571, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T25_U1 ( .a ({new_AGEMA_signal_5323, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_5322, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}), .c ({new_AGEMA_signal_5572, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T26_U1 ( .a ({new_AGEMA_signal_4955, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5153, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_5325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T27_U1 ( .a ({new_AGEMA_signal_4953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_4960, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_5156, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T1_U1 ( .a ({new_AGEMA_signal_4706, RoundKey[31]}), .b ({new_AGEMA_signal_4694, RoundKey[28]}), .c ({new_AGEMA_signal_4963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T2_U1 ( .a ({new_AGEMA_signal_4706, RoundKey[31]}), .b ({new_AGEMA_signal_4688, RoundKey[26]}), .c ({new_AGEMA_signal_4964, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T3_U1 ( .a ({new_AGEMA_signal_4706, RoundKey[31]}), .b ({new_AGEMA_signal_4685, RoundKey[25]}), .c ({new_AGEMA_signal_4965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T4_U1 ( .a ({new_AGEMA_signal_4694, RoundKey[28]}), .b ({new_AGEMA_signal_4688, RoundKey[26]}), .c ({new_AGEMA_signal_4966, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T5_U1 ( .a ({new_AGEMA_signal_4691, RoundKey[27]}), .b ({new_AGEMA_signal_4685, RoundKey[25]}), .c ({new_AGEMA_signal_4967, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T6_U1 ( .a ({new_AGEMA_signal_4963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_4967, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}), .c ({new_AGEMA_signal_5157, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T7_U1 ( .a ({new_AGEMA_signal_4703, RoundKey[30]}), .b ({new_AGEMA_signal_4697, RoundKey[29]}), .c ({new_AGEMA_signal_4968, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T8_U1 ( .a ({new_AGEMA_signal_4682, RoundKey[24]}), .b ({new_AGEMA_signal_5157, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .c ({new_AGEMA_signal_5332, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T9_U1 ( .a ({new_AGEMA_signal_4682, RoundKey[24]}), .b ({new_AGEMA_signal_4968, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_5158, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T10_U1 ( .a ({new_AGEMA_signal_5157, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_4968, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_5333, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T11_U1 ( .a ({new_AGEMA_signal_4703, RoundKey[30]}), .b ({new_AGEMA_signal_4688, RoundKey[26]}), .c ({new_AGEMA_signal_4969, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T12_U1 ( .a ({new_AGEMA_signal_4697, RoundKey[29]}), .b ({new_AGEMA_signal_4688, RoundKey[26]}), .c ({new_AGEMA_signal_4970, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T13_U1 ( .a ({new_AGEMA_signal_4965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_4966, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}), .c ({new_AGEMA_signal_5159, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T14_U1 ( .a ({new_AGEMA_signal_5157, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_4969, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_5334, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T15_U1 ( .a ({new_AGEMA_signal_4967, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_4969, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_5160, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T16_U1 ( .a ({new_AGEMA_signal_4967, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_4970, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_5161, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T17_U1 ( .a ({new_AGEMA_signal_5158, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}), .b ({new_AGEMA_signal_5161, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_5335, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T18_U1 ( .a ({new_AGEMA_signal_4694, RoundKey[28]}), .b ({new_AGEMA_signal_4682, RoundKey[24]}), .c ({new_AGEMA_signal_4971, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T19_U1 ( .a ({new_AGEMA_signal_4968, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_4971, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18}), .c ({new_AGEMA_signal_5162, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T20_U1 ( .a ({new_AGEMA_signal_4963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5162, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}), .c ({new_AGEMA_signal_5336, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T21_U1 ( .a ({new_AGEMA_signal_4685, RoundKey[25]}), .b ({new_AGEMA_signal_4682, RoundKey[24]}), .c ({new_AGEMA_signal_4972, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T22_U1 ( .a ({new_AGEMA_signal_4968, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_4972, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21}), .c ({new_AGEMA_signal_5163, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T23_U1 ( .a ({new_AGEMA_signal_4964, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_5163, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}), .c ({new_AGEMA_signal_5337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T24_U1 ( .a ({new_AGEMA_signal_4964, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_5333, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}), .c ({new_AGEMA_signal_5580, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T25_U1 ( .a ({new_AGEMA_signal_5336, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_5335, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}), .c ({new_AGEMA_signal_5581, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T26_U1 ( .a ({new_AGEMA_signal_4965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5161, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_5338, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T27_U1 ( .a ({new_AGEMA_signal_4963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_4970, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_5164, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27}) ) ;
    INV_X1 RoundCounterIns_U14 ( .A (RoundCounterIns_n13), .ZN (RoundCounterIns_n1) ) ;
    MUX2_X1 RoundCounterIns_U13 ( .S (RoundCounterIns_n5), .A (RoundCounterIns_n12), .B (RoundCounterIns_n11), .Z (RoundCounterIns_n13) ) ;
    NOR2_X1 RoundCounterIns_U12 ( .A1 (reset), .A2 (RoundCounterIns_n10), .ZN (RoundCounterIns_N8) ) ;
    XNOR2_X1 RoundCounterIns_U11 ( .A (RoundCounter[0]), .B (RoundCounter[1]), .ZN (RoundCounterIns_n10) ) ;
    MUX2_X1 RoundCounterIns_U10 ( .S (RoundCounter[3]), .A (RoundCounterIns_n9), .B (RoundCounterIns_n8), .Z (RoundCounterIns_N10) ) ;
    NAND2_X1 RoundCounterIns_U9 ( .A1 (RoundCounterIns_n12), .A2 (RoundCounterIns_n7), .ZN (RoundCounterIns_n8) ) ;
    NAND2_X1 RoundCounterIns_U8 ( .A1 (RoundCounterIns_n5), .A2 (RoundCounterIns_n2), .ZN (RoundCounterIns_n7) ) ;
    NOR2_X1 RoundCounterIns_U7 ( .A1 (RoundCounterIns_n4), .A2 (RoundCounterIns_N7), .ZN (RoundCounterIns_n12) ) ;
    NOR2_X1 RoundCounterIns_U6 ( .A1 (RoundCounter[1]), .A2 (reset), .ZN (RoundCounterIns_n4) ) ;
    NOR2_X1 RoundCounterIns_U5 ( .A1 (RoundCounterIns_n5), .A2 (RoundCounterIns_n11), .ZN (RoundCounterIns_n9) ) ;
    NAND2_X1 RoundCounterIns_U4 ( .A1 (RoundCounter[1]), .A2 (RoundCounterIns_n3), .ZN (RoundCounterIns_n11) ) ;
    NOR2_X1 RoundCounterIns_U3 ( .A1 (reset), .A2 (RoundCounterIns_n6), .ZN (RoundCounterIns_n3) ) ;
    NOR2_X1 RoundCounterIns_U2 ( .A1 (reset), .A2 (RoundCounter[0]), .ZN (RoundCounterIns_N7) ) ;
    INV_X1 RoundCounterIns_U1 ( .A (reset), .ZN (RoundCounterIns_n2) ) ;
    INV_X1 RoundCounterIns_count_reg_0__U1 ( .A (RoundCounter[0]), .ZN (RoundCounterIns_n6) ) ;
    INV_X1 RoundCounterIns_count_reg_2__U1 ( .A (RoundCounter[2]), .ZN (RoundCounterIns_n5) ) ;
    ClockGatingController #(9) ClockGatingInst ( .clk (clk), .rst (reset), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M1_U1 ( .a ({new_AGEMA_signal_5167, SubBytesIns_Inst_Sbox_0_T13}), .b ({new_AGEMA_signal_5165, SubBytesIns_Inst_Sbox_0_T6}), .clk (clk), .r (Fresh[0]), .c ({new_AGEMA_signal_5352, SubBytesIns_Inst_Sbox_0_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M2_U1 ( .a ({new_AGEMA_signal_5350, SubBytesIns_Inst_Sbox_0_T23}), .b ({new_AGEMA_signal_5345, SubBytesIns_Inst_Sbox_0_T8}), .clk (clk), .r (Fresh[1]), .c ({new_AGEMA_signal_5591, SubBytesIns_Inst_Sbox_0_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M3_U1 ( .a ({new_AGEMA_signal_5347, SubBytesIns_Inst_Sbox_0_T14}), .b ({new_AGEMA_signal_5352, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_5592, SubBytesIns_Inst_Sbox_0_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M4_U1 ( .a ({new_AGEMA_signal_5170, SubBytesIns_Inst_Sbox_0_T19}), .b ({ciphertext_s1[0], ciphertext_s0[0]}), .clk (clk), .r (Fresh[2]), .c ({new_AGEMA_signal_5353, SubBytesIns_Inst_Sbox_0_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M5_U1 ( .a ({new_AGEMA_signal_5353, SubBytesIns_Inst_Sbox_0_M4}), .b ({new_AGEMA_signal_5352, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_5593, SubBytesIns_Inst_Sbox_0_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M6_U1 ( .a ({new_AGEMA_signal_4975, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5169, SubBytesIns_Inst_Sbox_0_T16}), .clk (clk), .r (Fresh[3]), .c ({new_AGEMA_signal_5354, SubBytesIns_Inst_Sbox_0_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M7_U1 ( .a ({new_AGEMA_signal_5171, SubBytesIns_Inst_Sbox_0_T22}), .b ({new_AGEMA_signal_5166, SubBytesIns_Inst_Sbox_0_T9}), .clk (clk), .r (Fresh[4]), .c ({new_AGEMA_signal_5355, SubBytesIns_Inst_Sbox_0_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M8_U1 ( .a ({new_AGEMA_signal_5351, SubBytesIns_Inst_Sbox_0_T26}), .b ({new_AGEMA_signal_5354, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_5594, SubBytesIns_Inst_Sbox_0_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M9_U1 ( .a ({new_AGEMA_signal_5349, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_5348, SubBytesIns_Inst_Sbox_0_T17}), .clk (clk), .r (Fresh[5]), .c ({new_AGEMA_signal_5595, SubBytesIns_Inst_Sbox_0_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M10_U1 ( .a ({new_AGEMA_signal_5595, SubBytesIns_Inst_Sbox_0_M9}), .b ({new_AGEMA_signal_5354, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_5753, SubBytesIns_Inst_Sbox_0_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M11_U1 ( .a ({new_AGEMA_signal_4973, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5168, SubBytesIns_Inst_Sbox_0_T15}), .clk (clk), .r (Fresh[6]), .c ({new_AGEMA_signal_5356, SubBytesIns_Inst_Sbox_0_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M12_U1 ( .a ({new_AGEMA_signal_4976, SubBytesIns_Inst_Sbox_0_T4}), .b ({new_AGEMA_signal_5172, SubBytesIns_Inst_Sbox_0_T27}), .clk (clk), .r (Fresh[7]), .c ({new_AGEMA_signal_5357, SubBytesIns_Inst_Sbox_0_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M13_U1 ( .a ({new_AGEMA_signal_5357, SubBytesIns_Inst_Sbox_0_M12}), .b ({new_AGEMA_signal_5356, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_5596, SubBytesIns_Inst_Sbox_0_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M14_U1 ( .a ({new_AGEMA_signal_4974, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_5346, SubBytesIns_Inst_Sbox_0_T10}), .clk (clk), .r (Fresh[8]), .c ({new_AGEMA_signal_5597, SubBytesIns_Inst_Sbox_0_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M15_U1 ( .a ({new_AGEMA_signal_5597, SubBytesIns_Inst_Sbox_0_M14}), .b ({new_AGEMA_signal_5356, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_5754, SubBytesIns_Inst_Sbox_0_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M16_U1 ( .a ({new_AGEMA_signal_5592, SubBytesIns_Inst_Sbox_0_M3}), .b ({new_AGEMA_signal_5591, SubBytesIns_Inst_Sbox_0_M2}), .c ({new_AGEMA_signal_5755, SubBytesIns_Inst_Sbox_0_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M17_U1 ( .a ({new_AGEMA_signal_5593, SubBytesIns_Inst_Sbox_0_M5}), .b ({new_AGEMA_signal_5589, SubBytesIns_Inst_Sbox_0_T24}), .c ({new_AGEMA_signal_5756, SubBytesIns_Inst_Sbox_0_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M18_U1 ( .a ({new_AGEMA_signal_5594, SubBytesIns_Inst_Sbox_0_M8}), .b ({new_AGEMA_signal_5355, SubBytesIns_Inst_Sbox_0_M7}), .c ({new_AGEMA_signal_5757, SubBytesIns_Inst_Sbox_0_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M19_U1 ( .a ({new_AGEMA_signal_5753, SubBytesIns_Inst_Sbox_0_M10}), .b ({new_AGEMA_signal_5754, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_5849, SubBytesIns_Inst_Sbox_0_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M20_U1 ( .a ({new_AGEMA_signal_5755, SubBytesIns_Inst_Sbox_0_M16}), .b ({new_AGEMA_signal_5596, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_5850, SubBytesIns_Inst_Sbox_0_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M21_U1 ( .a ({new_AGEMA_signal_5756, SubBytesIns_Inst_Sbox_0_M17}), .b ({new_AGEMA_signal_5754, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_0_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M22_U1 ( .a ({new_AGEMA_signal_5757, SubBytesIns_Inst_Sbox_0_M18}), .b ({new_AGEMA_signal_5596, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_5852, SubBytesIns_Inst_Sbox_0_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M23_U1 ( .a ({new_AGEMA_signal_5849, SubBytesIns_Inst_Sbox_0_M19}), .b ({new_AGEMA_signal_5590, SubBytesIns_Inst_Sbox_0_T25}), .c ({new_AGEMA_signal_5929, SubBytesIns_Inst_Sbox_0_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M24_U1 ( .a ({new_AGEMA_signal_5852, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_5929, SubBytesIns_Inst_Sbox_0_M23}), .c ({new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_0_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M27_U1 ( .a ({new_AGEMA_signal_5850, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_0_M21}), .c ({new_AGEMA_signal_5931, SubBytesIns_Inst_Sbox_0_M27}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M1_U1 ( .a ({new_AGEMA_signal_5175, SubBytesIns_Inst_Sbox_1_T13}), .b ({new_AGEMA_signal_5173, SubBytesIns_Inst_Sbox_1_T6}), .clk (clk), .r (Fresh[9]), .c ({new_AGEMA_signal_5365, SubBytesIns_Inst_Sbox_1_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M2_U1 ( .a ({new_AGEMA_signal_5363, SubBytesIns_Inst_Sbox_1_T23}), .b ({new_AGEMA_signal_5358, SubBytesIns_Inst_Sbox_1_T8}), .clk (clk), .r (Fresh[10]), .c ({new_AGEMA_signal_5600, SubBytesIns_Inst_Sbox_1_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M3_U1 ( .a ({new_AGEMA_signal_5360, SubBytesIns_Inst_Sbox_1_T14}), .b ({new_AGEMA_signal_5365, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_5601, SubBytesIns_Inst_Sbox_1_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M4_U1 ( .a ({new_AGEMA_signal_5178, SubBytesIns_Inst_Sbox_1_T19}), .b ({ciphertext_s1[8], ciphertext_s0[8]}), .clk (clk), .r (Fresh[11]), .c ({new_AGEMA_signal_5366, SubBytesIns_Inst_Sbox_1_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M5_U1 ( .a ({new_AGEMA_signal_5366, SubBytesIns_Inst_Sbox_1_M4}), .b ({new_AGEMA_signal_5365, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_5602, SubBytesIns_Inst_Sbox_1_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M6_U1 ( .a ({new_AGEMA_signal_4985, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5177, SubBytesIns_Inst_Sbox_1_T16}), .clk (clk), .r (Fresh[12]), .c ({new_AGEMA_signal_5367, SubBytesIns_Inst_Sbox_1_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M7_U1 ( .a ({new_AGEMA_signal_5179, SubBytesIns_Inst_Sbox_1_T22}), .b ({new_AGEMA_signal_5174, SubBytesIns_Inst_Sbox_1_T9}), .clk (clk), .r (Fresh[13]), .c ({new_AGEMA_signal_5368, SubBytesIns_Inst_Sbox_1_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M8_U1 ( .a ({new_AGEMA_signal_5364, SubBytesIns_Inst_Sbox_1_T26}), .b ({new_AGEMA_signal_5367, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_5603, SubBytesIns_Inst_Sbox_1_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M9_U1 ( .a ({new_AGEMA_signal_5362, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_5361, SubBytesIns_Inst_Sbox_1_T17}), .clk (clk), .r (Fresh[14]), .c ({new_AGEMA_signal_5604, SubBytesIns_Inst_Sbox_1_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M10_U1 ( .a ({new_AGEMA_signal_5604, SubBytesIns_Inst_Sbox_1_M9}), .b ({new_AGEMA_signal_5367, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_5758, SubBytesIns_Inst_Sbox_1_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M11_U1 ( .a ({new_AGEMA_signal_4983, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5176, SubBytesIns_Inst_Sbox_1_T15}), .clk (clk), .r (Fresh[15]), .c ({new_AGEMA_signal_5369, SubBytesIns_Inst_Sbox_1_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M12_U1 ( .a ({new_AGEMA_signal_4986, SubBytesIns_Inst_Sbox_1_T4}), .b ({new_AGEMA_signal_5180, SubBytesIns_Inst_Sbox_1_T27}), .clk (clk), .r (Fresh[16]), .c ({new_AGEMA_signal_5370, SubBytesIns_Inst_Sbox_1_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M13_U1 ( .a ({new_AGEMA_signal_5370, SubBytesIns_Inst_Sbox_1_M12}), .b ({new_AGEMA_signal_5369, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_5605, SubBytesIns_Inst_Sbox_1_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M14_U1 ( .a ({new_AGEMA_signal_4984, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_5359, SubBytesIns_Inst_Sbox_1_T10}), .clk (clk), .r (Fresh[17]), .c ({new_AGEMA_signal_5606, SubBytesIns_Inst_Sbox_1_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M15_U1 ( .a ({new_AGEMA_signal_5606, SubBytesIns_Inst_Sbox_1_M14}), .b ({new_AGEMA_signal_5369, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_5759, SubBytesIns_Inst_Sbox_1_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M16_U1 ( .a ({new_AGEMA_signal_5601, SubBytesIns_Inst_Sbox_1_M3}), .b ({new_AGEMA_signal_5600, SubBytesIns_Inst_Sbox_1_M2}), .c ({new_AGEMA_signal_5760, SubBytesIns_Inst_Sbox_1_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M17_U1 ( .a ({new_AGEMA_signal_5602, SubBytesIns_Inst_Sbox_1_M5}), .b ({new_AGEMA_signal_5598, SubBytesIns_Inst_Sbox_1_T24}), .c ({new_AGEMA_signal_5761, SubBytesIns_Inst_Sbox_1_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M18_U1 ( .a ({new_AGEMA_signal_5603, SubBytesIns_Inst_Sbox_1_M8}), .b ({new_AGEMA_signal_5368, SubBytesIns_Inst_Sbox_1_M7}), .c ({new_AGEMA_signal_5762, SubBytesIns_Inst_Sbox_1_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M19_U1 ( .a ({new_AGEMA_signal_5758, SubBytesIns_Inst_Sbox_1_M10}), .b ({new_AGEMA_signal_5759, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_5853, SubBytesIns_Inst_Sbox_1_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M20_U1 ( .a ({new_AGEMA_signal_5760, SubBytesIns_Inst_Sbox_1_M16}), .b ({new_AGEMA_signal_5605, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_5854, SubBytesIns_Inst_Sbox_1_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M21_U1 ( .a ({new_AGEMA_signal_5761, SubBytesIns_Inst_Sbox_1_M17}), .b ({new_AGEMA_signal_5759, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_5855, SubBytesIns_Inst_Sbox_1_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M22_U1 ( .a ({new_AGEMA_signal_5762, SubBytesIns_Inst_Sbox_1_M18}), .b ({new_AGEMA_signal_5605, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_5856, SubBytesIns_Inst_Sbox_1_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M23_U1 ( .a ({new_AGEMA_signal_5853, SubBytesIns_Inst_Sbox_1_M19}), .b ({new_AGEMA_signal_5599, SubBytesIns_Inst_Sbox_1_T25}), .c ({new_AGEMA_signal_5933, SubBytesIns_Inst_Sbox_1_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M24_U1 ( .a ({new_AGEMA_signal_5856, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_5933, SubBytesIns_Inst_Sbox_1_M23}), .c ({new_AGEMA_signal_6018, SubBytesIns_Inst_Sbox_1_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M27_U1 ( .a ({new_AGEMA_signal_5854, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_5855, SubBytesIns_Inst_Sbox_1_M21}), .c ({new_AGEMA_signal_5935, SubBytesIns_Inst_Sbox_1_M27}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M1_U1 ( .a ({new_AGEMA_signal_5183, SubBytesIns_Inst_Sbox_2_T13}), .b ({new_AGEMA_signal_5181, SubBytesIns_Inst_Sbox_2_T6}), .clk (clk), .r (Fresh[18]), .c ({new_AGEMA_signal_5378, SubBytesIns_Inst_Sbox_2_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M2_U1 ( .a ({new_AGEMA_signal_5376, SubBytesIns_Inst_Sbox_2_T23}), .b ({new_AGEMA_signal_5371, SubBytesIns_Inst_Sbox_2_T8}), .clk (clk), .r (Fresh[19]), .c ({new_AGEMA_signal_5609, SubBytesIns_Inst_Sbox_2_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M3_U1 ( .a ({new_AGEMA_signal_5373, SubBytesIns_Inst_Sbox_2_T14}), .b ({new_AGEMA_signal_5378, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_5610, SubBytesIns_Inst_Sbox_2_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M4_U1 ( .a ({new_AGEMA_signal_5186, SubBytesIns_Inst_Sbox_2_T19}), .b ({ciphertext_s1[16], ciphertext_s0[16]}), .clk (clk), .r (Fresh[20]), .c ({new_AGEMA_signal_5379, SubBytesIns_Inst_Sbox_2_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M5_U1 ( .a ({new_AGEMA_signal_5379, SubBytesIns_Inst_Sbox_2_M4}), .b ({new_AGEMA_signal_5378, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_5611, SubBytesIns_Inst_Sbox_2_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M6_U1 ( .a ({new_AGEMA_signal_4995, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5185, SubBytesIns_Inst_Sbox_2_T16}), .clk (clk), .r (Fresh[21]), .c ({new_AGEMA_signal_5380, SubBytesIns_Inst_Sbox_2_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M7_U1 ( .a ({new_AGEMA_signal_5187, SubBytesIns_Inst_Sbox_2_T22}), .b ({new_AGEMA_signal_5182, SubBytesIns_Inst_Sbox_2_T9}), .clk (clk), .r (Fresh[22]), .c ({new_AGEMA_signal_5381, SubBytesIns_Inst_Sbox_2_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M8_U1 ( .a ({new_AGEMA_signal_5377, SubBytesIns_Inst_Sbox_2_T26}), .b ({new_AGEMA_signal_5380, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_5612, SubBytesIns_Inst_Sbox_2_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M9_U1 ( .a ({new_AGEMA_signal_5375, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_5374, SubBytesIns_Inst_Sbox_2_T17}), .clk (clk), .r (Fresh[23]), .c ({new_AGEMA_signal_5613, SubBytesIns_Inst_Sbox_2_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M10_U1 ( .a ({new_AGEMA_signal_5613, SubBytesIns_Inst_Sbox_2_M9}), .b ({new_AGEMA_signal_5380, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_5763, SubBytesIns_Inst_Sbox_2_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M11_U1 ( .a ({new_AGEMA_signal_4993, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5184, SubBytesIns_Inst_Sbox_2_T15}), .clk (clk), .r (Fresh[24]), .c ({new_AGEMA_signal_5382, SubBytesIns_Inst_Sbox_2_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M12_U1 ( .a ({new_AGEMA_signal_4996, SubBytesIns_Inst_Sbox_2_T4}), .b ({new_AGEMA_signal_5188, SubBytesIns_Inst_Sbox_2_T27}), .clk (clk), .r (Fresh[25]), .c ({new_AGEMA_signal_5383, SubBytesIns_Inst_Sbox_2_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M13_U1 ( .a ({new_AGEMA_signal_5383, SubBytesIns_Inst_Sbox_2_M12}), .b ({new_AGEMA_signal_5382, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_5614, SubBytesIns_Inst_Sbox_2_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M14_U1 ( .a ({new_AGEMA_signal_4994, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_5372, SubBytesIns_Inst_Sbox_2_T10}), .clk (clk), .r (Fresh[26]), .c ({new_AGEMA_signal_5615, SubBytesIns_Inst_Sbox_2_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M15_U1 ( .a ({new_AGEMA_signal_5615, SubBytesIns_Inst_Sbox_2_M14}), .b ({new_AGEMA_signal_5382, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_5764, SubBytesIns_Inst_Sbox_2_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M16_U1 ( .a ({new_AGEMA_signal_5610, SubBytesIns_Inst_Sbox_2_M3}), .b ({new_AGEMA_signal_5609, SubBytesIns_Inst_Sbox_2_M2}), .c ({new_AGEMA_signal_5765, SubBytesIns_Inst_Sbox_2_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M17_U1 ( .a ({new_AGEMA_signal_5611, SubBytesIns_Inst_Sbox_2_M5}), .b ({new_AGEMA_signal_5607, SubBytesIns_Inst_Sbox_2_T24}), .c ({new_AGEMA_signal_5766, SubBytesIns_Inst_Sbox_2_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M18_U1 ( .a ({new_AGEMA_signal_5612, SubBytesIns_Inst_Sbox_2_M8}), .b ({new_AGEMA_signal_5381, SubBytesIns_Inst_Sbox_2_M7}), .c ({new_AGEMA_signal_5767, SubBytesIns_Inst_Sbox_2_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M19_U1 ( .a ({new_AGEMA_signal_5763, SubBytesIns_Inst_Sbox_2_M10}), .b ({new_AGEMA_signal_5764, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_2_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M20_U1 ( .a ({new_AGEMA_signal_5765, SubBytesIns_Inst_Sbox_2_M16}), .b ({new_AGEMA_signal_5614, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_5858, SubBytesIns_Inst_Sbox_2_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M21_U1 ( .a ({new_AGEMA_signal_5766, SubBytesIns_Inst_Sbox_2_M17}), .b ({new_AGEMA_signal_5764, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_5859, SubBytesIns_Inst_Sbox_2_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M22_U1 ( .a ({new_AGEMA_signal_5767, SubBytesIns_Inst_Sbox_2_M18}), .b ({new_AGEMA_signal_5614, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_5860, SubBytesIns_Inst_Sbox_2_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M23_U1 ( .a ({new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_2_M19}), .b ({new_AGEMA_signal_5608, SubBytesIns_Inst_Sbox_2_T25}), .c ({new_AGEMA_signal_5937, SubBytesIns_Inst_Sbox_2_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M24_U1 ( .a ({new_AGEMA_signal_5860, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_5937, SubBytesIns_Inst_Sbox_2_M23}), .c ({new_AGEMA_signal_6023, SubBytesIns_Inst_Sbox_2_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M27_U1 ( .a ({new_AGEMA_signal_5858, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_5859, SubBytesIns_Inst_Sbox_2_M21}), .c ({new_AGEMA_signal_5939, SubBytesIns_Inst_Sbox_2_M27}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M1_U1 ( .a ({new_AGEMA_signal_5191, SubBytesIns_Inst_Sbox_3_T13}), .b ({new_AGEMA_signal_5189, SubBytesIns_Inst_Sbox_3_T6}), .clk (clk), .r (Fresh[27]), .c ({new_AGEMA_signal_5391, SubBytesIns_Inst_Sbox_3_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M2_U1 ( .a ({new_AGEMA_signal_5389, SubBytesIns_Inst_Sbox_3_T23}), .b ({new_AGEMA_signal_5384, SubBytesIns_Inst_Sbox_3_T8}), .clk (clk), .r (Fresh[28]), .c ({new_AGEMA_signal_5618, SubBytesIns_Inst_Sbox_3_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M3_U1 ( .a ({new_AGEMA_signal_5386, SubBytesIns_Inst_Sbox_3_T14}), .b ({new_AGEMA_signal_5391, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_5619, SubBytesIns_Inst_Sbox_3_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M4_U1 ( .a ({new_AGEMA_signal_5194, SubBytesIns_Inst_Sbox_3_T19}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .clk (clk), .r (Fresh[29]), .c ({new_AGEMA_signal_5392, SubBytesIns_Inst_Sbox_3_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M5_U1 ( .a ({new_AGEMA_signal_5392, SubBytesIns_Inst_Sbox_3_M4}), .b ({new_AGEMA_signal_5391, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_5620, SubBytesIns_Inst_Sbox_3_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M6_U1 ( .a ({new_AGEMA_signal_5005, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5193, SubBytesIns_Inst_Sbox_3_T16}), .clk (clk), .r (Fresh[30]), .c ({new_AGEMA_signal_5393, SubBytesIns_Inst_Sbox_3_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M7_U1 ( .a ({new_AGEMA_signal_5195, SubBytesIns_Inst_Sbox_3_T22}), .b ({new_AGEMA_signal_5190, SubBytesIns_Inst_Sbox_3_T9}), .clk (clk), .r (Fresh[31]), .c ({new_AGEMA_signal_5394, SubBytesIns_Inst_Sbox_3_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M8_U1 ( .a ({new_AGEMA_signal_5390, SubBytesIns_Inst_Sbox_3_T26}), .b ({new_AGEMA_signal_5393, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_5621, SubBytesIns_Inst_Sbox_3_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M9_U1 ( .a ({new_AGEMA_signal_5388, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_5387, SubBytesIns_Inst_Sbox_3_T17}), .clk (clk), .r (Fresh[32]), .c ({new_AGEMA_signal_5622, SubBytesIns_Inst_Sbox_3_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M10_U1 ( .a ({new_AGEMA_signal_5622, SubBytesIns_Inst_Sbox_3_M9}), .b ({new_AGEMA_signal_5393, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_5768, SubBytesIns_Inst_Sbox_3_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M11_U1 ( .a ({new_AGEMA_signal_5003, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5192, SubBytesIns_Inst_Sbox_3_T15}), .clk (clk), .r (Fresh[33]), .c ({new_AGEMA_signal_5395, SubBytesIns_Inst_Sbox_3_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M12_U1 ( .a ({new_AGEMA_signal_5006, SubBytesIns_Inst_Sbox_3_T4}), .b ({new_AGEMA_signal_5196, SubBytesIns_Inst_Sbox_3_T27}), .clk (clk), .r (Fresh[34]), .c ({new_AGEMA_signal_5396, SubBytesIns_Inst_Sbox_3_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M13_U1 ( .a ({new_AGEMA_signal_5396, SubBytesIns_Inst_Sbox_3_M12}), .b ({new_AGEMA_signal_5395, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_5623, SubBytesIns_Inst_Sbox_3_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M14_U1 ( .a ({new_AGEMA_signal_5004, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_5385, SubBytesIns_Inst_Sbox_3_T10}), .clk (clk), .r (Fresh[35]), .c ({new_AGEMA_signal_5624, SubBytesIns_Inst_Sbox_3_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M15_U1 ( .a ({new_AGEMA_signal_5624, SubBytesIns_Inst_Sbox_3_M14}), .b ({new_AGEMA_signal_5395, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_5769, SubBytesIns_Inst_Sbox_3_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M16_U1 ( .a ({new_AGEMA_signal_5619, SubBytesIns_Inst_Sbox_3_M3}), .b ({new_AGEMA_signal_5618, SubBytesIns_Inst_Sbox_3_M2}), .c ({new_AGEMA_signal_5770, SubBytesIns_Inst_Sbox_3_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M17_U1 ( .a ({new_AGEMA_signal_5620, SubBytesIns_Inst_Sbox_3_M5}), .b ({new_AGEMA_signal_5616, SubBytesIns_Inst_Sbox_3_T24}), .c ({new_AGEMA_signal_5771, SubBytesIns_Inst_Sbox_3_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M18_U1 ( .a ({new_AGEMA_signal_5621, SubBytesIns_Inst_Sbox_3_M8}), .b ({new_AGEMA_signal_5394, SubBytesIns_Inst_Sbox_3_M7}), .c ({new_AGEMA_signal_5772, SubBytesIns_Inst_Sbox_3_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M19_U1 ( .a ({new_AGEMA_signal_5768, SubBytesIns_Inst_Sbox_3_M10}), .b ({new_AGEMA_signal_5769, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_5861, SubBytesIns_Inst_Sbox_3_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M20_U1 ( .a ({new_AGEMA_signal_5770, SubBytesIns_Inst_Sbox_3_M16}), .b ({new_AGEMA_signal_5623, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_5862, SubBytesIns_Inst_Sbox_3_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M21_U1 ( .a ({new_AGEMA_signal_5771, SubBytesIns_Inst_Sbox_3_M17}), .b ({new_AGEMA_signal_5769, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_3_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M22_U1 ( .a ({new_AGEMA_signal_5772, SubBytesIns_Inst_Sbox_3_M18}), .b ({new_AGEMA_signal_5623, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_5864, SubBytesIns_Inst_Sbox_3_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M23_U1 ( .a ({new_AGEMA_signal_5861, SubBytesIns_Inst_Sbox_3_M19}), .b ({new_AGEMA_signal_5617, SubBytesIns_Inst_Sbox_3_T25}), .c ({new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_3_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M24_U1 ( .a ({new_AGEMA_signal_5864, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_3_M23}), .c ({new_AGEMA_signal_6028, SubBytesIns_Inst_Sbox_3_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M27_U1 ( .a ({new_AGEMA_signal_5862, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_3_M21}), .c ({new_AGEMA_signal_5943, SubBytesIns_Inst_Sbox_3_M27}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M1_U1 ( .a ({new_AGEMA_signal_5199, SubBytesIns_Inst_Sbox_4_T13}), .b ({new_AGEMA_signal_5197, SubBytesIns_Inst_Sbox_4_T6}), .clk (clk), .r (Fresh[36]), .c ({new_AGEMA_signal_5404, SubBytesIns_Inst_Sbox_4_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M2_U1 ( .a ({new_AGEMA_signal_5402, SubBytesIns_Inst_Sbox_4_T23}), .b ({new_AGEMA_signal_5397, SubBytesIns_Inst_Sbox_4_T8}), .clk (clk), .r (Fresh[37]), .c ({new_AGEMA_signal_5627, SubBytesIns_Inst_Sbox_4_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M3_U1 ( .a ({new_AGEMA_signal_5399, SubBytesIns_Inst_Sbox_4_T14}), .b ({new_AGEMA_signal_5404, SubBytesIns_Inst_Sbox_4_M1}), .c ({new_AGEMA_signal_5628, SubBytesIns_Inst_Sbox_4_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M4_U1 ( .a ({new_AGEMA_signal_5202, SubBytesIns_Inst_Sbox_4_T19}), .b ({ciphertext_s1[32], ciphertext_s0[32]}), .clk (clk), .r (Fresh[38]), .c ({new_AGEMA_signal_5405, SubBytesIns_Inst_Sbox_4_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M5_U1 ( .a ({new_AGEMA_signal_5405, SubBytesIns_Inst_Sbox_4_M4}), .b ({new_AGEMA_signal_5404, SubBytesIns_Inst_Sbox_4_M1}), .c ({new_AGEMA_signal_5629, SubBytesIns_Inst_Sbox_4_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M6_U1 ( .a ({new_AGEMA_signal_5015, SubBytesIns_Inst_Sbox_4_T3}), .b ({new_AGEMA_signal_5201, SubBytesIns_Inst_Sbox_4_T16}), .clk (clk), .r (Fresh[39]), .c ({new_AGEMA_signal_5406, SubBytesIns_Inst_Sbox_4_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M7_U1 ( .a ({new_AGEMA_signal_5203, SubBytesIns_Inst_Sbox_4_T22}), .b ({new_AGEMA_signal_5198, SubBytesIns_Inst_Sbox_4_T9}), .clk (clk), .r (Fresh[40]), .c ({new_AGEMA_signal_5407, SubBytesIns_Inst_Sbox_4_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M8_U1 ( .a ({new_AGEMA_signal_5403, SubBytesIns_Inst_Sbox_4_T26}), .b ({new_AGEMA_signal_5406, SubBytesIns_Inst_Sbox_4_M6}), .c ({new_AGEMA_signal_5630, SubBytesIns_Inst_Sbox_4_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M9_U1 ( .a ({new_AGEMA_signal_5401, SubBytesIns_Inst_Sbox_4_T20}), .b ({new_AGEMA_signal_5400, SubBytesIns_Inst_Sbox_4_T17}), .clk (clk), .r (Fresh[41]), .c ({new_AGEMA_signal_5631, SubBytesIns_Inst_Sbox_4_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M10_U1 ( .a ({new_AGEMA_signal_5631, SubBytesIns_Inst_Sbox_4_M9}), .b ({new_AGEMA_signal_5406, SubBytesIns_Inst_Sbox_4_M6}), .c ({new_AGEMA_signal_5773, SubBytesIns_Inst_Sbox_4_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M11_U1 ( .a ({new_AGEMA_signal_5013, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5200, SubBytesIns_Inst_Sbox_4_T15}), .clk (clk), .r (Fresh[42]), .c ({new_AGEMA_signal_5408, SubBytesIns_Inst_Sbox_4_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M12_U1 ( .a ({new_AGEMA_signal_5016, SubBytesIns_Inst_Sbox_4_T4}), .b ({new_AGEMA_signal_5204, SubBytesIns_Inst_Sbox_4_T27}), .clk (clk), .r (Fresh[43]), .c ({new_AGEMA_signal_5409, SubBytesIns_Inst_Sbox_4_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M13_U1 ( .a ({new_AGEMA_signal_5409, SubBytesIns_Inst_Sbox_4_M12}), .b ({new_AGEMA_signal_5408, SubBytesIns_Inst_Sbox_4_M11}), .c ({new_AGEMA_signal_5632, SubBytesIns_Inst_Sbox_4_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M14_U1 ( .a ({new_AGEMA_signal_5014, SubBytesIns_Inst_Sbox_4_T2}), .b ({new_AGEMA_signal_5398, SubBytesIns_Inst_Sbox_4_T10}), .clk (clk), .r (Fresh[44]), .c ({new_AGEMA_signal_5633, SubBytesIns_Inst_Sbox_4_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M15_U1 ( .a ({new_AGEMA_signal_5633, SubBytesIns_Inst_Sbox_4_M14}), .b ({new_AGEMA_signal_5408, SubBytesIns_Inst_Sbox_4_M11}), .c ({new_AGEMA_signal_5774, SubBytesIns_Inst_Sbox_4_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M16_U1 ( .a ({new_AGEMA_signal_5628, SubBytesIns_Inst_Sbox_4_M3}), .b ({new_AGEMA_signal_5627, SubBytesIns_Inst_Sbox_4_M2}), .c ({new_AGEMA_signal_5775, SubBytesIns_Inst_Sbox_4_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M17_U1 ( .a ({new_AGEMA_signal_5629, SubBytesIns_Inst_Sbox_4_M5}), .b ({new_AGEMA_signal_5625, SubBytesIns_Inst_Sbox_4_T24}), .c ({new_AGEMA_signal_5776, SubBytesIns_Inst_Sbox_4_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M18_U1 ( .a ({new_AGEMA_signal_5630, SubBytesIns_Inst_Sbox_4_M8}), .b ({new_AGEMA_signal_5407, SubBytesIns_Inst_Sbox_4_M7}), .c ({new_AGEMA_signal_5777, SubBytesIns_Inst_Sbox_4_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M19_U1 ( .a ({new_AGEMA_signal_5773, SubBytesIns_Inst_Sbox_4_M10}), .b ({new_AGEMA_signal_5774, SubBytesIns_Inst_Sbox_4_M15}), .c ({new_AGEMA_signal_5865, SubBytesIns_Inst_Sbox_4_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M20_U1 ( .a ({new_AGEMA_signal_5775, SubBytesIns_Inst_Sbox_4_M16}), .b ({new_AGEMA_signal_5632, SubBytesIns_Inst_Sbox_4_M13}), .c ({new_AGEMA_signal_5866, SubBytesIns_Inst_Sbox_4_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M21_U1 ( .a ({new_AGEMA_signal_5776, SubBytesIns_Inst_Sbox_4_M17}), .b ({new_AGEMA_signal_5774, SubBytesIns_Inst_Sbox_4_M15}), .c ({new_AGEMA_signal_5867, SubBytesIns_Inst_Sbox_4_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M22_U1 ( .a ({new_AGEMA_signal_5777, SubBytesIns_Inst_Sbox_4_M18}), .b ({new_AGEMA_signal_5632, SubBytesIns_Inst_Sbox_4_M13}), .c ({new_AGEMA_signal_5868, SubBytesIns_Inst_Sbox_4_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M23_U1 ( .a ({new_AGEMA_signal_5865, SubBytesIns_Inst_Sbox_4_M19}), .b ({new_AGEMA_signal_5626, SubBytesIns_Inst_Sbox_4_T25}), .c ({new_AGEMA_signal_5945, SubBytesIns_Inst_Sbox_4_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M24_U1 ( .a ({new_AGEMA_signal_5868, SubBytesIns_Inst_Sbox_4_M22}), .b ({new_AGEMA_signal_5945, SubBytesIns_Inst_Sbox_4_M23}), .c ({new_AGEMA_signal_6033, SubBytesIns_Inst_Sbox_4_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M27_U1 ( .a ({new_AGEMA_signal_5866, SubBytesIns_Inst_Sbox_4_M20}), .b ({new_AGEMA_signal_5867, SubBytesIns_Inst_Sbox_4_M21}), .c ({new_AGEMA_signal_5947, SubBytesIns_Inst_Sbox_4_M27}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M1_U1 ( .a ({new_AGEMA_signal_5207, SubBytesIns_Inst_Sbox_5_T13}), .b ({new_AGEMA_signal_5205, SubBytesIns_Inst_Sbox_5_T6}), .clk (clk), .r (Fresh[45]), .c ({new_AGEMA_signal_5417, SubBytesIns_Inst_Sbox_5_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M2_U1 ( .a ({new_AGEMA_signal_5415, SubBytesIns_Inst_Sbox_5_T23}), .b ({new_AGEMA_signal_5410, SubBytesIns_Inst_Sbox_5_T8}), .clk (clk), .r (Fresh[46]), .c ({new_AGEMA_signal_5636, SubBytesIns_Inst_Sbox_5_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M3_U1 ( .a ({new_AGEMA_signal_5412, SubBytesIns_Inst_Sbox_5_T14}), .b ({new_AGEMA_signal_5417, SubBytesIns_Inst_Sbox_5_M1}), .c ({new_AGEMA_signal_5637, SubBytesIns_Inst_Sbox_5_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M4_U1 ( .a ({new_AGEMA_signal_5210, SubBytesIns_Inst_Sbox_5_T19}), .b ({ciphertext_s1[40], ciphertext_s0[40]}), .clk (clk), .r (Fresh[47]), .c ({new_AGEMA_signal_5418, SubBytesIns_Inst_Sbox_5_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M5_U1 ( .a ({new_AGEMA_signal_5418, SubBytesIns_Inst_Sbox_5_M4}), .b ({new_AGEMA_signal_5417, SubBytesIns_Inst_Sbox_5_M1}), .c ({new_AGEMA_signal_5638, SubBytesIns_Inst_Sbox_5_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M6_U1 ( .a ({new_AGEMA_signal_5025, SubBytesIns_Inst_Sbox_5_T3}), .b ({new_AGEMA_signal_5209, SubBytesIns_Inst_Sbox_5_T16}), .clk (clk), .r (Fresh[48]), .c ({new_AGEMA_signal_5419, SubBytesIns_Inst_Sbox_5_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M7_U1 ( .a ({new_AGEMA_signal_5211, SubBytesIns_Inst_Sbox_5_T22}), .b ({new_AGEMA_signal_5206, SubBytesIns_Inst_Sbox_5_T9}), .clk (clk), .r (Fresh[49]), .c ({new_AGEMA_signal_5420, SubBytesIns_Inst_Sbox_5_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M8_U1 ( .a ({new_AGEMA_signal_5416, SubBytesIns_Inst_Sbox_5_T26}), .b ({new_AGEMA_signal_5419, SubBytesIns_Inst_Sbox_5_M6}), .c ({new_AGEMA_signal_5639, SubBytesIns_Inst_Sbox_5_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M9_U1 ( .a ({new_AGEMA_signal_5414, SubBytesIns_Inst_Sbox_5_T20}), .b ({new_AGEMA_signal_5413, SubBytesIns_Inst_Sbox_5_T17}), .clk (clk), .r (Fresh[50]), .c ({new_AGEMA_signal_5640, SubBytesIns_Inst_Sbox_5_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M10_U1 ( .a ({new_AGEMA_signal_5640, SubBytesIns_Inst_Sbox_5_M9}), .b ({new_AGEMA_signal_5419, SubBytesIns_Inst_Sbox_5_M6}), .c ({new_AGEMA_signal_5778, SubBytesIns_Inst_Sbox_5_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M11_U1 ( .a ({new_AGEMA_signal_5023, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5208, SubBytesIns_Inst_Sbox_5_T15}), .clk (clk), .r (Fresh[51]), .c ({new_AGEMA_signal_5421, SubBytesIns_Inst_Sbox_5_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M12_U1 ( .a ({new_AGEMA_signal_5026, SubBytesIns_Inst_Sbox_5_T4}), .b ({new_AGEMA_signal_5212, SubBytesIns_Inst_Sbox_5_T27}), .clk (clk), .r (Fresh[52]), .c ({new_AGEMA_signal_5422, SubBytesIns_Inst_Sbox_5_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M13_U1 ( .a ({new_AGEMA_signal_5422, SubBytesIns_Inst_Sbox_5_M12}), .b ({new_AGEMA_signal_5421, SubBytesIns_Inst_Sbox_5_M11}), .c ({new_AGEMA_signal_5641, SubBytesIns_Inst_Sbox_5_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M14_U1 ( .a ({new_AGEMA_signal_5024, SubBytesIns_Inst_Sbox_5_T2}), .b ({new_AGEMA_signal_5411, SubBytesIns_Inst_Sbox_5_T10}), .clk (clk), .r (Fresh[53]), .c ({new_AGEMA_signal_5642, SubBytesIns_Inst_Sbox_5_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M15_U1 ( .a ({new_AGEMA_signal_5642, SubBytesIns_Inst_Sbox_5_M14}), .b ({new_AGEMA_signal_5421, SubBytesIns_Inst_Sbox_5_M11}), .c ({new_AGEMA_signal_5779, SubBytesIns_Inst_Sbox_5_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M16_U1 ( .a ({new_AGEMA_signal_5637, SubBytesIns_Inst_Sbox_5_M3}), .b ({new_AGEMA_signal_5636, SubBytesIns_Inst_Sbox_5_M2}), .c ({new_AGEMA_signal_5780, SubBytesIns_Inst_Sbox_5_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M17_U1 ( .a ({new_AGEMA_signal_5638, SubBytesIns_Inst_Sbox_5_M5}), .b ({new_AGEMA_signal_5634, SubBytesIns_Inst_Sbox_5_T24}), .c ({new_AGEMA_signal_5781, SubBytesIns_Inst_Sbox_5_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M18_U1 ( .a ({new_AGEMA_signal_5639, SubBytesIns_Inst_Sbox_5_M8}), .b ({new_AGEMA_signal_5420, SubBytesIns_Inst_Sbox_5_M7}), .c ({new_AGEMA_signal_5782, SubBytesIns_Inst_Sbox_5_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M19_U1 ( .a ({new_AGEMA_signal_5778, SubBytesIns_Inst_Sbox_5_M10}), .b ({new_AGEMA_signal_5779, SubBytesIns_Inst_Sbox_5_M15}), .c ({new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_5_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M20_U1 ( .a ({new_AGEMA_signal_5780, SubBytesIns_Inst_Sbox_5_M16}), .b ({new_AGEMA_signal_5641, SubBytesIns_Inst_Sbox_5_M13}), .c ({new_AGEMA_signal_5870, SubBytesIns_Inst_Sbox_5_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M21_U1 ( .a ({new_AGEMA_signal_5781, SubBytesIns_Inst_Sbox_5_M17}), .b ({new_AGEMA_signal_5779, SubBytesIns_Inst_Sbox_5_M15}), .c ({new_AGEMA_signal_5871, SubBytesIns_Inst_Sbox_5_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M22_U1 ( .a ({new_AGEMA_signal_5782, SubBytesIns_Inst_Sbox_5_M18}), .b ({new_AGEMA_signal_5641, SubBytesIns_Inst_Sbox_5_M13}), .c ({new_AGEMA_signal_5872, SubBytesIns_Inst_Sbox_5_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M23_U1 ( .a ({new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_5_M19}), .b ({new_AGEMA_signal_5635, SubBytesIns_Inst_Sbox_5_T25}), .c ({new_AGEMA_signal_5949, SubBytesIns_Inst_Sbox_5_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M24_U1 ( .a ({new_AGEMA_signal_5872, SubBytesIns_Inst_Sbox_5_M22}), .b ({new_AGEMA_signal_5949, SubBytesIns_Inst_Sbox_5_M23}), .c ({new_AGEMA_signal_6038, SubBytesIns_Inst_Sbox_5_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M27_U1 ( .a ({new_AGEMA_signal_5870, SubBytesIns_Inst_Sbox_5_M20}), .b ({new_AGEMA_signal_5871, SubBytesIns_Inst_Sbox_5_M21}), .c ({new_AGEMA_signal_5951, SubBytesIns_Inst_Sbox_5_M27}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M1_U1 ( .a ({new_AGEMA_signal_5215, SubBytesIns_Inst_Sbox_6_T13}), .b ({new_AGEMA_signal_5213, SubBytesIns_Inst_Sbox_6_T6}), .clk (clk), .r (Fresh[54]), .c ({new_AGEMA_signal_5430, SubBytesIns_Inst_Sbox_6_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M2_U1 ( .a ({new_AGEMA_signal_5428, SubBytesIns_Inst_Sbox_6_T23}), .b ({new_AGEMA_signal_5423, SubBytesIns_Inst_Sbox_6_T8}), .clk (clk), .r (Fresh[55]), .c ({new_AGEMA_signal_5645, SubBytesIns_Inst_Sbox_6_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M3_U1 ( .a ({new_AGEMA_signal_5425, SubBytesIns_Inst_Sbox_6_T14}), .b ({new_AGEMA_signal_5430, SubBytesIns_Inst_Sbox_6_M1}), .c ({new_AGEMA_signal_5646, SubBytesIns_Inst_Sbox_6_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M4_U1 ( .a ({new_AGEMA_signal_5218, SubBytesIns_Inst_Sbox_6_T19}), .b ({ciphertext_s1[48], ciphertext_s0[48]}), .clk (clk), .r (Fresh[56]), .c ({new_AGEMA_signal_5431, SubBytesIns_Inst_Sbox_6_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M5_U1 ( .a ({new_AGEMA_signal_5431, SubBytesIns_Inst_Sbox_6_M4}), .b ({new_AGEMA_signal_5430, SubBytesIns_Inst_Sbox_6_M1}), .c ({new_AGEMA_signal_5647, SubBytesIns_Inst_Sbox_6_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M6_U1 ( .a ({new_AGEMA_signal_5035, SubBytesIns_Inst_Sbox_6_T3}), .b ({new_AGEMA_signal_5217, SubBytesIns_Inst_Sbox_6_T16}), .clk (clk), .r (Fresh[57]), .c ({new_AGEMA_signal_5432, SubBytesIns_Inst_Sbox_6_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M7_U1 ( .a ({new_AGEMA_signal_5219, SubBytesIns_Inst_Sbox_6_T22}), .b ({new_AGEMA_signal_5214, SubBytesIns_Inst_Sbox_6_T9}), .clk (clk), .r (Fresh[58]), .c ({new_AGEMA_signal_5433, SubBytesIns_Inst_Sbox_6_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M8_U1 ( .a ({new_AGEMA_signal_5429, SubBytesIns_Inst_Sbox_6_T26}), .b ({new_AGEMA_signal_5432, SubBytesIns_Inst_Sbox_6_M6}), .c ({new_AGEMA_signal_5648, SubBytesIns_Inst_Sbox_6_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M9_U1 ( .a ({new_AGEMA_signal_5427, SubBytesIns_Inst_Sbox_6_T20}), .b ({new_AGEMA_signal_5426, SubBytesIns_Inst_Sbox_6_T17}), .clk (clk), .r (Fresh[59]), .c ({new_AGEMA_signal_5649, SubBytesIns_Inst_Sbox_6_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M10_U1 ( .a ({new_AGEMA_signal_5649, SubBytesIns_Inst_Sbox_6_M9}), .b ({new_AGEMA_signal_5432, SubBytesIns_Inst_Sbox_6_M6}), .c ({new_AGEMA_signal_5783, SubBytesIns_Inst_Sbox_6_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M11_U1 ( .a ({new_AGEMA_signal_5033, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_5216, SubBytesIns_Inst_Sbox_6_T15}), .clk (clk), .r (Fresh[60]), .c ({new_AGEMA_signal_5434, SubBytesIns_Inst_Sbox_6_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M12_U1 ( .a ({new_AGEMA_signal_5036, SubBytesIns_Inst_Sbox_6_T4}), .b ({new_AGEMA_signal_5220, SubBytesIns_Inst_Sbox_6_T27}), .clk (clk), .r (Fresh[61]), .c ({new_AGEMA_signal_5435, SubBytesIns_Inst_Sbox_6_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M13_U1 ( .a ({new_AGEMA_signal_5435, SubBytesIns_Inst_Sbox_6_M12}), .b ({new_AGEMA_signal_5434, SubBytesIns_Inst_Sbox_6_M11}), .c ({new_AGEMA_signal_5650, SubBytesIns_Inst_Sbox_6_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M14_U1 ( .a ({new_AGEMA_signal_5034, SubBytesIns_Inst_Sbox_6_T2}), .b ({new_AGEMA_signal_5424, SubBytesIns_Inst_Sbox_6_T10}), .clk (clk), .r (Fresh[62]), .c ({new_AGEMA_signal_5651, SubBytesIns_Inst_Sbox_6_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M15_U1 ( .a ({new_AGEMA_signal_5651, SubBytesIns_Inst_Sbox_6_M14}), .b ({new_AGEMA_signal_5434, SubBytesIns_Inst_Sbox_6_M11}), .c ({new_AGEMA_signal_5784, SubBytesIns_Inst_Sbox_6_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M16_U1 ( .a ({new_AGEMA_signal_5646, SubBytesIns_Inst_Sbox_6_M3}), .b ({new_AGEMA_signal_5645, SubBytesIns_Inst_Sbox_6_M2}), .c ({new_AGEMA_signal_5785, SubBytesIns_Inst_Sbox_6_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M17_U1 ( .a ({new_AGEMA_signal_5647, SubBytesIns_Inst_Sbox_6_M5}), .b ({new_AGEMA_signal_5643, SubBytesIns_Inst_Sbox_6_T24}), .c ({new_AGEMA_signal_5786, SubBytesIns_Inst_Sbox_6_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M18_U1 ( .a ({new_AGEMA_signal_5648, SubBytesIns_Inst_Sbox_6_M8}), .b ({new_AGEMA_signal_5433, SubBytesIns_Inst_Sbox_6_M7}), .c ({new_AGEMA_signal_5787, SubBytesIns_Inst_Sbox_6_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M19_U1 ( .a ({new_AGEMA_signal_5783, SubBytesIns_Inst_Sbox_6_M10}), .b ({new_AGEMA_signal_5784, SubBytesIns_Inst_Sbox_6_M15}), .c ({new_AGEMA_signal_5873, SubBytesIns_Inst_Sbox_6_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M20_U1 ( .a ({new_AGEMA_signal_5785, SubBytesIns_Inst_Sbox_6_M16}), .b ({new_AGEMA_signal_5650, SubBytesIns_Inst_Sbox_6_M13}), .c ({new_AGEMA_signal_5874, SubBytesIns_Inst_Sbox_6_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M21_U1 ( .a ({new_AGEMA_signal_5786, SubBytesIns_Inst_Sbox_6_M17}), .b ({new_AGEMA_signal_5784, SubBytesIns_Inst_Sbox_6_M15}), .c ({new_AGEMA_signal_5875, SubBytesIns_Inst_Sbox_6_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M22_U1 ( .a ({new_AGEMA_signal_5787, SubBytesIns_Inst_Sbox_6_M18}), .b ({new_AGEMA_signal_5650, SubBytesIns_Inst_Sbox_6_M13}), .c ({new_AGEMA_signal_5876, SubBytesIns_Inst_Sbox_6_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M23_U1 ( .a ({new_AGEMA_signal_5873, SubBytesIns_Inst_Sbox_6_M19}), .b ({new_AGEMA_signal_5644, SubBytesIns_Inst_Sbox_6_T25}), .c ({new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_6_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M24_U1 ( .a ({new_AGEMA_signal_5876, SubBytesIns_Inst_Sbox_6_M22}), .b ({new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_6_M23}), .c ({new_AGEMA_signal_6043, SubBytesIns_Inst_Sbox_6_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M27_U1 ( .a ({new_AGEMA_signal_5874, SubBytesIns_Inst_Sbox_6_M20}), .b ({new_AGEMA_signal_5875, SubBytesIns_Inst_Sbox_6_M21}), .c ({new_AGEMA_signal_5955, SubBytesIns_Inst_Sbox_6_M27}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M1_U1 ( .a ({new_AGEMA_signal_5223, SubBytesIns_Inst_Sbox_7_T13}), .b ({new_AGEMA_signal_5221, SubBytesIns_Inst_Sbox_7_T6}), .clk (clk), .r (Fresh[63]), .c ({new_AGEMA_signal_5443, SubBytesIns_Inst_Sbox_7_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M2_U1 ( .a ({new_AGEMA_signal_5441, SubBytesIns_Inst_Sbox_7_T23}), .b ({new_AGEMA_signal_5436, SubBytesIns_Inst_Sbox_7_T8}), .clk (clk), .r (Fresh[64]), .c ({new_AGEMA_signal_5654, SubBytesIns_Inst_Sbox_7_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M3_U1 ( .a ({new_AGEMA_signal_5438, SubBytesIns_Inst_Sbox_7_T14}), .b ({new_AGEMA_signal_5443, SubBytesIns_Inst_Sbox_7_M1}), .c ({new_AGEMA_signal_5655, SubBytesIns_Inst_Sbox_7_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M4_U1 ( .a ({new_AGEMA_signal_5226, SubBytesIns_Inst_Sbox_7_T19}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .clk (clk), .r (Fresh[65]), .c ({new_AGEMA_signal_5444, SubBytesIns_Inst_Sbox_7_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M5_U1 ( .a ({new_AGEMA_signal_5444, SubBytesIns_Inst_Sbox_7_M4}), .b ({new_AGEMA_signal_5443, SubBytesIns_Inst_Sbox_7_M1}), .c ({new_AGEMA_signal_5656, SubBytesIns_Inst_Sbox_7_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M6_U1 ( .a ({new_AGEMA_signal_5045, SubBytesIns_Inst_Sbox_7_T3}), .b ({new_AGEMA_signal_5225, SubBytesIns_Inst_Sbox_7_T16}), .clk (clk), .r (Fresh[66]), .c ({new_AGEMA_signal_5445, SubBytesIns_Inst_Sbox_7_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M7_U1 ( .a ({new_AGEMA_signal_5227, SubBytesIns_Inst_Sbox_7_T22}), .b ({new_AGEMA_signal_5222, SubBytesIns_Inst_Sbox_7_T9}), .clk (clk), .r (Fresh[67]), .c ({new_AGEMA_signal_5446, SubBytesIns_Inst_Sbox_7_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M8_U1 ( .a ({new_AGEMA_signal_5442, SubBytesIns_Inst_Sbox_7_T26}), .b ({new_AGEMA_signal_5445, SubBytesIns_Inst_Sbox_7_M6}), .c ({new_AGEMA_signal_5657, SubBytesIns_Inst_Sbox_7_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M9_U1 ( .a ({new_AGEMA_signal_5440, SubBytesIns_Inst_Sbox_7_T20}), .b ({new_AGEMA_signal_5439, SubBytesIns_Inst_Sbox_7_T17}), .clk (clk), .r (Fresh[68]), .c ({new_AGEMA_signal_5658, SubBytesIns_Inst_Sbox_7_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M10_U1 ( .a ({new_AGEMA_signal_5658, SubBytesIns_Inst_Sbox_7_M9}), .b ({new_AGEMA_signal_5445, SubBytesIns_Inst_Sbox_7_M6}), .c ({new_AGEMA_signal_5788, SubBytesIns_Inst_Sbox_7_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M11_U1 ( .a ({new_AGEMA_signal_5043, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_5224, SubBytesIns_Inst_Sbox_7_T15}), .clk (clk), .r (Fresh[69]), .c ({new_AGEMA_signal_5447, SubBytesIns_Inst_Sbox_7_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M12_U1 ( .a ({new_AGEMA_signal_5046, SubBytesIns_Inst_Sbox_7_T4}), .b ({new_AGEMA_signal_5228, SubBytesIns_Inst_Sbox_7_T27}), .clk (clk), .r (Fresh[70]), .c ({new_AGEMA_signal_5448, SubBytesIns_Inst_Sbox_7_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M13_U1 ( .a ({new_AGEMA_signal_5448, SubBytesIns_Inst_Sbox_7_M12}), .b ({new_AGEMA_signal_5447, SubBytesIns_Inst_Sbox_7_M11}), .c ({new_AGEMA_signal_5659, SubBytesIns_Inst_Sbox_7_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M14_U1 ( .a ({new_AGEMA_signal_5044, SubBytesIns_Inst_Sbox_7_T2}), .b ({new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_7_T10}), .clk (clk), .r (Fresh[71]), .c ({new_AGEMA_signal_5660, SubBytesIns_Inst_Sbox_7_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M15_U1 ( .a ({new_AGEMA_signal_5660, SubBytesIns_Inst_Sbox_7_M14}), .b ({new_AGEMA_signal_5447, SubBytesIns_Inst_Sbox_7_M11}), .c ({new_AGEMA_signal_5789, SubBytesIns_Inst_Sbox_7_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M16_U1 ( .a ({new_AGEMA_signal_5655, SubBytesIns_Inst_Sbox_7_M3}), .b ({new_AGEMA_signal_5654, SubBytesIns_Inst_Sbox_7_M2}), .c ({new_AGEMA_signal_5790, SubBytesIns_Inst_Sbox_7_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M17_U1 ( .a ({new_AGEMA_signal_5656, SubBytesIns_Inst_Sbox_7_M5}), .b ({new_AGEMA_signal_5652, SubBytesIns_Inst_Sbox_7_T24}), .c ({new_AGEMA_signal_5791, SubBytesIns_Inst_Sbox_7_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M18_U1 ( .a ({new_AGEMA_signal_5657, SubBytesIns_Inst_Sbox_7_M8}), .b ({new_AGEMA_signal_5446, SubBytesIns_Inst_Sbox_7_M7}), .c ({new_AGEMA_signal_5792, SubBytesIns_Inst_Sbox_7_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M19_U1 ( .a ({new_AGEMA_signal_5788, SubBytesIns_Inst_Sbox_7_M10}), .b ({new_AGEMA_signal_5789, SubBytesIns_Inst_Sbox_7_M15}), .c ({new_AGEMA_signal_5877, SubBytesIns_Inst_Sbox_7_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M20_U1 ( .a ({new_AGEMA_signal_5790, SubBytesIns_Inst_Sbox_7_M16}), .b ({new_AGEMA_signal_5659, SubBytesIns_Inst_Sbox_7_M13}), .c ({new_AGEMA_signal_5878, SubBytesIns_Inst_Sbox_7_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M21_U1 ( .a ({new_AGEMA_signal_5791, SubBytesIns_Inst_Sbox_7_M17}), .b ({new_AGEMA_signal_5789, SubBytesIns_Inst_Sbox_7_M15}), .c ({new_AGEMA_signal_5879, SubBytesIns_Inst_Sbox_7_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M22_U1 ( .a ({new_AGEMA_signal_5792, SubBytesIns_Inst_Sbox_7_M18}), .b ({new_AGEMA_signal_5659, SubBytesIns_Inst_Sbox_7_M13}), .c ({new_AGEMA_signal_5880, SubBytesIns_Inst_Sbox_7_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M23_U1 ( .a ({new_AGEMA_signal_5877, SubBytesIns_Inst_Sbox_7_M19}), .b ({new_AGEMA_signal_5653, SubBytesIns_Inst_Sbox_7_T25}), .c ({new_AGEMA_signal_5957, SubBytesIns_Inst_Sbox_7_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M24_U1 ( .a ({new_AGEMA_signal_5880, SubBytesIns_Inst_Sbox_7_M22}), .b ({new_AGEMA_signal_5957, SubBytesIns_Inst_Sbox_7_M23}), .c ({new_AGEMA_signal_6048, SubBytesIns_Inst_Sbox_7_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M27_U1 ( .a ({new_AGEMA_signal_5878, SubBytesIns_Inst_Sbox_7_M20}), .b ({new_AGEMA_signal_5879, SubBytesIns_Inst_Sbox_7_M21}), .c ({new_AGEMA_signal_5959, SubBytesIns_Inst_Sbox_7_M27}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M1_U1 ( .a ({new_AGEMA_signal_5231, SubBytesIns_Inst_Sbox_8_T13}), .b ({new_AGEMA_signal_5229, SubBytesIns_Inst_Sbox_8_T6}), .clk (clk), .r (Fresh[72]), .c ({new_AGEMA_signal_5456, SubBytesIns_Inst_Sbox_8_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M2_U1 ( .a ({new_AGEMA_signal_5454, SubBytesIns_Inst_Sbox_8_T23}), .b ({new_AGEMA_signal_5449, SubBytesIns_Inst_Sbox_8_T8}), .clk (clk), .r (Fresh[73]), .c ({new_AGEMA_signal_5663, SubBytesIns_Inst_Sbox_8_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M3_U1 ( .a ({new_AGEMA_signal_5451, SubBytesIns_Inst_Sbox_8_T14}), .b ({new_AGEMA_signal_5456, SubBytesIns_Inst_Sbox_8_M1}), .c ({new_AGEMA_signal_5664, SubBytesIns_Inst_Sbox_8_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M4_U1 ( .a ({new_AGEMA_signal_5234, SubBytesIns_Inst_Sbox_8_T19}), .b ({ciphertext_s1[64], ciphertext_s0[64]}), .clk (clk), .r (Fresh[74]), .c ({new_AGEMA_signal_5457, SubBytesIns_Inst_Sbox_8_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M5_U1 ( .a ({new_AGEMA_signal_5457, SubBytesIns_Inst_Sbox_8_M4}), .b ({new_AGEMA_signal_5456, SubBytesIns_Inst_Sbox_8_M1}), .c ({new_AGEMA_signal_5665, SubBytesIns_Inst_Sbox_8_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M6_U1 ( .a ({new_AGEMA_signal_5055, SubBytesIns_Inst_Sbox_8_T3}), .b ({new_AGEMA_signal_5233, SubBytesIns_Inst_Sbox_8_T16}), .clk (clk), .r (Fresh[75]), .c ({new_AGEMA_signal_5458, SubBytesIns_Inst_Sbox_8_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M7_U1 ( .a ({new_AGEMA_signal_5235, SubBytesIns_Inst_Sbox_8_T22}), .b ({new_AGEMA_signal_5230, SubBytesIns_Inst_Sbox_8_T9}), .clk (clk), .r (Fresh[76]), .c ({new_AGEMA_signal_5459, SubBytesIns_Inst_Sbox_8_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M8_U1 ( .a ({new_AGEMA_signal_5455, SubBytesIns_Inst_Sbox_8_T26}), .b ({new_AGEMA_signal_5458, SubBytesIns_Inst_Sbox_8_M6}), .c ({new_AGEMA_signal_5666, SubBytesIns_Inst_Sbox_8_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M9_U1 ( .a ({new_AGEMA_signal_5453, SubBytesIns_Inst_Sbox_8_T20}), .b ({new_AGEMA_signal_5452, SubBytesIns_Inst_Sbox_8_T17}), .clk (clk), .r (Fresh[77]), .c ({new_AGEMA_signal_5667, SubBytesIns_Inst_Sbox_8_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M10_U1 ( .a ({new_AGEMA_signal_5667, SubBytesIns_Inst_Sbox_8_M9}), .b ({new_AGEMA_signal_5458, SubBytesIns_Inst_Sbox_8_M6}), .c ({new_AGEMA_signal_5793, SubBytesIns_Inst_Sbox_8_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M11_U1 ( .a ({new_AGEMA_signal_5053, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_5232, SubBytesIns_Inst_Sbox_8_T15}), .clk (clk), .r (Fresh[78]), .c ({new_AGEMA_signal_5460, SubBytesIns_Inst_Sbox_8_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M12_U1 ( .a ({new_AGEMA_signal_5056, SubBytesIns_Inst_Sbox_8_T4}), .b ({new_AGEMA_signal_5236, SubBytesIns_Inst_Sbox_8_T27}), .clk (clk), .r (Fresh[79]), .c ({new_AGEMA_signal_5461, SubBytesIns_Inst_Sbox_8_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M13_U1 ( .a ({new_AGEMA_signal_5461, SubBytesIns_Inst_Sbox_8_M12}), .b ({new_AGEMA_signal_5460, SubBytesIns_Inst_Sbox_8_M11}), .c ({new_AGEMA_signal_5668, SubBytesIns_Inst_Sbox_8_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M14_U1 ( .a ({new_AGEMA_signal_5054, SubBytesIns_Inst_Sbox_8_T2}), .b ({new_AGEMA_signal_5450, SubBytesIns_Inst_Sbox_8_T10}), .clk (clk), .r (Fresh[80]), .c ({new_AGEMA_signal_5669, SubBytesIns_Inst_Sbox_8_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M15_U1 ( .a ({new_AGEMA_signal_5669, SubBytesIns_Inst_Sbox_8_M14}), .b ({new_AGEMA_signal_5460, SubBytesIns_Inst_Sbox_8_M11}), .c ({new_AGEMA_signal_5794, SubBytesIns_Inst_Sbox_8_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M16_U1 ( .a ({new_AGEMA_signal_5664, SubBytesIns_Inst_Sbox_8_M3}), .b ({new_AGEMA_signal_5663, SubBytesIns_Inst_Sbox_8_M2}), .c ({new_AGEMA_signal_5795, SubBytesIns_Inst_Sbox_8_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M17_U1 ( .a ({new_AGEMA_signal_5665, SubBytesIns_Inst_Sbox_8_M5}), .b ({new_AGEMA_signal_5661, SubBytesIns_Inst_Sbox_8_T24}), .c ({new_AGEMA_signal_5796, SubBytesIns_Inst_Sbox_8_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M18_U1 ( .a ({new_AGEMA_signal_5666, SubBytesIns_Inst_Sbox_8_M8}), .b ({new_AGEMA_signal_5459, SubBytesIns_Inst_Sbox_8_M7}), .c ({new_AGEMA_signal_5797, SubBytesIns_Inst_Sbox_8_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M19_U1 ( .a ({new_AGEMA_signal_5793, SubBytesIns_Inst_Sbox_8_M10}), .b ({new_AGEMA_signal_5794, SubBytesIns_Inst_Sbox_8_M15}), .c ({new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_8_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M20_U1 ( .a ({new_AGEMA_signal_5795, SubBytesIns_Inst_Sbox_8_M16}), .b ({new_AGEMA_signal_5668, SubBytesIns_Inst_Sbox_8_M13}), .c ({new_AGEMA_signal_5882, SubBytesIns_Inst_Sbox_8_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M21_U1 ( .a ({new_AGEMA_signal_5796, SubBytesIns_Inst_Sbox_8_M17}), .b ({new_AGEMA_signal_5794, SubBytesIns_Inst_Sbox_8_M15}), .c ({new_AGEMA_signal_5883, SubBytesIns_Inst_Sbox_8_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M22_U1 ( .a ({new_AGEMA_signal_5797, SubBytesIns_Inst_Sbox_8_M18}), .b ({new_AGEMA_signal_5668, SubBytesIns_Inst_Sbox_8_M13}), .c ({new_AGEMA_signal_5884, SubBytesIns_Inst_Sbox_8_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M23_U1 ( .a ({new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_8_M19}), .b ({new_AGEMA_signal_5662, SubBytesIns_Inst_Sbox_8_T25}), .c ({new_AGEMA_signal_5961, SubBytesIns_Inst_Sbox_8_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M24_U1 ( .a ({new_AGEMA_signal_5884, SubBytesIns_Inst_Sbox_8_M22}), .b ({new_AGEMA_signal_5961, SubBytesIns_Inst_Sbox_8_M23}), .c ({new_AGEMA_signal_6053, SubBytesIns_Inst_Sbox_8_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M27_U1 ( .a ({new_AGEMA_signal_5882, SubBytesIns_Inst_Sbox_8_M20}), .b ({new_AGEMA_signal_5883, SubBytesIns_Inst_Sbox_8_M21}), .c ({new_AGEMA_signal_5963, SubBytesIns_Inst_Sbox_8_M27}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M1_U1 ( .a ({new_AGEMA_signal_5239, SubBytesIns_Inst_Sbox_9_T13}), .b ({new_AGEMA_signal_5237, SubBytesIns_Inst_Sbox_9_T6}), .clk (clk), .r (Fresh[81]), .c ({new_AGEMA_signal_5469, SubBytesIns_Inst_Sbox_9_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M2_U1 ( .a ({new_AGEMA_signal_5467, SubBytesIns_Inst_Sbox_9_T23}), .b ({new_AGEMA_signal_5462, SubBytesIns_Inst_Sbox_9_T8}), .clk (clk), .r (Fresh[82]), .c ({new_AGEMA_signal_5672, SubBytesIns_Inst_Sbox_9_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M3_U1 ( .a ({new_AGEMA_signal_5464, SubBytesIns_Inst_Sbox_9_T14}), .b ({new_AGEMA_signal_5469, SubBytesIns_Inst_Sbox_9_M1}), .c ({new_AGEMA_signal_5673, SubBytesIns_Inst_Sbox_9_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M4_U1 ( .a ({new_AGEMA_signal_5242, SubBytesIns_Inst_Sbox_9_T19}), .b ({ciphertext_s1[72], ciphertext_s0[72]}), .clk (clk), .r (Fresh[83]), .c ({new_AGEMA_signal_5470, SubBytesIns_Inst_Sbox_9_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M5_U1 ( .a ({new_AGEMA_signal_5470, SubBytesIns_Inst_Sbox_9_M4}), .b ({new_AGEMA_signal_5469, SubBytesIns_Inst_Sbox_9_M1}), .c ({new_AGEMA_signal_5674, SubBytesIns_Inst_Sbox_9_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M6_U1 ( .a ({new_AGEMA_signal_5065, SubBytesIns_Inst_Sbox_9_T3}), .b ({new_AGEMA_signal_5241, SubBytesIns_Inst_Sbox_9_T16}), .clk (clk), .r (Fresh[84]), .c ({new_AGEMA_signal_5471, SubBytesIns_Inst_Sbox_9_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M7_U1 ( .a ({new_AGEMA_signal_5243, SubBytesIns_Inst_Sbox_9_T22}), .b ({new_AGEMA_signal_5238, SubBytesIns_Inst_Sbox_9_T9}), .clk (clk), .r (Fresh[85]), .c ({new_AGEMA_signal_5472, SubBytesIns_Inst_Sbox_9_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M8_U1 ( .a ({new_AGEMA_signal_5468, SubBytesIns_Inst_Sbox_9_T26}), .b ({new_AGEMA_signal_5471, SubBytesIns_Inst_Sbox_9_M6}), .c ({new_AGEMA_signal_5675, SubBytesIns_Inst_Sbox_9_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M9_U1 ( .a ({new_AGEMA_signal_5466, SubBytesIns_Inst_Sbox_9_T20}), .b ({new_AGEMA_signal_5465, SubBytesIns_Inst_Sbox_9_T17}), .clk (clk), .r (Fresh[86]), .c ({new_AGEMA_signal_5676, SubBytesIns_Inst_Sbox_9_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M10_U1 ( .a ({new_AGEMA_signal_5676, SubBytesIns_Inst_Sbox_9_M9}), .b ({new_AGEMA_signal_5471, SubBytesIns_Inst_Sbox_9_M6}), .c ({new_AGEMA_signal_5798, SubBytesIns_Inst_Sbox_9_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M11_U1 ( .a ({new_AGEMA_signal_5063, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_5240, SubBytesIns_Inst_Sbox_9_T15}), .clk (clk), .r (Fresh[87]), .c ({new_AGEMA_signal_5473, SubBytesIns_Inst_Sbox_9_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M12_U1 ( .a ({new_AGEMA_signal_5066, SubBytesIns_Inst_Sbox_9_T4}), .b ({new_AGEMA_signal_5244, SubBytesIns_Inst_Sbox_9_T27}), .clk (clk), .r (Fresh[88]), .c ({new_AGEMA_signal_5474, SubBytesIns_Inst_Sbox_9_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M13_U1 ( .a ({new_AGEMA_signal_5474, SubBytesIns_Inst_Sbox_9_M12}), .b ({new_AGEMA_signal_5473, SubBytesIns_Inst_Sbox_9_M11}), .c ({new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_9_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M14_U1 ( .a ({new_AGEMA_signal_5064, SubBytesIns_Inst_Sbox_9_T2}), .b ({new_AGEMA_signal_5463, SubBytesIns_Inst_Sbox_9_T10}), .clk (clk), .r (Fresh[89]), .c ({new_AGEMA_signal_5678, SubBytesIns_Inst_Sbox_9_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M15_U1 ( .a ({new_AGEMA_signal_5678, SubBytesIns_Inst_Sbox_9_M14}), .b ({new_AGEMA_signal_5473, SubBytesIns_Inst_Sbox_9_M11}), .c ({new_AGEMA_signal_5799, SubBytesIns_Inst_Sbox_9_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M16_U1 ( .a ({new_AGEMA_signal_5673, SubBytesIns_Inst_Sbox_9_M3}), .b ({new_AGEMA_signal_5672, SubBytesIns_Inst_Sbox_9_M2}), .c ({new_AGEMA_signal_5800, SubBytesIns_Inst_Sbox_9_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M17_U1 ( .a ({new_AGEMA_signal_5674, SubBytesIns_Inst_Sbox_9_M5}), .b ({new_AGEMA_signal_5670, SubBytesIns_Inst_Sbox_9_T24}), .c ({new_AGEMA_signal_5801, SubBytesIns_Inst_Sbox_9_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M18_U1 ( .a ({new_AGEMA_signal_5675, SubBytesIns_Inst_Sbox_9_M8}), .b ({new_AGEMA_signal_5472, SubBytesIns_Inst_Sbox_9_M7}), .c ({new_AGEMA_signal_5802, SubBytesIns_Inst_Sbox_9_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M19_U1 ( .a ({new_AGEMA_signal_5798, SubBytesIns_Inst_Sbox_9_M10}), .b ({new_AGEMA_signal_5799, SubBytesIns_Inst_Sbox_9_M15}), .c ({new_AGEMA_signal_5885, SubBytesIns_Inst_Sbox_9_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M20_U1 ( .a ({new_AGEMA_signal_5800, SubBytesIns_Inst_Sbox_9_M16}), .b ({new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_9_M13}), .c ({new_AGEMA_signal_5886, SubBytesIns_Inst_Sbox_9_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M21_U1 ( .a ({new_AGEMA_signal_5801, SubBytesIns_Inst_Sbox_9_M17}), .b ({new_AGEMA_signal_5799, SubBytesIns_Inst_Sbox_9_M15}), .c ({new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_9_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M22_U1 ( .a ({new_AGEMA_signal_5802, SubBytesIns_Inst_Sbox_9_M18}), .b ({new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_9_M13}), .c ({new_AGEMA_signal_5888, SubBytesIns_Inst_Sbox_9_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M23_U1 ( .a ({new_AGEMA_signal_5885, SubBytesIns_Inst_Sbox_9_M19}), .b ({new_AGEMA_signal_5671, SubBytesIns_Inst_Sbox_9_T25}), .c ({new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_9_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M24_U1 ( .a ({new_AGEMA_signal_5888, SubBytesIns_Inst_Sbox_9_M22}), .b ({new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_9_M23}), .c ({new_AGEMA_signal_6058, SubBytesIns_Inst_Sbox_9_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M27_U1 ( .a ({new_AGEMA_signal_5886, SubBytesIns_Inst_Sbox_9_M20}), .b ({new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_9_M21}), .c ({new_AGEMA_signal_5967, SubBytesIns_Inst_Sbox_9_M27}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M1_U1 ( .a ({new_AGEMA_signal_5247, SubBytesIns_Inst_Sbox_10_T13}), .b ({new_AGEMA_signal_5245, SubBytesIns_Inst_Sbox_10_T6}), .clk (clk), .r (Fresh[90]), .c ({new_AGEMA_signal_5482, SubBytesIns_Inst_Sbox_10_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M2_U1 ( .a ({new_AGEMA_signal_5480, SubBytesIns_Inst_Sbox_10_T23}), .b ({new_AGEMA_signal_5475, SubBytesIns_Inst_Sbox_10_T8}), .clk (clk), .r (Fresh[91]), .c ({new_AGEMA_signal_5681, SubBytesIns_Inst_Sbox_10_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M3_U1 ( .a ({new_AGEMA_signal_5477, SubBytesIns_Inst_Sbox_10_T14}), .b ({new_AGEMA_signal_5482, SubBytesIns_Inst_Sbox_10_M1}), .c ({new_AGEMA_signal_5682, SubBytesIns_Inst_Sbox_10_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M4_U1 ( .a ({new_AGEMA_signal_5250, SubBytesIns_Inst_Sbox_10_T19}), .b ({ciphertext_s1[80], ciphertext_s0[80]}), .clk (clk), .r (Fresh[92]), .c ({new_AGEMA_signal_5483, SubBytesIns_Inst_Sbox_10_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M5_U1 ( .a ({new_AGEMA_signal_5483, SubBytesIns_Inst_Sbox_10_M4}), .b ({new_AGEMA_signal_5482, SubBytesIns_Inst_Sbox_10_M1}), .c ({new_AGEMA_signal_5683, SubBytesIns_Inst_Sbox_10_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M6_U1 ( .a ({new_AGEMA_signal_5075, SubBytesIns_Inst_Sbox_10_T3}), .b ({new_AGEMA_signal_5249, SubBytesIns_Inst_Sbox_10_T16}), .clk (clk), .r (Fresh[93]), .c ({new_AGEMA_signal_5484, SubBytesIns_Inst_Sbox_10_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M7_U1 ( .a ({new_AGEMA_signal_5251, SubBytesIns_Inst_Sbox_10_T22}), .b ({new_AGEMA_signal_5246, SubBytesIns_Inst_Sbox_10_T9}), .clk (clk), .r (Fresh[94]), .c ({new_AGEMA_signal_5485, SubBytesIns_Inst_Sbox_10_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M8_U1 ( .a ({new_AGEMA_signal_5481, SubBytesIns_Inst_Sbox_10_T26}), .b ({new_AGEMA_signal_5484, SubBytesIns_Inst_Sbox_10_M6}), .c ({new_AGEMA_signal_5684, SubBytesIns_Inst_Sbox_10_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M9_U1 ( .a ({new_AGEMA_signal_5479, SubBytesIns_Inst_Sbox_10_T20}), .b ({new_AGEMA_signal_5478, SubBytesIns_Inst_Sbox_10_T17}), .clk (clk), .r (Fresh[95]), .c ({new_AGEMA_signal_5685, SubBytesIns_Inst_Sbox_10_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M10_U1 ( .a ({new_AGEMA_signal_5685, SubBytesIns_Inst_Sbox_10_M9}), .b ({new_AGEMA_signal_5484, SubBytesIns_Inst_Sbox_10_M6}), .c ({new_AGEMA_signal_5803, SubBytesIns_Inst_Sbox_10_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M11_U1 ( .a ({new_AGEMA_signal_5073, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_5248, SubBytesIns_Inst_Sbox_10_T15}), .clk (clk), .r (Fresh[96]), .c ({new_AGEMA_signal_5486, SubBytesIns_Inst_Sbox_10_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M12_U1 ( .a ({new_AGEMA_signal_5076, SubBytesIns_Inst_Sbox_10_T4}), .b ({new_AGEMA_signal_5252, SubBytesIns_Inst_Sbox_10_T27}), .clk (clk), .r (Fresh[97]), .c ({new_AGEMA_signal_5487, SubBytesIns_Inst_Sbox_10_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M13_U1 ( .a ({new_AGEMA_signal_5487, SubBytesIns_Inst_Sbox_10_M12}), .b ({new_AGEMA_signal_5486, SubBytesIns_Inst_Sbox_10_M11}), .c ({new_AGEMA_signal_5686, SubBytesIns_Inst_Sbox_10_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M14_U1 ( .a ({new_AGEMA_signal_5074, SubBytesIns_Inst_Sbox_10_T2}), .b ({new_AGEMA_signal_5476, SubBytesIns_Inst_Sbox_10_T10}), .clk (clk), .r (Fresh[98]), .c ({new_AGEMA_signal_5687, SubBytesIns_Inst_Sbox_10_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M15_U1 ( .a ({new_AGEMA_signal_5687, SubBytesIns_Inst_Sbox_10_M14}), .b ({new_AGEMA_signal_5486, SubBytesIns_Inst_Sbox_10_M11}), .c ({new_AGEMA_signal_5804, SubBytesIns_Inst_Sbox_10_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M16_U1 ( .a ({new_AGEMA_signal_5682, SubBytesIns_Inst_Sbox_10_M3}), .b ({new_AGEMA_signal_5681, SubBytesIns_Inst_Sbox_10_M2}), .c ({new_AGEMA_signal_5805, SubBytesIns_Inst_Sbox_10_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M17_U1 ( .a ({new_AGEMA_signal_5683, SubBytesIns_Inst_Sbox_10_M5}), .b ({new_AGEMA_signal_5679, SubBytesIns_Inst_Sbox_10_T24}), .c ({new_AGEMA_signal_5806, SubBytesIns_Inst_Sbox_10_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M18_U1 ( .a ({new_AGEMA_signal_5684, SubBytesIns_Inst_Sbox_10_M8}), .b ({new_AGEMA_signal_5485, SubBytesIns_Inst_Sbox_10_M7}), .c ({new_AGEMA_signal_5807, SubBytesIns_Inst_Sbox_10_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M19_U1 ( .a ({new_AGEMA_signal_5803, SubBytesIns_Inst_Sbox_10_M10}), .b ({new_AGEMA_signal_5804, SubBytesIns_Inst_Sbox_10_M15}), .c ({new_AGEMA_signal_5889, SubBytesIns_Inst_Sbox_10_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M20_U1 ( .a ({new_AGEMA_signal_5805, SubBytesIns_Inst_Sbox_10_M16}), .b ({new_AGEMA_signal_5686, SubBytesIns_Inst_Sbox_10_M13}), .c ({new_AGEMA_signal_5890, SubBytesIns_Inst_Sbox_10_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M21_U1 ( .a ({new_AGEMA_signal_5806, SubBytesIns_Inst_Sbox_10_M17}), .b ({new_AGEMA_signal_5804, SubBytesIns_Inst_Sbox_10_M15}), .c ({new_AGEMA_signal_5891, SubBytesIns_Inst_Sbox_10_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M22_U1 ( .a ({new_AGEMA_signal_5807, SubBytesIns_Inst_Sbox_10_M18}), .b ({new_AGEMA_signal_5686, SubBytesIns_Inst_Sbox_10_M13}), .c ({new_AGEMA_signal_5892, SubBytesIns_Inst_Sbox_10_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M23_U1 ( .a ({new_AGEMA_signal_5889, SubBytesIns_Inst_Sbox_10_M19}), .b ({new_AGEMA_signal_5680, SubBytesIns_Inst_Sbox_10_T25}), .c ({new_AGEMA_signal_5969, SubBytesIns_Inst_Sbox_10_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M24_U1 ( .a ({new_AGEMA_signal_5892, SubBytesIns_Inst_Sbox_10_M22}), .b ({new_AGEMA_signal_5969, SubBytesIns_Inst_Sbox_10_M23}), .c ({new_AGEMA_signal_6063, SubBytesIns_Inst_Sbox_10_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M27_U1 ( .a ({new_AGEMA_signal_5890, SubBytesIns_Inst_Sbox_10_M20}), .b ({new_AGEMA_signal_5891, SubBytesIns_Inst_Sbox_10_M21}), .c ({new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_10_M27}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M1_U1 ( .a ({new_AGEMA_signal_5255, SubBytesIns_Inst_Sbox_11_T13}), .b ({new_AGEMA_signal_5253, SubBytesIns_Inst_Sbox_11_T6}), .clk (clk), .r (Fresh[99]), .c ({new_AGEMA_signal_5495, SubBytesIns_Inst_Sbox_11_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M2_U1 ( .a ({new_AGEMA_signal_5493, SubBytesIns_Inst_Sbox_11_T23}), .b ({new_AGEMA_signal_5488, SubBytesIns_Inst_Sbox_11_T8}), .clk (clk), .r (Fresh[100]), .c ({new_AGEMA_signal_5690, SubBytesIns_Inst_Sbox_11_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M3_U1 ( .a ({new_AGEMA_signal_5490, SubBytesIns_Inst_Sbox_11_T14}), .b ({new_AGEMA_signal_5495, SubBytesIns_Inst_Sbox_11_M1}), .c ({new_AGEMA_signal_5691, SubBytesIns_Inst_Sbox_11_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M4_U1 ( .a ({new_AGEMA_signal_5258, SubBytesIns_Inst_Sbox_11_T19}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .clk (clk), .r (Fresh[101]), .c ({new_AGEMA_signal_5496, SubBytesIns_Inst_Sbox_11_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M5_U1 ( .a ({new_AGEMA_signal_5496, SubBytesIns_Inst_Sbox_11_M4}), .b ({new_AGEMA_signal_5495, SubBytesIns_Inst_Sbox_11_M1}), .c ({new_AGEMA_signal_5692, SubBytesIns_Inst_Sbox_11_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M6_U1 ( .a ({new_AGEMA_signal_5085, SubBytesIns_Inst_Sbox_11_T3}), .b ({new_AGEMA_signal_5257, SubBytesIns_Inst_Sbox_11_T16}), .clk (clk), .r (Fresh[102]), .c ({new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_11_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M7_U1 ( .a ({new_AGEMA_signal_5259, SubBytesIns_Inst_Sbox_11_T22}), .b ({new_AGEMA_signal_5254, SubBytesIns_Inst_Sbox_11_T9}), .clk (clk), .r (Fresh[103]), .c ({new_AGEMA_signal_5498, SubBytesIns_Inst_Sbox_11_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M8_U1 ( .a ({new_AGEMA_signal_5494, SubBytesIns_Inst_Sbox_11_T26}), .b ({new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_11_M6}), .c ({new_AGEMA_signal_5693, SubBytesIns_Inst_Sbox_11_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M9_U1 ( .a ({new_AGEMA_signal_5492, SubBytesIns_Inst_Sbox_11_T20}), .b ({new_AGEMA_signal_5491, SubBytesIns_Inst_Sbox_11_T17}), .clk (clk), .r (Fresh[104]), .c ({new_AGEMA_signal_5694, SubBytesIns_Inst_Sbox_11_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M10_U1 ( .a ({new_AGEMA_signal_5694, SubBytesIns_Inst_Sbox_11_M9}), .b ({new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_11_M6}), .c ({new_AGEMA_signal_5808, SubBytesIns_Inst_Sbox_11_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M11_U1 ( .a ({new_AGEMA_signal_5083, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_5256, SubBytesIns_Inst_Sbox_11_T15}), .clk (clk), .r (Fresh[105]), .c ({new_AGEMA_signal_5499, SubBytesIns_Inst_Sbox_11_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M12_U1 ( .a ({new_AGEMA_signal_5086, SubBytesIns_Inst_Sbox_11_T4}), .b ({new_AGEMA_signal_5260, SubBytesIns_Inst_Sbox_11_T27}), .clk (clk), .r (Fresh[106]), .c ({new_AGEMA_signal_5500, SubBytesIns_Inst_Sbox_11_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M13_U1 ( .a ({new_AGEMA_signal_5500, SubBytesIns_Inst_Sbox_11_M12}), .b ({new_AGEMA_signal_5499, SubBytesIns_Inst_Sbox_11_M11}), .c ({new_AGEMA_signal_5695, SubBytesIns_Inst_Sbox_11_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M14_U1 ( .a ({new_AGEMA_signal_5084, SubBytesIns_Inst_Sbox_11_T2}), .b ({new_AGEMA_signal_5489, SubBytesIns_Inst_Sbox_11_T10}), .clk (clk), .r (Fresh[107]), .c ({new_AGEMA_signal_5696, SubBytesIns_Inst_Sbox_11_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M15_U1 ( .a ({new_AGEMA_signal_5696, SubBytesIns_Inst_Sbox_11_M14}), .b ({new_AGEMA_signal_5499, SubBytesIns_Inst_Sbox_11_M11}), .c ({new_AGEMA_signal_5809, SubBytesIns_Inst_Sbox_11_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M16_U1 ( .a ({new_AGEMA_signal_5691, SubBytesIns_Inst_Sbox_11_M3}), .b ({new_AGEMA_signal_5690, SubBytesIns_Inst_Sbox_11_M2}), .c ({new_AGEMA_signal_5810, SubBytesIns_Inst_Sbox_11_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M17_U1 ( .a ({new_AGEMA_signal_5692, SubBytesIns_Inst_Sbox_11_M5}), .b ({new_AGEMA_signal_5688, SubBytesIns_Inst_Sbox_11_T24}), .c ({new_AGEMA_signal_5811, SubBytesIns_Inst_Sbox_11_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M18_U1 ( .a ({new_AGEMA_signal_5693, SubBytesIns_Inst_Sbox_11_M8}), .b ({new_AGEMA_signal_5498, SubBytesIns_Inst_Sbox_11_M7}), .c ({new_AGEMA_signal_5812, SubBytesIns_Inst_Sbox_11_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M19_U1 ( .a ({new_AGEMA_signal_5808, SubBytesIns_Inst_Sbox_11_M10}), .b ({new_AGEMA_signal_5809, SubBytesIns_Inst_Sbox_11_M15}), .c ({new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_11_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M20_U1 ( .a ({new_AGEMA_signal_5810, SubBytesIns_Inst_Sbox_11_M16}), .b ({new_AGEMA_signal_5695, SubBytesIns_Inst_Sbox_11_M13}), .c ({new_AGEMA_signal_5894, SubBytesIns_Inst_Sbox_11_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M21_U1 ( .a ({new_AGEMA_signal_5811, SubBytesIns_Inst_Sbox_11_M17}), .b ({new_AGEMA_signal_5809, SubBytesIns_Inst_Sbox_11_M15}), .c ({new_AGEMA_signal_5895, SubBytesIns_Inst_Sbox_11_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M22_U1 ( .a ({new_AGEMA_signal_5812, SubBytesIns_Inst_Sbox_11_M18}), .b ({new_AGEMA_signal_5695, SubBytesIns_Inst_Sbox_11_M13}), .c ({new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_11_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M23_U1 ( .a ({new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_11_M19}), .b ({new_AGEMA_signal_5689, SubBytesIns_Inst_Sbox_11_T25}), .c ({new_AGEMA_signal_5973, SubBytesIns_Inst_Sbox_11_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M24_U1 ( .a ({new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_11_M22}), .b ({new_AGEMA_signal_5973, SubBytesIns_Inst_Sbox_11_M23}), .c ({new_AGEMA_signal_6068, SubBytesIns_Inst_Sbox_11_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M27_U1 ( .a ({new_AGEMA_signal_5894, SubBytesIns_Inst_Sbox_11_M20}), .b ({new_AGEMA_signal_5895, SubBytesIns_Inst_Sbox_11_M21}), .c ({new_AGEMA_signal_5975, SubBytesIns_Inst_Sbox_11_M27}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M1_U1 ( .a ({new_AGEMA_signal_5263, SubBytesIns_Inst_Sbox_12_T13}), .b ({new_AGEMA_signal_5261, SubBytesIns_Inst_Sbox_12_T6}), .clk (clk), .r (Fresh[108]), .c ({new_AGEMA_signal_5508, SubBytesIns_Inst_Sbox_12_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M2_U1 ( .a ({new_AGEMA_signal_5506, SubBytesIns_Inst_Sbox_12_T23}), .b ({new_AGEMA_signal_5501, SubBytesIns_Inst_Sbox_12_T8}), .clk (clk), .r (Fresh[109]), .c ({new_AGEMA_signal_5699, SubBytesIns_Inst_Sbox_12_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M3_U1 ( .a ({new_AGEMA_signal_5503, SubBytesIns_Inst_Sbox_12_T14}), .b ({new_AGEMA_signal_5508, SubBytesIns_Inst_Sbox_12_M1}), .c ({new_AGEMA_signal_5700, SubBytesIns_Inst_Sbox_12_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M4_U1 ( .a ({new_AGEMA_signal_5266, SubBytesIns_Inst_Sbox_12_T19}), .b ({ciphertext_s1[96], ciphertext_s0[96]}), .clk (clk), .r (Fresh[110]), .c ({new_AGEMA_signal_5509, SubBytesIns_Inst_Sbox_12_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M5_U1 ( .a ({new_AGEMA_signal_5509, SubBytesIns_Inst_Sbox_12_M4}), .b ({new_AGEMA_signal_5508, SubBytesIns_Inst_Sbox_12_M1}), .c ({new_AGEMA_signal_5701, SubBytesIns_Inst_Sbox_12_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M6_U1 ( .a ({new_AGEMA_signal_5095, SubBytesIns_Inst_Sbox_12_T3}), .b ({new_AGEMA_signal_5265, SubBytesIns_Inst_Sbox_12_T16}), .clk (clk), .r (Fresh[111]), .c ({new_AGEMA_signal_5510, SubBytesIns_Inst_Sbox_12_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M7_U1 ( .a ({new_AGEMA_signal_5267, SubBytesIns_Inst_Sbox_12_T22}), .b ({new_AGEMA_signal_5262, SubBytesIns_Inst_Sbox_12_T9}), .clk (clk), .r (Fresh[112]), .c ({new_AGEMA_signal_5511, SubBytesIns_Inst_Sbox_12_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M8_U1 ( .a ({new_AGEMA_signal_5507, SubBytesIns_Inst_Sbox_12_T26}), .b ({new_AGEMA_signal_5510, SubBytesIns_Inst_Sbox_12_M6}), .c ({new_AGEMA_signal_5702, SubBytesIns_Inst_Sbox_12_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M9_U1 ( .a ({new_AGEMA_signal_5505, SubBytesIns_Inst_Sbox_12_T20}), .b ({new_AGEMA_signal_5504, SubBytesIns_Inst_Sbox_12_T17}), .clk (clk), .r (Fresh[113]), .c ({new_AGEMA_signal_5703, SubBytesIns_Inst_Sbox_12_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M10_U1 ( .a ({new_AGEMA_signal_5703, SubBytesIns_Inst_Sbox_12_M9}), .b ({new_AGEMA_signal_5510, SubBytesIns_Inst_Sbox_12_M6}), .c ({new_AGEMA_signal_5813, SubBytesIns_Inst_Sbox_12_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M11_U1 ( .a ({new_AGEMA_signal_5093, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_5264, SubBytesIns_Inst_Sbox_12_T15}), .clk (clk), .r (Fresh[114]), .c ({new_AGEMA_signal_5512, SubBytesIns_Inst_Sbox_12_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M12_U1 ( .a ({new_AGEMA_signal_5096, SubBytesIns_Inst_Sbox_12_T4}), .b ({new_AGEMA_signal_5268, SubBytesIns_Inst_Sbox_12_T27}), .clk (clk), .r (Fresh[115]), .c ({new_AGEMA_signal_5513, SubBytesIns_Inst_Sbox_12_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M13_U1 ( .a ({new_AGEMA_signal_5513, SubBytesIns_Inst_Sbox_12_M12}), .b ({new_AGEMA_signal_5512, SubBytesIns_Inst_Sbox_12_M11}), .c ({new_AGEMA_signal_5704, SubBytesIns_Inst_Sbox_12_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M14_U1 ( .a ({new_AGEMA_signal_5094, SubBytesIns_Inst_Sbox_12_T2}), .b ({new_AGEMA_signal_5502, SubBytesIns_Inst_Sbox_12_T10}), .clk (clk), .r (Fresh[116]), .c ({new_AGEMA_signal_5705, SubBytesIns_Inst_Sbox_12_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M15_U1 ( .a ({new_AGEMA_signal_5705, SubBytesIns_Inst_Sbox_12_M14}), .b ({new_AGEMA_signal_5512, SubBytesIns_Inst_Sbox_12_M11}), .c ({new_AGEMA_signal_5814, SubBytesIns_Inst_Sbox_12_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M16_U1 ( .a ({new_AGEMA_signal_5700, SubBytesIns_Inst_Sbox_12_M3}), .b ({new_AGEMA_signal_5699, SubBytesIns_Inst_Sbox_12_M2}), .c ({new_AGEMA_signal_5815, SubBytesIns_Inst_Sbox_12_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M17_U1 ( .a ({new_AGEMA_signal_5701, SubBytesIns_Inst_Sbox_12_M5}), .b ({new_AGEMA_signal_5697, SubBytesIns_Inst_Sbox_12_T24}), .c ({new_AGEMA_signal_5816, SubBytesIns_Inst_Sbox_12_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M18_U1 ( .a ({new_AGEMA_signal_5702, SubBytesIns_Inst_Sbox_12_M8}), .b ({new_AGEMA_signal_5511, SubBytesIns_Inst_Sbox_12_M7}), .c ({new_AGEMA_signal_5817, SubBytesIns_Inst_Sbox_12_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M19_U1 ( .a ({new_AGEMA_signal_5813, SubBytesIns_Inst_Sbox_12_M10}), .b ({new_AGEMA_signal_5814, SubBytesIns_Inst_Sbox_12_M15}), .c ({new_AGEMA_signal_5897, SubBytesIns_Inst_Sbox_12_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M20_U1 ( .a ({new_AGEMA_signal_5815, SubBytesIns_Inst_Sbox_12_M16}), .b ({new_AGEMA_signal_5704, SubBytesIns_Inst_Sbox_12_M13}), .c ({new_AGEMA_signal_5898, SubBytesIns_Inst_Sbox_12_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M21_U1 ( .a ({new_AGEMA_signal_5816, SubBytesIns_Inst_Sbox_12_M17}), .b ({new_AGEMA_signal_5814, SubBytesIns_Inst_Sbox_12_M15}), .c ({new_AGEMA_signal_5899, SubBytesIns_Inst_Sbox_12_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M22_U1 ( .a ({new_AGEMA_signal_5817, SubBytesIns_Inst_Sbox_12_M18}), .b ({new_AGEMA_signal_5704, SubBytesIns_Inst_Sbox_12_M13}), .c ({new_AGEMA_signal_5900, SubBytesIns_Inst_Sbox_12_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M23_U1 ( .a ({new_AGEMA_signal_5897, SubBytesIns_Inst_Sbox_12_M19}), .b ({new_AGEMA_signal_5698, SubBytesIns_Inst_Sbox_12_T25}), .c ({new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_12_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M24_U1 ( .a ({new_AGEMA_signal_5900, SubBytesIns_Inst_Sbox_12_M22}), .b ({new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_12_M23}), .c ({new_AGEMA_signal_6073, SubBytesIns_Inst_Sbox_12_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M27_U1 ( .a ({new_AGEMA_signal_5898, SubBytesIns_Inst_Sbox_12_M20}), .b ({new_AGEMA_signal_5899, SubBytesIns_Inst_Sbox_12_M21}), .c ({new_AGEMA_signal_5979, SubBytesIns_Inst_Sbox_12_M27}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M1_U1 ( .a ({new_AGEMA_signal_5271, SubBytesIns_Inst_Sbox_13_T13}), .b ({new_AGEMA_signal_5269, SubBytesIns_Inst_Sbox_13_T6}), .clk (clk), .r (Fresh[117]), .c ({new_AGEMA_signal_5521, SubBytesIns_Inst_Sbox_13_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M2_U1 ( .a ({new_AGEMA_signal_5519, SubBytesIns_Inst_Sbox_13_T23}), .b ({new_AGEMA_signal_5514, SubBytesIns_Inst_Sbox_13_T8}), .clk (clk), .r (Fresh[118]), .c ({new_AGEMA_signal_5708, SubBytesIns_Inst_Sbox_13_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M3_U1 ( .a ({new_AGEMA_signal_5516, SubBytesIns_Inst_Sbox_13_T14}), .b ({new_AGEMA_signal_5521, SubBytesIns_Inst_Sbox_13_M1}), .c ({new_AGEMA_signal_5709, SubBytesIns_Inst_Sbox_13_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M4_U1 ( .a ({new_AGEMA_signal_5274, SubBytesIns_Inst_Sbox_13_T19}), .b ({ciphertext_s1[104], ciphertext_s0[104]}), .clk (clk), .r (Fresh[119]), .c ({new_AGEMA_signal_5522, SubBytesIns_Inst_Sbox_13_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M5_U1 ( .a ({new_AGEMA_signal_5522, SubBytesIns_Inst_Sbox_13_M4}), .b ({new_AGEMA_signal_5521, SubBytesIns_Inst_Sbox_13_M1}), .c ({new_AGEMA_signal_5710, SubBytesIns_Inst_Sbox_13_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M6_U1 ( .a ({new_AGEMA_signal_5105, SubBytesIns_Inst_Sbox_13_T3}), .b ({new_AGEMA_signal_5273, SubBytesIns_Inst_Sbox_13_T16}), .clk (clk), .r (Fresh[120]), .c ({new_AGEMA_signal_5523, SubBytesIns_Inst_Sbox_13_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M7_U1 ( .a ({new_AGEMA_signal_5275, SubBytesIns_Inst_Sbox_13_T22}), .b ({new_AGEMA_signal_5270, SubBytesIns_Inst_Sbox_13_T9}), .clk (clk), .r (Fresh[121]), .c ({new_AGEMA_signal_5524, SubBytesIns_Inst_Sbox_13_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M8_U1 ( .a ({new_AGEMA_signal_5520, SubBytesIns_Inst_Sbox_13_T26}), .b ({new_AGEMA_signal_5523, SubBytesIns_Inst_Sbox_13_M6}), .c ({new_AGEMA_signal_5711, SubBytesIns_Inst_Sbox_13_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M9_U1 ( .a ({new_AGEMA_signal_5518, SubBytesIns_Inst_Sbox_13_T20}), .b ({new_AGEMA_signal_5517, SubBytesIns_Inst_Sbox_13_T17}), .clk (clk), .r (Fresh[122]), .c ({new_AGEMA_signal_5712, SubBytesIns_Inst_Sbox_13_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M10_U1 ( .a ({new_AGEMA_signal_5712, SubBytesIns_Inst_Sbox_13_M9}), .b ({new_AGEMA_signal_5523, SubBytesIns_Inst_Sbox_13_M6}), .c ({new_AGEMA_signal_5818, SubBytesIns_Inst_Sbox_13_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M11_U1 ( .a ({new_AGEMA_signal_5103, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_5272, SubBytesIns_Inst_Sbox_13_T15}), .clk (clk), .r (Fresh[123]), .c ({new_AGEMA_signal_5525, SubBytesIns_Inst_Sbox_13_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M12_U1 ( .a ({new_AGEMA_signal_5106, SubBytesIns_Inst_Sbox_13_T4}), .b ({new_AGEMA_signal_5276, SubBytesIns_Inst_Sbox_13_T27}), .clk (clk), .r (Fresh[124]), .c ({new_AGEMA_signal_5526, SubBytesIns_Inst_Sbox_13_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M13_U1 ( .a ({new_AGEMA_signal_5526, SubBytesIns_Inst_Sbox_13_M12}), .b ({new_AGEMA_signal_5525, SubBytesIns_Inst_Sbox_13_M11}), .c ({new_AGEMA_signal_5713, SubBytesIns_Inst_Sbox_13_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M14_U1 ( .a ({new_AGEMA_signal_5104, SubBytesIns_Inst_Sbox_13_T2}), .b ({new_AGEMA_signal_5515, SubBytesIns_Inst_Sbox_13_T10}), .clk (clk), .r (Fresh[125]), .c ({new_AGEMA_signal_5714, SubBytesIns_Inst_Sbox_13_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M15_U1 ( .a ({new_AGEMA_signal_5714, SubBytesIns_Inst_Sbox_13_M14}), .b ({new_AGEMA_signal_5525, SubBytesIns_Inst_Sbox_13_M11}), .c ({new_AGEMA_signal_5819, SubBytesIns_Inst_Sbox_13_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M16_U1 ( .a ({new_AGEMA_signal_5709, SubBytesIns_Inst_Sbox_13_M3}), .b ({new_AGEMA_signal_5708, SubBytesIns_Inst_Sbox_13_M2}), .c ({new_AGEMA_signal_5820, SubBytesIns_Inst_Sbox_13_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M17_U1 ( .a ({new_AGEMA_signal_5710, SubBytesIns_Inst_Sbox_13_M5}), .b ({new_AGEMA_signal_5706, SubBytesIns_Inst_Sbox_13_T24}), .c ({new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_13_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M18_U1 ( .a ({new_AGEMA_signal_5711, SubBytesIns_Inst_Sbox_13_M8}), .b ({new_AGEMA_signal_5524, SubBytesIns_Inst_Sbox_13_M7}), .c ({new_AGEMA_signal_5822, SubBytesIns_Inst_Sbox_13_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M19_U1 ( .a ({new_AGEMA_signal_5818, SubBytesIns_Inst_Sbox_13_M10}), .b ({new_AGEMA_signal_5819, SubBytesIns_Inst_Sbox_13_M15}), .c ({new_AGEMA_signal_5901, SubBytesIns_Inst_Sbox_13_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M20_U1 ( .a ({new_AGEMA_signal_5820, SubBytesIns_Inst_Sbox_13_M16}), .b ({new_AGEMA_signal_5713, SubBytesIns_Inst_Sbox_13_M13}), .c ({new_AGEMA_signal_5902, SubBytesIns_Inst_Sbox_13_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M21_U1 ( .a ({new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_13_M17}), .b ({new_AGEMA_signal_5819, SubBytesIns_Inst_Sbox_13_M15}), .c ({new_AGEMA_signal_5903, SubBytesIns_Inst_Sbox_13_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M22_U1 ( .a ({new_AGEMA_signal_5822, SubBytesIns_Inst_Sbox_13_M18}), .b ({new_AGEMA_signal_5713, SubBytesIns_Inst_Sbox_13_M13}), .c ({new_AGEMA_signal_5904, SubBytesIns_Inst_Sbox_13_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M23_U1 ( .a ({new_AGEMA_signal_5901, SubBytesIns_Inst_Sbox_13_M19}), .b ({new_AGEMA_signal_5707, SubBytesIns_Inst_Sbox_13_T25}), .c ({new_AGEMA_signal_5981, SubBytesIns_Inst_Sbox_13_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M24_U1 ( .a ({new_AGEMA_signal_5904, SubBytesIns_Inst_Sbox_13_M22}), .b ({new_AGEMA_signal_5981, SubBytesIns_Inst_Sbox_13_M23}), .c ({new_AGEMA_signal_6078, SubBytesIns_Inst_Sbox_13_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M27_U1 ( .a ({new_AGEMA_signal_5902, SubBytesIns_Inst_Sbox_13_M20}), .b ({new_AGEMA_signal_5903, SubBytesIns_Inst_Sbox_13_M21}), .c ({new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_13_M27}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M1_U1 ( .a ({new_AGEMA_signal_5279, SubBytesIns_Inst_Sbox_14_T13}), .b ({new_AGEMA_signal_5277, SubBytesIns_Inst_Sbox_14_T6}), .clk (clk), .r (Fresh[126]), .c ({new_AGEMA_signal_5534, SubBytesIns_Inst_Sbox_14_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M2_U1 ( .a ({new_AGEMA_signal_5532, SubBytesIns_Inst_Sbox_14_T23}), .b ({new_AGEMA_signal_5527, SubBytesIns_Inst_Sbox_14_T8}), .clk (clk), .r (Fresh[127]), .c ({new_AGEMA_signal_5717, SubBytesIns_Inst_Sbox_14_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M3_U1 ( .a ({new_AGEMA_signal_5529, SubBytesIns_Inst_Sbox_14_T14}), .b ({new_AGEMA_signal_5534, SubBytesIns_Inst_Sbox_14_M1}), .c ({new_AGEMA_signal_5718, SubBytesIns_Inst_Sbox_14_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M4_U1 ( .a ({new_AGEMA_signal_5282, SubBytesIns_Inst_Sbox_14_T19}), .b ({ciphertext_s1[112], ciphertext_s0[112]}), .clk (clk), .r (Fresh[128]), .c ({new_AGEMA_signal_5535, SubBytesIns_Inst_Sbox_14_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M5_U1 ( .a ({new_AGEMA_signal_5535, SubBytesIns_Inst_Sbox_14_M4}), .b ({new_AGEMA_signal_5534, SubBytesIns_Inst_Sbox_14_M1}), .c ({new_AGEMA_signal_5719, SubBytesIns_Inst_Sbox_14_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M6_U1 ( .a ({new_AGEMA_signal_5115, SubBytesIns_Inst_Sbox_14_T3}), .b ({new_AGEMA_signal_5281, SubBytesIns_Inst_Sbox_14_T16}), .clk (clk), .r (Fresh[129]), .c ({new_AGEMA_signal_5536, SubBytesIns_Inst_Sbox_14_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M7_U1 ( .a ({new_AGEMA_signal_5283, SubBytesIns_Inst_Sbox_14_T22}), .b ({new_AGEMA_signal_5278, SubBytesIns_Inst_Sbox_14_T9}), .clk (clk), .r (Fresh[130]), .c ({new_AGEMA_signal_5537, SubBytesIns_Inst_Sbox_14_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M8_U1 ( .a ({new_AGEMA_signal_5533, SubBytesIns_Inst_Sbox_14_T26}), .b ({new_AGEMA_signal_5536, SubBytesIns_Inst_Sbox_14_M6}), .c ({new_AGEMA_signal_5720, SubBytesIns_Inst_Sbox_14_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M9_U1 ( .a ({new_AGEMA_signal_5531, SubBytesIns_Inst_Sbox_14_T20}), .b ({new_AGEMA_signal_5530, SubBytesIns_Inst_Sbox_14_T17}), .clk (clk), .r (Fresh[131]), .c ({new_AGEMA_signal_5721, SubBytesIns_Inst_Sbox_14_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M10_U1 ( .a ({new_AGEMA_signal_5721, SubBytesIns_Inst_Sbox_14_M9}), .b ({new_AGEMA_signal_5536, SubBytesIns_Inst_Sbox_14_M6}), .c ({new_AGEMA_signal_5823, SubBytesIns_Inst_Sbox_14_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M11_U1 ( .a ({new_AGEMA_signal_5113, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_5280, SubBytesIns_Inst_Sbox_14_T15}), .clk (clk), .r (Fresh[132]), .c ({new_AGEMA_signal_5538, SubBytesIns_Inst_Sbox_14_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M12_U1 ( .a ({new_AGEMA_signal_5116, SubBytesIns_Inst_Sbox_14_T4}), .b ({new_AGEMA_signal_5284, SubBytesIns_Inst_Sbox_14_T27}), .clk (clk), .r (Fresh[133]), .c ({new_AGEMA_signal_5539, SubBytesIns_Inst_Sbox_14_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M13_U1 ( .a ({new_AGEMA_signal_5539, SubBytesIns_Inst_Sbox_14_M12}), .b ({new_AGEMA_signal_5538, SubBytesIns_Inst_Sbox_14_M11}), .c ({new_AGEMA_signal_5722, SubBytesIns_Inst_Sbox_14_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M14_U1 ( .a ({new_AGEMA_signal_5114, SubBytesIns_Inst_Sbox_14_T2}), .b ({new_AGEMA_signal_5528, SubBytesIns_Inst_Sbox_14_T10}), .clk (clk), .r (Fresh[134]), .c ({new_AGEMA_signal_5723, SubBytesIns_Inst_Sbox_14_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M15_U1 ( .a ({new_AGEMA_signal_5723, SubBytesIns_Inst_Sbox_14_M14}), .b ({new_AGEMA_signal_5538, SubBytesIns_Inst_Sbox_14_M11}), .c ({new_AGEMA_signal_5824, SubBytesIns_Inst_Sbox_14_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M16_U1 ( .a ({new_AGEMA_signal_5718, SubBytesIns_Inst_Sbox_14_M3}), .b ({new_AGEMA_signal_5717, SubBytesIns_Inst_Sbox_14_M2}), .c ({new_AGEMA_signal_5825, SubBytesIns_Inst_Sbox_14_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M17_U1 ( .a ({new_AGEMA_signal_5719, SubBytesIns_Inst_Sbox_14_M5}), .b ({new_AGEMA_signal_5715, SubBytesIns_Inst_Sbox_14_T24}), .c ({new_AGEMA_signal_5826, SubBytesIns_Inst_Sbox_14_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M18_U1 ( .a ({new_AGEMA_signal_5720, SubBytesIns_Inst_Sbox_14_M8}), .b ({new_AGEMA_signal_5537, SubBytesIns_Inst_Sbox_14_M7}), .c ({new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_14_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M19_U1 ( .a ({new_AGEMA_signal_5823, SubBytesIns_Inst_Sbox_14_M10}), .b ({new_AGEMA_signal_5824, SubBytesIns_Inst_Sbox_14_M15}), .c ({new_AGEMA_signal_5905, SubBytesIns_Inst_Sbox_14_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M20_U1 ( .a ({new_AGEMA_signal_5825, SubBytesIns_Inst_Sbox_14_M16}), .b ({new_AGEMA_signal_5722, SubBytesIns_Inst_Sbox_14_M13}), .c ({new_AGEMA_signal_5906, SubBytesIns_Inst_Sbox_14_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M21_U1 ( .a ({new_AGEMA_signal_5826, SubBytesIns_Inst_Sbox_14_M17}), .b ({new_AGEMA_signal_5824, SubBytesIns_Inst_Sbox_14_M15}), .c ({new_AGEMA_signal_5907, SubBytesIns_Inst_Sbox_14_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M22_U1 ( .a ({new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_14_M18}), .b ({new_AGEMA_signal_5722, SubBytesIns_Inst_Sbox_14_M13}), .c ({new_AGEMA_signal_5908, SubBytesIns_Inst_Sbox_14_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M23_U1 ( .a ({new_AGEMA_signal_5905, SubBytesIns_Inst_Sbox_14_M19}), .b ({new_AGEMA_signal_5716, SubBytesIns_Inst_Sbox_14_T25}), .c ({new_AGEMA_signal_5985, SubBytesIns_Inst_Sbox_14_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M24_U1 ( .a ({new_AGEMA_signal_5908, SubBytesIns_Inst_Sbox_14_M22}), .b ({new_AGEMA_signal_5985, SubBytesIns_Inst_Sbox_14_M23}), .c ({new_AGEMA_signal_6083, SubBytesIns_Inst_Sbox_14_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M27_U1 ( .a ({new_AGEMA_signal_5906, SubBytesIns_Inst_Sbox_14_M20}), .b ({new_AGEMA_signal_5907, SubBytesIns_Inst_Sbox_14_M21}), .c ({new_AGEMA_signal_5987, SubBytesIns_Inst_Sbox_14_M27}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M1_U1 ( .a ({new_AGEMA_signal_5287, SubBytesIns_Inst_Sbox_15_T13}), .b ({new_AGEMA_signal_5285, SubBytesIns_Inst_Sbox_15_T6}), .clk (clk), .r (Fresh[135]), .c ({new_AGEMA_signal_5547, SubBytesIns_Inst_Sbox_15_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M2_U1 ( .a ({new_AGEMA_signal_5545, SubBytesIns_Inst_Sbox_15_T23}), .b ({new_AGEMA_signal_5540, SubBytesIns_Inst_Sbox_15_T8}), .clk (clk), .r (Fresh[136]), .c ({new_AGEMA_signal_5726, SubBytesIns_Inst_Sbox_15_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M3_U1 ( .a ({new_AGEMA_signal_5542, SubBytesIns_Inst_Sbox_15_T14}), .b ({new_AGEMA_signal_5547, SubBytesIns_Inst_Sbox_15_M1}), .c ({new_AGEMA_signal_5727, SubBytesIns_Inst_Sbox_15_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M4_U1 ( .a ({new_AGEMA_signal_5290, SubBytesIns_Inst_Sbox_15_T19}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .clk (clk), .r (Fresh[137]), .c ({new_AGEMA_signal_5548, SubBytesIns_Inst_Sbox_15_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M5_U1 ( .a ({new_AGEMA_signal_5548, SubBytesIns_Inst_Sbox_15_M4}), .b ({new_AGEMA_signal_5547, SubBytesIns_Inst_Sbox_15_M1}), .c ({new_AGEMA_signal_5728, SubBytesIns_Inst_Sbox_15_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M6_U1 ( .a ({new_AGEMA_signal_5125, SubBytesIns_Inst_Sbox_15_T3}), .b ({new_AGEMA_signal_5289, SubBytesIns_Inst_Sbox_15_T16}), .clk (clk), .r (Fresh[138]), .c ({new_AGEMA_signal_5549, SubBytesIns_Inst_Sbox_15_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M7_U1 ( .a ({new_AGEMA_signal_5291, SubBytesIns_Inst_Sbox_15_T22}), .b ({new_AGEMA_signal_5286, SubBytesIns_Inst_Sbox_15_T9}), .clk (clk), .r (Fresh[139]), .c ({new_AGEMA_signal_5550, SubBytesIns_Inst_Sbox_15_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M8_U1 ( .a ({new_AGEMA_signal_5546, SubBytesIns_Inst_Sbox_15_T26}), .b ({new_AGEMA_signal_5549, SubBytesIns_Inst_Sbox_15_M6}), .c ({new_AGEMA_signal_5729, SubBytesIns_Inst_Sbox_15_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M9_U1 ( .a ({new_AGEMA_signal_5544, SubBytesIns_Inst_Sbox_15_T20}), .b ({new_AGEMA_signal_5543, SubBytesIns_Inst_Sbox_15_T17}), .clk (clk), .r (Fresh[140]), .c ({new_AGEMA_signal_5730, SubBytesIns_Inst_Sbox_15_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M10_U1 ( .a ({new_AGEMA_signal_5730, SubBytesIns_Inst_Sbox_15_M9}), .b ({new_AGEMA_signal_5549, SubBytesIns_Inst_Sbox_15_M6}), .c ({new_AGEMA_signal_5828, SubBytesIns_Inst_Sbox_15_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M11_U1 ( .a ({new_AGEMA_signal_5123, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_5288, SubBytesIns_Inst_Sbox_15_T15}), .clk (clk), .r (Fresh[141]), .c ({new_AGEMA_signal_5551, SubBytesIns_Inst_Sbox_15_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M12_U1 ( .a ({new_AGEMA_signal_5126, SubBytesIns_Inst_Sbox_15_T4}), .b ({new_AGEMA_signal_5292, SubBytesIns_Inst_Sbox_15_T27}), .clk (clk), .r (Fresh[142]), .c ({new_AGEMA_signal_5552, SubBytesIns_Inst_Sbox_15_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M13_U1 ( .a ({new_AGEMA_signal_5552, SubBytesIns_Inst_Sbox_15_M12}), .b ({new_AGEMA_signal_5551, SubBytesIns_Inst_Sbox_15_M11}), .c ({new_AGEMA_signal_5731, SubBytesIns_Inst_Sbox_15_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M14_U1 ( .a ({new_AGEMA_signal_5124, SubBytesIns_Inst_Sbox_15_T2}), .b ({new_AGEMA_signal_5541, SubBytesIns_Inst_Sbox_15_T10}), .clk (clk), .r (Fresh[143]), .c ({new_AGEMA_signal_5732, SubBytesIns_Inst_Sbox_15_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M15_U1 ( .a ({new_AGEMA_signal_5732, SubBytesIns_Inst_Sbox_15_M14}), .b ({new_AGEMA_signal_5551, SubBytesIns_Inst_Sbox_15_M11}), .c ({new_AGEMA_signal_5829, SubBytesIns_Inst_Sbox_15_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M16_U1 ( .a ({new_AGEMA_signal_5727, SubBytesIns_Inst_Sbox_15_M3}), .b ({new_AGEMA_signal_5726, SubBytesIns_Inst_Sbox_15_M2}), .c ({new_AGEMA_signal_5830, SubBytesIns_Inst_Sbox_15_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M17_U1 ( .a ({new_AGEMA_signal_5728, SubBytesIns_Inst_Sbox_15_M5}), .b ({new_AGEMA_signal_5724, SubBytesIns_Inst_Sbox_15_T24}), .c ({new_AGEMA_signal_5831, SubBytesIns_Inst_Sbox_15_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M18_U1 ( .a ({new_AGEMA_signal_5729, SubBytesIns_Inst_Sbox_15_M8}), .b ({new_AGEMA_signal_5550, SubBytesIns_Inst_Sbox_15_M7}), .c ({new_AGEMA_signal_5832, SubBytesIns_Inst_Sbox_15_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M19_U1 ( .a ({new_AGEMA_signal_5828, SubBytesIns_Inst_Sbox_15_M10}), .b ({new_AGEMA_signal_5829, SubBytesIns_Inst_Sbox_15_M15}), .c ({new_AGEMA_signal_5909, SubBytesIns_Inst_Sbox_15_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M20_U1 ( .a ({new_AGEMA_signal_5830, SubBytesIns_Inst_Sbox_15_M16}), .b ({new_AGEMA_signal_5731, SubBytesIns_Inst_Sbox_15_M13}), .c ({new_AGEMA_signal_5910, SubBytesIns_Inst_Sbox_15_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M21_U1 ( .a ({new_AGEMA_signal_5831, SubBytesIns_Inst_Sbox_15_M17}), .b ({new_AGEMA_signal_5829, SubBytesIns_Inst_Sbox_15_M15}), .c ({new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_15_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M22_U1 ( .a ({new_AGEMA_signal_5832, SubBytesIns_Inst_Sbox_15_M18}), .b ({new_AGEMA_signal_5731, SubBytesIns_Inst_Sbox_15_M13}), .c ({new_AGEMA_signal_5912, SubBytesIns_Inst_Sbox_15_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M23_U1 ( .a ({new_AGEMA_signal_5909, SubBytesIns_Inst_Sbox_15_M19}), .b ({new_AGEMA_signal_5725, SubBytesIns_Inst_Sbox_15_T25}), .c ({new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_15_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M24_U1 ( .a ({new_AGEMA_signal_5912, SubBytesIns_Inst_Sbox_15_M22}), .b ({new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_15_M23}), .c ({new_AGEMA_signal_6088, SubBytesIns_Inst_Sbox_15_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M27_U1 ( .a ({new_AGEMA_signal_5910, SubBytesIns_Inst_Sbox_15_M20}), .b ({new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_15_M21}), .c ({new_AGEMA_signal_5991, SubBytesIns_Inst_Sbox_15_M27}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M1_U1 ( .a ({new_AGEMA_signal_5135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13}), .b ({new_AGEMA_signal_5133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .clk (clk), .r (Fresh[144]), .c ({new_AGEMA_signal_5300, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M2_U1 ( .a ({new_AGEMA_signal_5298, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23}), .b ({new_AGEMA_signal_5293, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8}), .clk (clk), .r (Fresh[145]), .c ({new_AGEMA_signal_5555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M3_U1 ( .a ({new_AGEMA_signal_5295, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14}), .b ({new_AGEMA_signal_5300, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_5556, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M4_U1 ( .a ({new_AGEMA_signal_5138, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}), .b ({new_AGEMA_signal_4655, RoundKey[16]}), .clk (clk), .r (Fresh[146]), .c ({new_AGEMA_signal_5301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M5_U1 ( .a ({new_AGEMA_signal_5301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4}), .b ({new_AGEMA_signal_5300, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_5557, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M6_U1 ( .a ({new_AGEMA_signal_4935, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .clk (clk), .r (Fresh[147]), .c ({new_AGEMA_signal_5302, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M7_U1 ( .a ({new_AGEMA_signal_5139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}), .b ({new_AGEMA_signal_5134, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}), .clk (clk), .r (Fresh[148]), .c ({new_AGEMA_signal_5303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M8_U1 ( .a ({new_AGEMA_signal_5299, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26}), .b ({new_AGEMA_signal_5302, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_5558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M9_U1 ( .a ({new_AGEMA_signal_5297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_5296, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}), .clk (clk), .r (Fresh[149]), .c ({new_AGEMA_signal_5559, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M10_U1 ( .a ({new_AGEMA_signal_5559, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9}), .b ({new_AGEMA_signal_5302, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_5733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M11_U1 ( .a ({new_AGEMA_signal_4933, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5136, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15}), .clk (clk), .r (Fresh[150]), .c ({new_AGEMA_signal_5304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M12_U1 ( .a ({new_AGEMA_signal_4936, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}), .b ({new_AGEMA_signal_5140, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27}), .clk (clk), .r (Fresh[151]), .c ({new_AGEMA_signal_5305, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M13_U1 ( .a ({new_AGEMA_signal_5305, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12}), .b ({new_AGEMA_signal_5304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_5560, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M14_U1 ( .a ({new_AGEMA_signal_4934, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_5294, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}), .clk (clk), .r (Fresh[152]), .c ({new_AGEMA_signal_5561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M15_U1 ( .a ({new_AGEMA_signal_5561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14}), .b ({new_AGEMA_signal_5304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_5734, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M16_U1 ( .a ({new_AGEMA_signal_5556, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3}), .b ({new_AGEMA_signal_5555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2}), .c ({new_AGEMA_signal_5735, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M17_U1 ( .a ({new_AGEMA_signal_5557, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5}), .b ({new_AGEMA_signal_5553, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24}), .c ({new_AGEMA_signal_5736, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M18_U1 ( .a ({new_AGEMA_signal_5558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8}), .b ({new_AGEMA_signal_5303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7}), .c ({new_AGEMA_signal_5737, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M19_U1 ( .a ({new_AGEMA_signal_5733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10}), .b ({new_AGEMA_signal_5734, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_5833, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M20_U1 ( .a ({new_AGEMA_signal_5735, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16}), .b ({new_AGEMA_signal_5560, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_5834, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M21_U1 ( .a ({new_AGEMA_signal_5736, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17}), .b ({new_AGEMA_signal_5734, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_5835, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M22_U1 ( .a ({new_AGEMA_signal_5737, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18}), .b ({new_AGEMA_signal_5560, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_5836, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M23_U1 ( .a ({new_AGEMA_signal_5833, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19}), .b ({new_AGEMA_signal_5554, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25}), .c ({new_AGEMA_signal_5913, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M24_U1 ( .a ({new_AGEMA_signal_5836, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_5913, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}), .c ({new_AGEMA_signal_5993, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M27_U1 ( .a ({new_AGEMA_signal_5834, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_5835, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}), .c ({new_AGEMA_signal_5915, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M1_U1 ( .a ({new_AGEMA_signal_5143, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13}), .b ({new_AGEMA_signal_5141, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .clk (clk), .r (Fresh[153]), .c ({new_AGEMA_signal_5313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M2_U1 ( .a ({new_AGEMA_signal_5311, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23}), .b ({new_AGEMA_signal_5306, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8}), .clk (clk), .r (Fresh[154]), .c ({new_AGEMA_signal_5564, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M3_U1 ( .a ({new_AGEMA_signal_5308, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14}), .b ({new_AGEMA_signal_5313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_5565, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M4_U1 ( .a ({new_AGEMA_signal_5146, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}), .b ({new_AGEMA_signal_4898, RoundKey[8]}), .clk (clk), .r (Fresh[155]), .c ({new_AGEMA_signal_5314, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M5_U1 ( .a ({new_AGEMA_signal_5314, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4}), .b ({new_AGEMA_signal_5313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_5566, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M6_U1 ( .a ({new_AGEMA_signal_4945, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .clk (clk), .r (Fresh[156]), .c ({new_AGEMA_signal_5315, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M7_U1 ( .a ({new_AGEMA_signal_5147, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}), .b ({new_AGEMA_signal_5142, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}), .clk (clk), .r (Fresh[157]), .c ({new_AGEMA_signal_5316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M8_U1 ( .a ({new_AGEMA_signal_5312, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26}), .b ({new_AGEMA_signal_5315, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_5567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M9_U1 ( .a ({new_AGEMA_signal_5310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_5309, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}), .clk (clk), .r (Fresh[158]), .c ({new_AGEMA_signal_5568, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M10_U1 ( .a ({new_AGEMA_signal_5568, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9}), .b ({new_AGEMA_signal_5315, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_5738, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M11_U1 ( .a ({new_AGEMA_signal_4943, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5144, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15}), .clk (clk), .r (Fresh[159]), .c ({new_AGEMA_signal_5317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M12_U1 ( .a ({new_AGEMA_signal_4946, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}), .b ({new_AGEMA_signal_5148, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27}), .clk (clk), .r (Fresh[160]), .c ({new_AGEMA_signal_5318, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M13_U1 ( .a ({new_AGEMA_signal_5318, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12}), .b ({new_AGEMA_signal_5317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_5569, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M14_U1 ( .a ({new_AGEMA_signal_4944, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_5307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}), .clk (clk), .r (Fresh[161]), .c ({new_AGEMA_signal_5570, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M15_U1 ( .a ({new_AGEMA_signal_5570, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14}), .b ({new_AGEMA_signal_5317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_5739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M16_U1 ( .a ({new_AGEMA_signal_5565, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3}), .b ({new_AGEMA_signal_5564, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2}), .c ({new_AGEMA_signal_5740, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M17_U1 ( .a ({new_AGEMA_signal_5566, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5}), .b ({new_AGEMA_signal_5562, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24}), .c ({new_AGEMA_signal_5741, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M18_U1 ( .a ({new_AGEMA_signal_5567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8}), .b ({new_AGEMA_signal_5316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7}), .c ({new_AGEMA_signal_5742, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M19_U1 ( .a ({new_AGEMA_signal_5738, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10}), .b ({new_AGEMA_signal_5739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_5837, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M20_U1 ( .a ({new_AGEMA_signal_5740, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16}), .b ({new_AGEMA_signal_5569, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_5838, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M21_U1 ( .a ({new_AGEMA_signal_5741, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17}), .b ({new_AGEMA_signal_5739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_5839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M22_U1 ( .a ({new_AGEMA_signal_5742, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18}), .b ({new_AGEMA_signal_5569, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_5840, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M23_U1 ( .a ({new_AGEMA_signal_5837, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19}), .b ({new_AGEMA_signal_5563, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25}), .c ({new_AGEMA_signal_5917, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M24_U1 ( .a ({new_AGEMA_signal_5840, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_5917, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}), .c ({new_AGEMA_signal_5998, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M27_U1 ( .a ({new_AGEMA_signal_5838, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_5839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}), .c ({new_AGEMA_signal_5919, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M1_U1 ( .a ({new_AGEMA_signal_5151, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13}), .b ({new_AGEMA_signal_5149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .clk (clk), .r (Fresh[162]), .c ({new_AGEMA_signal_5326, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M2_U1 ( .a ({new_AGEMA_signal_5324, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23}), .b ({new_AGEMA_signal_5319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8}), .clk (clk), .r (Fresh[163]), .c ({new_AGEMA_signal_5573, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M3_U1 ( .a ({new_AGEMA_signal_5321, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14}), .b ({new_AGEMA_signal_5326, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_5574, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M4_U1 ( .a ({new_AGEMA_signal_5154, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}), .b ({new_AGEMA_signal_4550, RoundKey[0]}), .clk (clk), .r (Fresh[164]), .c ({new_AGEMA_signal_5327, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M5_U1 ( .a ({new_AGEMA_signal_5327, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4}), .b ({new_AGEMA_signal_5326, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_5575, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M6_U1 ( .a ({new_AGEMA_signal_4955, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5153, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .clk (clk), .r (Fresh[165]), .c ({new_AGEMA_signal_5328, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M7_U1 ( .a ({new_AGEMA_signal_5155, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}), .b ({new_AGEMA_signal_5150, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}), .clk (clk), .r (Fresh[166]), .c ({new_AGEMA_signal_5329, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M8_U1 ( .a ({new_AGEMA_signal_5325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26}), .b ({new_AGEMA_signal_5328, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_5576, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M9_U1 ( .a ({new_AGEMA_signal_5323, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_5322, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}), .clk (clk), .r (Fresh[167]), .c ({new_AGEMA_signal_5577, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M10_U1 ( .a ({new_AGEMA_signal_5577, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9}), .b ({new_AGEMA_signal_5328, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_5743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M11_U1 ( .a ({new_AGEMA_signal_4953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5152, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15}), .clk (clk), .r (Fresh[168]), .c ({new_AGEMA_signal_5330, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M12_U1 ( .a ({new_AGEMA_signal_4956, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}), .b ({new_AGEMA_signal_5156, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27}), .clk (clk), .r (Fresh[169]), .c ({new_AGEMA_signal_5331, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M13_U1 ( .a ({new_AGEMA_signal_5331, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12}), .b ({new_AGEMA_signal_5330, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_5578, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M14_U1 ( .a ({new_AGEMA_signal_4954, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_5320, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}), .clk (clk), .r (Fresh[170]), .c ({new_AGEMA_signal_5579, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M15_U1 ( .a ({new_AGEMA_signal_5579, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14}), .b ({new_AGEMA_signal_5330, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_5744, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M16_U1 ( .a ({new_AGEMA_signal_5574, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3}), .b ({new_AGEMA_signal_5573, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2}), .c ({new_AGEMA_signal_5745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M17_U1 ( .a ({new_AGEMA_signal_5575, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5}), .b ({new_AGEMA_signal_5571, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24}), .c ({new_AGEMA_signal_5746, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M18_U1 ( .a ({new_AGEMA_signal_5576, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8}), .b ({new_AGEMA_signal_5329, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7}), .c ({new_AGEMA_signal_5747, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M19_U1 ( .a ({new_AGEMA_signal_5743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10}), .b ({new_AGEMA_signal_5744, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_5841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M20_U1 ( .a ({new_AGEMA_signal_5745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16}), .b ({new_AGEMA_signal_5578, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_5842, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M21_U1 ( .a ({new_AGEMA_signal_5746, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17}), .b ({new_AGEMA_signal_5744, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_5843, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M22_U1 ( .a ({new_AGEMA_signal_5747, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18}), .b ({new_AGEMA_signal_5578, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_5844, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M23_U1 ( .a ({new_AGEMA_signal_5841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19}), .b ({new_AGEMA_signal_5572, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25}), .c ({new_AGEMA_signal_5921, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M24_U1 ( .a ({new_AGEMA_signal_5844, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_5921, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}), .c ({new_AGEMA_signal_6003, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M27_U1 ( .a ({new_AGEMA_signal_5842, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_5843, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}), .c ({new_AGEMA_signal_5923, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M1_U1 ( .a ({new_AGEMA_signal_5159, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13}), .b ({new_AGEMA_signal_5157, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .clk (clk), .r (Fresh[171]), .c ({new_AGEMA_signal_5339, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M2_U1 ( .a ({new_AGEMA_signal_5337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23}), .b ({new_AGEMA_signal_5332, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8}), .clk (clk), .r (Fresh[172]), .c ({new_AGEMA_signal_5582, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M3_U1 ( .a ({new_AGEMA_signal_5334, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14}), .b ({new_AGEMA_signal_5339, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_5583, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M4_U1 ( .a ({new_AGEMA_signal_5162, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}), .b ({new_AGEMA_signal_4682, RoundKey[24]}), .clk (clk), .r (Fresh[173]), .c ({new_AGEMA_signal_5340, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M5_U1 ( .a ({new_AGEMA_signal_5340, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4}), .b ({new_AGEMA_signal_5339, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_5584, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M6_U1 ( .a ({new_AGEMA_signal_4965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5161, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .clk (clk), .r (Fresh[174]), .c ({new_AGEMA_signal_5341, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M7_U1 ( .a ({new_AGEMA_signal_5163, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}), .b ({new_AGEMA_signal_5158, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}), .clk (clk), .r (Fresh[175]), .c ({new_AGEMA_signal_5342, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M8_U1 ( .a ({new_AGEMA_signal_5338, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26}), .b ({new_AGEMA_signal_5341, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_5585, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M9_U1 ( .a ({new_AGEMA_signal_5336, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_5335, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}), .clk (clk), .r (Fresh[176]), .c ({new_AGEMA_signal_5586, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M10_U1 ( .a ({new_AGEMA_signal_5586, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9}), .b ({new_AGEMA_signal_5341, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_5748, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M11_U1 ( .a ({new_AGEMA_signal_4963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5160, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15}), .clk (clk), .r (Fresh[177]), .c ({new_AGEMA_signal_5343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M12_U1 ( .a ({new_AGEMA_signal_4966, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}), .b ({new_AGEMA_signal_5164, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27}), .clk (clk), .r (Fresh[178]), .c ({new_AGEMA_signal_5344, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M13_U1 ( .a ({new_AGEMA_signal_5344, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12}), .b ({new_AGEMA_signal_5343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_5587, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M14_U1 ( .a ({new_AGEMA_signal_4964, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_5333, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}), .clk (clk), .r (Fresh[179]), .c ({new_AGEMA_signal_5588, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M15_U1 ( .a ({new_AGEMA_signal_5588, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14}), .b ({new_AGEMA_signal_5343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M16_U1 ( .a ({new_AGEMA_signal_5583, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3}), .b ({new_AGEMA_signal_5582, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2}), .c ({new_AGEMA_signal_5750, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M17_U1 ( .a ({new_AGEMA_signal_5584, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5}), .b ({new_AGEMA_signal_5580, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24}), .c ({new_AGEMA_signal_5751, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M18_U1 ( .a ({new_AGEMA_signal_5585, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8}), .b ({new_AGEMA_signal_5342, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7}), .c ({new_AGEMA_signal_5752, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M19_U1 ( .a ({new_AGEMA_signal_5748, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10}), .b ({new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_5845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M20_U1 ( .a ({new_AGEMA_signal_5750, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16}), .b ({new_AGEMA_signal_5587, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_5846, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M21_U1 ( .a ({new_AGEMA_signal_5751, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17}), .b ({new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_5847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M22_U1 ( .a ({new_AGEMA_signal_5752, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18}), .b ({new_AGEMA_signal_5587, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_5848, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M23_U1 ( .a ({new_AGEMA_signal_5845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19}), .b ({new_AGEMA_signal_5581, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25}), .c ({new_AGEMA_signal_5925, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M24_U1 ( .a ({new_AGEMA_signal_5848, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_5925, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}), .c ({new_AGEMA_signal_6008, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M27_U1 ( .a ({new_AGEMA_signal_5846, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_5847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}), .c ({new_AGEMA_signal_5927, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M25_U1 ( .a ({new_AGEMA_signal_5852, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_5850, SubBytesIns_Inst_Sbox_0_M20}), .clk (clk), .r (Fresh[180]), .c ({new_AGEMA_signal_5930, SubBytesIns_Inst_Sbox_0_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M26_U1 ( .a ({new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_5930, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_6014, SubBytesIns_Inst_Sbox_0_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M28_U1 ( .a ({new_AGEMA_signal_5929, SubBytesIns_Inst_Sbox_0_M23}), .b ({new_AGEMA_signal_5930, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_6015, SubBytesIns_Inst_Sbox_0_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M31_U1 ( .a ({new_AGEMA_signal_5850, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_5929, SubBytesIns_Inst_Sbox_0_M23}), .clk (clk), .r (Fresh[181]), .c ({new_AGEMA_signal_6016, SubBytesIns_Inst_Sbox_0_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M33_U1 ( .a ({new_AGEMA_signal_5931, SubBytesIns_Inst_Sbox_0_M27}), .b ({new_AGEMA_signal_5930, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_6017, SubBytesIns_Inst_Sbox_0_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M34_U1 ( .a ({new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_5852, SubBytesIns_Inst_Sbox_0_M22}), .clk (clk), .r (Fresh[182]), .c ({new_AGEMA_signal_5932, SubBytesIns_Inst_Sbox_0_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M36_U1 ( .a ({new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_0_M24}), .b ({new_AGEMA_signal_5930, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_6117, SubBytesIns_Inst_Sbox_0_M36}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M25_U1 ( .a ({new_AGEMA_signal_5856, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_5854, SubBytesIns_Inst_Sbox_1_M20}), .clk (clk), .r (Fresh[183]), .c ({new_AGEMA_signal_5934, SubBytesIns_Inst_Sbox_1_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M26_U1 ( .a ({new_AGEMA_signal_5855, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_5934, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_6019, SubBytesIns_Inst_Sbox_1_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M28_U1 ( .a ({new_AGEMA_signal_5933, SubBytesIns_Inst_Sbox_1_M23}), .b ({new_AGEMA_signal_5934, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_6020, SubBytesIns_Inst_Sbox_1_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M31_U1 ( .a ({new_AGEMA_signal_5854, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_5933, SubBytesIns_Inst_Sbox_1_M23}), .clk (clk), .r (Fresh[184]), .c ({new_AGEMA_signal_6021, SubBytesIns_Inst_Sbox_1_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M33_U1 ( .a ({new_AGEMA_signal_5935, SubBytesIns_Inst_Sbox_1_M27}), .b ({new_AGEMA_signal_5934, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_6022, SubBytesIns_Inst_Sbox_1_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M34_U1 ( .a ({new_AGEMA_signal_5855, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_5856, SubBytesIns_Inst_Sbox_1_M22}), .clk (clk), .r (Fresh[185]), .c ({new_AGEMA_signal_5936, SubBytesIns_Inst_Sbox_1_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M36_U1 ( .a ({new_AGEMA_signal_6018, SubBytesIns_Inst_Sbox_1_M24}), .b ({new_AGEMA_signal_5934, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_6122, SubBytesIns_Inst_Sbox_1_M36}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M25_U1 ( .a ({new_AGEMA_signal_5860, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_5858, SubBytesIns_Inst_Sbox_2_M20}), .clk (clk), .r (Fresh[186]), .c ({new_AGEMA_signal_5938, SubBytesIns_Inst_Sbox_2_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M26_U1 ( .a ({new_AGEMA_signal_5859, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_5938, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_6024, SubBytesIns_Inst_Sbox_2_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M28_U1 ( .a ({new_AGEMA_signal_5937, SubBytesIns_Inst_Sbox_2_M23}), .b ({new_AGEMA_signal_5938, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_6025, SubBytesIns_Inst_Sbox_2_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M31_U1 ( .a ({new_AGEMA_signal_5858, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_5937, SubBytesIns_Inst_Sbox_2_M23}), .clk (clk), .r (Fresh[187]), .c ({new_AGEMA_signal_6026, SubBytesIns_Inst_Sbox_2_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M33_U1 ( .a ({new_AGEMA_signal_5939, SubBytesIns_Inst_Sbox_2_M27}), .b ({new_AGEMA_signal_5938, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_6027, SubBytesIns_Inst_Sbox_2_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M34_U1 ( .a ({new_AGEMA_signal_5859, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_5860, SubBytesIns_Inst_Sbox_2_M22}), .clk (clk), .r (Fresh[188]), .c ({new_AGEMA_signal_5940, SubBytesIns_Inst_Sbox_2_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M36_U1 ( .a ({new_AGEMA_signal_6023, SubBytesIns_Inst_Sbox_2_M24}), .b ({new_AGEMA_signal_5938, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_6127, SubBytesIns_Inst_Sbox_2_M36}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M25_U1 ( .a ({new_AGEMA_signal_5864, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_5862, SubBytesIns_Inst_Sbox_3_M20}), .clk (clk), .r (Fresh[189]), .c ({new_AGEMA_signal_5942, SubBytesIns_Inst_Sbox_3_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M26_U1 ( .a ({new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_5942, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_6029, SubBytesIns_Inst_Sbox_3_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M28_U1 ( .a ({new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_3_M23}), .b ({new_AGEMA_signal_5942, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_6030, SubBytesIns_Inst_Sbox_3_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M31_U1 ( .a ({new_AGEMA_signal_5862, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_3_M23}), .clk (clk), .r (Fresh[190]), .c ({new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_3_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M33_U1 ( .a ({new_AGEMA_signal_5943, SubBytesIns_Inst_Sbox_3_M27}), .b ({new_AGEMA_signal_5942, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_6032, SubBytesIns_Inst_Sbox_3_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M34_U1 ( .a ({new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_5864, SubBytesIns_Inst_Sbox_3_M22}), .clk (clk), .r (Fresh[191]), .c ({new_AGEMA_signal_5944, SubBytesIns_Inst_Sbox_3_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M36_U1 ( .a ({new_AGEMA_signal_6028, SubBytesIns_Inst_Sbox_3_M24}), .b ({new_AGEMA_signal_5942, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_6132, SubBytesIns_Inst_Sbox_3_M36}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M25_U1 ( .a ({new_AGEMA_signal_5868, SubBytesIns_Inst_Sbox_4_M22}), .b ({new_AGEMA_signal_5866, SubBytesIns_Inst_Sbox_4_M20}), .clk (clk), .r (Fresh[192]), .c ({new_AGEMA_signal_5946, SubBytesIns_Inst_Sbox_4_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M26_U1 ( .a ({new_AGEMA_signal_5867, SubBytesIns_Inst_Sbox_4_M21}), .b ({new_AGEMA_signal_5946, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_6034, SubBytesIns_Inst_Sbox_4_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M28_U1 ( .a ({new_AGEMA_signal_5945, SubBytesIns_Inst_Sbox_4_M23}), .b ({new_AGEMA_signal_5946, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_6035, SubBytesIns_Inst_Sbox_4_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M31_U1 ( .a ({new_AGEMA_signal_5866, SubBytesIns_Inst_Sbox_4_M20}), .b ({new_AGEMA_signal_5945, SubBytesIns_Inst_Sbox_4_M23}), .clk (clk), .r (Fresh[193]), .c ({new_AGEMA_signal_6036, SubBytesIns_Inst_Sbox_4_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M33_U1 ( .a ({new_AGEMA_signal_5947, SubBytesIns_Inst_Sbox_4_M27}), .b ({new_AGEMA_signal_5946, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_6037, SubBytesIns_Inst_Sbox_4_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M34_U1 ( .a ({new_AGEMA_signal_5867, SubBytesIns_Inst_Sbox_4_M21}), .b ({new_AGEMA_signal_5868, SubBytesIns_Inst_Sbox_4_M22}), .clk (clk), .r (Fresh[194]), .c ({new_AGEMA_signal_5948, SubBytesIns_Inst_Sbox_4_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M36_U1 ( .a ({new_AGEMA_signal_6033, SubBytesIns_Inst_Sbox_4_M24}), .b ({new_AGEMA_signal_5946, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_6137, SubBytesIns_Inst_Sbox_4_M36}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M25_U1 ( .a ({new_AGEMA_signal_5872, SubBytesIns_Inst_Sbox_5_M22}), .b ({new_AGEMA_signal_5870, SubBytesIns_Inst_Sbox_5_M20}), .clk (clk), .r (Fresh[195]), .c ({new_AGEMA_signal_5950, SubBytesIns_Inst_Sbox_5_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M26_U1 ( .a ({new_AGEMA_signal_5871, SubBytesIns_Inst_Sbox_5_M21}), .b ({new_AGEMA_signal_5950, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_6039, SubBytesIns_Inst_Sbox_5_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M28_U1 ( .a ({new_AGEMA_signal_5949, SubBytesIns_Inst_Sbox_5_M23}), .b ({new_AGEMA_signal_5950, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_6040, SubBytesIns_Inst_Sbox_5_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M31_U1 ( .a ({new_AGEMA_signal_5870, SubBytesIns_Inst_Sbox_5_M20}), .b ({new_AGEMA_signal_5949, SubBytesIns_Inst_Sbox_5_M23}), .clk (clk), .r (Fresh[196]), .c ({new_AGEMA_signal_6041, SubBytesIns_Inst_Sbox_5_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M33_U1 ( .a ({new_AGEMA_signal_5951, SubBytesIns_Inst_Sbox_5_M27}), .b ({new_AGEMA_signal_5950, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_6042, SubBytesIns_Inst_Sbox_5_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M34_U1 ( .a ({new_AGEMA_signal_5871, SubBytesIns_Inst_Sbox_5_M21}), .b ({new_AGEMA_signal_5872, SubBytesIns_Inst_Sbox_5_M22}), .clk (clk), .r (Fresh[197]), .c ({new_AGEMA_signal_5952, SubBytesIns_Inst_Sbox_5_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M36_U1 ( .a ({new_AGEMA_signal_6038, SubBytesIns_Inst_Sbox_5_M24}), .b ({new_AGEMA_signal_5950, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_6142, SubBytesIns_Inst_Sbox_5_M36}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M25_U1 ( .a ({new_AGEMA_signal_5876, SubBytesIns_Inst_Sbox_6_M22}), .b ({new_AGEMA_signal_5874, SubBytesIns_Inst_Sbox_6_M20}), .clk (clk), .r (Fresh[198]), .c ({new_AGEMA_signal_5954, SubBytesIns_Inst_Sbox_6_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M26_U1 ( .a ({new_AGEMA_signal_5875, SubBytesIns_Inst_Sbox_6_M21}), .b ({new_AGEMA_signal_5954, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_6044, SubBytesIns_Inst_Sbox_6_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M28_U1 ( .a ({new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_6_M23}), .b ({new_AGEMA_signal_5954, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_6045, SubBytesIns_Inst_Sbox_6_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M31_U1 ( .a ({new_AGEMA_signal_5874, SubBytesIns_Inst_Sbox_6_M20}), .b ({new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_6_M23}), .clk (clk), .r (Fresh[199]), .c ({new_AGEMA_signal_6046, SubBytesIns_Inst_Sbox_6_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M33_U1 ( .a ({new_AGEMA_signal_5955, SubBytesIns_Inst_Sbox_6_M27}), .b ({new_AGEMA_signal_5954, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_6047, SubBytesIns_Inst_Sbox_6_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M34_U1 ( .a ({new_AGEMA_signal_5875, SubBytesIns_Inst_Sbox_6_M21}), .b ({new_AGEMA_signal_5876, SubBytesIns_Inst_Sbox_6_M22}), .clk (clk), .r (Fresh[200]), .c ({new_AGEMA_signal_5956, SubBytesIns_Inst_Sbox_6_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M36_U1 ( .a ({new_AGEMA_signal_6043, SubBytesIns_Inst_Sbox_6_M24}), .b ({new_AGEMA_signal_5954, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_6147, SubBytesIns_Inst_Sbox_6_M36}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M25_U1 ( .a ({new_AGEMA_signal_5880, SubBytesIns_Inst_Sbox_7_M22}), .b ({new_AGEMA_signal_5878, SubBytesIns_Inst_Sbox_7_M20}), .clk (clk), .r (Fresh[201]), .c ({new_AGEMA_signal_5958, SubBytesIns_Inst_Sbox_7_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M26_U1 ( .a ({new_AGEMA_signal_5879, SubBytesIns_Inst_Sbox_7_M21}), .b ({new_AGEMA_signal_5958, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_6049, SubBytesIns_Inst_Sbox_7_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M28_U1 ( .a ({new_AGEMA_signal_5957, SubBytesIns_Inst_Sbox_7_M23}), .b ({new_AGEMA_signal_5958, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_6050, SubBytesIns_Inst_Sbox_7_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M31_U1 ( .a ({new_AGEMA_signal_5878, SubBytesIns_Inst_Sbox_7_M20}), .b ({new_AGEMA_signal_5957, SubBytesIns_Inst_Sbox_7_M23}), .clk (clk), .r (Fresh[202]), .c ({new_AGEMA_signal_6051, SubBytesIns_Inst_Sbox_7_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M33_U1 ( .a ({new_AGEMA_signal_5959, SubBytesIns_Inst_Sbox_7_M27}), .b ({new_AGEMA_signal_5958, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_6052, SubBytesIns_Inst_Sbox_7_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M34_U1 ( .a ({new_AGEMA_signal_5879, SubBytesIns_Inst_Sbox_7_M21}), .b ({new_AGEMA_signal_5880, SubBytesIns_Inst_Sbox_7_M22}), .clk (clk), .r (Fresh[203]), .c ({new_AGEMA_signal_5960, SubBytesIns_Inst_Sbox_7_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M36_U1 ( .a ({new_AGEMA_signal_6048, SubBytesIns_Inst_Sbox_7_M24}), .b ({new_AGEMA_signal_5958, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_6152, SubBytesIns_Inst_Sbox_7_M36}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M25_U1 ( .a ({new_AGEMA_signal_5884, SubBytesIns_Inst_Sbox_8_M22}), .b ({new_AGEMA_signal_5882, SubBytesIns_Inst_Sbox_8_M20}), .clk (clk), .r (Fresh[204]), .c ({new_AGEMA_signal_5962, SubBytesIns_Inst_Sbox_8_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M26_U1 ( .a ({new_AGEMA_signal_5883, SubBytesIns_Inst_Sbox_8_M21}), .b ({new_AGEMA_signal_5962, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_6054, SubBytesIns_Inst_Sbox_8_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M28_U1 ( .a ({new_AGEMA_signal_5961, SubBytesIns_Inst_Sbox_8_M23}), .b ({new_AGEMA_signal_5962, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_6055, SubBytesIns_Inst_Sbox_8_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M31_U1 ( .a ({new_AGEMA_signal_5882, SubBytesIns_Inst_Sbox_8_M20}), .b ({new_AGEMA_signal_5961, SubBytesIns_Inst_Sbox_8_M23}), .clk (clk), .r (Fresh[205]), .c ({new_AGEMA_signal_6056, SubBytesIns_Inst_Sbox_8_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M33_U1 ( .a ({new_AGEMA_signal_5963, SubBytesIns_Inst_Sbox_8_M27}), .b ({new_AGEMA_signal_5962, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_6057, SubBytesIns_Inst_Sbox_8_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M34_U1 ( .a ({new_AGEMA_signal_5883, SubBytesIns_Inst_Sbox_8_M21}), .b ({new_AGEMA_signal_5884, SubBytesIns_Inst_Sbox_8_M22}), .clk (clk), .r (Fresh[206]), .c ({new_AGEMA_signal_5964, SubBytesIns_Inst_Sbox_8_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M36_U1 ( .a ({new_AGEMA_signal_6053, SubBytesIns_Inst_Sbox_8_M24}), .b ({new_AGEMA_signal_5962, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_6157, SubBytesIns_Inst_Sbox_8_M36}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M25_U1 ( .a ({new_AGEMA_signal_5888, SubBytesIns_Inst_Sbox_9_M22}), .b ({new_AGEMA_signal_5886, SubBytesIns_Inst_Sbox_9_M20}), .clk (clk), .r (Fresh[207]), .c ({new_AGEMA_signal_5966, SubBytesIns_Inst_Sbox_9_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M26_U1 ( .a ({new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_9_M21}), .b ({new_AGEMA_signal_5966, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_6059, SubBytesIns_Inst_Sbox_9_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M28_U1 ( .a ({new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_9_M23}), .b ({new_AGEMA_signal_5966, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_6060, SubBytesIns_Inst_Sbox_9_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M31_U1 ( .a ({new_AGEMA_signal_5886, SubBytesIns_Inst_Sbox_9_M20}), .b ({new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_9_M23}), .clk (clk), .r (Fresh[208]), .c ({new_AGEMA_signal_6061, SubBytesIns_Inst_Sbox_9_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M33_U1 ( .a ({new_AGEMA_signal_5967, SubBytesIns_Inst_Sbox_9_M27}), .b ({new_AGEMA_signal_5966, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_6062, SubBytesIns_Inst_Sbox_9_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M34_U1 ( .a ({new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_9_M21}), .b ({new_AGEMA_signal_5888, SubBytesIns_Inst_Sbox_9_M22}), .clk (clk), .r (Fresh[209]), .c ({new_AGEMA_signal_5968, SubBytesIns_Inst_Sbox_9_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M36_U1 ( .a ({new_AGEMA_signal_6058, SubBytesIns_Inst_Sbox_9_M24}), .b ({new_AGEMA_signal_5966, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_6162, SubBytesIns_Inst_Sbox_9_M36}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M25_U1 ( .a ({new_AGEMA_signal_5892, SubBytesIns_Inst_Sbox_10_M22}), .b ({new_AGEMA_signal_5890, SubBytesIns_Inst_Sbox_10_M20}), .clk (clk), .r (Fresh[210]), .c ({new_AGEMA_signal_5970, SubBytesIns_Inst_Sbox_10_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M26_U1 ( .a ({new_AGEMA_signal_5891, SubBytesIns_Inst_Sbox_10_M21}), .b ({new_AGEMA_signal_5970, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_6064, SubBytesIns_Inst_Sbox_10_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M28_U1 ( .a ({new_AGEMA_signal_5969, SubBytesIns_Inst_Sbox_10_M23}), .b ({new_AGEMA_signal_5970, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_6065, SubBytesIns_Inst_Sbox_10_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M31_U1 ( .a ({new_AGEMA_signal_5890, SubBytesIns_Inst_Sbox_10_M20}), .b ({new_AGEMA_signal_5969, SubBytesIns_Inst_Sbox_10_M23}), .clk (clk), .r (Fresh[211]), .c ({new_AGEMA_signal_6066, SubBytesIns_Inst_Sbox_10_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M33_U1 ( .a ({new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_10_M27}), .b ({new_AGEMA_signal_5970, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_6067, SubBytesIns_Inst_Sbox_10_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M34_U1 ( .a ({new_AGEMA_signal_5891, SubBytesIns_Inst_Sbox_10_M21}), .b ({new_AGEMA_signal_5892, SubBytesIns_Inst_Sbox_10_M22}), .clk (clk), .r (Fresh[212]), .c ({new_AGEMA_signal_5972, SubBytesIns_Inst_Sbox_10_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M36_U1 ( .a ({new_AGEMA_signal_6063, SubBytesIns_Inst_Sbox_10_M24}), .b ({new_AGEMA_signal_5970, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_6167, SubBytesIns_Inst_Sbox_10_M36}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M25_U1 ( .a ({new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_11_M22}), .b ({new_AGEMA_signal_5894, SubBytesIns_Inst_Sbox_11_M20}), .clk (clk), .r (Fresh[213]), .c ({new_AGEMA_signal_5974, SubBytesIns_Inst_Sbox_11_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M26_U1 ( .a ({new_AGEMA_signal_5895, SubBytesIns_Inst_Sbox_11_M21}), .b ({new_AGEMA_signal_5974, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_6069, SubBytesIns_Inst_Sbox_11_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M28_U1 ( .a ({new_AGEMA_signal_5973, SubBytesIns_Inst_Sbox_11_M23}), .b ({new_AGEMA_signal_5974, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_6070, SubBytesIns_Inst_Sbox_11_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M31_U1 ( .a ({new_AGEMA_signal_5894, SubBytesIns_Inst_Sbox_11_M20}), .b ({new_AGEMA_signal_5973, SubBytesIns_Inst_Sbox_11_M23}), .clk (clk), .r (Fresh[214]), .c ({new_AGEMA_signal_6071, SubBytesIns_Inst_Sbox_11_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M33_U1 ( .a ({new_AGEMA_signal_5975, SubBytesIns_Inst_Sbox_11_M27}), .b ({new_AGEMA_signal_5974, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_6072, SubBytesIns_Inst_Sbox_11_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M34_U1 ( .a ({new_AGEMA_signal_5895, SubBytesIns_Inst_Sbox_11_M21}), .b ({new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_11_M22}), .clk (clk), .r (Fresh[215]), .c ({new_AGEMA_signal_5976, SubBytesIns_Inst_Sbox_11_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M36_U1 ( .a ({new_AGEMA_signal_6068, SubBytesIns_Inst_Sbox_11_M24}), .b ({new_AGEMA_signal_5974, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_6172, SubBytesIns_Inst_Sbox_11_M36}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M25_U1 ( .a ({new_AGEMA_signal_5900, SubBytesIns_Inst_Sbox_12_M22}), .b ({new_AGEMA_signal_5898, SubBytesIns_Inst_Sbox_12_M20}), .clk (clk), .r (Fresh[216]), .c ({new_AGEMA_signal_5978, SubBytesIns_Inst_Sbox_12_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M26_U1 ( .a ({new_AGEMA_signal_5899, SubBytesIns_Inst_Sbox_12_M21}), .b ({new_AGEMA_signal_5978, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_6074, SubBytesIns_Inst_Sbox_12_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M28_U1 ( .a ({new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_12_M23}), .b ({new_AGEMA_signal_5978, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_6075, SubBytesIns_Inst_Sbox_12_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M31_U1 ( .a ({new_AGEMA_signal_5898, SubBytesIns_Inst_Sbox_12_M20}), .b ({new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_12_M23}), .clk (clk), .r (Fresh[217]), .c ({new_AGEMA_signal_6076, SubBytesIns_Inst_Sbox_12_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M33_U1 ( .a ({new_AGEMA_signal_5979, SubBytesIns_Inst_Sbox_12_M27}), .b ({new_AGEMA_signal_5978, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_6077, SubBytesIns_Inst_Sbox_12_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M34_U1 ( .a ({new_AGEMA_signal_5899, SubBytesIns_Inst_Sbox_12_M21}), .b ({new_AGEMA_signal_5900, SubBytesIns_Inst_Sbox_12_M22}), .clk (clk), .r (Fresh[218]), .c ({new_AGEMA_signal_5980, SubBytesIns_Inst_Sbox_12_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M36_U1 ( .a ({new_AGEMA_signal_6073, SubBytesIns_Inst_Sbox_12_M24}), .b ({new_AGEMA_signal_5978, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_6177, SubBytesIns_Inst_Sbox_12_M36}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M25_U1 ( .a ({new_AGEMA_signal_5904, SubBytesIns_Inst_Sbox_13_M22}), .b ({new_AGEMA_signal_5902, SubBytesIns_Inst_Sbox_13_M20}), .clk (clk), .r (Fresh[219]), .c ({new_AGEMA_signal_5982, SubBytesIns_Inst_Sbox_13_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M26_U1 ( .a ({new_AGEMA_signal_5903, SubBytesIns_Inst_Sbox_13_M21}), .b ({new_AGEMA_signal_5982, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_6079, SubBytesIns_Inst_Sbox_13_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M28_U1 ( .a ({new_AGEMA_signal_5981, SubBytesIns_Inst_Sbox_13_M23}), .b ({new_AGEMA_signal_5982, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_6080, SubBytesIns_Inst_Sbox_13_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M31_U1 ( .a ({new_AGEMA_signal_5902, SubBytesIns_Inst_Sbox_13_M20}), .b ({new_AGEMA_signal_5981, SubBytesIns_Inst_Sbox_13_M23}), .clk (clk), .r (Fresh[220]), .c ({new_AGEMA_signal_6081, SubBytesIns_Inst_Sbox_13_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M33_U1 ( .a ({new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_13_M27}), .b ({new_AGEMA_signal_5982, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_6082, SubBytesIns_Inst_Sbox_13_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M34_U1 ( .a ({new_AGEMA_signal_5903, SubBytesIns_Inst_Sbox_13_M21}), .b ({new_AGEMA_signal_5904, SubBytesIns_Inst_Sbox_13_M22}), .clk (clk), .r (Fresh[221]), .c ({new_AGEMA_signal_5984, SubBytesIns_Inst_Sbox_13_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M36_U1 ( .a ({new_AGEMA_signal_6078, SubBytesIns_Inst_Sbox_13_M24}), .b ({new_AGEMA_signal_5982, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_6182, SubBytesIns_Inst_Sbox_13_M36}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M25_U1 ( .a ({new_AGEMA_signal_5908, SubBytesIns_Inst_Sbox_14_M22}), .b ({new_AGEMA_signal_5906, SubBytesIns_Inst_Sbox_14_M20}), .clk (clk), .r (Fresh[222]), .c ({new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_14_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M26_U1 ( .a ({new_AGEMA_signal_5907, SubBytesIns_Inst_Sbox_14_M21}), .b ({new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_6084, SubBytesIns_Inst_Sbox_14_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M28_U1 ( .a ({new_AGEMA_signal_5985, SubBytesIns_Inst_Sbox_14_M23}), .b ({new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_6085, SubBytesIns_Inst_Sbox_14_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M31_U1 ( .a ({new_AGEMA_signal_5906, SubBytesIns_Inst_Sbox_14_M20}), .b ({new_AGEMA_signal_5985, SubBytesIns_Inst_Sbox_14_M23}), .clk (clk), .r (Fresh[223]), .c ({new_AGEMA_signal_6086, SubBytesIns_Inst_Sbox_14_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M33_U1 ( .a ({new_AGEMA_signal_5987, SubBytesIns_Inst_Sbox_14_M27}), .b ({new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_6087, SubBytesIns_Inst_Sbox_14_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M34_U1 ( .a ({new_AGEMA_signal_5907, SubBytesIns_Inst_Sbox_14_M21}), .b ({new_AGEMA_signal_5908, SubBytesIns_Inst_Sbox_14_M22}), .clk (clk), .r (Fresh[224]), .c ({new_AGEMA_signal_5988, SubBytesIns_Inst_Sbox_14_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M36_U1 ( .a ({new_AGEMA_signal_6083, SubBytesIns_Inst_Sbox_14_M24}), .b ({new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_6187, SubBytesIns_Inst_Sbox_14_M36}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M25_U1 ( .a ({new_AGEMA_signal_5912, SubBytesIns_Inst_Sbox_15_M22}), .b ({new_AGEMA_signal_5910, SubBytesIns_Inst_Sbox_15_M20}), .clk (clk), .r (Fresh[225]), .c ({new_AGEMA_signal_5990, SubBytesIns_Inst_Sbox_15_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M26_U1 ( .a ({new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_15_M21}), .b ({new_AGEMA_signal_5990, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_6089, SubBytesIns_Inst_Sbox_15_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M28_U1 ( .a ({new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_15_M23}), .b ({new_AGEMA_signal_5990, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_6090, SubBytesIns_Inst_Sbox_15_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M31_U1 ( .a ({new_AGEMA_signal_5910, SubBytesIns_Inst_Sbox_15_M20}), .b ({new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_15_M23}), .clk (clk), .r (Fresh[226]), .c ({new_AGEMA_signal_6091, SubBytesIns_Inst_Sbox_15_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M33_U1 ( .a ({new_AGEMA_signal_5991, SubBytesIns_Inst_Sbox_15_M27}), .b ({new_AGEMA_signal_5990, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_6092, SubBytesIns_Inst_Sbox_15_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M34_U1 ( .a ({new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_15_M21}), .b ({new_AGEMA_signal_5912, SubBytesIns_Inst_Sbox_15_M22}), .clk (clk), .r (Fresh[227]), .c ({new_AGEMA_signal_5992, SubBytesIns_Inst_Sbox_15_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M36_U1 ( .a ({new_AGEMA_signal_6088, SubBytesIns_Inst_Sbox_15_M24}), .b ({new_AGEMA_signal_5990, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_6192, SubBytesIns_Inst_Sbox_15_M36}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M25_U1 ( .a ({new_AGEMA_signal_5836, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_5834, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}), .clk (clk), .r (Fresh[228]), .c ({new_AGEMA_signal_5914, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M26_U1 ( .a ({new_AGEMA_signal_5835, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_5914, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_5994, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M28_U1 ( .a ({new_AGEMA_signal_5913, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}), .b ({new_AGEMA_signal_5914, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_5995, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M31_U1 ( .a ({new_AGEMA_signal_5834, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_5913, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}), .clk (clk), .r (Fresh[229]), .c ({new_AGEMA_signal_5996, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M33_U1 ( .a ({new_AGEMA_signal_5915, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27}), .b ({new_AGEMA_signal_5914, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_5997, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M34_U1 ( .a ({new_AGEMA_signal_5835, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_5836, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}), .clk (clk), .r (Fresh[230]), .c ({new_AGEMA_signal_5916, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M36_U1 ( .a ({new_AGEMA_signal_5993, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24}), .b ({new_AGEMA_signal_5914, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_6097, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M25_U1 ( .a ({new_AGEMA_signal_5840, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_5838, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}), .clk (clk), .r (Fresh[231]), .c ({new_AGEMA_signal_5918, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M26_U1 ( .a ({new_AGEMA_signal_5839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_5918, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_5999, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M28_U1 ( .a ({new_AGEMA_signal_5917, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}), .b ({new_AGEMA_signal_5918, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_6000, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M31_U1 ( .a ({new_AGEMA_signal_5838, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_5917, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}), .clk (clk), .r (Fresh[232]), .c ({new_AGEMA_signal_6001, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M33_U1 ( .a ({new_AGEMA_signal_5919, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27}), .b ({new_AGEMA_signal_5918, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_6002, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M34_U1 ( .a ({new_AGEMA_signal_5839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_5840, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}), .clk (clk), .r (Fresh[233]), .c ({new_AGEMA_signal_5920, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M36_U1 ( .a ({new_AGEMA_signal_5998, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24}), .b ({new_AGEMA_signal_5918, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_6102, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M25_U1 ( .a ({new_AGEMA_signal_5844, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_5842, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}), .clk (clk), .r (Fresh[234]), .c ({new_AGEMA_signal_5922, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M26_U1 ( .a ({new_AGEMA_signal_5843, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_5922, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_6004, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M28_U1 ( .a ({new_AGEMA_signal_5921, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}), .b ({new_AGEMA_signal_5922, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_6005, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M31_U1 ( .a ({new_AGEMA_signal_5842, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_5921, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}), .clk (clk), .r (Fresh[235]), .c ({new_AGEMA_signal_6006, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M33_U1 ( .a ({new_AGEMA_signal_5923, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27}), .b ({new_AGEMA_signal_5922, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_6007, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M34_U1 ( .a ({new_AGEMA_signal_5843, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_5844, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}), .clk (clk), .r (Fresh[236]), .c ({new_AGEMA_signal_5924, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M36_U1 ( .a ({new_AGEMA_signal_6003, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24}), .b ({new_AGEMA_signal_5922, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_6107, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M25_U1 ( .a ({new_AGEMA_signal_5848, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_5846, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}), .clk (clk), .r (Fresh[237]), .c ({new_AGEMA_signal_5926, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M26_U1 ( .a ({new_AGEMA_signal_5847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_5926, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_6009, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M28_U1 ( .a ({new_AGEMA_signal_5925, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}), .b ({new_AGEMA_signal_5926, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_6010, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M31_U1 ( .a ({new_AGEMA_signal_5846, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_5925, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}), .clk (clk), .r (Fresh[238]), .c ({new_AGEMA_signal_6011, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M33_U1 ( .a ({new_AGEMA_signal_5927, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27}), .b ({new_AGEMA_signal_5926, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_6012, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M34_U1 ( .a ({new_AGEMA_signal_5847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_5848, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}), .clk (clk), .r (Fresh[239]), .c ({new_AGEMA_signal_5928, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M36_U1 ( .a ({new_AGEMA_signal_6008, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24}), .b ({new_AGEMA_signal_5926, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_6112, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M29_U1 ( .a ({new_AGEMA_signal_6015, SubBytesIns_Inst_Sbox_0_M28}), .b ({new_AGEMA_signal_5931, SubBytesIns_Inst_Sbox_0_M27}), .clk (clk), .r (Fresh[240]), .c ({new_AGEMA_signal_6113, SubBytesIns_Inst_Sbox_0_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M30_U1 ( .a ({new_AGEMA_signal_6014, SubBytesIns_Inst_Sbox_0_M26}), .b ({new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_0_M24}), .clk (clk), .r (Fresh[241]), .c ({new_AGEMA_signal_6114, SubBytesIns_Inst_Sbox_0_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M32_U1 ( .a ({new_AGEMA_signal_5931, SubBytesIns_Inst_Sbox_0_M27}), .b ({new_AGEMA_signal_6016, SubBytesIns_Inst_Sbox_0_M31}), .clk (clk), .r (Fresh[242]), .c ({new_AGEMA_signal_6115, SubBytesIns_Inst_Sbox_0_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M35_U1 ( .a ({new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_0_M24}), .b ({new_AGEMA_signal_5932, SubBytesIns_Inst_Sbox_0_M34}), .clk (clk), .r (Fresh[243]), .c ({new_AGEMA_signal_6116, SubBytesIns_Inst_Sbox_0_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M37_U1 ( .a ({new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_6113, SubBytesIns_Inst_Sbox_0_M29}), .c ({new_AGEMA_signal_6209, SubBytesIns_Inst_Sbox_0_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M38_U1 ( .a ({new_AGEMA_signal_6115, SubBytesIns_Inst_Sbox_0_M32}), .b ({new_AGEMA_signal_6017, SubBytesIns_Inst_Sbox_0_M33}), .c ({new_AGEMA_signal_6210, SubBytesIns_Inst_Sbox_0_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M39_U1 ( .a ({new_AGEMA_signal_5929, SubBytesIns_Inst_Sbox_0_M23}), .b ({new_AGEMA_signal_6114, SubBytesIns_Inst_Sbox_0_M30}), .c ({new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_0_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M40_U1 ( .a ({new_AGEMA_signal_6116, SubBytesIns_Inst_Sbox_0_M35}), .b ({new_AGEMA_signal_6117, SubBytesIns_Inst_Sbox_0_M36}), .c ({new_AGEMA_signal_6212, SubBytesIns_Inst_Sbox_0_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M41_U1 ( .a ({new_AGEMA_signal_6210, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_6212, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_6321, SubBytesIns_Inst_Sbox_0_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M42_U1 ( .a ({new_AGEMA_signal_6209, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_0_M39}), .c ({new_AGEMA_signal_6322, SubBytesIns_Inst_Sbox_0_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M43_U1 ( .a ({new_AGEMA_signal_6209, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_6210, SubBytesIns_Inst_Sbox_0_M38}), .c ({new_AGEMA_signal_6323, SubBytesIns_Inst_Sbox_0_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M44_U1 ( .a ({new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_6212, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_6324, SubBytesIns_Inst_Sbox_0_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M45_U1 ( .a ({new_AGEMA_signal_6322, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_6321, SubBytesIns_Inst_Sbox_0_M41}), .c ({new_AGEMA_signal_6561, SubBytesIns_Inst_Sbox_0_M45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M29_U1 ( .a ({new_AGEMA_signal_6020, SubBytesIns_Inst_Sbox_1_M28}), .b ({new_AGEMA_signal_5935, SubBytesIns_Inst_Sbox_1_M27}), .clk (clk), .r (Fresh[244]), .c ({new_AGEMA_signal_6118, SubBytesIns_Inst_Sbox_1_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M30_U1 ( .a ({new_AGEMA_signal_6019, SubBytesIns_Inst_Sbox_1_M26}), .b ({new_AGEMA_signal_6018, SubBytesIns_Inst_Sbox_1_M24}), .clk (clk), .r (Fresh[245]), .c ({new_AGEMA_signal_6119, SubBytesIns_Inst_Sbox_1_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M32_U1 ( .a ({new_AGEMA_signal_5935, SubBytesIns_Inst_Sbox_1_M27}), .b ({new_AGEMA_signal_6021, SubBytesIns_Inst_Sbox_1_M31}), .clk (clk), .r (Fresh[246]), .c ({new_AGEMA_signal_6120, SubBytesIns_Inst_Sbox_1_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M35_U1 ( .a ({new_AGEMA_signal_6018, SubBytesIns_Inst_Sbox_1_M24}), .b ({new_AGEMA_signal_5936, SubBytesIns_Inst_Sbox_1_M34}), .clk (clk), .r (Fresh[247]), .c ({new_AGEMA_signal_6121, SubBytesIns_Inst_Sbox_1_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M37_U1 ( .a ({new_AGEMA_signal_5855, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_6118, SubBytesIns_Inst_Sbox_1_M29}), .c ({new_AGEMA_signal_6213, SubBytesIns_Inst_Sbox_1_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M38_U1 ( .a ({new_AGEMA_signal_6120, SubBytesIns_Inst_Sbox_1_M32}), .b ({new_AGEMA_signal_6022, SubBytesIns_Inst_Sbox_1_M33}), .c ({new_AGEMA_signal_6214, SubBytesIns_Inst_Sbox_1_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M39_U1 ( .a ({new_AGEMA_signal_5933, SubBytesIns_Inst_Sbox_1_M23}), .b ({new_AGEMA_signal_6119, SubBytesIns_Inst_Sbox_1_M30}), .c ({new_AGEMA_signal_6215, SubBytesIns_Inst_Sbox_1_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M40_U1 ( .a ({new_AGEMA_signal_6121, SubBytesIns_Inst_Sbox_1_M35}), .b ({new_AGEMA_signal_6122, SubBytesIns_Inst_Sbox_1_M36}), .c ({new_AGEMA_signal_6216, SubBytesIns_Inst_Sbox_1_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M41_U1 ( .a ({new_AGEMA_signal_6214, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_6216, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_6333, SubBytesIns_Inst_Sbox_1_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M42_U1 ( .a ({new_AGEMA_signal_6213, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_6215, SubBytesIns_Inst_Sbox_1_M39}), .c ({new_AGEMA_signal_6334, SubBytesIns_Inst_Sbox_1_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M43_U1 ( .a ({new_AGEMA_signal_6213, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_6214, SubBytesIns_Inst_Sbox_1_M38}), .c ({new_AGEMA_signal_6335, SubBytesIns_Inst_Sbox_1_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M44_U1 ( .a ({new_AGEMA_signal_6215, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_6216, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_6336, SubBytesIns_Inst_Sbox_1_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M45_U1 ( .a ({new_AGEMA_signal_6334, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_6333, SubBytesIns_Inst_Sbox_1_M41}), .c ({new_AGEMA_signal_6573, SubBytesIns_Inst_Sbox_1_M45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M29_U1 ( .a ({new_AGEMA_signal_6025, SubBytesIns_Inst_Sbox_2_M28}), .b ({new_AGEMA_signal_5939, SubBytesIns_Inst_Sbox_2_M27}), .clk (clk), .r (Fresh[248]), .c ({new_AGEMA_signal_6123, SubBytesIns_Inst_Sbox_2_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M30_U1 ( .a ({new_AGEMA_signal_6024, SubBytesIns_Inst_Sbox_2_M26}), .b ({new_AGEMA_signal_6023, SubBytesIns_Inst_Sbox_2_M24}), .clk (clk), .r (Fresh[249]), .c ({new_AGEMA_signal_6124, SubBytesIns_Inst_Sbox_2_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M32_U1 ( .a ({new_AGEMA_signal_5939, SubBytesIns_Inst_Sbox_2_M27}), .b ({new_AGEMA_signal_6026, SubBytesIns_Inst_Sbox_2_M31}), .clk (clk), .r (Fresh[250]), .c ({new_AGEMA_signal_6125, SubBytesIns_Inst_Sbox_2_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M35_U1 ( .a ({new_AGEMA_signal_6023, SubBytesIns_Inst_Sbox_2_M24}), .b ({new_AGEMA_signal_5940, SubBytesIns_Inst_Sbox_2_M34}), .clk (clk), .r (Fresh[251]), .c ({new_AGEMA_signal_6126, SubBytesIns_Inst_Sbox_2_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M37_U1 ( .a ({new_AGEMA_signal_5859, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_6123, SubBytesIns_Inst_Sbox_2_M29}), .c ({new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_2_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M38_U1 ( .a ({new_AGEMA_signal_6125, SubBytesIns_Inst_Sbox_2_M32}), .b ({new_AGEMA_signal_6027, SubBytesIns_Inst_Sbox_2_M33}), .c ({new_AGEMA_signal_6218, SubBytesIns_Inst_Sbox_2_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M39_U1 ( .a ({new_AGEMA_signal_5937, SubBytesIns_Inst_Sbox_2_M23}), .b ({new_AGEMA_signal_6124, SubBytesIns_Inst_Sbox_2_M30}), .c ({new_AGEMA_signal_6219, SubBytesIns_Inst_Sbox_2_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M40_U1 ( .a ({new_AGEMA_signal_6126, SubBytesIns_Inst_Sbox_2_M35}), .b ({new_AGEMA_signal_6127, SubBytesIns_Inst_Sbox_2_M36}), .c ({new_AGEMA_signal_6220, SubBytesIns_Inst_Sbox_2_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M41_U1 ( .a ({new_AGEMA_signal_6218, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_6220, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_6345, SubBytesIns_Inst_Sbox_2_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M42_U1 ( .a ({new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_6219, SubBytesIns_Inst_Sbox_2_M39}), .c ({new_AGEMA_signal_6346, SubBytesIns_Inst_Sbox_2_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M43_U1 ( .a ({new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_6218, SubBytesIns_Inst_Sbox_2_M38}), .c ({new_AGEMA_signal_6347, SubBytesIns_Inst_Sbox_2_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M44_U1 ( .a ({new_AGEMA_signal_6219, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_6220, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_6348, SubBytesIns_Inst_Sbox_2_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M45_U1 ( .a ({new_AGEMA_signal_6346, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_6345, SubBytesIns_Inst_Sbox_2_M41}), .c ({new_AGEMA_signal_6585, SubBytesIns_Inst_Sbox_2_M45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M29_U1 ( .a ({new_AGEMA_signal_6030, SubBytesIns_Inst_Sbox_3_M28}), .b ({new_AGEMA_signal_5943, SubBytesIns_Inst_Sbox_3_M27}), .clk (clk), .r (Fresh[252]), .c ({new_AGEMA_signal_6128, SubBytesIns_Inst_Sbox_3_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M30_U1 ( .a ({new_AGEMA_signal_6029, SubBytesIns_Inst_Sbox_3_M26}), .b ({new_AGEMA_signal_6028, SubBytesIns_Inst_Sbox_3_M24}), .clk (clk), .r (Fresh[253]), .c ({new_AGEMA_signal_6129, SubBytesIns_Inst_Sbox_3_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M32_U1 ( .a ({new_AGEMA_signal_5943, SubBytesIns_Inst_Sbox_3_M27}), .b ({new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_3_M31}), .clk (clk), .r (Fresh[254]), .c ({new_AGEMA_signal_6130, SubBytesIns_Inst_Sbox_3_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M35_U1 ( .a ({new_AGEMA_signal_6028, SubBytesIns_Inst_Sbox_3_M24}), .b ({new_AGEMA_signal_5944, SubBytesIns_Inst_Sbox_3_M34}), .clk (clk), .r (Fresh[255]), .c ({new_AGEMA_signal_6131, SubBytesIns_Inst_Sbox_3_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M37_U1 ( .a ({new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_6128, SubBytesIns_Inst_Sbox_3_M29}), .c ({new_AGEMA_signal_6221, SubBytesIns_Inst_Sbox_3_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M38_U1 ( .a ({new_AGEMA_signal_6130, SubBytesIns_Inst_Sbox_3_M32}), .b ({new_AGEMA_signal_6032, SubBytesIns_Inst_Sbox_3_M33}), .c ({new_AGEMA_signal_6222, SubBytesIns_Inst_Sbox_3_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M39_U1 ( .a ({new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_3_M23}), .b ({new_AGEMA_signal_6129, SubBytesIns_Inst_Sbox_3_M30}), .c ({new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_3_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M40_U1 ( .a ({new_AGEMA_signal_6131, SubBytesIns_Inst_Sbox_3_M35}), .b ({new_AGEMA_signal_6132, SubBytesIns_Inst_Sbox_3_M36}), .c ({new_AGEMA_signal_6224, SubBytesIns_Inst_Sbox_3_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M41_U1 ( .a ({new_AGEMA_signal_6222, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_6224, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_6357, SubBytesIns_Inst_Sbox_3_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M42_U1 ( .a ({new_AGEMA_signal_6221, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_3_M39}), .c ({new_AGEMA_signal_6358, SubBytesIns_Inst_Sbox_3_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M43_U1 ( .a ({new_AGEMA_signal_6221, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_6222, SubBytesIns_Inst_Sbox_3_M38}), .c ({new_AGEMA_signal_6359, SubBytesIns_Inst_Sbox_3_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M44_U1 ( .a ({new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_6224, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_6360, SubBytesIns_Inst_Sbox_3_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M45_U1 ( .a ({new_AGEMA_signal_6358, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_6357, SubBytesIns_Inst_Sbox_3_M41}), .c ({new_AGEMA_signal_6597, SubBytesIns_Inst_Sbox_3_M45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M29_U1 ( .a ({new_AGEMA_signal_6035, SubBytesIns_Inst_Sbox_4_M28}), .b ({new_AGEMA_signal_5947, SubBytesIns_Inst_Sbox_4_M27}), .clk (clk), .r (Fresh[256]), .c ({new_AGEMA_signal_6133, SubBytesIns_Inst_Sbox_4_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M30_U1 ( .a ({new_AGEMA_signal_6034, SubBytesIns_Inst_Sbox_4_M26}), .b ({new_AGEMA_signal_6033, SubBytesIns_Inst_Sbox_4_M24}), .clk (clk), .r (Fresh[257]), .c ({new_AGEMA_signal_6134, SubBytesIns_Inst_Sbox_4_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M32_U1 ( .a ({new_AGEMA_signal_5947, SubBytesIns_Inst_Sbox_4_M27}), .b ({new_AGEMA_signal_6036, SubBytesIns_Inst_Sbox_4_M31}), .clk (clk), .r (Fresh[258]), .c ({new_AGEMA_signal_6135, SubBytesIns_Inst_Sbox_4_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M35_U1 ( .a ({new_AGEMA_signal_6033, SubBytesIns_Inst_Sbox_4_M24}), .b ({new_AGEMA_signal_5948, SubBytesIns_Inst_Sbox_4_M34}), .clk (clk), .r (Fresh[259]), .c ({new_AGEMA_signal_6136, SubBytesIns_Inst_Sbox_4_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M37_U1 ( .a ({new_AGEMA_signal_5867, SubBytesIns_Inst_Sbox_4_M21}), .b ({new_AGEMA_signal_6133, SubBytesIns_Inst_Sbox_4_M29}), .c ({new_AGEMA_signal_6225, SubBytesIns_Inst_Sbox_4_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M38_U1 ( .a ({new_AGEMA_signal_6135, SubBytesIns_Inst_Sbox_4_M32}), .b ({new_AGEMA_signal_6037, SubBytesIns_Inst_Sbox_4_M33}), .c ({new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_4_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M39_U1 ( .a ({new_AGEMA_signal_5945, SubBytesIns_Inst_Sbox_4_M23}), .b ({new_AGEMA_signal_6134, SubBytesIns_Inst_Sbox_4_M30}), .c ({new_AGEMA_signal_6227, SubBytesIns_Inst_Sbox_4_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M40_U1 ( .a ({new_AGEMA_signal_6136, SubBytesIns_Inst_Sbox_4_M35}), .b ({new_AGEMA_signal_6137, SubBytesIns_Inst_Sbox_4_M36}), .c ({new_AGEMA_signal_6228, SubBytesIns_Inst_Sbox_4_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M41_U1 ( .a ({new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_4_M38}), .b ({new_AGEMA_signal_6228, SubBytesIns_Inst_Sbox_4_M40}), .c ({new_AGEMA_signal_6369, SubBytesIns_Inst_Sbox_4_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M42_U1 ( .a ({new_AGEMA_signal_6225, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_6227, SubBytesIns_Inst_Sbox_4_M39}), .c ({new_AGEMA_signal_6370, SubBytesIns_Inst_Sbox_4_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M43_U1 ( .a ({new_AGEMA_signal_6225, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_4_M38}), .c ({new_AGEMA_signal_6371, SubBytesIns_Inst_Sbox_4_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M44_U1 ( .a ({new_AGEMA_signal_6227, SubBytesIns_Inst_Sbox_4_M39}), .b ({new_AGEMA_signal_6228, SubBytesIns_Inst_Sbox_4_M40}), .c ({new_AGEMA_signal_6372, SubBytesIns_Inst_Sbox_4_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M45_U1 ( .a ({new_AGEMA_signal_6370, SubBytesIns_Inst_Sbox_4_M42}), .b ({new_AGEMA_signal_6369, SubBytesIns_Inst_Sbox_4_M41}), .c ({new_AGEMA_signal_6609, SubBytesIns_Inst_Sbox_4_M45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M29_U1 ( .a ({new_AGEMA_signal_6040, SubBytesIns_Inst_Sbox_5_M28}), .b ({new_AGEMA_signal_5951, SubBytesIns_Inst_Sbox_5_M27}), .clk (clk), .r (Fresh[260]), .c ({new_AGEMA_signal_6138, SubBytesIns_Inst_Sbox_5_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M30_U1 ( .a ({new_AGEMA_signal_6039, SubBytesIns_Inst_Sbox_5_M26}), .b ({new_AGEMA_signal_6038, SubBytesIns_Inst_Sbox_5_M24}), .clk (clk), .r (Fresh[261]), .c ({new_AGEMA_signal_6139, SubBytesIns_Inst_Sbox_5_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M32_U1 ( .a ({new_AGEMA_signal_5951, SubBytesIns_Inst_Sbox_5_M27}), .b ({new_AGEMA_signal_6041, SubBytesIns_Inst_Sbox_5_M31}), .clk (clk), .r (Fresh[262]), .c ({new_AGEMA_signal_6140, SubBytesIns_Inst_Sbox_5_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M35_U1 ( .a ({new_AGEMA_signal_6038, SubBytesIns_Inst_Sbox_5_M24}), .b ({new_AGEMA_signal_5952, SubBytesIns_Inst_Sbox_5_M34}), .clk (clk), .r (Fresh[263]), .c ({new_AGEMA_signal_6141, SubBytesIns_Inst_Sbox_5_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M37_U1 ( .a ({new_AGEMA_signal_5871, SubBytesIns_Inst_Sbox_5_M21}), .b ({new_AGEMA_signal_6138, SubBytesIns_Inst_Sbox_5_M29}), .c ({new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_5_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M38_U1 ( .a ({new_AGEMA_signal_6140, SubBytesIns_Inst_Sbox_5_M32}), .b ({new_AGEMA_signal_6042, SubBytesIns_Inst_Sbox_5_M33}), .c ({new_AGEMA_signal_6230, SubBytesIns_Inst_Sbox_5_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M39_U1 ( .a ({new_AGEMA_signal_5949, SubBytesIns_Inst_Sbox_5_M23}), .b ({new_AGEMA_signal_6139, SubBytesIns_Inst_Sbox_5_M30}), .c ({new_AGEMA_signal_6231, SubBytesIns_Inst_Sbox_5_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M40_U1 ( .a ({new_AGEMA_signal_6141, SubBytesIns_Inst_Sbox_5_M35}), .b ({new_AGEMA_signal_6142, SubBytesIns_Inst_Sbox_5_M36}), .c ({new_AGEMA_signal_6232, SubBytesIns_Inst_Sbox_5_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M41_U1 ( .a ({new_AGEMA_signal_6230, SubBytesIns_Inst_Sbox_5_M38}), .b ({new_AGEMA_signal_6232, SubBytesIns_Inst_Sbox_5_M40}), .c ({new_AGEMA_signal_6381, SubBytesIns_Inst_Sbox_5_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M42_U1 ( .a ({new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_6231, SubBytesIns_Inst_Sbox_5_M39}), .c ({new_AGEMA_signal_6382, SubBytesIns_Inst_Sbox_5_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M43_U1 ( .a ({new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_6230, SubBytesIns_Inst_Sbox_5_M38}), .c ({new_AGEMA_signal_6383, SubBytesIns_Inst_Sbox_5_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M44_U1 ( .a ({new_AGEMA_signal_6231, SubBytesIns_Inst_Sbox_5_M39}), .b ({new_AGEMA_signal_6232, SubBytesIns_Inst_Sbox_5_M40}), .c ({new_AGEMA_signal_6384, SubBytesIns_Inst_Sbox_5_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M45_U1 ( .a ({new_AGEMA_signal_6382, SubBytesIns_Inst_Sbox_5_M42}), .b ({new_AGEMA_signal_6381, SubBytesIns_Inst_Sbox_5_M41}), .c ({new_AGEMA_signal_6621, SubBytesIns_Inst_Sbox_5_M45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M29_U1 ( .a ({new_AGEMA_signal_6045, SubBytesIns_Inst_Sbox_6_M28}), .b ({new_AGEMA_signal_5955, SubBytesIns_Inst_Sbox_6_M27}), .clk (clk), .r (Fresh[264]), .c ({new_AGEMA_signal_6143, SubBytesIns_Inst_Sbox_6_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M30_U1 ( .a ({new_AGEMA_signal_6044, SubBytesIns_Inst_Sbox_6_M26}), .b ({new_AGEMA_signal_6043, SubBytesIns_Inst_Sbox_6_M24}), .clk (clk), .r (Fresh[265]), .c ({new_AGEMA_signal_6144, SubBytesIns_Inst_Sbox_6_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M32_U1 ( .a ({new_AGEMA_signal_5955, SubBytesIns_Inst_Sbox_6_M27}), .b ({new_AGEMA_signal_6046, SubBytesIns_Inst_Sbox_6_M31}), .clk (clk), .r (Fresh[266]), .c ({new_AGEMA_signal_6145, SubBytesIns_Inst_Sbox_6_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M35_U1 ( .a ({new_AGEMA_signal_6043, SubBytesIns_Inst_Sbox_6_M24}), .b ({new_AGEMA_signal_5956, SubBytesIns_Inst_Sbox_6_M34}), .clk (clk), .r (Fresh[267]), .c ({new_AGEMA_signal_6146, SubBytesIns_Inst_Sbox_6_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M37_U1 ( .a ({new_AGEMA_signal_5875, SubBytesIns_Inst_Sbox_6_M21}), .b ({new_AGEMA_signal_6143, SubBytesIns_Inst_Sbox_6_M29}), .c ({new_AGEMA_signal_6233, SubBytesIns_Inst_Sbox_6_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M38_U1 ( .a ({new_AGEMA_signal_6145, SubBytesIns_Inst_Sbox_6_M32}), .b ({new_AGEMA_signal_6047, SubBytesIns_Inst_Sbox_6_M33}), .c ({new_AGEMA_signal_6234, SubBytesIns_Inst_Sbox_6_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M39_U1 ( .a ({new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_6_M23}), .b ({new_AGEMA_signal_6144, SubBytesIns_Inst_Sbox_6_M30}), .c ({new_AGEMA_signal_6235, SubBytesIns_Inst_Sbox_6_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M40_U1 ( .a ({new_AGEMA_signal_6146, SubBytesIns_Inst_Sbox_6_M35}), .b ({new_AGEMA_signal_6147, SubBytesIns_Inst_Sbox_6_M36}), .c ({new_AGEMA_signal_6236, SubBytesIns_Inst_Sbox_6_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M41_U1 ( .a ({new_AGEMA_signal_6234, SubBytesIns_Inst_Sbox_6_M38}), .b ({new_AGEMA_signal_6236, SubBytesIns_Inst_Sbox_6_M40}), .c ({new_AGEMA_signal_6393, SubBytesIns_Inst_Sbox_6_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M42_U1 ( .a ({new_AGEMA_signal_6233, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_6235, SubBytesIns_Inst_Sbox_6_M39}), .c ({new_AGEMA_signal_6394, SubBytesIns_Inst_Sbox_6_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M43_U1 ( .a ({new_AGEMA_signal_6233, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_6234, SubBytesIns_Inst_Sbox_6_M38}), .c ({new_AGEMA_signal_6395, SubBytesIns_Inst_Sbox_6_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M44_U1 ( .a ({new_AGEMA_signal_6235, SubBytesIns_Inst_Sbox_6_M39}), .b ({new_AGEMA_signal_6236, SubBytesIns_Inst_Sbox_6_M40}), .c ({new_AGEMA_signal_6396, SubBytesIns_Inst_Sbox_6_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M45_U1 ( .a ({new_AGEMA_signal_6394, SubBytesIns_Inst_Sbox_6_M42}), .b ({new_AGEMA_signal_6393, SubBytesIns_Inst_Sbox_6_M41}), .c ({new_AGEMA_signal_6633, SubBytesIns_Inst_Sbox_6_M45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M29_U1 ( .a ({new_AGEMA_signal_6050, SubBytesIns_Inst_Sbox_7_M28}), .b ({new_AGEMA_signal_5959, SubBytesIns_Inst_Sbox_7_M27}), .clk (clk), .r (Fresh[268]), .c ({new_AGEMA_signal_6148, SubBytesIns_Inst_Sbox_7_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M30_U1 ( .a ({new_AGEMA_signal_6049, SubBytesIns_Inst_Sbox_7_M26}), .b ({new_AGEMA_signal_6048, SubBytesIns_Inst_Sbox_7_M24}), .clk (clk), .r (Fresh[269]), .c ({new_AGEMA_signal_6149, SubBytesIns_Inst_Sbox_7_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M32_U1 ( .a ({new_AGEMA_signal_5959, SubBytesIns_Inst_Sbox_7_M27}), .b ({new_AGEMA_signal_6051, SubBytesIns_Inst_Sbox_7_M31}), .clk (clk), .r (Fresh[270]), .c ({new_AGEMA_signal_6150, SubBytesIns_Inst_Sbox_7_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M35_U1 ( .a ({new_AGEMA_signal_6048, SubBytesIns_Inst_Sbox_7_M24}), .b ({new_AGEMA_signal_5960, SubBytesIns_Inst_Sbox_7_M34}), .clk (clk), .r (Fresh[271]), .c ({new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_7_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M37_U1 ( .a ({new_AGEMA_signal_5879, SubBytesIns_Inst_Sbox_7_M21}), .b ({new_AGEMA_signal_6148, SubBytesIns_Inst_Sbox_7_M29}), .c ({new_AGEMA_signal_6237, SubBytesIns_Inst_Sbox_7_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M38_U1 ( .a ({new_AGEMA_signal_6150, SubBytesIns_Inst_Sbox_7_M32}), .b ({new_AGEMA_signal_6052, SubBytesIns_Inst_Sbox_7_M33}), .c ({new_AGEMA_signal_6238, SubBytesIns_Inst_Sbox_7_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M39_U1 ( .a ({new_AGEMA_signal_5957, SubBytesIns_Inst_Sbox_7_M23}), .b ({new_AGEMA_signal_6149, SubBytesIns_Inst_Sbox_7_M30}), .c ({new_AGEMA_signal_6239, SubBytesIns_Inst_Sbox_7_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M40_U1 ( .a ({new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_7_M35}), .b ({new_AGEMA_signal_6152, SubBytesIns_Inst_Sbox_7_M36}), .c ({new_AGEMA_signal_6240, SubBytesIns_Inst_Sbox_7_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M41_U1 ( .a ({new_AGEMA_signal_6238, SubBytesIns_Inst_Sbox_7_M38}), .b ({new_AGEMA_signal_6240, SubBytesIns_Inst_Sbox_7_M40}), .c ({new_AGEMA_signal_6405, SubBytesIns_Inst_Sbox_7_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M42_U1 ( .a ({new_AGEMA_signal_6237, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_6239, SubBytesIns_Inst_Sbox_7_M39}), .c ({new_AGEMA_signal_6406, SubBytesIns_Inst_Sbox_7_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M43_U1 ( .a ({new_AGEMA_signal_6237, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_6238, SubBytesIns_Inst_Sbox_7_M38}), .c ({new_AGEMA_signal_6407, SubBytesIns_Inst_Sbox_7_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M44_U1 ( .a ({new_AGEMA_signal_6239, SubBytesIns_Inst_Sbox_7_M39}), .b ({new_AGEMA_signal_6240, SubBytesIns_Inst_Sbox_7_M40}), .c ({new_AGEMA_signal_6408, SubBytesIns_Inst_Sbox_7_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M45_U1 ( .a ({new_AGEMA_signal_6406, SubBytesIns_Inst_Sbox_7_M42}), .b ({new_AGEMA_signal_6405, SubBytesIns_Inst_Sbox_7_M41}), .c ({new_AGEMA_signal_6645, SubBytesIns_Inst_Sbox_7_M45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M29_U1 ( .a ({new_AGEMA_signal_6055, SubBytesIns_Inst_Sbox_8_M28}), .b ({new_AGEMA_signal_5963, SubBytesIns_Inst_Sbox_8_M27}), .clk (clk), .r (Fresh[272]), .c ({new_AGEMA_signal_6153, SubBytesIns_Inst_Sbox_8_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M30_U1 ( .a ({new_AGEMA_signal_6054, SubBytesIns_Inst_Sbox_8_M26}), .b ({new_AGEMA_signal_6053, SubBytesIns_Inst_Sbox_8_M24}), .clk (clk), .r (Fresh[273]), .c ({new_AGEMA_signal_6154, SubBytesIns_Inst_Sbox_8_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M32_U1 ( .a ({new_AGEMA_signal_5963, SubBytesIns_Inst_Sbox_8_M27}), .b ({new_AGEMA_signal_6056, SubBytesIns_Inst_Sbox_8_M31}), .clk (clk), .r (Fresh[274]), .c ({new_AGEMA_signal_6155, SubBytesIns_Inst_Sbox_8_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M35_U1 ( .a ({new_AGEMA_signal_6053, SubBytesIns_Inst_Sbox_8_M24}), .b ({new_AGEMA_signal_5964, SubBytesIns_Inst_Sbox_8_M34}), .clk (clk), .r (Fresh[275]), .c ({new_AGEMA_signal_6156, SubBytesIns_Inst_Sbox_8_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M37_U1 ( .a ({new_AGEMA_signal_5883, SubBytesIns_Inst_Sbox_8_M21}), .b ({new_AGEMA_signal_6153, SubBytesIns_Inst_Sbox_8_M29}), .c ({new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_8_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M38_U1 ( .a ({new_AGEMA_signal_6155, SubBytesIns_Inst_Sbox_8_M32}), .b ({new_AGEMA_signal_6057, SubBytesIns_Inst_Sbox_8_M33}), .c ({new_AGEMA_signal_6242, SubBytesIns_Inst_Sbox_8_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M39_U1 ( .a ({new_AGEMA_signal_5961, SubBytesIns_Inst_Sbox_8_M23}), .b ({new_AGEMA_signal_6154, SubBytesIns_Inst_Sbox_8_M30}), .c ({new_AGEMA_signal_6243, SubBytesIns_Inst_Sbox_8_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M40_U1 ( .a ({new_AGEMA_signal_6156, SubBytesIns_Inst_Sbox_8_M35}), .b ({new_AGEMA_signal_6157, SubBytesIns_Inst_Sbox_8_M36}), .c ({new_AGEMA_signal_6244, SubBytesIns_Inst_Sbox_8_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M41_U1 ( .a ({new_AGEMA_signal_6242, SubBytesIns_Inst_Sbox_8_M38}), .b ({new_AGEMA_signal_6244, SubBytesIns_Inst_Sbox_8_M40}), .c ({new_AGEMA_signal_6417, SubBytesIns_Inst_Sbox_8_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M42_U1 ( .a ({new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_6243, SubBytesIns_Inst_Sbox_8_M39}), .c ({new_AGEMA_signal_6418, SubBytesIns_Inst_Sbox_8_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M43_U1 ( .a ({new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_6242, SubBytesIns_Inst_Sbox_8_M38}), .c ({new_AGEMA_signal_6419, SubBytesIns_Inst_Sbox_8_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M44_U1 ( .a ({new_AGEMA_signal_6243, SubBytesIns_Inst_Sbox_8_M39}), .b ({new_AGEMA_signal_6244, SubBytesIns_Inst_Sbox_8_M40}), .c ({new_AGEMA_signal_6420, SubBytesIns_Inst_Sbox_8_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M45_U1 ( .a ({new_AGEMA_signal_6418, SubBytesIns_Inst_Sbox_8_M42}), .b ({new_AGEMA_signal_6417, SubBytesIns_Inst_Sbox_8_M41}), .c ({new_AGEMA_signal_6657, SubBytesIns_Inst_Sbox_8_M45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M29_U1 ( .a ({new_AGEMA_signal_6060, SubBytesIns_Inst_Sbox_9_M28}), .b ({new_AGEMA_signal_5967, SubBytesIns_Inst_Sbox_9_M27}), .clk (clk), .r (Fresh[276]), .c ({new_AGEMA_signal_6158, SubBytesIns_Inst_Sbox_9_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M30_U1 ( .a ({new_AGEMA_signal_6059, SubBytesIns_Inst_Sbox_9_M26}), .b ({new_AGEMA_signal_6058, SubBytesIns_Inst_Sbox_9_M24}), .clk (clk), .r (Fresh[277]), .c ({new_AGEMA_signal_6159, SubBytesIns_Inst_Sbox_9_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M32_U1 ( .a ({new_AGEMA_signal_5967, SubBytesIns_Inst_Sbox_9_M27}), .b ({new_AGEMA_signal_6061, SubBytesIns_Inst_Sbox_9_M31}), .clk (clk), .r (Fresh[278]), .c ({new_AGEMA_signal_6160, SubBytesIns_Inst_Sbox_9_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M35_U1 ( .a ({new_AGEMA_signal_6058, SubBytesIns_Inst_Sbox_9_M24}), .b ({new_AGEMA_signal_5968, SubBytesIns_Inst_Sbox_9_M34}), .clk (clk), .r (Fresh[279]), .c ({new_AGEMA_signal_6161, SubBytesIns_Inst_Sbox_9_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M37_U1 ( .a ({new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_9_M21}), .b ({new_AGEMA_signal_6158, SubBytesIns_Inst_Sbox_9_M29}), .c ({new_AGEMA_signal_6245, SubBytesIns_Inst_Sbox_9_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M38_U1 ( .a ({new_AGEMA_signal_6160, SubBytesIns_Inst_Sbox_9_M32}), .b ({new_AGEMA_signal_6062, SubBytesIns_Inst_Sbox_9_M33}), .c ({new_AGEMA_signal_6246, SubBytesIns_Inst_Sbox_9_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M39_U1 ( .a ({new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_9_M23}), .b ({new_AGEMA_signal_6159, SubBytesIns_Inst_Sbox_9_M30}), .c ({new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_9_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M40_U1 ( .a ({new_AGEMA_signal_6161, SubBytesIns_Inst_Sbox_9_M35}), .b ({new_AGEMA_signal_6162, SubBytesIns_Inst_Sbox_9_M36}), .c ({new_AGEMA_signal_6248, SubBytesIns_Inst_Sbox_9_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M41_U1 ( .a ({new_AGEMA_signal_6246, SubBytesIns_Inst_Sbox_9_M38}), .b ({new_AGEMA_signal_6248, SubBytesIns_Inst_Sbox_9_M40}), .c ({new_AGEMA_signal_6429, SubBytesIns_Inst_Sbox_9_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M42_U1 ( .a ({new_AGEMA_signal_6245, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_9_M39}), .c ({new_AGEMA_signal_6430, SubBytesIns_Inst_Sbox_9_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M43_U1 ( .a ({new_AGEMA_signal_6245, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_6246, SubBytesIns_Inst_Sbox_9_M38}), .c ({new_AGEMA_signal_6431, SubBytesIns_Inst_Sbox_9_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M44_U1 ( .a ({new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_9_M39}), .b ({new_AGEMA_signal_6248, SubBytesIns_Inst_Sbox_9_M40}), .c ({new_AGEMA_signal_6432, SubBytesIns_Inst_Sbox_9_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M45_U1 ( .a ({new_AGEMA_signal_6430, SubBytesIns_Inst_Sbox_9_M42}), .b ({new_AGEMA_signal_6429, SubBytesIns_Inst_Sbox_9_M41}), .c ({new_AGEMA_signal_6669, SubBytesIns_Inst_Sbox_9_M45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M29_U1 ( .a ({new_AGEMA_signal_6065, SubBytesIns_Inst_Sbox_10_M28}), .b ({new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_10_M27}), .clk (clk), .r (Fresh[280]), .c ({new_AGEMA_signal_6163, SubBytesIns_Inst_Sbox_10_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M30_U1 ( .a ({new_AGEMA_signal_6064, SubBytesIns_Inst_Sbox_10_M26}), .b ({new_AGEMA_signal_6063, SubBytesIns_Inst_Sbox_10_M24}), .clk (clk), .r (Fresh[281]), .c ({new_AGEMA_signal_6164, SubBytesIns_Inst_Sbox_10_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M32_U1 ( .a ({new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_10_M27}), .b ({new_AGEMA_signal_6066, SubBytesIns_Inst_Sbox_10_M31}), .clk (clk), .r (Fresh[282]), .c ({new_AGEMA_signal_6165, SubBytesIns_Inst_Sbox_10_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M35_U1 ( .a ({new_AGEMA_signal_6063, SubBytesIns_Inst_Sbox_10_M24}), .b ({new_AGEMA_signal_5972, SubBytesIns_Inst_Sbox_10_M34}), .clk (clk), .r (Fresh[283]), .c ({new_AGEMA_signal_6166, SubBytesIns_Inst_Sbox_10_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M37_U1 ( .a ({new_AGEMA_signal_5891, SubBytesIns_Inst_Sbox_10_M21}), .b ({new_AGEMA_signal_6163, SubBytesIns_Inst_Sbox_10_M29}), .c ({new_AGEMA_signal_6249, SubBytesIns_Inst_Sbox_10_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M38_U1 ( .a ({new_AGEMA_signal_6165, SubBytesIns_Inst_Sbox_10_M32}), .b ({new_AGEMA_signal_6067, SubBytesIns_Inst_Sbox_10_M33}), .c ({new_AGEMA_signal_6250, SubBytesIns_Inst_Sbox_10_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M39_U1 ( .a ({new_AGEMA_signal_5969, SubBytesIns_Inst_Sbox_10_M23}), .b ({new_AGEMA_signal_6164, SubBytesIns_Inst_Sbox_10_M30}), .c ({new_AGEMA_signal_6251, SubBytesIns_Inst_Sbox_10_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M40_U1 ( .a ({new_AGEMA_signal_6166, SubBytesIns_Inst_Sbox_10_M35}), .b ({new_AGEMA_signal_6167, SubBytesIns_Inst_Sbox_10_M36}), .c ({new_AGEMA_signal_6252, SubBytesIns_Inst_Sbox_10_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M41_U1 ( .a ({new_AGEMA_signal_6250, SubBytesIns_Inst_Sbox_10_M38}), .b ({new_AGEMA_signal_6252, SubBytesIns_Inst_Sbox_10_M40}), .c ({new_AGEMA_signal_6441, SubBytesIns_Inst_Sbox_10_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M42_U1 ( .a ({new_AGEMA_signal_6249, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_6251, SubBytesIns_Inst_Sbox_10_M39}), .c ({new_AGEMA_signal_6442, SubBytesIns_Inst_Sbox_10_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M43_U1 ( .a ({new_AGEMA_signal_6249, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_6250, SubBytesIns_Inst_Sbox_10_M38}), .c ({new_AGEMA_signal_6443, SubBytesIns_Inst_Sbox_10_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M44_U1 ( .a ({new_AGEMA_signal_6251, SubBytesIns_Inst_Sbox_10_M39}), .b ({new_AGEMA_signal_6252, SubBytesIns_Inst_Sbox_10_M40}), .c ({new_AGEMA_signal_6444, SubBytesIns_Inst_Sbox_10_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M45_U1 ( .a ({new_AGEMA_signal_6442, SubBytesIns_Inst_Sbox_10_M42}), .b ({new_AGEMA_signal_6441, SubBytesIns_Inst_Sbox_10_M41}), .c ({new_AGEMA_signal_6681, SubBytesIns_Inst_Sbox_10_M45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M29_U1 ( .a ({new_AGEMA_signal_6070, SubBytesIns_Inst_Sbox_11_M28}), .b ({new_AGEMA_signal_5975, SubBytesIns_Inst_Sbox_11_M27}), .clk (clk), .r (Fresh[284]), .c ({new_AGEMA_signal_6168, SubBytesIns_Inst_Sbox_11_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M30_U1 ( .a ({new_AGEMA_signal_6069, SubBytesIns_Inst_Sbox_11_M26}), .b ({new_AGEMA_signal_6068, SubBytesIns_Inst_Sbox_11_M24}), .clk (clk), .r (Fresh[285]), .c ({new_AGEMA_signal_6169, SubBytesIns_Inst_Sbox_11_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M32_U1 ( .a ({new_AGEMA_signal_5975, SubBytesIns_Inst_Sbox_11_M27}), .b ({new_AGEMA_signal_6071, SubBytesIns_Inst_Sbox_11_M31}), .clk (clk), .r (Fresh[286]), .c ({new_AGEMA_signal_6170, SubBytesIns_Inst_Sbox_11_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M35_U1 ( .a ({new_AGEMA_signal_6068, SubBytesIns_Inst_Sbox_11_M24}), .b ({new_AGEMA_signal_5976, SubBytesIns_Inst_Sbox_11_M34}), .clk (clk), .r (Fresh[287]), .c ({new_AGEMA_signal_6171, SubBytesIns_Inst_Sbox_11_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M37_U1 ( .a ({new_AGEMA_signal_5895, SubBytesIns_Inst_Sbox_11_M21}), .b ({new_AGEMA_signal_6168, SubBytesIns_Inst_Sbox_11_M29}), .c ({new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_11_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M38_U1 ( .a ({new_AGEMA_signal_6170, SubBytesIns_Inst_Sbox_11_M32}), .b ({new_AGEMA_signal_6072, SubBytesIns_Inst_Sbox_11_M33}), .c ({new_AGEMA_signal_6254, SubBytesIns_Inst_Sbox_11_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M39_U1 ( .a ({new_AGEMA_signal_5973, SubBytesIns_Inst_Sbox_11_M23}), .b ({new_AGEMA_signal_6169, SubBytesIns_Inst_Sbox_11_M30}), .c ({new_AGEMA_signal_6255, SubBytesIns_Inst_Sbox_11_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M40_U1 ( .a ({new_AGEMA_signal_6171, SubBytesIns_Inst_Sbox_11_M35}), .b ({new_AGEMA_signal_6172, SubBytesIns_Inst_Sbox_11_M36}), .c ({new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_11_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M41_U1 ( .a ({new_AGEMA_signal_6254, SubBytesIns_Inst_Sbox_11_M38}), .b ({new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_11_M40}), .c ({new_AGEMA_signal_6453, SubBytesIns_Inst_Sbox_11_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M42_U1 ( .a ({new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_6255, SubBytesIns_Inst_Sbox_11_M39}), .c ({new_AGEMA_signal_6454, SubBytesIns_Inst_Sbox_11_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M43_U1 ( .a ({new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_6254, SubBytesIns_Inst_Sbox_11_M38}), .c ({new_AGEMA_signal_6455, SubBytesIns_Inst_Sbox_11_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M44_U1 ( .a ({new_AGEMA_signal_6255, SubBytesIns_Inst_Sbox_11_M39}), .b ({new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_11_M40}), .c ({new_AGEMA_signal_6456, SubBytesIns_Inst_Sbox_11_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M45_U1 ( .a ({new_AGEMA_signal_6454, SubBytesIns_Inst_Sbox_11_M42}), .b ({new_AGEMA_signal_6453, SubBytesIns_Inst_Sbox_11_M41}), .c ({new_AGEMA_signal_6693, SubBytesIns_Inst_Sbox_11_M45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M29_U1 ( .a ({new_AGEMA_signal_6075, SubBytesIns_Inst_Sbox_12_M28}), .b ({new_AGEMA_signal_5979, SubBytesIns_Inst_Sbox_12_M27}), .clk (clk), .r (Fresh[288]), .c ({new_AGEMA_signal_6173, SubBytesIns_Inst_Sbox_12_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M30_U1 ( .a ({new_AGEMA_signal_6074, SubBytesIns_Inst_Sbox_12_M26}), .b ({new_AGEMA_signal_6073, SubBytesIns_Inst_Sbox_12_M24}), .clk (clk), .r (Fresh[289]), .c ({new_AGEMA_signal_6174, SubBytesIns_Inst_Sbox_12_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M32_U1 ( .a ({new_AGEMA_signal_5979, SubBytesIns_Inst_Sbox_12_M27}), .b ({new_AGEMA_signal_6076, SubBytesIns_Inst_Sbox_12_M31}), .clk (clk), .r (Fresh[290]), .c ({new_AGEMA_signal_6175, SubBytesIns_Inst_Sbox_12_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M35_U1 ( .a ({new_AGEMA_signal_6073, SubBytesIns_Inst_Sbox_12_M24}), .b ({new_AGEMA_signal_5980, SubBytesIns_Inst_Sbox_12_M34}), .clk (clk), .r (Fresh[291]), .c ({new_AGEMA_signal_6176, SubBytesIns_Inst_Sbox_12_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M37_U1 ( .a ({new_AGEMA_signal_5899, SubBytesIns_Inst_Sbox_12_M21}), .b ({new_AGEMA_signal_6173, SubBytesIns_Inst_Sbox_12_M29}), .c ({new_AGEMA_signal_6257, SubBytesIns_Inst_Sbox_12_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M38_U1 ( .a ({new_AGEMA_signal_6175, SubBytesIns_Inst_Sbox_12_M32}), .b ({new_AGEMA_signal_6077, SubBytesIns_Inst_Sbox_12_M33}), .c ({new_AGEMA_signal_6258, SubBytesIns_Inst_Sbox_12_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M39_U1 ( .a ({new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_12_M23}), .b ({new_AGEMA_signal_6174, SubBytesIns_Inst_Sbox_12_M30}), .c ({new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_12_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M40_U1 ( .a ({new_AGEMA_signal_6176, SubBytesIns_Inst_Sbox_12_M35}), .b ({new_AGEMA_signal_6177, SubBytesIns_Inst_Sbox_12_M36}), .c ({new_AGEMA_signal_6260, SubBytesIns_Inst_Sbox_12_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M41_U1 ( .a ({new_AGEMA_signal_6258, SubBytesIns_Inst_Sbox_12_M38}), .b ({new_AGEMA_signal_6260, SubBytesIns_Inst_Sbox_12_M40}), .c ({new_AGEMA_signal_6465, SubBytesIns_Inst_Sbox_12_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M42_U1 ( .a ({new_AGEMA_signal_6257, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_12_M39}), .c ({new_AGEMA_signal_6466, SubBytesIns_Inst_Sbox_12_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M43_U1 ( .a ({new_AGEMA_signal_6257, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_6258, SubBytesIns_Inst_Sbox_12_M38}), .c ({new_AGEMA_signal_6467, SubBytesIns_Inst_Sbox_12_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M44_U1 ( .a ({new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_12_M39}), .b ({new_AGEMA_signal_6260, SubBytesIns_Inst_Sbox_12_M40}), .c ({new_AGEMA_signal_6468, SubBytesIns_Inst_Sbox_12_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M45_U1 ( .a ({new_AGEMA_signal_6466, SubBytesIns_Inst_Sbox_12_M42}), .b ({new_AGEMA_signal_6465, SubBytesIns_Inst_Sbox_12_M41}), .c ({new_AGEMA_signal_6705, SubBytesIns_Inst_Sbox_12_M45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M29_U1 ( .a ({new_AGEMA_signal_6080, SubBytesIns_Inst_Sbox_13_M28}), .b ({new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_13_M27}), .clk (clk), .r (Fresh[292]), .c ({new_AGEMA_signal_6178, SubBytesIns_Inst_Sbox_13_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M30_U1 ( .a ({new_AGEMA_signal_6079, SubBytesIns_Inst_Sbox_13_M26}), .b ({new_AGEMA_signal_6078, SubBytesIns_Inst_Sbox_13_M24}), .clk (clk), .r (Fresh[293]), .c ({new_AGEMA_signal_6179, SubBytesIns_Inst_Sbox_13_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M32_U1 ( .a ({new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_13_M27}), .b ({new_AGEMA_signal_6081, SubBytesIns_Inst_Sbox_13_M31}), .clk (clk), .r (Fresh[294]), .c ({new_AGEMA_signal_6180, SubBytesIns_Inst_Sbox_13_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M35_U1 ( .a ({new_AGEMA_signal_6078, SubBytesIns_Inst_Sbox_13_M24}), .b ({new_AGEMA_signal_5984, SubBytesIns_Inst_Sbox_13_M34}), .clk (clk), .r (Fresh[295]), .c ({new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_13_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M37_U1 ( .a ({new_AGEMA_signal_5903, SubBytesIns_Inst_Sbox_13_M21}), .b ({new_AGEMA_signal_6178, SubBytesIns_Inst_Sbox_13_M29}), .c ({new_AGEMA_signal_6261, SubBytesIns_Inst_Sbox_13_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M38_U1 ( .a ({new_AGEMA_signal_6180, SubBytesIns_Inst_Sbox_13_M32}), .b ({new_AGEMA_signal_6082, SubBytesIns_Inst_Sbox_13_M33}), .c ({new_AGEMA_signal_6262, SubBytesIns_Inst_Sbox_13_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M39_U1 ( .a ({new_AGEMA_signal_5981, SubBytesIns_Inst_Sbox_13_M23}), .b ({new_AGEMA_signal_6179, SubBytesIns_Inst_Sbox_13_M30}), .c ({new_AGEMA_signal_6263, SubBytesIns_Inst_Sbox_13_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M40_U1 ( .a ({new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_13_M35}), .b ({new_AGEMA_signal_6182, SubBytesIns_Inst_Sbox_13_M36}), .c ({new_AGEMA_signal_6264, SubBytesIns_Inst_Sbox_13_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M41_U1 ( .a ({new_AGEMA_signal_6262, SubBytesIns_Inst_Sbox_13_M38}), .b ({new_AGEMA_signal_6264, SubBytesIns_Inst_Sbox_13_M40}), .c ({new_AGEMA_signal_6477, SubBytesIns_Inst_Sbox_13_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M42_U1 ( .a ({new_AGEMA_signal_6261, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_6263, SubBytesIns_Inst_Sbox_13_M39}), .c ({new_AGEMA_signal_6478, SubBytesIns_Inst_Sbox_13_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M43_U1 ( .a ({new_AGEMA_signal_6261, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_6262, SubBytesIns_Inst_Sbox_13_M38}), .c ({new_AGEMA_signal_6479, SubBytesIns_Inst_Sbox_13_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M44_U1 ( .a ({new_AGEMA_signal_6263, SubBytesIns_Inst_Sbox_13_M39}), .b ({new_AGEMA_signal_6264, SubBytesIns_Inst_Sbox_13_M40}), .c ({new_AGEMA_signal_6480, SubBytesIns_Inst_Sbox_13_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M45_U1 ( .a ({new_AGEMA_signal_6478, SubBytesIns_Inst_Sbox_13_M42}), .b ({new_AGEMA_signal_6477, SubBytesIns_Inst_Sbox_13_M41}), .c ({new_AGEMA_signal_6717, SubBytesIns_Inst_Sbox_13_M45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M29_U1 ( .a ({new_AGEMA_signal_6085, SubBytesIns_Inst_Sbox_14_M28}), .b ({new_AGEMA_signal_5987, SubBytesIns_Inst_Sbox_14_M27}), .clk (clk), .r (Fresh[296]), .c ({new_AGEMA_signal_6183, SubBytesIns_Inst_Sbox_14_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M30_U1 ( .a ({new_AGEMA_signal_6084, SubBytesIns_Inst_Sbox_14_M26}), .b ({new_AGEMA_signal_6083, SubBytesIns_Inst_Sbox_14_M24}), .clk (clk), .r (Fresh[297]), .c ({new_AGEMA_signal_6184, SubBytesIns_Inst_Sbox_14_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M32_U1 ( .a ({new_AGEMA_signal_5987, SubBytesIns_Inst_Sbox_14_M27}), .b ({new_AGEMA_signal_6086, SubBytesIns_Inst_Sbox_14_M31}), .clk (clk), .r (Fresh[298]), .c ({new_AGEMA_signal_6185, SubBytesIns_Inst_Sbox_14_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M35_U1 ( .a ({new_AGEMA_signal_6083, SubBytesIns_Inst_Sbox_14_M24}), .b ({new_AGEMA_signal_5988, SubBytesIns_Inst_Sbox_14_M34}), .clk (clk), .r (Fresh[299]), .c ({new_AGEMA_signal_6186, SubBytesIns_Inst_Sbox_14_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M37_U1 ( .a ({new_AGEMA_signal_5907, SubBytesIns_Inst_Sbox_14_M21}), .b ({new_AGEMA_signal_6183, SubBytesIns_Inst_Sbox_14_M29}), .c ({new_AGEMA_signal_6265, SubBytesIns_Inst_Sbox_14_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M38_U1 ( .a ({new_AGEMA_signal_6185, SubBytesIns_Inst_Sbox_14_M32}), .b ({new_AGEMA_signal_6087, SubBytesIns_Inst_Sbox_14_M33}), .c ({new_AGEMA_signal_6266, SubBytesIns_Inst_Sbox_14_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M39_U1 ( .a ({new_AGEMA_signal_5985, SubBytesIns_Inst_Sbox_14_M23}), .b ({new_AGEMA_signal_6184, SubBytesIns_Inst_Sbox_14_M30}), .c ({new_AGEMA_signal_6267, SubBytesIns_Inst_Sbox_14_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M40_U1 ( .a ({new_AGEMA_signal_6186, SubBytesIns_Inst_Sbox_14_M35}), .b ({new_AGEMA_signal_6187, SubBytesIns_Inst_Sbox_14_M36}), .c ({new_AGEMA_signal_6268, SubBytesIns_Inst_Sbox_14_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M41_U1 ( .a ({new_AGEMA_signal_6266, SubBytesIns_Inst_Sbox_14_M38}), .b ({new_AGEMA_signal_6268, SubBytesIns_Inst_Sbox_14_M40}), .c ({new_AGEMA_signal_6489, SubBytesIns_Inst_Sbox_14_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M42_U1 ( .a ({new_AGEMA_signal_6265, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_6267, SubBytesIns_Inst_Sbox_14_M39}), .c ({new_AGEMA_signal_6490, SubBytesIns_Inst_Sbox_14_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M43_U1 ( .a ({new_AGEMA_signal_6265, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_6266, SubBytesIns_Inst_Sbox_14_M38}), .c ({new_AGEMA_signal_6491, SubBytesIns_Inst_Sbox_14_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M44_U1 ( .a ({new_AGEMA_signal_6267, SubBytesIns_Inst_Sbox_14_M39}), .b ({new_AGEMA_signal_6268, SubBytesIns_Inst_Sbox_14_M40}), .c ({new_AGEMA_signal_6492, SubBytesIns_Inst_Sbox_14_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M45_U1 ( .a ({new_AGEMA_signal_6490, SubBytesIns_Inst_Sbox_14_M42}), .b ({new_AGEMA_signal_6489, SubBytesIns_Inst_Sbox_14_M41}), .c ({new_AGEMA_signal_6729, SubBytesIns_Inst_Sbox_14_M45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M29_U1 ( .a ({new_AGEMA_signal_6090, SubBytesIns_Inst_Sbox_15_M28}), .b ({new_AGEMA_signal_5991, SubBytesIns_Inst_Sbox_15_M27}), .clk (clk), .r (Fresh[300]), .c ({new_AGEMA_signal_6188, SubBytesIns_Inst_Sbox_15_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M30_U1 ( .a ({new_AGEMA_signal_6089, SubBytesIns_Inst_Sbox_15_M26}), .b ({new_AGEMA_signal_6088, SubBytesIns_Inst_Sbox_15_M24}), .clk (clk), .r (Fresh[301]), .c ({new_AGEMA_signal_6189, SubBytesIns_Inst_Sbox_15_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M32_U1 ( .a ({new_AGEMA_signal_5991, SubBytesIns_Inst_Sbox_15_M27}), .b ({new_AGEMA_signal_6091, SubBytesIns_Inst_Sbox_15_M31}), .clk (clk), .r (Fresh[302]), .c ({new_AGEMA_signal_6190, SubBytesIns_Inst_Sbox_15_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M35_U1 ( .a ({new_AGEMA_signal_6088, SubBytesIns_Inst_Sbox_15_M24}), .b ({new_AGEMA_signal_5992, SubBytesIns_Inst_Sbox_15_M34}), .clk (clk), .r (Fresh[303]), .c ({new_AGEMA_signal_6191, SubBytesIns_Inst_Sbox_15_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M37_U1 ( .a ({new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_15_M21}), .b ({new_AGEMA_signal_6188, SubBytesIns_Inst_Sbox_15_M29}), .c ({new_AGEMA_signal_6269, SubBytesIns_Inst_Sbox_15_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M38_U1 ( .a ({new_AGEMA_signal_6190, SubBytesIns_Inst_Sbox_15_M32}), .b ({new_AGEMA_signal_6092, SubBytesIns_Inst_Sbox_15_M33}), .c ({new_AGEMA_signal_6270, SubBytesIns_Inst_Sbox_15_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M39_U1 ( .a ({new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_15_M23}), .b ({new_AGEMA_signal_6189, SubBytesIns_Inst_Sbox_15_M30}), .c ({new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M40_U1 ( .a ({new_AGEMA_signal_6191, SubBytesIns_Inst_Sbox_15_M35}), .b ({new_AGEMA_signal_6192, SubBytesIns_Inst_Sbox_15_M36}), .c ({new_AGEMA_signal_6272, SubBytesIns_Inst_Sbox_15_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M41_U1 ( .a ({new_AGEMA_signal_6270, SubBytesIns_Inst_Sbox_15_M38}), .b ({new_AGEMA_signal_6272, SubBytesIns_Inst_Sbox_15_M40}), .c ({new_AGEMA_signal_6501, SubBytesIns_Inst_Sbox_15_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M42_U1 ( .a ({new_AGEMA_signal_6269, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_M39}), .c ({new_AGEMA_signal_6502, SubBytesIns_Inst_Sbox_15_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M43_U1 ( .a ({new_AGEMA_signal_6269, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_6270, SubBytesIns_Inst_Sbox_15_M38}), .c ({new_AGEMA_signal_6503, SubBytesIns_Inst_Sbox_15_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M44_U1 ( .a ({new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_M39}), .b ({new_AGEMA_signal_6272, SubBytesIns_Inst_Sbox_15_M40}), .c ({new_AGEMA_signal_6504, SubBytesIns_Inst_Sbox_15_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M45_U1 ( .a ({new_AGEMA_signal_6502, SubBytesIns_Inst_Sbox_15_M42}), .b ({new_AGEMA_signal_6501, SubBytesIns_Inst_Sbox_15_M41}), .c ({new_AGEMA_signal_6741, SubBytesIns_Inst_Sbox_15_M45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M29_U1 ( .a ({new_AGEMA_signal_5995, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28}), .b ({new_AGEMA_signal_5915, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27}), .clk (clk), .r (Fresh[304]), .c ({new_AGEMA_signal_6093, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M30_U1 ( .a ({new_AGEMA_signal_5994, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26}), .b ({new_AGEMA_signal_5993, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24}), .clk (clk), .r (Fresh[305]), .c ({new_AGEMA_signal_6094, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M32_U1 ( .a ({new_AGEMA_signal_5915, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27}), .b ({new_AGEMA_signal_5996, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31}), .clk (clk), .r (Fresh[306]), .c ({new_AGEMA_signal_6095, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M35_U1 ( .a ({new_AGEMA_signal_5993, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24}), .b ({new_AGEMA_signal_5916, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34}), .clk (clk), .r (Fresh[307]), .c ({new_AGEMA_signal_6096, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M37_U1 ( .a ({new_AGEMA_signal_5835, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_6093, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29}), .c ({new_AGEMA_signal_6193, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M38_U1 ( .a ({new_AGEMA_signal_6095, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32}), .b ({new_AGEMA_signal_5997, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33}), .c ({new_AGEMA_signal_6194, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M39_U1 ( .a ({new_AGEMA_signal_5913, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}), .b ({new_AGEMA_signal_6094, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30}), .c ({new_AGEMA_signal_6195, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M40_U1 ( .a ({new_AGEMA_signal_6096, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35}), .b ({new_AGEMA_signal_6097, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36}), .c ({new_AGEMA_signal_6196, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M41_U1 ( .a ({new_AGEMA_signal_6194, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_6196, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_6273, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M42_U1 ( .a ({new_AGEMA_signal_6193, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_6195, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .c ({new_AGEMA_signal_6274, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M43_U1 ( .a ({new_AGEMA_signal_6193, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_6194, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .c ({new_AGEMA_signal_6275, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M44_U1 ( .a ({new_AGEMA_signal_6195, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_6196, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_6276, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M45_U1 ( .a ({new_AGEMA_signal_6274, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_6273, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}), .c ({new_AGEMA_signal_6513, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M29_U1 ( .a ({new_AGEMA_signal_6000, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28}), .b ({new_AGEMA_signal_5919, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27}), .clk (clk), .r (Fresh[308]), .c ({new_AGEMA_signal_6098, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M30_U1 ( .a ({new_AGEMA_signal_5999, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26}), .b ({new_AGEMA_signal_5998, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24}), .clk (clk), .r (Fresh[309]), .c ({new_AGEMA_signal_6099, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M32_U1 ( .a ({new_AGEMA_signal_5919, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27}), .b ({new_AGEMA_signal_6001, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31}), .clk (clk), .r (Fresh[310]), .c ({new_AGEMA_signal_6100, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M35_U1 ( .a ({new_AGEMA_signal_5998, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24}), .b ({new_AGEMA_signal_5920, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34}), .clk (clk), .r (Fresh[311]), .c ({new_AGEMA_signal_6101, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M37_U1 ( .a ({new_AGEMA_signal_5839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_6098, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29}), .c ({new_AGEMA_signal_6197, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M38_U1 ( .a ({new_AGEMA_signal_6100, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32}), .b ({new_AGEMA_signal_6002, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33}), .c ({new_AGEMA_signal_6198, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M39_U1 ( .a ({new_AGEMA_signal_5917, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}), .b ({new_AGEMA_signal_6099, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30}), .c ({new_AGEMA_signal_6199, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M40_U1 ( .a ({new_AGEMA_signal_6101, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35}), .b ({new_AGEMA_signal_6102, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36}), .c ({new_AGEMA_signal_6200, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M41_U1 ( .a ({new_AGEMA_signal_6198, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_6200, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_6285, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M42_U1 ( .a ({new_AGEMA_signal_6197, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_6199, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .c ({new_AGEMA_signal_6286, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M43_U1 ( .a ({new_AGEMA_signal_6197, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_6198, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .c ({new_AGEMA_signal_6287, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M44_U1 ( .a ({new_AGEMA_signal_6199, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_6200, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_6288, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M45_U1 ( .a ({new_AGEMA_signal_6286, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_6285, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}), .c ({new_AGEMA_signal_6525, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M29_U1 ( .a ({new_AGEMA_signal_6005, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28}), .b ({new_AGEMA_signal_5923, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27}), .clk (clk), .r (Fresh[312]), .c ({new_AGEMA_signal_6103, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M30_U1 ( .a ({new_AGEMA_signal_6004, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26}), .b ({new_AGEMA_signal_6003, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24}), .clk (clk), .r (Fresh[313]), .c ({new_AGEMA_signal_6104, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M32_U1 ( .a ({new_AGEMA_signal_5923, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27}), .b ({new_AGEMA_signal_6006, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31}), .clk (clk), .r (Fresh[314]), .c ({new_AGEMA_signal_6105, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M35_U1 ( .a ({new_AGEMA_signal_6003, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24}), .b ({new_AGEMA_signal_5924, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34}), .clk (clk), .r (Fresh[315]), .c ({new_AGEMA_signal_6106, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M37_U1 ( .a ({new_AGEMA_signal_5843, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_6103, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29}), .c ({new_AGEMA_signal_6201, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M38_U1 ( .a ({new_AGEMA_signal_6105, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32}), .b ({new_AGEMA_signal_6007, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33}), .c ({new_AGEMA_signal_6202, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M39_U1 ( .a ({new_AGEMA_signal_5921, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}), .b ({new_AGEMA_signal_6104, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30}), .c ({new_AGEMA_signal_6203, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M40_U1 ( .a ({new_AGEMA_signal_6106, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35}), .b ({new_AGEMA_signal_6107, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36}), .c ({new_AGEMA_signal_6204, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M41_U1 ( .a ({new_AGEMA_signal_6202, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_6204, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_6297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M42_U1 ( .a ({new_AGEMA_signal_6201, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_6203, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .c ({new_AGEMA_signal_6298, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M43_U1 ( .a ({new_AGEMA_signal_6201, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_6202, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .c ({new_AGEMA_signal_6299, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M44_U1 ( .a ({new_AGEMA_signal_6203, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_6204, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_6300, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M45_U1 ( .a ({new_AGEMA_signal_6298, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_6297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}), .c ({new_AGEMA_signal_6537, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M29_U1 ( .a ({new_AGEMA_signal_6010, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28}), .b ({new_AGEMA_signal_5927, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27}), .clk (clk), .r (Fresh[316]), .c ({new_AGEMA_signal_6108, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M30_U1 ( .a ({new_AGEMA_signal_6009, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26}), .b ({new_AGEMA_signal_6008, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24}), .clk (clk), .r (Fresh[317]), .c ({new_AGEMA_signal_6109, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M32_U1 ( .a ({new_AGEMA_signal_5927, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27}), .b ({new_AGEMA_signal_6011, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31}), .clk (clk), .r (Fresh[318]), .c ({new_AGEMA_signal_6110, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M35_U1 ( .a ({new_AGEMA_signal_6008, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24}), .b ({new_AGEMA_signal_5928, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34}), .clk (clk), .r (Fresh[319]), .c ({new_AGEMA_signal_6111, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M37_U1 ( .a ({new_AGEMA_signal_5847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_6108, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29}), .c ({new_AGEMA_signal_6205, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M38_U1 ( .a ({new_AGEMA_signal_6110, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32}), .b ({new_AGEMA_signal_6012, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33}), .c ({new_AGEMA_signal_6206, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M39_U1 ( .a ({new_AGEMA_signal_5925, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}), .b ({new_AGEMA_signal_6109, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30}), .c ({new_AGEMA_signal_6207, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M40_U1 ( .a ({new_AGEMA_signal_6111, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35}), .b ({new_AGEMA_signal_6112, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36}), .c ({new_AGEMA_signal_6208, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M41_U1 ( .a ({new_AGEMA_signal_6206, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_6208, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_6309, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M42_U1 ( .a ({new_AGEMA_signal_6205, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_6207, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .c ({new_AGEMA_signal_6310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M43_U1 ( .a ({new_AGEMA_signal_6205, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_6206, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .c ({new_AGEMA_signal_6311, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M44_U1 ( .a ({new_AGEMA_signal_6207, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_6208, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_6312, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M45_U1 ( .a ({new_AGEMA_signal_6310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_6309, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}), .c ({new_AGEMA_signal_6549, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_masked #(.security_order(1), .pipeline(0)) U858 ( .s (n321), .b ({new_AGEMA_signal_7231, MixColumnsInput[0]}), .a ({new_AGEMA_signal_8096, MixColumnsOutput[0]}), .c ({new_AGEMA_signal_8190, RoundOutput[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U859 ( .s (n321), .b ({new_AGEMA_signal_7388, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .a ({new_AGEMA_signal_8271, MixColumnsOutput[100]}), .c ({new_AGEMA_signal_8383, RoundOutput[100]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U860 ( .s (n321), .b ({new_AGEMA_signal_7387, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .a ({new_AGEMA_signal_7973, MixColumnsOutput[101]}), .c ({new_AGEMA_signal_8191, RoundOutput[101]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U861 ( .s (n321), .b ({new_AGEMA_signal_7386, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .a ({new_AGEMA_signal_7972, MixColumnsOutput[102]}), .c ({new_AGEMA_signal_8192, RoundOutput[102]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U862 ( .s (n321), .b ({new_AGEMA_signal_7385, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .a ({new_AGEMA_signal_7971, MixColumnsOutput[103]}), .c ({new_AGEMA_signal_8193, RoundOutput[103]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U863 ( .s (n321), .b ({new_AGEMA_signal_7242, MixColumnsInput[104]}), .a ({new_AGEMA_signal_7970, MixColumnsOutput[104]}), .c ({new_AGEMA_signal_8194, RoundOutput[104]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U864 ( .s (n321), .b ({new_AGEMA_signal_7426, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .a ({new_AGEMA_signal_8270, MixColumnsOutput[105]}), .c ({new_AGEMA_signal_8384, RoundOutput[105]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U865 ( .s (n321), .b ({new_AGEMA_signal_7425, MixColumnsInput[106]}), .a ({new_AGEMA_signal_7999, MixColumnsOutput[106]}), .c ({new_AGEMA_signal_8195, RoundOutput[106]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U866 ( .s (n315), .b ({new_AGEMA_signal_7424, MixColumnsInput[107]}), .a ({new_AGEMA_signal_8281, MixColumnsOutput[107]}), .c ({new_AGEMA_signal_8385, RoundOutput[107]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U867 ( .s (n316), .b ({new_AGEMA_signal_7423, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .a ({new_AGEMA_signal_8280, MixColumnsOutput[108]}), .c ({new_AGEMA_signal_8386, RoundOutput[108]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U868 ( .s (n317), .b ({new_AGEMA_signal_7422, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .a ({new_AGEMA_signal_7996, MixColumnsOutput[109]}), .c ({new_AGEMA_signal_8196, RoundOutput[109]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U869 ( .s (n318), .b ({new_AGEMA_signal_7453, MixColumnsInput[10]}), .a ({new_AGEMA_signal_8095, MixColumnsOutput[10]}), .c ({new_AGEMA_signal_8197, RoundOutput[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U870 ( .s (n319), .b ({new_AGEMA_signal_7421, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .a ({new_AGEMA_signal_7995, MixColumnsOutput[110]}), .c ({new_AGEMA_signal_8198, RoundOutput[110]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U871 ( .s (n320), .b ({new_AGEMA_signal_7420, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .a ({new_AGEMA_signal_7994, MixColumnsOutput[111]}), .c ({new_AGEMA_signal_8199, RoundOutput[111]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U872 ( .s (n319), .b ({new_AGEMA_signal_7297, MixColumnsInput[112]}), .a ({new_AGEMA_signal_7993, MixColumnsOutput[112]}), .c ({new_AGEMA_signal_8200, RoundOutput[112]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U873 ( .s (n318), .b ({new_AGEMA_signal_7461, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .a ({new_AGEMA_signal_8279, MixColumnsOutput[113]}), .c ({new_AGEMA_signal_8387, RoundOutput[113]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U874 ( .s (n318), .b ({new_AGEMA_signal_7460, MixColumnsInput[114]}), .a ({new_AGEMA_signal_7991, MixColumnsOutput[114]}), .c ({new_AGEMA_signal_8201, RoundOutput[114]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U875 ( .s (n315), .b ({new_AGEMA_signal_7459, MixColumnsInput[115]}), .a ({new_AGEMA_signal_8278, MixColumnsOutput[115]}), .c ({new_AGEMA_signal_8388, RoundOutput[115]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U876 ( .s (n316), .b ({new_AGEMA_signal_7458, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .a ({new_AGEMA_signal_8276, MixColumnsOutput[116]}), .c ({new_AGEMA_signal_8389, RoundOutput[116]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U877 ( .s (n317), .b ({new_AGEMA_signal_7457, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .a ({new_AGEMA_signal_7987, MixColumnsOutput[117]}), .c ({new_AGEMA_signal_8202, RoundOutput[117]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U878 ( .s (n319), .b ({new_AGEMA_signal_7456, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .a ({new_AGEMA_signal_7986, MixColumnsOutput[118]}), .c ({new_AGEMA_signal_8203, RoundOutput[118]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U879 ( .s (n320), .b ({new_AGEMA_signal_7455, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .a ({new_AGEMA_signal_7985, MixColumnsOutput[119]}), .c ({new_AGEMA_signal_8204, RoundOutput[119]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U880 ( .s (n320), .b ({new_AGEMA_signal_7452, MixColumnsInput[11]}), .a ({new_AGEMA_signal_8317, MixColumnsOutput[11]}), .c ({new_AGEMA_signal_8390, RoundOutput[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U881 ( .s (n319), .b ({new_AGEMA_signal_7352, MixColumnsInput[120]}), .a ({new_AGEMA_signal_7984, MixColumnsOutput[120]}), .c ({new_AGEMA_signal_8205, RoundOutput[120]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U882 ( .s (n318), .b ({new_AGEMA_signal_7496, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .a ({new_AGEMA_signal_8275, MixColumnsOutput[121]}), .c ({new_AGEMA_signal_8391, RoundOutput[121]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U883 ( .s (n319), .b ({new_AGEMA_signal_7495, MixColumnsInput[122]}), .a ({new_AGEMA_signal_7982, MixColumnsOutput[122]}), .c ({new_AGEMA_signal_8206, RoundOutput[122]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U884 ( .s (n320), .b ({new_AGEMA_signal_7494, MixColumnsInput[123]}), .a ({new_AGEMA_signal_8274, MixColumnsOutput[123]}), .c ({new_AGEMA_signal_8392, RoundOutput[123]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U885 ( .s (n316), .b ({new_AGEMA_signal_7493, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .a ({new_AGEMA_signal_8273, MixColumnsOutput[124]}), .c ({new_AGEMA_signal_8393, RoundOutput[124]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U886 ( .s (n320), .b ({new_AGEMA_signal_7492, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .a ({new_AGEMA_signal_7979, MixColumnsOutput[125]}), .c ({new_AGEMA_signal_8207, RoundOutput[125]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U887 ( .s (n316), .b ({new_AGEMA_signal_7491, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .a ({new_AGEMA_signal_7977, MixColumnsOutput[126]}), .c ({new_AGEMA_signal_8208, RoundOutput[126]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U888 ( .s (n317), .b ({new_AGEMA_signal_7490, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .a ({new_AGEMA_signal_7976, MixColumnsOutput[127]}), .c ({new_AGEMA_signal_8209, RoundOutput[127]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U889 ( .s (n315), .b ({new_AGEMA_signal_7451, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .a ({new_AGEMA_signal_8316, MixColumnsOutput[12]}), .c ({new_AGEMA_signal_8394, RoundOutput[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U890 ( .s (n317), .b ({new_AGEMA_signal_7450, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .a ({new_AGEMA_signal_8092, MixColumnsOutput[13]}), .c ({new_AGEMA_signal_8210, RoundOutput[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U891 ( .s (n316), .b ({new_AGEMA_signal_7449, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .a ({new_AGEMA_signal_8091, MixColumnsOutput[14]}), .c ({new_AGEMA_signal_8211, RoundOutput[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U892 ( .s (n317), .b ({new_AGEMA_signal_7448, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .a ({new_AGEMA_signal_8090, MixColumnsOutput[15]}), .c ({new_AGEMA_signal_8212, RoundOutput[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U893 ( .s (n315), .b ({new_AGEMA_signal_7341, MixColumnsInput[16]}), .a ({new_AGEMA_signal_8089, MixColumnsOutput[16]}), .c ({new_AGEMA_signal_8213, RoundOutput[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U894 ( .s (n318), .b ({new_AGEMA_signal_7489, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .a ({new_AGEMA_signal_8315, MixColumnsOutput[17]}), .c ({new_AGEMA_signal_8395, RoundOutput[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U895 ( .s (n319), .b ({new_AGEMA_signal_7488, MixColumnsInput[18]}), .a ({new_AGEMA_signal_8087, MixColumnsOutput[18]}), .c ({new_AGEMA_signal_8214, RoundOutput[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U896 ( .s (n320), .b ({new_AGEMA_signal_7487, MixColumnsInput[19]}), .a ({new_AGEMA_signal_8314, MixColumnsOutput[19]}), .c ({new_AGEMA_signal_8396, RoundOutput[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U897 ( .s (n318), .b ({new_AGEMA_signal_7419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .a ({new_AGEMA_signal_8313, MixColumnsOutput[1]}), .c ({new_AGEMA_signal_8397, RoundOutput[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U898 ( .s (n319), .b ({new_AGEMA_signal_7486, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .a ({new_AGEMA_signal_8312, MixColumnsOutput[20]}), .c ({new_AGEMA_signal_8398, RoundOutput[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U899 ( .s (n316), .b ({new_AGEMA_signal_7485, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .a ({new_AGEMA_signal_8083, MixColumnsOutput[21]}), .c ({new_AGEMA_signal_8215, RoundOutput[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U900 ( .s (n317), .b ({new_AGEMA_signal_7484, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .a ({new_AGEMA_signal_8082, MixColumnsOutput[22]}), .c ({new_AGEMA_signal_8216, RoundOutput[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U901 ( .s (n315), .b ({new_AGEMA_signal_7483, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .a ({new_AGEMA_signal_8081, MixColumnsOutput[23]}), .c ({new_AGEMA_signal_8217, RoundOutput[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U902 ( .s (n320), .b ({new_AGEMA_signal_7220, MixColumnsInput[24]}), .a ({new_AGEMA_signal_8080, MixColumnsOutput[24]}), .c ({new_AGEMA_signal_8218, RoundOutput[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U903 ( .s (n318), .b ({new_AGEMA_signal_7412, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .a ({new_AGEMA_signal_8311, MixColumnsOutput[25]}), .c ({new_AGEMA_signal_8399, RoundOutput[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U904 ( .s (n316), .b ({new_AGEMA_signal_7411, MixColumnsInput[26]}), .a ({new_AGEMA_signal_8078, MixColumnsOutput[26]}), .c ({new_AGEMA_signal_8219, RoundOutput[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U905 ( .s (n317), .b ({new_AGEMA_signal_7410, MixColumnsInput[27]}), .a ({new_AGEMA_signal_8310, MixColumnsOutput[27]}), .c ({new_AGEMA_signal_8400, RoundOutput[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U906 ( .s (n315), .b ({new_AGEMA_signal_7409, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .a ({new_AGEMA_signal_8309, MixColumnsOutput[28]}), .c ({new_AGEMA_signal_8401, RoundOutput[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U907 ( .s (n319), .b ({new_AGEMA_signal_7408, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .a ({new_AGEMA_signal_8075, MixColumnsOutput[29]}), .c ({new_AGEMA_signal_8220, RoundOutput[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U908 ( .s (n315), .b ({new_AGEMA_signal_7418, MixColumnsInput[2]}), .a ({new_AGEMA_signal_8074, MixColumnsOutput[2]}), .c ({new_AGEMA_signal_8221, RoundOutput[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U909 ( .s (n320), .b ({new_AGEMA_signal_7407, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .a ({new_AGEMA_signal_8073, MixColumnsOutput[30]}), .c ({new_AGEMA_signal_8222, RoundOutput[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U910 ( .s (n318), .b ({new_AGEMA_signal_7406, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .a ({new_AGEMA_signal_8072, MixColumnsOutput[31]}), .c ({new_AGEMA_signal_8223, RoundOutput[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U911 ( .s (n316), .b ({new_AGEMA_signal_7275, MixColumnsInput[32]}), .a ({new_AGEMA_signal_8064, MixColumnsOutput[32]}), .c ({new_AGEMA_signal_8224, RoundOutput[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U912 ( .s (n317), .b ({new_AGEMA_signal_7447, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .a ({new_AGEMA_signal_8301, MixColumnsOutput[33]}), .c ({new_AGEMA_signal_8402, RoundOutput[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U913 ( .s (n315), .b ({new_AGEMA_signal_7446, MixColumnsInput[34]}), .a ({new_AGEMA_signal_8042, MixColumnsOutput[34]}), .c ({new_AGEMA_signal_8225, RoundOutput[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U914 ( .s (n320), .b ({new_AGEMA_signal_7445, MixColumnsInput[35]}), .a ({new_AGEMA_signal_8296, MixColumnsOutput[35]}), .c ({new_AGEMA_signal_8403, RoundOutput[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U915 ( .s (n320), .b ({new_AGEMA_signal_7444, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .a ({new_AGEMA_signal_8295, MixColumnsOutput[36]}), .c ({new_AGEMA_signal_8404, RoundOutput[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U916 ( .s (n320), .b ({new_AGEMA_signal_7443, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .a ({new_AGEMA_signal_8037, MixColumnsOutput[37]}), .c ({new_AGEMA_signal_8226, RoundOutput[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U917 ( .s (n320), .b ({new_AGEMA_signal_7442, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .a ({new_AGEMA_signal_8036, MixColumnsOutput[38]}), .c ({new_AGEMA_signal_8227, RoundOutput[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U918 ( .s (n320), .b ({new_AGEMA_signal_7441, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .a ({new_AGEMA_signal_8035, MixColumnsOutput[39]}), .c ({new_AGEMA_signal_8228, RoundOutput[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U919 ( .s (n320), .b ({new_AGEMA_signal_7417, MixColumnsInput[3]}), .a ({new_AGEMA_signal_8308, MixColumnsOutput[3]}), .c ({new_AGEMA_signal_8405, RoundOutput[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U920 ( .s (n320), .b ({new_AGEMA_signal_7330, MixColumnsInput[40]}), .a ({new_AGEMA_signal_8034, MixColumnsOutput[40]}), .c ({new_AGEMA_signal_8229, RoundOutput[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U921 ( .s (n320), .b ({new_AGEMA_signal_7482, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .a ({new_AGEMA_signal_8294, MixColumnsOutput[41]}), .c ({new_AGEMA_signal_8406, RoundOutput[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U922 ( .s (n320), .b ({new_AGEMA_signal_7481, MixColumnsInput[42]}), .a ({new_AGEMA_signal_8063, MixColumnsOutput[42]}), .c ({new_AGEMA_signal_8230, RoundOutput[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U923 ( .s (n320), .b ({new_AGEMA_signal_7480, MixColumnsInput[43]}), .a ({new_AGEMA_signal_8305, MixColumnsOutput[43]}), .c ({new_AGEMA_signal_8407, RoundOutput[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U924 ( .s (n320), .b ({new_AGEMA_signal_7479, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .a ({new_AGEMA_signal_8304, MixColumnsOutput[44]}), .c ({new_AGEMA_signal_8408, RoundOutput[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U925 ( .s (n320), .b ({new_AGEMA_signal_7478, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .a ({new_AGEMA_signal_8060, MixColumnsOutput[45]}), .c ({new_AGEMA_signal_8231, RoundOutput[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U926 ( .s (n319), .b ({new_AGEMA_signal_7477, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .a ({new_AGEMA_signal_8059, MixColumnsOutput[46]}), .c ({new_AGEMA_signal_8232, RoundOutput[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U927 ( .s (n319), .b ({new_AGEMA_signal_7476, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .a ({new_AGEMA_signal_8058, MixColumnsOutput[47]}), .c ({new_AGEMA_signal_8233, RoundOutput[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U928 ( .s (n319), .b ({new_AGEMA_signal_7209, MixColumnsInput[48]}), .a ({new_AGEMA_signal_8057, MixColumnsOutput[48]}), .c ({new_AGEMA_signal_8234, RoundOutput[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U929 ( .s (n319), .b ({new_AGEMA_signal_7405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .a ({new_AGEMA_signal_8303, MixColumnsOutput[49]}), .c ({new_AGEMA_signal_8409, RoundOutput[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U930 ( .s (n319), .b ({new_AGEMA_signal_7416, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .a ({new_AGEMA_signal_8307, MixColumnsOutput[4]}), .c ({new_AGEMA_signal_8410, RoundOutput[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U931 ( .s (n319), .b ({new_AGEMA_signal_7404, MixColumnsInput[50]}), .a ({new_AGEMA_signal_8055, MixColumnsOutput[50]}), .c ({new_AGEMA_signal_8235, RoundOutput[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U932 ( .s (n319), .b ({new_AGEMA_signal_7403, MixColumnsInput[51]}), .a ({new_AGEMA_signal_8302, MixColumnsOutput[51]}), .c ({new_AGEMA_signal_8411, RoundOutput[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U933 ( .s (n319), .b ({new_AGEMA_signal_7402, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .a ({new_AGEMA_signal_8300, MixColumnsOutput[52]}), .c ({new_AGEMA_signal_8412, RoundOutput[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U934 ( .s (n319), .b ({new_AGEMA_signal_7401, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .a ({new_AGEMA_signal_8051, MixColumnsOutput[53]}), .c ({new_AGEMA_signal_8236, RoundOutput[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U935 ( .s (n319), .b ({new_AGEMA_signal_7400, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .a ({new_AGEMA_signal_8050, MixColumnsOutput[54]}), .c ({new_AGEMA_signal_8237, RoundOutput[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U936 ( .s (n319), .b ({new_AGEMA_signal_7399, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .a ({new_AGEMA_signal_8049, MixColumnsOutput[55]}), .c ({new_AGEMA_signal_8238, RoundOutput[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U937 ( .s (n319), .b ({new_AGEMA_signal_7264, MixColumnsInput[56]}), .a ({new_AGEMA_signal_8048, MixColumnsOutput[56]}), .c ({new_AGEMA_signal_8239, RoundOutput[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U938 ( .s (n318), .b ({new_AGEMA_signal_7440, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .a ({new_AGEMA_signal_8299, MixColumnsOutput[57]}), .c ({new_AGEMA_signal_8413, RoundOutput[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U939 ( .s (n318), .b ({new_AGEMA_signal_7439, MixColumnsInput[58]}), .a ({new_AGEMA_signal_8046, MixColumnsOutput[58]}), .c ({new_AGEMA_signal_8240, RoundOutput[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U940 ( .s (n318), .b ({new_AGEMA_signal_7438, MixColumnsInput[59]}), .a ({new_AGEMA_signal_8298, MixColumnsOutput[59]}), .c ({new_AGEMA_signal_8414, RoundOutput[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U941 ( .s (n318), .b ({new_AGEMA_signal_7415, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .a ({new_AGEMA_signal_8069, MixColumnsOutput[5]}), .c ({new_AGEMA_signal_8241, RoundOutput[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U942 ( .s (n318), .b ({new_AGEMA_signal_7437, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .a ({new_AGEMA_signal_8297, MixColumnsOutput[60]}), .c ({new_AGEMA_signal_8415, RoundOutput[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U943 ( .s (n318), .b ({new_AGEMA_signal_7436, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .a ({new_AGEMA_signal_8043, MixColumnsOutput[61]}), .c ({new_AGEMA_signal_8242, RoundOutput[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U944 ( .s (n318), .b ({new_AGEMA_signal_7435, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .a ({new_AGEMA_signal_8041, MixColumnsOutput[62]}), .c ({new_AGEMA_signal_8243, RoundOutput[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U945 ( .s (n318), .b ({new_AGEMA_signal_7434, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .a ({new_AGEMA_signal_8040, MixColumnsOutput[63]}), .c ({new_AGEMA_signal_8244, RoundOutput[63]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U946 ( .s (n318), .b ({new_AGEMA_signal_7319, MixColumnsInput[64]}), .a ({new_AGEMA_signal_8032, MixColumnsOutput[64]}), .c ({new_AGEMA_signal_8245, RoundOutput[64]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U947 ( .s (n318), .b ({new_AGEMA_signal_7475, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .a ({new_AGEMA_signal_8289, MixColumnsOutput[65]}), .c ({new_AGEMA_signal_8416, RoundOutput[65]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U948 ( .s (n318), .b ({new_AGEMA_signal_7474, MixColumnsInput[66]}), .a ({new_AGEMA_signal_8010, MixColumnsOutput[66]}), .c ({new_AGEMA_signal_8246, RoundOutput[66]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U949 ( .s (n318), .b ({new_AGEMA_signal_7473, MixColumnsInput[67]}), .a ({new_AGEMA_signal_8284, MixColumnsOutput[67]}), .c ({new_AGEMA_signal_8417, RoundOutput[67]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U950 ( .s (n317), .b ({new_AGEMA_signal_7472, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .a ({new_AGEMA_signal_8283, MixColumnsOutput[68]}), .c ({new_AGEMA_signal_8418, RoundOutput[68]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U951 ( .s (n317), .b ({new_AGEMA_signal_7471, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .a ({new_AGEMA_signal_8005, MixColumnsOutput[69]}), .c ({new_AGEMA_signal_8247, RoundOutput[69]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U952 ( .s (n317), .b ({new_AGEMA_signal_7414, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .a ({new_AGEMA_signal_8068, MixColumnsOutput[6]}), .c ({new_AGEMA_signal_8248, RoundOutput[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U953 ( .s (n317), .b ({new_AGEMA_signal_7470, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .a ({new_AGEMA_signal_8004, MixColumnsOutput[70]}), .c ({new_AGEMA_signal_8249, RoundOutput[70]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U954 ( .s (n317), .b ({new_AGEMA_signal_7469, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .a ({new_AGEMA_signal_8003, MixColumnsOutput[71]}), .c ({new_AGEMA_signal_8250, RoundOutput[71]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U955 ( .s (n317), .b ({new_AGEMA_signal_7198, MixColumnsInput[72]}), .a ({new_AGEMA_signal_8002, MixColumnsOutput[72]}), .c ({new_AGEMA_signal_8251, RoundOutput[72]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U956 ( .s (n317), .b ({new_AGEMA_signal_7398, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .a ({new_AGEMA_signal_8282, MixColumnsOutput[73]}), .c ({new_AGEMA_signal_8419, RoundOutput[73]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U957 ( .s (n317), .b ({new_AGEMA_signal_7397, MixColumnsInput[74]}), .a ({new_AGEMA_signal_8031, MixColumnsOutput[74]}), .c ({new_AGEMA_signal_8252, RoundOutput[74]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U958 ( .s (n317), .b ({new_AGEMA_signal_7396, MixColumnsInput[75]}), .a ({new_AGEMA_signal_8293, MixColumnsOutput[75]}), .c ({new_AGEMA_signal_8420, RoundOutput[75]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U959 ( .s (n317), .b ({new_AGEMA_signal_7395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .a ({new_AGEMA_signal_8292, MixColumnsOutput[76]}), .c ({new_AGEMA_signal_8421, RoundOutput[76]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U960 ( .s (n317), .b ({new_AGEMA_signal_7394, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .a ({new_AGEMA_signal_8028, MixColumnsOutput[77]}), .c ({new_AGEMA_signal_8253, RoundOutput[77]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U961 ( .s (n317), .b ({new_AGEMA_signal_7393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .a ({new_AGEMA_signal_8027, MixColumnsOutput[78]}), .c ({new_AGEMA_signal_8254, RoundOutput[78]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U962 ( .s (n316), .b ({new_AGEMA_signal_7392, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .a ({new_AGEMA_signal_8026, MixColumnsOutput[79]}), .c ({new_AGEMA_signal_8255, RoundOutput[79]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U963 ( .s (n316), .b ({new_AGEMA_signal_7413, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .a ({new_AGEMA_signal_8067, MixColumnsOutput[7]}), .c ({new_AGEMA_signal_8256, RoundOutput[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U964 ( .s (n316), .b ({new_AGEMA_signal_7253, MixColumnsInput[80]}), .a ({new_AGEMA_signal_8025, MixColumnsOutput[80]}), .c ({new_AGEMA_signal_8257, RoundOutput[80]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U965 ( .s (n316), .b ({new_AGEMA_signal_7433, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .a ({new_AGEMA_signal_8291, MixColumnsOutput[81]}), .c ({new_AGEMA_signal_8422, RoundOutput[81]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U966 ( .s (n316), .b ({new_AGEMA_signal_7432, MixColumnsInput[82]}), .a ({new_AGEMA_signal_8023, MixColumnsOutput[82]}), .c ({new_AGEMA_signal_8258, RoundOutput[82]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U967 ( .s (n316), .b ({new_AGEMA_signal_7431, MixColumnsInput[83]}), .a ({new_AGEMA_signal_8290, MixColumnsOutput[83]}), .c ({new_AGEMA_signal_8423, RoundOutput[83]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U968 ( .s (n316), .b ({new_AGEMA_signal_7430, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .a ({new_AGEMA_signal_8288, MixColumnsOutput[84]}), .c ({new_AGEMA_signal_8424, RoundOutput[84]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U969 ( .s (n316), .b ({new_AGEMA_signal_7429, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .a ({new_AGEMA_signal_8019, MixColumnsOutput[85]}), .c ({new_AGEMA_signal_8259, RoundOutput[85]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U970 ( .s (n316), .b ({new_AGEMA_signal_7428, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .a ({new_AGEMA_signal_8018, MixColumnsOutput[86]}), .c ({new_AGEMA_signal_8260, RoundOutput[86]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U971 ( .s (n316), .b ({new_AGEMA_signal_7427, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .a ({new_AGEMA_signal_8017, MixColumnsOutput[87]}), .c ({new_AGEMA_signal_8261, RoundOutput[87]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U972 ( .s (n316), .b ({new_AGEMA_signal_7308, MixColumnsInput[88]}), .a ({new_AGEMA_signal_8016, MixColumnsOutput[88]}), .c ({new_AGEMA_signal_8262, RoundOutput[88]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U973 ( .s (n316), .b ({new_AGEMA_signal_7468, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .a ({new_AGEMA_signal_8287, MixColumnsOutput[89]}), .c ({new_AGEMA_signal_8425, RoundOutput[89]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U974 ( .s (n315), .b ({new_AGEMA_signal_7286, MixColumnsInput[8]}), .a ({new_AGEMA_signal_8066, MixColumnsOutput[8]}), .c ({new_AGEMA_signal_8263, RoundOutput[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U975 ( .s (n315), .b ({new_AGEMA_signal_7467, MixColumnsInput[90]}), .a ({new_AGEMA_signal_8014, MixColumnsOutput[90]}), .c ({new_AGEMA_signal_8264, RoundOutput[90]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U976 ( .s (n315), .b ({new_AGEMA_signal_7466, MixColumnsInput[91]}), .a ({new_AGEMA_signal_8286, MixColumnsOutput[91]}), .c ({new_AGEMA_signal_8426, RoundOutput[91]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U977 ( .s (n315), .b ({new_AGEMA_signal_7465, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .a ({new_AGEMA_signal_8285, MixColumnsOutput[92]}), .c ({new_AGEMA_signal_8427, RoundOutput[92]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U978 ( .s (n315), .b ({new_AGEMA_signal_7464, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .a ({new_AGEMA_signal_8011, MixColumnsOutput[93]}), .c ({new_AGEMA_signal_8265, RoundOutput[93]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U979 ( .s (n315), .b ({new_AGEMA_signal_7463, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .a ({new_AGEMA_signal_8009, MixColumnsOutput[94]}), .c ({new_AGEMA_signal_8266, RoundOutput[94]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U980 ( .s (n315), .b ({new_AGEMA_signal_7462, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .a ({new_AGEMA_signal_8008, MixColumnsOutput[95]}), .c ({new_AGEMA_signal_8267, RoundOutput[95]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U981 ( .s (n315), .b ({new_AGEMA_signal_7187, MixColumnsInput[96]}), .a ({new_AGEMA_signal_8000, MixColumnsOutput[96]}), .c ({new_AGEMA_signal_8268, RoundOutput[96]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U982 ( .s (n315), .b ({new_AGEMA_signal_7391, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .a ({new_AGEMA_signal_8277, MixColumnsOutput[97]}), .c ({new_AGEMA_signal_8428, RoundOutput[97]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U983 ( .s (n315), .b ({new_AGEMA_signal_7390, MixColumnsInput[98]}), .a ({new_AGEMA_signal_7978, MixColumnsOutput[98]}), .c ({new_AGEMA_signal_8269, RoundOutput[98]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U984 ( .s (n315), .b ({new_AGEMA_signal_7389, MixColumnsInput[99]}), .a ({new_AGEMA_signal_8272, MixColumnsOutput[99]}), .c ({new_AGEMA_signal_8429, RoundOutput[99]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) U985 ( .s (n315), .b ({new_AGEMA_signal_7454, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .a ({new_AGEMA_signal_8306, MixColumnsOutput[9]}), .c ({new_AGEMA_signal_8430, RoundOutput[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8190, RoundOutput[0]}), .a ({plaintext_s1[0], plaintext_s0[0]}), .c ({new_AGEMA_signal_8432, RoundReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8397, RoundOutput[1]}), .a ({plaintext_s1[1], plaintext_s0[1]}), .c ({new_AGEMA_signal_8606, RoundReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8221, RoundOutput[2]}), .a ({plaintext_s1[2], plaintext_s0[2]}), .c ({new_AGEMA_signal_8434, RoundReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8405, RoundOutput[3]}), .a ({plaintext_s1[3], plaintext_s0[3]}), .c ({new_AGEMA_signal_8608, RoundReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8410, RoundOutput[4]}), .a ({plaintext_s1[4], plaintext_s0[4]}), .c ({new_AGEMA_signal_8610, RoundReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8241, RoundOutput[5]}), .a ({plaintext_s1[5], plaintext_s0[5]}), .c ({new_AGEMA_signal_8436, RoundReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8248, RoundOutput[6]}), .a ({plaintext_s1[6], plaintext_s0[6]}), .c ({new_AGEMA_signal_8438, RoundReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8256, RoundOutput[7]}), .a ({plaintext_s1[7], plaintext_s0[7]}), .c ({new_AGEMA_signal_8440, RoundReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8263, RoundOutput[8]}), .a ({plaintext_s1[8], plaintext_s0[8]}), .c ({new_AGEMA_signal_8442, RoundReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8430, RoundOutput[9]}), .a ({plaintext_s1[9], plaintext_s0[9]}), .c ({new_AGEMA_signal_8612, RoundReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8197, RoundOutput[10]}), .a ({plaintext_s1[10], plaintext_s0[10]}), .c ({new_AGEMA_signal_8444, RoundReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8390, RoundOutput[11]}), .a ({plaintext_s1[11], plaintext_s0[11]}), .c ({new_AGEMA_signal_8614, RoundReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8394, RoundOutput[12]}), .a ({plaintext_s1[12], plaintext_s0[12]}), .c ({new_AGEMA_signal_8616, RoundReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8210, RoundOutput[13]}), .a ({plaintext_s1[13], plaintext_s0[13]}), .c ({new_AGEMA_signal_8446, RoundReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8211, RoundOutput[14]}), .a ({plaintext_s1[14], plaintext_s0[14]}), .c ({new_AGEMA_signal_8448, RoundReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8212, RoundOutput[15]}), .a ({plaintext_s1[15], plaintext_s0[15]}), .c ({new_AGEMA_signal_8450, RoundReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8213, RoundOutput[16]}), .a ({plaintext_s1[16], plaintext_s0[16]}), .c ({new_AGEMA_signal_8452, RoundReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8395, RoundOutput[17]}), .a ({plaintext_s1[17], plaintext_s0[17]}), .c ({new_AGEMA_signal_8618, RoundReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8214, RoundOutput[18]}), .a ({plaintext_s1[18], plaintext_s0[18]}), .c ({new_AGEMA_signal_8454, RoundReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8396, RoundOutput[19]}), .a ({plaintext_s1[19], plaintext_s0[19]}), .c ({new_AGEMA_signal_8620, RoundReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8398, RoundOutput[20]}), .a ({plaintext_s1[20], plaintext_s0[20]}), .c ({new_AGEMA_signal_8622, RoundReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8215, RoundOutput[21]}), .a ({plaintext_s1[21], plaintext_s0[21]}), .c ({new_AGEMA_signal_8456, RoundReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8216, RoundOutput[22]}), .a ({plaintext_s1[22], plaintext_s0[22]}), .c ({new_AGEMA_signal_8458, RoundReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8217, RoundOutput[23]}), .a ({plaintext_s1[23], plaintext_s0[23]}), .c ({new_AGEMA_signal_8460, RoundReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8218, RoundOutput[24]}), .a ({plaintext_s1[24], plaintext_s0[24]}), .c ({new_AGEMA_signal_8462, RoundReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8399, RoundOutput[25]}), .a ({plaintext_s1[25], plaintext_s0[25]}), .c ({new_AGEMA_signal_8624, RoundReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8219, RoundOutput[26]}), .a ({plaintext_s1[26], plaintext_s0[26]}), .c ({new_AGEMA_signal_8464, RoundReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8400, RoundOutput[27]}), .a ({plaintext_s1[27], plaintext_s0[27]}), .c ({new_AGEMA_signal_8626, RoundReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8401, RoundOutput[28]}), .a ({plaintext_s1[28], plaintext_s0[28]}), .c ({new_AGEMA_signal_8628, RoundReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8220, RoundOutput[29]}), .a ({plaintext_s1[29], plaintext_s0[29]}), .c ({new_AGEMA_signal_8466, RoundReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8222, RoundOutput[30]}), .a ({plaintext_s1[30], plaintext_s0[30]}), .c ({new_AGEMA_signal_8468, RoundReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8223, RoundOutput[31]}), .a ({plaintext_s1[31], plaintext_s0[31]}), .c ({new_AGEMA_signal_8470, RoundReg_Inst_ff_SDE_31_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8224, RoundOutput[32]}), .a ({plaintext_s1[32], plaintext_s0[32]}), .c ({new_AGEMA_signal_8472, RoundReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8402, RoundOutput[33]}), .a ({plaintext_s1[33], plaintext_s0[33]}), .c ({new_AGEMA_signal_8630, RoundReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8225, RoundOutput[34]}), .a ({plaintext_s1[34], plaintext_s0[34]}), .c ({new_AGEMA_signal_8474, RoundReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8403, RoundOutput[35]}), .a ({plaintext_s1[35], plaintext_s0[35]}), .c ({new_AGEMA_signal_8632, RoundReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8404, RoundOutput[36]}), .a ({plaintext_s1[36], plaintext_s0[36]}), .c ({new_AGEMA_signal_8634, RoundReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8226, RoundOutput[37]}), .a ({plaintext_s1[37], plaintext_s0[37]}), .c ({new_AGEMA_signal_8476, RoundReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8227, RoundOutput[38]}), .a ({plaintext_s1[38], plaintext_s0[38]}), .c ({new_AGEMA_signal_8478, RoundReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8228, RoundOutput[39]}), .a ({plaintext_s1[39], plaintext_s0[39]}), .c ({new_AGEMA_signal_8480, RoundReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8229, RoundOutput[40]}), .a ({plaintext_s1[40], plaintext_s0[40]}), .c ({new_AGEMA_signal_8482, RoundReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8406, RoundOutput[41]}), .a ({plaintext_s1[41], plaintext_s0[41]}), .c ({new_AGEMA_signal_8636, RoundReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8230, RoundOutput[42]}), .a ({plaintext_s1[42], plaintext_s0[42]}), .c ({new_AGEMA_signal_8484, RoundReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8407, RoundOutput[43]}), .a ({plaintext_s1[43], plaintext_s0[43]}), .c ({new_AGEMA_signal_8638, RoundReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8408, RoundOutput[44]}), .a ({plaintext_s1[44], plaintext_s0[44]}), .c ({new_AGEMA_signal_8640, RoundReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8231, RoundOutput[45]}), .a ({plaintext_s1[45], plaintext_s0[45]}), .c ({new_AGEMA_signal_8486, RoundReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8232, RoundOutput[46]}), .a ({plaintext_s1[46], plaintext_s0[46]}), .c ({new_AGEMA_signal_8488, RoundReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8233, RoundOutput[47]}), .a ({plaintext_s1[47], plaintext_s0[47]}), .c ({new_AGEMA_signal_8490, RoundReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8234, RoundOutput[48]}), .a ({plaintext_s1[48], plaintext_s0[48]}), .c ({new_AGEMA_signal_8492, RoundReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8409, RoundOutput[49]}), .a ({plaintext_s1[49], plaintext_s0[49]}), .c ({new_AGEMA_signal_8642, RoundReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8235, RoundOutput[50]}), .a ({plaintext_s1[50], plaintext_s0[50]}), .c ({new_AGEMA_signal_8494, RoundReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8411, RoundOutput[51]}), .a ({plaintext_s1[51], plaintext_s0[51]}), .c ({new_AGEMA_signal_8644, RoundReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8412, RoundOutput[52]}), .a ({plaintext_s1[52], plaintext_s0[52]}), .c ({new_AGEMA_signal_8646, RoundReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8236, RoundOutput[53]}), .a ({plaintext_s1[53], plaintext_s0[53]}), .c ({new_AGEMA_signal_8496, RoundReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8237, RoundOutput[54]}), .a ({plaintext_s1[54], plaintext_s0[54]}), .c ({new_AGEMA_signal_8498, RoundReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8238, RoundOutput[55]}), .a ({plaintext_s1[55], plaintext_s0[55]}), .c ({new_AGEMA_signal_8500, RoundReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8239, RoundOutput[56]}), .a ({plaintext_s1[56], plaintext_s0[56]}), .c ({new_AGEMA_signal_8502, RoundReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8413, RoundOutput[57]}), .a ({plaintext_s1[57], plaintext_s0[57]}), .c ({new_AGEMA_signal_8648, RoundReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8240, RoundOutput[58]}), .a ({plaintext_s1[58], plaintext_s0[58]}), .c ({new_AGEMA_signal_8504, RoundReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8414, RoundOutput[59]}), .a ({plaintext_s1[59], plaintext_s0[59]}), .c ({new_AGEMA_signal_8650, RoundReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8415, RoundOutput[60]}), .a ({plaintext_s1[60], plaintext_s0[60]}), .c ({new_AGEMA_signal_8652, RoundReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8242, RoundOutput[61]}), .a ({plaintext_s1[61], plaintext_s0[61]}), .c ({new_AGEMA_signal_8506, RoundReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8243, RoundOutput[62]}), .a ({plaintext_s1[62], plaintext_s0[62]}), .c ({new_AGEMA_signal_8508, RoundReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8244, RoundOutput[63]}), .a ({plaintext_s1[63], plaintext_s0[63]}), .c ({new_AGEMA_signal_8510, RoundReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8245, RoundOutput[64]}), .a ({plaintext_s1[64], plaintext_s0[64]}), .c ({new_AGEMA_signal_8512, RoundReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8416, RoundOutput[65]}), .a ({plaintext_s1[65], plaintext_s0[65]}), .c ({new_AGEMA_signal_8654, RoundReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8246, RoundOutput[66]}), .a ({plaintext_s1[66], plaintext_s0[66]}), .c ({new_AGEMA_signal_8514, RoundReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8417, RoundOutput[67]}), .a ({plaintext_s1[67], plaintext_s0[67]}), .c ({new_AGEMA_signal_8656, RoundReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8418, RoundOutput[68]}), .a ({plaintext_s1[68], plaintext_s0[68]}), .c ({new_AGEMA_signal_8658, RoundReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8247, RoundOutput[69]}), .a ({plaintext_s1[69], plaintext_s0[69]}), .c ({new_AGEMA_signal_8516, RoundReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8249, RoundOutput[70]}), .a ({plaintext_s1[70], plaintext_s0[70]}), .c ({new_AGEMA_signal_8518, RoundReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8250, RoundOutput[71]}), .a ({plaintext_s1[71], plaintext_s0[71]}), .c ({new_AGEMA_signal_8520, RoundReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8251, RoundOutput[72]}), .a ({plaintext_s1[72], plaintext_s0[72]}), .c ({new_AGEMA_signal_8522, RoundReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8419, RoundOutput[73]}), .a ({plaintext_s1[73], plaintext_s0[73]}), .c ({new_AGEMA_signal_8660, RoundReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8252, RoundOutput[74]}), .a ({plaintext_s1[74], plaintext_s0[74]}), .c ({new_AGEMA_signal_8524, RoundReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8420, RoundOutput[75]}), .a ({plaintext_s1[75], plaintext_s0[75]}), .c ({new_AGEMA_signal_8662, RoundReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8421, RoundOutput[76]}), .a ({plaintext_s1[76], plaintext_s0[76]}), .c ({new_AGEMA_signal_8664, RoundReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8253, RoundOutput[77]}), .a ({plaintext_s1[77], plaintext_s0[77]}), .c ({new_AGEMA_signal_8526, RoundReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8254, RoundOutput[78]}), .a ({plaintext_s1[78], plaintext_s0[78]}), .c ({new_AGEMA_signal_8528, RoundReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8255, RoundOutput[79]}), .a ({plaintext_s1[79], plaintext_s0[79]}), .c ({new_AGEMA_signal_8530, RoundReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8257, RoundOutput[80]}), .a ({plaintext_s1[80], plaintext_s0[80]}), .c ({new_AGEMA_signal_8532, RoundReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8422, RoundOutput[81]}), .a ({plaintext_s1[81], plaintext_s0[81]}), .c ({new_AGEMA_signal_8666, RoundReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8258, RoundOutput[82]}), .a ({plaintext_s1[82], plaintext_s0[82]}), .c ({new_AGEMA_signal_8534, RoundReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8423, RoundOutput[83]}), .a ({plaintext_s1[83], plaintext_s0[83]}), .c ({new_AGEMA_signal_8668, RoundReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8424, RoundOutput[84]}), .a ({plaintext_s1[84], plaintext_s0[84]}), .c ({new_AGEMA_signal_8670, RoundReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8259, RoundOutput[85]}), .a ({plaintext_s1[85], plaintext_s0[85]}), .c ({new_AGEMA_signal_8536, RoundReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8260, RoundOutput[86]}), .a ({plaintext_s1[86], plaintext_s0[86]}), .c ({new_AGEMA_signal_8538, RoundReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8261, RoundOutput[87]}), .a ({plaintext_s1[87], plaintext_s0[87]}), .c ({new_AGEMA_signal_8540, RoundReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8262, RoundOutput[88]}), .a ({plaintext_s1[88], plaintext_s0[88]}), .c ({new_AGEMA_signal_8542, RoundReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8425, RoundOutput[89]}), .a ({plaintext_s1[89], plaintext_s0[89]}), .c ({new_AGEMA_signal_8672, RoundReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8264, RoundOutput[90]}), .a ({plaintext_s1[90], plaintext_s0[90]}), .c ({new_AGEMA_signal_8544, RoundReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8426, RoundOutput[91]}), .a ({plaintext_s1[91], plaintext_s0[91]}), .c ({new_AGEMA_signal_8674, RoundReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8427, RoundOutput[92]}), .a ({plaintext_s1[92], plaintext_s0[92]}), .c ({new_AGEMA_signal_8676, RoundReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8265, RoundOutput[93]}), .a ({plaintext_s1[93], plaintext_s0[93]}), .c ({new_AGEMA_signal_8546, RoundReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8266, RoundOutput[94]}), .a ({plaintext_s1[94], plaintext_s0[94]}), .c ({new_AGEMA_signal_8548, RoundReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8267, RoundOutput[95]}), .a ({plaintext_s1[95], plaintext_s0[95]}), .c ({new_AGEMA_signal_8550, RoundReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8268, RoundOutput[96]}), .a ({plaintext_s1[96], plaintext_s0[96]}), .c ({new_AGEMA_signal_8552, RoundReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8428, RoundOutput[97]}), .a ({plaintext_s1[97], plaintext_s0[97]}), .c ({new_AGEMA_signal_8678, RoundReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8269, RoundOutput[98]}), .a ({plaintext_s1[98], plaintext_s0[98]}), .c ({new_AGEMA_signal_8554, RoundReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8429, RoundOutput[99]}), .a ({plaintext_s1[99], plaintext_s0[99]}), .c ({new_AGEMA_signal_8680, RoundReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8383, RoundOutput[100]}), .a ({plaintext_s1[100], plaintext_s0[100]}), .c ({new_AGEMA_signal_8682, RoundReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8191, RoundOutput[101]}), .a ({plaintext_s1[101], plaintext_s0[101]}), .c ({new_AGEMA_signal_8556, RoundReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8192, RoundOutput[102]}), .a ({plaintext_s1[102], plaintext_s0[102]}), .c ({new_AGEMA_signal_8558, RoundReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8193, RoundOutput[103]}), .a ({plaintext_s1[103], plaintext_s0[103]}), .c ({new_AGEMA_signal_8560, RoundReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8194, RoundOutput[104]}), .a ({plaintext_s1[104], plaintext_s0[104]}), .c ({new_AGEMA_signal_8562, RoundReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8384, RoundOutput[105]}), .a ({plaintext_s1[105], plaintext_s0[105]}), .c ({new_AGEMA_signal_8684, RoundReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8195, RoundOutput[106]}), .a ({plaintext_s1[106], plaintext_s0[106]}), .c ({new_AGEMA_signal_8564, RoundReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8385, RoundOutput[107]}), .a ({plaintext_s1[107], plaintext_s0[107]}), .c ({new_AGEMA_signal_8686, RoundReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8386, RoundOutput[108]}), .a ({plaintext_s1[108], plaintext_s0[108]}), .c ({new_AGEMA_signal_8688, RoundReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8196, RoundOutput[109]}), .a ({plaintext_s1[109], plaintext_s0[109]}), .c ({new_AGEMA_signal_8566, RoundReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8198, RoundOutput[110]}), .a ({plaintext_s1[110], plaintext_s0[110]}), .c ({new_AGEMA_signal_8568, RoundReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8199, RoundOutput[111]}), .a ({plaintext_s1[111], plaintext_s0[111]}), .c ({new_AGEMA_signal_8570, RoundReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8200, RoundOutput[112]}), .a ({plaintext_s1[112], plaintext_s0[112]}), .c ({new_AGEMA_signal_8572, RoundReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8387, RoundOutput[113]}), .a ({plaintext_s1[113], plaintext_s0[113]}), .c ({new_AGEMA_signal_8690, RoundReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8201, RoundOutput[114]}), .a ({plaintext_s1[114], plaintext_s0[114]}), .c ({new_AGEMA_signal_8574, RoundReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8388, RoundOutput[115]}), .a ({plaintext_s1[115], plaintext_s0[115]}), .c ({new_AGEMA_signal_8692, RoundReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8389, RoundOutput[116]}), .a ({plaintext_s1[116], plaintext_s0[116]}), .c ({new_AGEMA_signal_8694, RoundReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8202, RoundOutput[117]}), .a ({plaintext_s1[117], plaintext_s0[117]}), .c ({new_AGEMA_signal_8576, RoundReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8203, RoundOutput[118]}), .a ({plaintext_s1[118], plaintext_s0[118]}), .c ({new_AGEMA_signal_8578, RoundReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8204, RoundOutput[119]}), .a ({plaintext_s1[119], plaintext_s0[119]}), .c ({new_AGEMA_signal_8580, RoundReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8205, RoundOutput[120]}), .a ({plaintext_s1[120], plaintext_s0[120]}), .c ({new_AGEMA_signal_8582, RoundReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8391, RoundOutput[121]}), .a ({plaintext_s1[121], plaintext_s0[121]}), .c ({new_AGEMA_signal_8696, RoundReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8206, RoundOutput[122]}), .a ({plaintext_s1[122], plaintext_s0[122]}), .c ({new_AGEMA_signal_8584, RoundReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8392, RoundOutput[123]}), .a ({plaintext_s1[123], plaintext_s0[123]}), .c ({new_AGEMA_signal_8698, RoundReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8393, RoundOutput[124]}), .a ({plaintext_s1[124], plaintext_s0[124]}), .c ({new_AGEMA_signal_8700, RoundReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8207, RoundOutput[125]}), .a ({plaintext_s1[125], plaintext_s0[125]}), .c ({new_AGEMA_signal_8586, RoundReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8208, RoundOutput[126]}), .a ({plaintext_s1[126], plaintext_s0[126]}), .c ({new_AGEMA_signal_8588, RoundReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8209, RoundOutput[127]}), .a ({plaintext_s1[127], plaintext_s0[127]}), .c ({new_AGEMA_signal_8590, RoundReg_Inst_ff_SDE_127_next_state}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M46_U1 ( .a ({new_AGEMA_signal_6324, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_5165, SubBytesIns_Inst_Sbox_0_T6}), .clk (clk), .r (Fresh[320]), .c ({new_AGEMA_signal_6562, SubBytesIns_Inst_Sbox_0_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M47_U1 ( .a ({new_AGEMA_signal_6212, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_5345, SubBytesIns_Inst_Sbox_0_T8}), .clk (clk), .r (Fresh[321]), .c ({new_AGEMA_signal_6325, SubBytesIns_Inst_Sbox_0_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M48_U1 ( .a ({new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_0_M39}), .b ({ciphertext_s1[0], ciphertext_s0[0]}), .clk (clk), .r (Fresh[322]), .c ({new_AGEMA_signal_6326, SubBytesIns_Inst_Sbox_0_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M49_U1 ( .a ({new_AGEMA_signal_6323, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_5169, SubBytesIns_Inst_Sbox_0_T16}), .clk (clk), .r (Fresh[323]), .c ({new_AGEMA_signal_6563, SubBytesIns_Inst_Sbox_0_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M50_U1 ( .a ({new_AGEMA_signal_6210, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_5166, SubBytesIns_Inst_Sbox_0_T9}), .clk (clk), .r (Fresh[324]), .c ({new_AGEMA_signal_6327, SubBytesIns_Inst_Sbox_0_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M51_U1 ( .a ({new_AGEMA_signal_6209, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_5348, SubBytesIns_Inst_Sbox_0_T17}), .clk (clk), .r (Fresh[325]), .c ({new_AGEMA_signal_6328, SubBytesIns_Inst_Sbox_0_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M52_U1 ( .a ({new_AGEMA_signal_6322, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_5168, SubBytesIns_Inst_Sbox_0_T15}), .clk (clk), .r (Fresh[326]), .c ({new_AGEMA_signal_6564, SubBytesIns_Inst_Sbox_0_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M53_U1 ( .a ({new_AGEMA_signal_6561, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_5172, SubBytesIns_Inst_Sbox_0_T27}), .clk (clk), .r (Fresh[327]), .c ({new_AGEMA_signal_6793, SubBytesIns_Inst_Sbox_0_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M54_U1 ( .a ({new_AGEMA_signal_6321, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_5346, SubBytesIns_Inst_Sbox_0_T10}), .clk (clk), .r (Fresh[328]), .c ({new_AGEMA_signal_6565, SubBytesIns_Inst_Sbox_0_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M55_U1 ( .a ({new_AGEMA_signal_6324, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_5167, SubBytesIns_Inst_Sbox_0_T13}), .clk (clk), .r (Fresh[329]), .c ({new_AGEMA_signal_6566, SubBytesIns_Inst_Sbox_0_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M56_U1 ( .a ({new_AGEMA_signal_6212, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_5350, SubBytesIns_Inst_Sbox_0_T23}), .clk (clk), .r (Fresh[330]), .c ({new_AGEMA_signal_6329, SubBytesIns_Inst_Sbox_0_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M57_U1 ( .a ({new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_5170, SubBytesIns_Inst_Sbox_0_T19}), .clk (clk), .r (Fresh[331]), .c ({new_AGEMA_signal_6330, SubBytesIns_Inst_Sbox_0_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M58_U1 ( .a ({new_AGEMA_signal_6323, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_4975, SubBytesIns_Inst_Sbox_0_T3}), .clk (clk), .r (Fresh[332]), .c ({new_AGEMA_signal_6567, SubBytesIns_Inst_Sbox_0_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M59_U1 ( .a ({new_AGEMA_signal_6210, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_5171, SubBytesIns_Inst_Sbox_0_T22}), .clk (clk), .r (Fresh[333]), .c ({new_AGEMA_signal_6331, SubBytesIns_Inst_Sbox_0_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M60_U1 ( .a ({new_AGEMA_signal_6209, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_5349, SubBytesIns_Inst_Sbox_0_T20}), .clk (clk), .r (Fresh[334]), .c ({new_AGEMA_signal_6332, SubBytesIns_Inst_Sbox_0_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M61_U1 ( .a ({new_AGEMA_signal_6322, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_4973, SubBytesIns_Inst_Sbox_0_T1}), .clk (clk), .r (Fresh[335]), .c ({new_AGEMA_signal_6568, SubBytesIns_Inst_Sbox_0_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M62_U1 ( .a ({new_AGEMA_signal_6561, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_4976, SubBytesIns_Inst_Sbox_0_T4}), .clk (clk), .r (Fresh[336]), .c ({new_AGEMA_signal_6794, SubBytesIns_Inst_Sbox_0_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M63_U1 ( .a ({new_AGEMA_signal_6321, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_4974, SubBytesIns_Inst_Sbox_0_T2}), .clk (clk), .r (Fresh[337]), .c ({new_AGEMA_signal_6569, SubBytesIns_Inst_Sbox_0_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L0_U1 ( .a ({new_AGEMA_signal_6568, SubBytesIns_Inst_Sbox_0_M61}), .b ({new_AGEMA_signal_6794, SubBytesIns_Inst_Sbox_0_M62}), .c ({new_AGEMA_signal_6989, SubBytesIns_Inst_Sbox_0_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L1_U1 ( .a ({new_AGEMA_signal_6327, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_6329, SubBytesIns_Inst_Sbox_0_M56}), .c ({new_AGEMA_signal_6570, SubBytesIns_Inst_Sbox_0_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L2_U1 ( .a ({new_AGEMA_signal_6562, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_6326, SubBytesIns_Inst_Sbox_0_M48}), .c ({new_AGEMA_signal_6795, SubBytesIns_Inst_Sbox_0_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L3_U1 ( .a ({new_AGEMA_signal_6325, SubBytesIns_Inst_Sbox_0_M47}), .b ({new_AGEMA_signal_6566, SubBytesIns_Inst_Sbox_0_M55}), .c ({new_AGEMA_signal_6796, SubBytesIns_Inst_Sbox_0_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L4_U1 ( .a ({new_AGEMA_signal_6565, SubBytesIns_Inst_Sbox_0_M54}), .b ({new_AGEMA_signal_6567, SubBytesIns_Inst_Sbox_0_M58}), .c ({new_AGEMA_signal_6797, SubBytesIns_Inst_Sbox_0_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L5_U1 ( .a ({new_AGEMA_signal_6563, SubBytesIns_Inst_Sbox_0_M49}), .b ({new_AGEMA_signal_6568, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_6798, SubBytesIns_Inst_Sbox_0_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L6_U1 ( .a ({new_AGEMA_signal_6794, SubBytesIns_Inst_Sbox_0_M62}), .b ({new_AGEMA_signal_6798, SubBytesIns_Inst_Sbox_0_L5}), .c ({new_AGEMA_signal_6990, SubBytesIns_Inst_Sbox_0_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L7_U1 ( .a ({new_AGEMA_signal_6562, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_6796, SubBytesIns_Inst_Sbox_0_L3}), .c ({new_AGEMA_signal_6991, SubBytesIns_Inst_Sbox_0_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L8_U1 ( .a ({new_AGEMA_signal_6328, SubBytesIns_Inst_Sbox_0_M51}), .b ({new_AGEMA_signal_6331, SubBytesIns_Inst_Sbox_0_M59}), .c ({new_AGEMA_signal_6571, SubBytesIns_Inst_Sbox_0_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L9_U1 ( .a ({new_AGEMA_signal_6564, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_6793, SubBytesIns_Inst_Sbox_0_M53}), .c ({new_AGEMA_signal_6992, SubBytesIns_Inst_Sbox_0_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L10_U1 ( .a ({new_AGEMA_signal_6793, SubBytesIns_Inst_Sbox_0_M53}), .b ({new_AGEMA_signal_6797, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_6993, SubBytesIns_Inst_Sbox_0_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L11_U1 ( .a ({new_AGEMA_signal_6332, SubBytesIns_Inst_Sbox_0_M60}), .b ({new_AGEMA_signal_6795, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_6994, SubBytesIns_Inst_Sbox_0_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L12_U1 ( .a ({new_AGEMA_signal_6326, SubBytesIns_Inst_Sbox_0_M48}), .b ({new_AGEMA_signal_6328, SubBytesIns_Inst_Sbox_0_M51}), .c ({new_AGEMA_signal_6572, SubBytesIns_Inst_Sbox_0_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L13_U1 ( .a ({new_AGEMA_signal_6327, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_6989, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_7177, SubBytesIns_Inst_Sbox_0_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L14_U1 ( .a ({new_AGEMA_signal_6564, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_6568, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_6799, SubBytesIns_Inst_Sbox_0_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L15_U1 ( .a ({new_AGEMA_signal_6566, SubBytesIns_Inst_Sbox_0_M55}), .b ({new_AGEMA_signal_6570, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_6800, SubBytesIns_Inst_Sbox_0_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L16_U1 ( .a ({new_AGEMA_signal_6329, SubBytesIns_Inst_Sbox_0_M56}), .b ({new_AGEMA_signal_6989, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_7178, SubBytesIns_Inst_Sbox_0_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L17_U1 ( .a ({new_AGEMA_signal_6330, SubBytesIns_Inst_Sbox_0_M57}), .b ({new_AGEMA_signal_6570, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_6801, SubBytesIns_Inst_Sbox_0_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L18_U1 ( .a ({new_AGEMA_signal_6567, SubBytesIns_Inst_Sbox_0_M58}), .b ({new_AGEMA_signal_6571, SubBytesIns_Inst_Sbox_0_L8}), .c ({new_AGEMA_signal_6802, SubBytesIns_Inst_Sbox_0_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L19_U1 ( .a ({new_AGEMA_signal_6569, SubBytesIns_Inst_Sbox_0_M63}), .b ({new_AGEMA_signal_6797, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_6995, SubBytesIns_Inst_Sbox_0_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L20_U1 ( .a ({new_AGEMA_signal_6989, SubBytesIns_Inst_Sbox_0_L0}), .b ({new_AGEMA_signal_6570, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_7179, SubBytesIns_Inst_Sbox_0_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L21_U1 ( .a ({new_AGEMA_signal_6570, SubBytesIns_Inst_Sbox_0_L1}), .b ({new_AGEMA_signal_6991, SubBytesIns_Inst_Sbox_0_L7}), .c ({new_AGEMA_signal_7180, SubBytesIns_Inst_Sbox_0_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L22_U1 ( .a ({new_AGEMA_signal_6796, SubBytesIns_Inst_Sbox_0_L3}), .b ({new_AGEMA_signal_6572, SubBytesIns_Inst_Sbox_0_L12}), .c ({new_AGEMA_signal_6996, SubBytesIns_Inst_Sbox_0_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L23_U1 ( .a ({new_AGEMA_signal_6802, SubBytesIns_Inst_Sbox_0_L18}), .b ({new_AGEMA_signal_6795, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_6997, SubBytesIns_Inst_Sbox_0_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L24_U1 ( .a ({new_AGEMA_signal_6800, SubBytesIns_Inst_Sbox_0_L15}), .b ({new_AGEMA_signal_6992, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_7181, SubBytesIns_Inst_Sbox_0_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L25_U1 ( .a ({new_AGEMA_signal_6990, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_6993, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_7182, SubBytesIns_Inst_Sbox_0_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L26_U1 ( .a ({new_AGEMA_signal_6991, SubBytesIns_Inst_Sbox_0_L7}), .b ({new_AGEMA_signal_6992, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_7183, SubBytesIns_Inst_Sbox_0_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L27_U1 ( .a ({new_AGEMA_signal_6571, SubBytesIns_Inst_Sbox_0_L8}), .b ({new_AGEMA_signal_6993, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_7184, SubBytesIns_Inst_Sbox_0_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L28_U1 ( .a ({new_AGEMA_signal_6994, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_6799, SubBytesIns_Inst_Sbox_0_L14}), .c ({new_AGEMA_signal_7185, SubBytesIns_Inst_Sbox_0_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L29_U1 ( .a ({new_AGEMA_signal_6994, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_6801, SubBytesIns_Inst_Sbox_0_L17}), .c ({new_AGEMA_signal_7186, SubBytesIns_Inst_Sbox_0_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S0_U1 ( .a ({new_AGEMA_signal_6990, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_7181, SubBytesIns_Inst_Sbox_0_L24}), .c ({new_AGEMA_signal_7385, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S1_U1 ( .a ({new_AGEMA_signal_7178, SubBytesIns_Inst_Sbox_0_L16}), .b ({new_AGEMA_signal_7183, SubBytesIns_Inst_Sbox_0_L26}), .c ({new_AGEMA_signal_7386, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S2_U1 ( .a ({new_AGEMA_signal_6995, SubBytesIns_Inst_Sbox_0_L19}), .b ({new_AGEMA_signal_7185, SubBytesIns_Inst_Sbox_0_L28}), .c ({new_AGEMA_signal_7387, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S3_U1 ( .a ({new_AGEMA_signal_6990, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_7180, SubBytesIns_Inst_Sbox_0_L21}), .c ({new_AGEMA_signal_7388, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S4_U1 ( .a ({new_AGEMA_signal_7179, SubBytesIns_Inst_Sbox_0_L20}), .b ({new_AGEMA_signal_6996, SubBytesIns_Inst_Sbox_0_L22}), .c ({new_AGEMA_signal_7389, MixColumnsInput[99]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S5_U1 ( .a ({new_AGEMA_signal_7182, SubBytesIns_Inst_Sbox_0_L25}), .b ({new_AGEMA_signal_7186, SubBytesIns_Inst_Sbox_0_L29}), .c ({new_AGEMA_signal_7390, MixColumnsInput[98]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S6_U1 ( .a ({new_AGEMA_signal_7177, SubBytesIns_Inst_Sbox_0_L13}), .b ({new_AGEMA_signal_7184, SubBytesIns_Inst_Sbox_0_L27}), .c ({new_AGEMA_signal_7391, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S7_U1 ( .a ({new_AGEMA_signal_6990, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_6997, SubBytesIns_Inst_Sbox_0_L23}), .c ({new_AGEMA_signal_7187, MixColumnsInput[96]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M46_U1 ( .a ({new_AGEMA_signal_6336, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_5173, SubBytesIns_Inst_Sbox_1_T6}), .clk (clk), .r (Fresh[338]), .c ({new_AGEMA_signal_6574, SubBytesIns_Inst_Sbox_1_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M47_U1 ( .a ({new_AGEMA_signal_6216, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_5358, SubBytesIns_Inst_Sbox_1_T8}), .clk (clk), .r (Fresh[339]), .c ({new_AGEMA_signal_6337, SubBytesIns_Inst_Sbox_1_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M48_U1 ( .a ({new_AGEMA_signal_6215, SubBytesIns_Inst_Sbox_1_M39}), .b ({ciphertext_s1[8], ciphertext_s0[8]}), .clk (clk), .r (Fresh[340]), .c ({new_AGEMA_signal_6338, SubBytesIns_Inst_Sbox_1_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M49_U1 ( .a ({new_AGEMA_signal_6335, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_5177, SubBytesIns_Inst_Sbox_1_T16}), .clk (clk), .r (Fresh[341]), .c ({new_AGEMA_signal_6575, SubBytesIns_Inst_Sbox_1_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M50_U1 ( .a ({new_AGEMA_signal_6214, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_5174, SubBytesIns_Inst_Sbox_1_T9}), .clk (clk), .r (Fresh[342]), .c ({new_AGEMA_signal_6339, SubBytesIns_Inst_Sbox_1_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M51_U1 ( .a ({new_AGEMA_signal_6213, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_5361, SubBytesIns_Inst_Sbox_1_T17}), .clk (clk), .r (Fresh[343]), .c ({new_AGEMA_signal_6340, SubBytesIns_Inst_Sbox_1_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M52_U1 ( .a ({new_AGEMA_signal_6334, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_5176, SubBytesIns_Inst_Sbox_1_T15}), .clk (clk), .r (Fresh[344]), .c ({new_AGEMA_signal_6576, SubBytesIns_Inst_Sbox_1_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M53_U1 ( .a ({new_AGEMA_signal_6573, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_5180, SubBytesIns_Inst_Sbox_1_T27}), .clk (clk), .r (Fresh[345]), .c ({new_AGEMA_signal_6803, SubBytesIns_Inst_Sbox_1_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M54_U1 ( .a ({new_AGEMA_signal_6333, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_5359, SubBytesIns_Inst_Sbox_1_T10}), .clk (clk), .r (Fresh[346]), .c ({new_AGEMA_signal_6577, SubBytesIns_Inst_Sbox_1_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M55_U1 ( .a ({new_AGEMA_signal_6336, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_5175, SubBytesIns_Inst_Sbox_1_T13}), .clk (clk), .r (Fresh[347]), .c ({new_AGEMA_signal_6578, SubBytesIns_Inst_Sbox_1_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M56_U1 ( .a ({new_AGEMA_signal_6216, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_5363, SubBytesIns_Inst_Sbox_1_T23}), .clk (clk), .r (Fresh[348]), .c ({new_AGEMA_signal_6341, SubBytesIns_Inst_Sbox_1_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M57_U1 ( .a ({new_AGEMA_signal_6215, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_5178, SubBytesIns_Inst_Sbox_1_T19}), .clk (clk), .r (Fresh[349]), .c ({new_AGEMA_signal_6342, SubBytesIns_Inst_Sbox_1_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M58_U1 ( .a ({new_AGEMA_signal_6335, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_4985, SubBytesIns_Inst_Sbox_1_T3}), .clk (clk), .r (Fresh[350]), .c ({new_AGEMA_signal_6579, SubBytesIns_Inst_Sbox_1_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M59_U1 ( .a ({new_AGEMA_signal_6214, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_5179, SubBytesIns_Inst_Sbox_1_T22}), .clk (clk), .r (Fresh[351]), .c ({new_AGEMA_signal_6343, SubBytesIns_Inst_Sbox_1_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M60_U1 ( .a ({new_AGEMA_signal_6213, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_5362, SubBytesIns_Inst_Sbox_1_T20}), .clk (clk), .r (Fresh[352]), .c ({new_AGEMA_signal_6344, SubBytesIns_Inst_Sbox_1_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M61_U1 ( .a ({new_AGEMA_signal_6334, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_4983, SubBytesIns_Inst_Sbox_1_T1}), .clk (clk), .r (Fresh[353]), .c ({new_AGEMA_signal_6580, SubBytesIns_Inst_Sbox_1_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M62_U1 ( .a ({new_AGEMA_signal_6573, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_4986, SubBytesIns_Inst_Sbox_1_T4}), .clk (clk), .r (Fresh[354]), .c ({new_AGEMA_signal_6804, SubBytesIns_Inst_Sbox_1_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M63_U1 ( .a ({new_AGEMA_signal_6333, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_4984, SubBytesIns_Inst_Sbox_1_T2}), .clk (clk), .r (Fresh[355]), .c ({new_AGEMA_signal_6581, SubBytesIns_Inst_Sbox_1_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L0_U1 ( .a ({new_AGEMA_signal_6580, SubBytesIns_Inst_Sbox_1_M61}), .b ({new_AGEMA_signal_6804, SubBytesIns_Inst_Sbox_1_M62}), .c ({new_AGEMA_signal_6998, SubBytesIns_Inst_Sbox_1_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L1_U1 ( .a ({new_AGEMA_signal_6339, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_6341, SubBytesIns_Inst_Sbox_1_M56}), .c ({new_AGEMA_signal_6582, SubBytesIns_Inst_Sbox_1_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L2_U1 ( .a ({new_AGEMA_signal_6574, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_6338, SubBytesIns_Inst_Sbox_1_M48}), .c ({new_AGEMA_signal_6805, SubBytesIns_Inst_Sbox_1_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L3_U1 ( .a ({new_AGEMA_signal_6337, SubBytesIns_Inst_Sbox_1_M47}), .b ({new_AGEMA_signal_6578, SubBytesIns_Inst_Sbox_1_M55}), .c ({new_AGEMA_signal_6806, SubBytesIns_Inst_Sbox_1_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L4_U1 ( .a ({new_AGEMA_signal_6577, SubBytesIns_Inst_Sbox_1_M54}), .b ({new_AGEMA_signal_6579, SubBytesIns_Inst_Sbox_1_M58}), .c ({new_AGEMA_signal_6807, SubBytesIns_Inst_Sbox_1_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L5_U1 ( .a ({new_AGEMA_signal_6575, SubBytesIns_Inst_Sbox_1_M49}), .b ({new_AGEMA_signal_6580, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_6808, SubBytesIns_Inst_Sbox_1_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L6_U1 ( .a ({new_AGEMA_signal_6804, SubBytesIns_Inst_Sbox_1_M62}), .b ({new_AGEMA_signal_6808, SubBytesIns_Inst_Sbox_1_L5}), .c ({new_AGEMA_signal_6999, SubBytesIns_Inst_Sbox_1_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L7_U1 ( .a ({new_AGEMA_signal_6574, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_6806, SubBytesIns_Inst_Sbox_1_L3}), .c ({new_AGEMA_signal_7000, SubBytesIns_Inst_Sbox_1_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L8_U1 ( .a ({new_AGEMA_signal_6340, SubBytesIns_Inst_Sbox_1_M51}), .b ({new_AGEMA_signal_6343, SubBytesIns_Inst_Sbox_1_M59}), .c ({new_AGEMA_signal_6583, SubBytesIns_Inst_Sbox_1_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L9_U1 ( .a ({new_AGEMA_signal_6576, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_6803, SubBytesIns_Inst_Sbox_1_M53}), .c ({new_AGEMA_signal_7001, SubBytesIns_Inst_Sbox_1_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L10_U1 ( .a ({new_AGEMA_signal_6803, SubBytesIns_Inst_Sbox_1_M53}), .b ({new_AGEMA_signal_6807, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_7002, SubBytesIns_Inst_Sbox_1_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L11_U1 ( .a ({new_AGEMA_signal_6344, SubBytesIns_Inst_Sbox_1_M60}), .b ({new_AGEMA_signal_6805, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_7003, SubBytesIns_Inst_Sbox_1_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L12_U1 ( .a ({new_AGEMA_signal_6338, SubBytesIns_Inst_Sbox_1_M48}), .b ({new_AGEMA_signal_6340, SubBytesIns_Inst_Sbox_1_M51}), .c ({new_AGEMA_signal_6584, SubBytesIns_Inst_Sbox_1_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L13_U1 ( .a ({new_AGEMA_signal_6339, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_6998, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_7188, SubBytesIns_Inst_Sbox_1_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L14_U1 ( .a ({new_AGEMA_signal_6576, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_6580, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_6809, SubBytesIns_Inst_Sbox_1_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L15_U1 ( .a ({new_AGEMA_signal_6578, SubBytesIns_Inst_Sbox_1_M55}), .b ({new_AGEMA_signal_6582, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_6810, SubBytesIns_Inst_Sbox_1_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L16_U1 ( .a ({new_AGEMA_signal_6341, SubBytesIns_Inst_Sbox_1_M56}), .b ({new_AGEMA_signal_6998, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_7189, SubBytesIns_Inst_Sbox_1_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L17_U1 ( .a ({new_AGEMA_signal_6342, SubBytesIns_Inst_Sbox_1_M57}), .b ({new_AGEMA_signal_6582, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_6811, SubBytesIns_Inst_Sbox_1_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L18_U1 ( .a ({new_AGEMA_signal_6579, SubBytesIns_Inst_Sbox_1_M58}), .b ({new_AGEMA_signal_6583, SubBytesIns_Inst_Sbox_1_L8}), .c ({new_AGEMA_signal_6812, SubBytesIns_Inst_Sbox_1_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L19_U1 ( .a ({new_AGEMA_signal_6581, SubBytesIns_Inst_Sbox_1_M63}), .b ({new_AGEMA_signal_6807, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_7004, SubBytesIns_Inst_Sbox_1_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L20_U1 ( .a ({new_AGEMA_signal_6998, SubBytesIns_Inst_Sbox_1_L0}), .b ({new_AGEMA_signal_6582, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_7190, SubBytesIns_Inst_Sbox_1_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L21_U1 ( .a ({new_AGEMA_signal_6582, SubBytesIns_Inst_Sbox_1_L1}), .b ({new_AGEMA_signal_7000, SubBytesIns_Inst_Sbox_1_L7}), .c ({new_AGEMA_signal_7191, SubBytesIns_Inst_Sbox_1_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L22_U1 ( .a ({new_AGEMA_signal_6806, SubBytesIns_Inst_Sbox_1_L3}), .b ({new_AGEMA_signal_6584, SubBytesIns_Inst_Sbox_1_L12}), .c ({new_AGEMA_signal_7005, SubBytesIns_Inst_Sbox_1_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L23_U1 ( .a ({new_AGEMA_signal_6812, SubBytesIns_Inst_Sbox_1_L18}), .b ({new_AGEMA_signal_6805, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_7006, SubBytesIns_Inst_Sbox_1_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L24_U1 ( .a ({new_AGEMA_signal_6810, SubBytesIns_Inst_Sbox_1_L15}), .b ({new_AGEMA_signal_7001, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_7192, SubBytesIns_Inst_Sbox_1_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L25_U1 ( .a ({new_AGEMA_signal_6999, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_7002, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_7193, SubBytesIns_Inst_Sbox_1_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L26_U1 ( .a ({new_AGEMA_signal_7000, SubBytesIns_Inst_Sbox_1_L7}), .b ({new_AGEMA_signal_7001, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_7194, SubBytesIns_Inst_Sbox_1_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L27_U1 ( .a ({new_AGEMA_signal_6583, SubBytesIns_Inst_Sbox_1_L8}), .b ({new_AGEMA_signal_7002, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_7195, SubBytesIns_Inst_Sbox_1_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L28_U1 ( .a ({new_AGEMA_signal_7003, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_6809, SubBytesIns_Inst_Sbox_1_L14}), .c ({new_AGEMA_signal_7196, SubBytesIns_Inst_Sbox_1_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L29_U1 ( .a ({new_AGEMA_signal_7003, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_6811, SubBytesIns_Inst_Sbox_1_L17}), .c ({new_AGEMA_signal_7197, SubBytesIns_Inst_Sbox_1_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S0_U1 ( .a ({new_AGEMA_signal_6999, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_7192, SubBytesIns_Inst_Sbox_1_L24}), .c ({new_AGEMA_signal_7392, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S1_U1 ( .a ({new_AGEMA_signal_7189, SubBytesIns_Inst_Sbox_1_L16}), .b ({new_AGEMA_signal_7194, SubBytesIns_Inst_Sbox_1_L26}), .c ({new_AGEMA_signal_7393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S2_U1 ( .a ({new_AGEMA_signal_7004, SubBytesIns_Inst_Sbox_1_L19}), .b ({new_AGEMA_signal_7196, SubBytesIns_Inst_Sbox_1_L28}), .c ({new_AGEMA_signal_7394, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S3_U1 ( .a ({new_AGEMA_signal_6999, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_7191, SubBytesIns_Inst_Sbox_1_L21}), .c ({new_AGEMA_signal_7395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S4_U1 ( .a ({new_AGEMA_signal_7190, SubBytesIns_Inst_Sbox_1_L20}), .b ({new_AGEMA_signal_7005, SubBytesIns_Inst_Sbox_1_L22}), .c ({new_AGEMA_signal_7396, MixColumnsInput[75]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S5_U1 ( .a ({new_AGEMA_signal_7193, SubBytesIns_Inst_Sbox_1_L25}), .b ({new_AGEMA_signal_7197, SubBytesIns_Inst_Sbox_1_L29}), .c ({new_AGEMA_signal_7397, MixColumnsInput[74]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S6_U1 ( .a ({new_AGEMA_signal_7188, SubBytesIns_Inst_Sbox_1_L13}), .b ({new_AGEMA_signal_7195, SubBytesIns_Inst_Sbox_1_L27}), .c ({new_AGEMA_signal_7398, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S7_U1 ( .a ({new_AGEMA_signal_6999, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_7006, SubBytesIns_Inst_Sbox_1_L23}), .c ({new_AGEMA_signal_7198, MixColumnsInput[72]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M46_U1 ( .a ({new_AGEMA_signal_6348, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_5181, SubBytesIns_Inst_Sbox_2_T6}), .clk (clk), .r (Fresh[356]), .c ({new_AGEMA_signal_6586, SubBytesIns_Inst_Sbox_2_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M47_U1 ( .a ({new_AGEMA_signal_6220, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_5371, SubBytesIns_Inst_Sbox_2_T8}), .clk (clk), .r (Fresh[357]), .c ({new_AGEMA_signal_6349, SubBytesIns_Inst_Sbox_2_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M48_U1 ( .a ({new_AGEMA_signal_6219, SubBytesIns_Inst_Sbox_2_M39}), .b ({ciphertext_s1[16], ciphertext_s0[16]}), .clk (clk), .r (Fresh[358]), .c ({new_AGEMA_signal_6350, SubBytesIns_Inst_Sbox_2_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M49_U1 ( .a ({new_AGEMA_signal_6347, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_5185, SubBytesIns_Inst_Sbox_2_T16}), .clk (clk), .r (Fresh[359]), .c ({new_AGEMA_signal_6587, SubBytesIns_Inst_Sbox_2_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M50_U1 ( .a ({new_AGEMA_signal_6218, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_5182, SubBytesIns_Inst_Sbox_2_T9}), .clk (clk), .r (Fresh[360]), .c ({new_AGEMA_signal_6351, SubBytesIns_Inst_Sbox_2_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M51_U1 ( .a ({new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_5374, SubBytesIns_Inst_Sbox_2_T17}), .clk (clk), .r (Fresh[361]), .c ({new_AGEMA_signal_6352, SubBytesIns_Inst_Sbox_2_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M52_U1 ( .a ({new_AGEMA_signal_6346, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_5184, SubBytesIns_Inst_Sbox_2_T15}), .clk (clk), .r (Fresh[362]), .c ({new_AGEMA_signal_6588, SubBytesIns_Inst_Sbox_2_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M53_U1 ( .a ({new_AGEMA_signal_6585, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_5188, SubBytesIns_Inst_Sbox_2_T27}), .clk (clk), .r (Fresh[363]), .c ({new_AGEMA_signal_6813, SubBytesIns_Inst_Sbox_2_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M54_U1 ( .a ({new_AGEMA_signal_6345, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_5372, SubBytesIns_Inst_Sbox_2_T10}), .clk (clk), .r (Fresh[364]), .c ({new_AGEMA_signal_6589, SubBytesIns_Inst_Sbox_2_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M55_U1 ( .a ({new_AGEMA_signal_6348, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_5183, SubBytesIns_Inst_Sbox_2_T13}), .clk (clk), .r (Fresh[365]), .c ({new_AGEMA_signal_6590, SubBytesIns_Inst_Sbox_2_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M56_U1 ( .a ({new_AGEMA_signal_6220, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_5376, SubBytesIns_Inst_Sbox_2_T23}), .clk (clk), .r (Fresh[366]), .c ({new_AGEMA_signal_6353, SubBytesIns_Inst_Sbox_2_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M57_U1 ( .a ({new_AGEMA_signal_6219, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_5186, SubBytesIns_Inst_Sbox_2_T19}), .clk (clk), .r (Fresh[367]), .c ({new_AGEMA_signal_6354, SubBytesIns_Inst_Sbox_2_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M58_U1 ( .a ({new_AGEMA_signal_6347, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_4995, SubBytesIns_Inst_Sbox_2_T3}), .clk (clk), .r (Fresh[368]), .c ({new_AGEMA_signal_6591, SubBytesIns_Inst_Sbox_2_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M59_U1 ( .a ({new_AGEMA_signal_6218, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_5187, SubBytesIns_Inst_Sbox_2_T22}), .clk (clk), .r (Fresh[369]), .c ({new_AGEMA_signal_6355, SubBytesIns_Inst_Sbox_2_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M60_U1 ( .a ({new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_5375, SubBytesIns_Inst_Sbox_2_T20}), .clk (clk), .r (Fresh[370]), .c ({new_AGEMA_signal_6356, SubBytesIns_Inst_Sbox_2_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M61_U1 ( .a ({new_AGEMA_signal_6346, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_4993, SubBytesIns_Inst_Sbox_2_T1}), .clk (clk), .r (Fresh[371]), .c ({new_AGEMA_signal_6592, SubBytesIns_Inst_Sbox_2_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M62_U1 ( .a ({new_AGEMA_signal_6585, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_4996, SubBytesIns_Inst_Sbox_2_T4}), .clk (clk), .r (Fresh[372]), .c ({new_AGEMA_signal_6814, SubBytesIns_Inst_Sbox_2_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M63_U1 ( .a ({new_AGEMA_signal_6345, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_4994, SubBytesIns_Inst_Sbox_2_T2}), .clk (clk), .r (Fresh[373]), .c ({new_AGEMA_signal_6593, SubBytesIns_Inst_Sbox_2_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L0_U1 ( .a ({new_AGEMA_signal_6592, SubBytesIns_Inst_Sbox_2_M61}), .b ({new_AGEMA_signal_6814, SubBytesIns_Inst_Sbox_2_M62}), .c ({new_AGEMA_signal_7007, SubBytesIns_Inst_Sbox_2_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L1_U1 ( .a ({new_AGEMA_signal_6351, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_6353, SubBytesIns_Inst_Sbox_2_M56}), .c ({new_AGEMA_signal_6594, SubBytesIns_Inst_Sbox_2_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L2_U1 ( .a ({new_AGEMA_signal_6586, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_6350, SubBytesIns_Inst_Sbox_2_M48}), .c ({new_AGEMA_signal_6815, SubBytesIns_Inst_Sbox_2_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L3_U1 ( .a ({new_AGEMA_signal_6349, SubBytesIns_Inst_Sbox_2_M47}), .b ({new_AGEMA_signal_6590, SubBytesIns_Inst_Sbox_2_M55}), .c ({new_AGEMA_signal_6816, SubBytesIns_Inst_Sbox_2_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L4_U1 ( .a ({new_AGEMA_signal_6589, SubBytesIns_Inst_Sbox_2_M54}), .b ({new_AGEMA_signal_6591, SubBytesIns_Inst_Sbox_2_M58}), .c ({new_AGEMA_signal_6817, SubBytesIns_Inst_Sbox_2_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L5_U1 ( .a ({new_AGEMA_signal_6587, SubBytesIns_Inst_Sbox_2_M49}), .b ({new_AGEMA_signal_6592, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_6818, SubBytesIns_Inst_Sbox_2_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L6_U1 ( .a ({new_AGEMA_signal_6814, SubBytesIns_Inst_Sbox_2_M62}), .b ({new_AGEMA_signal_6818, SubBytesIns_Inst_Sbox_2_L5}), .c ({new_AGEMA_signal_7008, SubBytesIns_Inst_Sbox_2_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L7_U1 ( .a ({new_AGEMA_signal_6586, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_6816, SubBytesIns_Inst_Sbox_2_L3}), .c ({new_AGEMA_signal_7009, SubBytesIns_Inst_Sbox_2_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L8_U1 ( .a ({new_AGEMA_signal_6352, SubBytesIns_Inst_Sbox_2_M51}), .b ({new_AGEMA_signal_6355, SubBytesIns_Inst_Sbox_2_M59}), .c ({new_AGEMA_signal_6595, SubBytesIns_Inst_Sbox_2_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L9_U1 ( .a ({new_AGEMA_signal_6588, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_6813, SubBytesIns_Inst_Sbox_2_M53}), .c ({new_AGEMA_signal_7010, SubBytesIns_Inst_Sbox_2_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L10_U1 ( .a ({new_AGEMA_signal_6813, SubBytesIns_Inst_Sbox_2_M53}), .b ({new_AGEMA_signal_6817, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_7011, SubBytesIns_Inst_Sbox_2_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L11_U1 ( .a ({new_AGEMA_signal_6356, SubBytesIns_Inst_Sbox_2_M60}), .b ({new_AGEMA_signal_6815, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_7012, SubBytesIns_Inst_Sbox_2_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L12_U1 ( .a ({new_AGEMA_signal_6350, SubBytesIns_Inst_Sbox_2_M48}), .b ({new_AGEMA_signal_6352, SubBytesIns_Inst_Sbox_2_M51}), .c ({new_AGEMA_signal_6596, SubBytesIns_Inst_Sbox_2_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L13_U1 ( .a ({new_AGEMA_signal_6351, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_7007, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_7199, SubBytesIns_Inst_Sbox_2_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L14_U1 ( .a ({new_AGEMA_signal_6588, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_6592, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_6819, SubBytesIns_Inst_Sbox_2_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L15_U1 ( .a ({new_AGEMA_signal_6590, SubBytesIns_Inst_Sbox_2_M55}), .b ({new_AGEMA_signal_6594, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_6820, SubBytesIns_Inst_Sbox_2_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L16_U1 ( .a ({new_AGEMA_signal_6353, SubBytesIns_Inst_Sbox_2_M56}), .b ({new_AGEMA_signal_7007, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_7200, SubBytesIns_Inst_Sbox_2_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L17_U1 ( .a ({new_AGEMA_signal_6354, SubBytesIns_Inst_Sbox_2_M57}), .b ({new_AGEMA_signal_6594, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_6821, SubBytesIns_Inst_Sbox_2_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L18_U1 ( .a ({new_AGEMA_signal_6591, SubBytesIns_Inst_Sbox_2_M58}), .b ({new_AGEMA_signal_6595, SubBytesIns_Inst_Sbox_2_L8}), .c ({new_AGEMA_signal_6822, SubBytesIns_Inst_Sbox_2_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L19_U1 ( .a ({new_AGEMA_signal_6593, SubBytesIns_Inst_Sbox_2_M63}), .b ({new_AGEMA_signal_6817, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_7013, SubBytesIns_Inst_Sbox_2_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L20_U1 ( .a ({new_AGEMA_signal_7007, SubBytesIns_Inst_Sbox_2_L0}), .b ({new_AGEMA_signal_6594, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_7201, SubBytesIns_Inst_Sbox_2_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L21_U1 ( .a ({new_AGEMA_signal_6594, SubBytesIns_Inst_Sbox_2_L1}), .b ({new_AGEMA_signal_7009, SubBytesIns_Inst_Sbox_2_L7}), .c ({new_AGEMA_signal_7202, SubBytesIns_Inst_Sbox_2_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L22_U1 ( .a ({new_AGEMA_signal_6816, SubBytesIns_Inst_Sbox_2_L3}), .b ({new_AGEMA_signal_6596, SubBytesIns_Inst_Sbox_2_L12}), .c ({new_AGEMA_signal_7014, SubBytesIns_Inst_Sbox_2_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L23_U1 ( .a ({new_AGEMA_signal_6822, SubBytesIns_Inst_Sbox_2_L18}), .b ({new_AGEMA_signal_6815, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_7015, SubBytesIns_Inst_Sbox_2_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L24_U1 ( .a ({new_AGEMA_signal_6820, SubBytesIns_Inst_Sbox_2_L15}), .b ({new_AGEMA_signal_7010, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_7203, SubBytesIns_Inst_Sbox_2_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L25_U1 ( .a ({new_AGEMA_signal_7008, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_7011, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_7204, SubBytesIns_Inst_Sbox_2_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L26_U1 ( .a ({new_AGEMA_signal_7009, SubBytesIns_Inst_Sbox_2_L7}), .b ({new_AGEMA_signal_7010, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_7205, SubBytesIns_Inst_Sbox_2_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L27_U1 ( .a ({new_AGEMA_signal_6595, SubBytesIns_Inst_Sbox_2_L8}), .b ({new_AGEMA_signal_7011, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_7206, SubBytesIns_Inst_Sbox_2_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L28_U1 ( .a ({new_AGEMA_signal_7012, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_6819, SubBytesIns_Inst_Sbox_2_L14}), .c ({new_AGEMA_signal_7207, SubBytesIns_Inst_Sbox_2_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L29_U1 ( .a ({new_AGEMA_signal_7012, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_6821, SubBytesIns_Inst_Sbox_2_L17}), .c ({new_AGEMA_signal_7208, SubBytesIns_Inst_Sbox_2_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S0_U1 ( .a ({new_AGEMA_signal_7008, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_7203, SubBytesIns_Inst_Sbox_2_L24}), .c ({new_AGEMA_signal_7399, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S1_U1 ( .a ({new_AGEMA_signal_7200, SubBytesIns_Inst_Sbox_2_L16}), .b ({new_AGEMA_signal_7205, SubBytesIns_Inst_Sbox_2_L26}), .c ({new_AGEMA_signal_7400, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S2_U1 ( .a ({new_AGEMA_signal_7013, SubBytesIns_Inst_Sbox_2_L19}), .b ({new_AGEMA_signal_7207, SubBytesIns_Inst_Sbox_2_L28}), .c ({new_AGEMA_signal_7401, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S3_U1 ( .a ({new_AGEMA_signal_7008, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_7202, SubBytesIns_Inst_Sbox_2_L21}), .c ({new_AGEMA_signal_7402, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S4_U1 ( .a ({new_AGEMA_signal_7201, SubBytesIns_Inst_Sbox_2_L20}), .b ({new_AGEMA_signal_7014, SubBytesIns_Inst_Sbox_2_L22}), .c ({new_AGEMA_signal_7403, MixColumnsInput[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S5_U1 ( .a ({new_AGEMA_signal_7204, SubBytesIns_Inst_Sbox_2_L25}), .b ({new_AGEMA_signal_7208, SubBytesIns_Inst_Sbox_2_L29}), .c ({new_AGEMA_signal_7404, MixColumnsInput[50]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S6_U1 ( .a ({new_AGEMA_signal_7199, SubBytesIns_Inst_Sbox_2_L13}), .b ({new_AGEMA_signal_7206, SubBytesIns_Inst_Sbox_2_L27}), .c ({new_AGEMA_signal_7405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S7_U1 ( .a ({new_AGEMA_signal_7008, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_7015, SubBytesIns_Inst_Sbox_2_L23}), .c ({new_AGEMA_signal_7209, MixColumnsInput[48]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M46_U1 ( .a ({new_AGEMA_signal_6360, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_5189, SubBytesIns_Inst_Sbox_3_T6}), .clk (clk), .r (Fresh[374]), .c ({new_AGEMA_signal_6598, SubBytesIns_Inst_Sbox_3_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M47_U1 ( .a ({new_AGEMA_signal_6224, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_5384, SubBytesIns_Inst_Sbox_3_T8}), .clk (clk), .r (Fresh[375]), .c ({new_AGEMA_signal_6361, SubBytesIns_Inst_Sbox_3_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M48_U1 ( .a ({new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_3_M39}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .clk (clk), .r (Fresh[376]), .c ({new_AGEMA_signal_6362, SubBytesIns_Inst_Sbox_3_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M49_U1 ( .a ({new_AGEMA_signal_6359, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_5193, SubBytesIns_Inst_Sbox_3_T16}), .clk (clk), .r (Fresh[377]), .c ({new_AGEMA_signal_6599, SubBytesIns_Inst_Sbox_3_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M50_U1 ( .a ({new_AGEMA_signal_6222, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_5190, SubBytesIns_Inst_Sbox_3_T9}), .clk (clk), .r (Fresh[378]), .c ({new_AGEMA_signal_6363, SubBytesIns_Inst_Sbox_3_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M51_U1 ( .a ({new_AGEMA_signal_6221, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_5387, SubBytesIns_Inst_Sbox_3_T17}), .clk (clk), .r (Fresh[379]), .c ({new_AGEMA_signal_6364, SubBytesIns_Inst_Sbox_3_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M52_U1 ( .a ({new_AGEMA_signal_6358, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_5192, SubBytesIns_Inst_Sbox_3_T15}), .clk (clk), .r (Fresh[380]), .c ({new_AGEMA_signal_6600, SubBytesIns_Inst_Sbox_3_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M53_U1 ( .a ({new_AGEMA_signal_6597, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_5196, SubBytesIns_Inst_Sbox_3_T27}), .clk (clk), .r (Fresh[381]), .c ({new_AGEMA_signal_6823, SubBytesIns_Inst_Sbox_3_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M54_U1 ( .a ({new_AGEMA_signal_6357, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_5385, SubBytesIns_Inst_Sbox_3_T10}), .clk (clk), .r (Fresh[382]), .c ({new_AGEMA_signal_6601, SubBytesIns_Inst_Sbox_3_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M55_U1 ( .a ({new_AGEMA_signal_6360, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_5191, SubBytesIns_Inst_Sbox_3_T13}), .clk (clk), .r (Fresh[383]), .c ({new_AGEMA_signal_6602, SubBytesIns_Inst_Sbox_3_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M56_U1 ( .a ({new_AGEMA_signal_6224, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_5389, SubBytesIns_Inst_Sbox_3_T23}), .clk (clk), .r (Fresh[384]), .c ({new_AGEMA_signal_6365, SubBytesIns_Inst_Sbox_3_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M57_U1 ( .a ({new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_5194, SubBytesIns_Inst_Sbox_3_T19}), .clk (clk), .r (Fresh[385]), .c ({new_AGEMA_signal_6366, SubBytesIns_Inst_Sbox_3_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M58_U1 ( .a ({new_AGEMA_signal_6359, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_5005, SubBytesIns_Inst_Sbox_3_T3}), .clk (clk), .r (Fresh[386]), .c ({new_AGEMA_signal_6603, SubBytesIns_Inst_Sbox_3_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M59_U1 ( .a ({new_AGEMA_signal_6222, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_5195, SubBytesIns_Inst_Sbox_3_T22}), .clk (clk), .r (Fresh[387]), .c ({new_AGEMA_signal_6367, SubBytesIns_Inst_Sbox_3_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M60_U1 ( .a ({new_AGEMA_signal_6221, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_5388, SubBytesIns_Inst_Sbox_3_T20}), .clk (clk), .r (Fresh[388]), .c ({new_AGEMA_signal_6368, SubBytesIns_Inst_Sbox_3_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M61_U1 ( .a ({new_AGEMA_signal_6358, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_5003, SubBytesIns_Inst_Sbox_3_T1}), .clk (clk), .r (Fresh[389]), .c ({new_AGEMA_signal_6604, SubBytesIns_Inst_Sbox_3_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M62_U1 ( .a ({new_AGEMA_signal_6597, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_5006, SubBytesIns_Inst_Sbox_3_T4}), .clk (clk), .r (Fresh[390]), .c ({new_AGEMA_signal_6824, SubBytesIns_Inst_Sbox_3_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M63_U1 ( .a ({new_AGEMA_signal_6357, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_5004, SubBytesIns_Inst_Sbox_3_T2}), .clk (clk), .r (Fresh[391]), .c ({new_AGEMA_signal_6605, SubBytesIns_Inst_Sbox_3_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L0_U1 ( .a ({new_AGEMA_signal_6604, SubBytesIns_Inst_Sbox_3_M61}), .b ({new_AGEMA_signal_6824, SubBytesIns_Inst_Sbox_3_M62}), .c ({new_AGEMA_signal_7016, SubBytesIns_Inst_Sbox_3_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L1_U1 ( .a ({new_AGEMA_signal_6363, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_6365, SubBytesIns_Inst_Sbox_3_M56}), .c ({new_AGEMA_signal_6606, SubBytesIns_Inst_Sbox_3_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L2_U1 ( .a ({new_AGEMA_signal_6598, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_6362, SubBytesIns_Inst_Sbox_3_M48}), .c ({new_AGEMA_signal_6825, SubBytesIns_Inst_Sbox_3_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L3_U1 ( .a ({new_AGEMA_signal_6361, SubBytesIns_Inst_Sbox_3_M47}), .b ({new_AGEMA_signal_6602, SubBytesIns_Inst_Sbox_3_M55}), .c ({new_AGEMA_signal_6826, SubBytesIns_Inst_Sbox_3_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L4_U1 ( .a ({new_AGEMA_signal_6601, SubBytesIns_Inst_Sbox_3_M54}), .b ({new_AGEMA_signal_6603, SubBytesIns_Inst_Sbox_3_M58}), .c ({new_AGEMA_signal_6827, SubBytesIns_Inst_Sbox_3_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L5_U1 ( .a ({new_AGEMA_signal_6599, SubBytesIns_Inst_Sbox_3_M49}), .b ({new_AGEMA_signal_6604, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_6828, SubBytesIns_Inst_Sbox_3_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L6_U1 ( .a ({new_AGEMA_signal_6824, SubBytesIns_Inst_Sbox_3_M62}), .b ({new_AGEMA_signal_6828, SubBytesIns_Inst_Sbox_3_L5}), .c ({new_AGEMA_signal_7017, SubBytesIns_Inst_Sbox_3_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L7_U1 ( .a ({new_AGEMA_signal_6598, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_6826, SubBytesIns_Inst_Sbox_3_L3}), .c ({new_AGEMA_signal_7018, SubBytesIns_Inst_Sbox_3_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L8_U1 ( .a ({new_AGEMA_signal_6364, SubBytesIns_Inst_Sbox_3_M51}), .b ({new_AGEMA_signal_6367, SubBytesIns_Inst_Sbox_3_M59}), .c ({new_AGEMA_signal_6607, SubBytesIns_Inst_Sbox_3_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L9_U1 ( .a ({new_AGEMA_signal_6600, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_6823, SubBytesIns_Inst_Sbox_3_M53}), .c ({new_AGEMA_signal_7019, SubBytesIns_Inst_Sbox_3_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L10_U1 ( .a ({new_AGEMA_signal_6823, SubBytesIns_Inst_Sbox_3_M53}), .b ({new_AGEMA_signal_6827, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_7020, SubBytesIns_Inst_Sbox_3_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L11_U1 ( .a ({new_AGEMA_signal_6368, SubBytesIns_Inst_Sbox_3_M60}), .b ({new_AGEMA_signal_6825, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_7021, SubBytesIns_Inst_Sbox_3_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L12_U1 ( .a ({new_AGEMA_signal_6362, SubBytesIns_Inst_Sbox_3_M48}), .b ({new_AGEMA_signal_6364, SubBytesIns_Inst_Sbox_3_M51}), .c ({new_AGEMA_signal_6608, SubBytesIns_Inst_Sbox_3_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L13_U1 ( .a ({new_AGEMA_signal_6363, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_7016, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_7210, SubBytesIns_Inst_Sbox_3_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L14_U1 ( .a ({new_AGEMA_signal_6600, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_6604, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_6829, SubBytesIns_Inst_Sbox_3_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L15_U1 ( .a ({new_AGEMA_signal_6602, SubBytesIns_Inst_Sbox_3_M55}), .b ({new_AGEMA_signal_6606, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_6830, SubBytesIns_Inst_Sbox_3_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L16_U1 ( .a ({new_AGEMA_signal_6365, SubBytesIns_Inst_Sbox_3_M56}), .b ({new_AGEMA_signal_7016, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_7211, SubBytesIns_Inst_Sbox_3_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L17_U1 ( .a ({new_AGEMA_signal_6366, SubBytesIns_Inst_Sbox_3_M57}), .b ({new_AGEMA_signal_6606, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_6831, SubBytesIns_Inst_Sbox_3_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L18_U1 ( .a ({new_AGEMA_signal_6603, SubBytesIns_Inst_Sbox_3_M58}), .b ({new_AGEMA_signal_6607, SubBytesIns_Inst_Sbox_3_L8}), .c ({new_AGEMA_signal_6832, SubBytesIns_Inst_Sbox_3_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L19_U1 ( .a ({new_AGEMA_signal_6605, SubBytesIns_Inst_Sbox_3_M63}), .b ({new_AGEMA_signal_6827, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_7022, SubBytesIns_Inst_Sbox_3_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L20_U1 ( .a ({new_AGEMA_signal_7016, SubBytesIns_Inst_Sbox_3_L0}), .b ({new_AGEMA_signal_6606, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_7212, SubBytesIns_Inst_Sbox_3_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L21_U1 ( .a ({new_AGEMA_signal_6606, SubBytesIns_Inst_Sbox_3_L1}), .b ({new_AGEMA_signal_7018, SubBytesIns_Inst_Sbox_3_L7}), .c ({new_AGEMA_signal_7213, SubBytesIns_Inst_Sbox_3_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L22_U1 ( .a ({new_AGEMA_signal_6826, SubBytesIns_Inst_Sbox_3_L3}), .b ({new_AGEMA_signal_6608, SubBytesIns_Inst_Sbox_3_L12}), .c ({new_AGEMA_signal_7023, SubBytesIns_Inst_Sbox_3_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L23_U1 ( .a ({new_AGEMA_signal_6832, SubBytesIns_Inst_Sbox_3_L18}), .b ({new_AGEMA_signal_6825, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_7024, SubBytesIns_Inst_Sbox_3_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L24_U1 ( .a ({new_AGEMA_signal_6830, SubBytesIns_Inst_Sbox_3_L15}), .b ({new_AGEMA_signal_7019, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_7214, SubBytesIns_Inst_Sbox_3_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L25_U1 ( .a ({new_AGEMA_signal_7017, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_7020, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_7215, SubBytesIns_Inst_Sbox_3_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L26_U1 ( .a ({new_AGEMA_signal_7018, SubBytesIns_Inst_Sbox_3_L7}), .b ({new_AGEMA_signal_7019, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_7216, SubBytesIns_Inst_Sbox_3_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L27_U1 ( .a ({new_AGEMA_signal_6607, SubBytesIns_Inst_Sbox_3_L8}), .b ({new_AGEMA_signal_7020, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_7217, SubBytesIns_Inst_Sbox_3_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L28_U1 ( .a ({new_AGEMA_signal_7021, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_6829, SubBytesIns_Inst_Sbox_3_L14}), .c ({new_AGEMA_signal_7218, SubBytesIns_Inst_Sbox_3_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L29_U1 ( .a ({new_AGEMA_signal_7021, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_6831, SubBytesIns_Inst_Sbox_3_L17}), .c ({new_AGEMA_signal_7219, SubBytesIns_Inst_Sbox_3_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S0_U1 ( .a ({new_AGEMA_signal_7017, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_7214, SubBytesIns_Inst_Sbox_3_L24}), .c ({new_AGEMA_signal_7406, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S1_U1 ( .a ({new_AGEMA_signal_7211, SubBytesIns_Inst_Sbox_3_L16}), .b ({new_AGEMA_signal_7216, SubBytesIns_Inst_Sbox_3_L26}), .c ({new_AGEMA_signal_7407, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S2_U1 ( .a ({new_AGEMA_signal_7022, SubBytesIns_Inst_Sbox_3_L19}), .b ({new_AGEMA_signal_7218, SubBytesIns_Inst_Sbox_3_L28}), .c ({new_AGEMA_signal_7408, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S3_U1 ( .a ({new_AGEMA_signal_7017, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_7213, SubBytesIns_Inst_Sbox_3_L21}), .c ({new_AGEMA_signal_7409, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S4_U1 ( .a ({new_AGEMA_signal_7212, SubBytesIns_Inst_Sbox_3_L20}), .b ({new_AGEMA_signal_7023, SubBytesIns_Inst_Sbox_3_L22}), .c ({new_AGEMA_signal_7410, MixColumnsInput[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S5_U1 ( .a ({new_AGEMA_signal_7215, SubBytesIns_Inst_Sbox_3_L25}), .b ({new_AGEMA_signal_7219, SubBytesIns_Inst_Sbox_3_L29}), .c ({new_AGEMA_signal_7411, MixColumnsInput[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S6_U1 ( .a ({new_AGEMA_signal_7210, SubBytesIns_Inst_Sbox_3_L13}), .b ({new_AGEMA_signal_7217, SubBytesIns_Inst_Sbox_3_L27}), .c ({new_AGEMA_signal_7412, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S7_U1 ( .a ({new_AGEMA_signal_7017, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_7024, SubBytesIns_Inst_Sbox_3_L23}), .c ({new_AGEMA_signal_7220, MixColumnsInput[24]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M46_U1 ( .a ({new_AGEMA_signal_6372, SubBytesIns_Inst_Sbox_4_M44}), .b ({new_AGEMA_signal_5197, SubBytesIns_Inst_Sbox_4_T6}), .clk (clk), .r (Fresh[392]), .c ({new_AGEMA_signal_6610, SubBytesIns_Inst_Sbox_4_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M47_U1 ( .a ({new_AGEMA_signal_6228, SubBytesIns_Inst_Sbox_4_M40}), .b ({new_AGEMA_signal_5397, SubBytesIns_Inst_Sbox_4_T8}), .clk (clk), .r (Fresh[393]), .c ({new_AGEMA_signal_6373, SubBytesIns_Inst_Sbox_4_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M48_U1 ( .a ({new_AGEMA_signal_6227, SubBytesIns_Inst_Sbox_4_M39}), .b ({ciphertext_s1[32], ciphertext_s0[32]}), .clk (clk), .r (Fresh[394]), .c ({new_AGEMA_signal_6374, SubBytesIns_Inst_Sbox_4_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M49_U1 ( .a ({new_AGEMA_signal_6371, SubBytesIns_Inst_Sbox_4_M43}), .b ({new_AGEMA_signal_5201, SubBytesIns_Inst_Sbox_4_T16}), .clk (clk), .r (Fresh[395]), .c ({new_AGEMA_signal_6611, SubBytesIns_Inst_Sbox_4_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M50_U1 ( .a ({new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_4_M38}), .b ({new_AGEMA_signal_5198, SubBytesIns_Inst_Sbox_4_T9}), .clk (clk), .r (Fresh[396]), .c ({new_AGEMA_signal_6375, SubBytesIns_Inst_Sbox_4_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M51_U1 ( .a ({new_AGEMA_signal_6225, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_5400, SubBytesIns_Inst_Sbox_4_T17}), .clk (clk), .r (Fresh[397]), .c ({new_AGEMA_signal_6376, SubBytesIns_Inst_Sbox_4_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M52_U1 ( .a ({new_AGEMA_signal_6370, SubBytesIns_Inst_Sbox_4_M42}), .b ({new_AGEMA_signal_5200, SubBytesIns_Inst_Sbox_4_T15}), .clk (clk), .r (Fresh[398]), .c ({new_AGEMA_signal_6612, SubBytesIns_Inst_Sbox_4_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M53_U1 ( .a ({new_AGEMA_signal_6609, SubBytesIns_Inst_Sbox_4_M45}), .b ({new_AGEMA_signal_5204, SubBytesIns_Inst_Sbox_4_T27}), .clk (clk), .r (Fresh[399]), .c ({new_AGEMA_signal_6833, SubBytesIns_Inst_Sbox_4_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M54_U1 ( .a ({new_AGEMA_signal_6369, SubBytesIns_Inst_Sbox_4_M41}), .b ({new_AGEMA_signal_5398, SubBytesIns_Inst_Sbox_4_T10}), .clk (clk), .r (Fresh[400]), .c ({new_AGEMA_signal_6613, SubBytesIns_Inst_Sbox_4_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M55_U1 ( .a ({new_AGEMA_signal_6372, SubBytesIns_Inst_Sbox_4_M44}), .b ({new_AGEMA_signal_5199, SubBytesIns_Inst_Sbox_4_T13}), .clk (clk), .r (Fresh[401]), .c ({new_AGEMA_signal_6614, SubBytesIns_Inst_Sbox_4_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M56_U1 ( .a ({new_AGEMA_signal_6228, SubBytesIns_Inst_Sbox_4_M40}), .b ({new_AGEMA_signal_5402, SubBytesIns_Inst_Sbox_4_T23}), .clk (clk), .r (Fresh[402]), .c ({new_AGEMA_signal_6377, SubBytesIns_Inst_Sbox_4_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M57_U1 ( .a ({new_AGEMA_signal_6227, SubBytesIns_Inst_Sbox_4_M39}), .b ({new_AGEMA_signal_5202, SubBytesIns_Inst_Sbox_4_T19}), .clk (clk), .r (Fresh[403]), .c ({new_AGEMA_signal_6378, SubBytesIns_Inst_Sbox_4_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M58_U1 ( .a ({new_AGEMA_signal_6371, SubBytesIns_Inst_Sbox_4_M43}), .b ({new_AGEMA_signal_5015, SubBytesIns_Inst_Sbox_4_T3}), .clk (clk), .r (Fresh[404]), .c ({new_AGEMA_signal_6615, SubBytesIns_Inst_Sbox_4_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M59_U1 ( .a ({new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_4_M38}), .b ({new_AGEMA_signal_5203, SubBytesIns_Inst_Sbox_4_T22}), .clk (clk), .r (Fresh[405]), .c ({new_AGEMA_signal_6379, SubBytesIns_Inst_Sbox_4_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M60_U1 ( .a ({new_AGEMA_signal_6225, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_5401, SubBytesIns_Inst_Sbox_4_T20}), .clk (clk), .r (Fresh[406]), .c ({new_AGEMA_signal_6380, SubBytesIns_Inst_Sbox_4_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M61_U1 ( .a ({new_AGEMA_signal_6370, SubBytesIns_Inst_Sbox_4_M42}), .b ({new_AGEMA_signal_5013, SubBytesIns_Inst_Sbox_4_T1}), .clk (clk), .r (Fresh[407]), .c ({new_AGEMA_signal_6616, SubBytesIns_Inst_Sbox_4_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M62_U1 ( .a ({new_AGEMA_signal_6609, SubBytesIns_Inst_Sbox_4_M45}), .b ({new_AGEMA_signal_5016, SubBytesIns_Inst_Sbox_4_T4}), .clk (clk), .r (Fresh[408]), .c ({new_AGEMA_signal_6834, SubBytesIns_Inst_Sbox_4_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M63_U1 ( .a ({new_AGEMA_signal_6369, SubBytesIns_Inst_Sbox_4_M41}), .b ({new_AGEMA_signal_5014, SubBytesIns_Inst_Sbox_4_T2}), .clk (clk), .r (Fresh[409]), .c ({new_AGEMA_signal_6617, SubBytesIns_Inst_Sbox_4_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L0_U1 ( .a ({new_AGEMA_signal_6616, SubBytesIns_Inst_Sbox_4_M61}), .b ({new_AGEMA_signal_6834, SubBytesIns_Inst_Sbox_4_M62}), .c ({new_AGEMA_signal_7025, SubBytesIns_Inst_Sbox_4_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L1_U1 ( .a ({new_AGEMA_signal_6375, SubBytesIns_Inst_Sbox_4_M50}), .b ({new_AGEMA_signal_6377, SubBytesIns_Inst_Sbox_4_M56}), .c ({new_AGEMA_signal_6618, SubBytesIns_Inst_Sbox_4_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L2_U1 ( .a ({new_AGEMA_signal_6610, SubBytesIns_Inst_Sbox_4_M46}), .b ({new_AGEMA_signal_6374, SubBytesIns_Inst_Sbox_4_M48}), .c ({new_AGEMA_signal_6835, SubBytesIns_Inst_Sbox_4_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L3_U1 ( .a ({new_AGEMA_signal_6373, SubBytesIns_Inst_Sbox_4_M47}), .b ({new_AGEMA_signal_6614, SubBytesIns_Inst_Sbox_4_M55}), .c ({new_AGEMA_signal_6836, SubBytesIns_Inst_Sbox_4_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L4_U1 ( .a ({new_AGEMA_signal_6613, SubBytesIns_Inst_Sbox_4_M54}), .b ({new_AGEMA_signal_6615, SubBytesIns_Inst_Sbox_4_M58}), .c ({new_AGEMA_signal_6837, SubBytesIns_Inst_Sbox_4_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L5_U1 ( .a ({new_AGEMA_signal_6611, SubBytesIns_Inst_Sbox_4_M49}), .b ({new_AGEMA_signal_6616, SubBytesIns_Inst_Sbox_4_M61}), .c ({new_AGEMA_signal_6838, SubBytesIns_Inst_Sbox_4_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L6_U1 ( .a ({new_AGEMA_signal_6834, SubBytesIns_Inst_Sbox_4_M62}), .b ({new_AGEMA_signal_6838, SubBytesIns_Inst_Sbox_4_L5}), .c ({new_AGEMA_signal_7026, SubBytesIns_Inst_Sbox_4_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L7_U1 ( .a ({new_AGEMA_signal_6610, SubBytesIns_Inst_Sbox_4_M46}), .b ({new_AGEMA_signal_6836, SubBytesIns_Inst_Sbox_4_L3}), .c ({new_AGEMA_signal_7027, SubBytesIns_Inst_Sbox_4_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L8_U1 ( .a ({new_AGEMA_signal_6376, SubBytesIns_Inst_Sbox_4_M51}), .b ({new_AGEMA_signal_6379, SubBytesIns_Inst_Sbox_4_M59}), .c ({new_AGEMA_signal_6619, SubBytesIns_Inst_Sbox_4_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L9_U1 ( .a ({new_AGEMA_signal_6612, SubBytesIns_Inst_Sbox_4_M52}), .b ({new_AGEMA_signal_6833, SubBytesIns_Inst_Sbox_4_M53}), .c ({new_AGEMA_signal_7028, SubBytesIns_Inst_Sbox_4_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L10_U1 ( .a ({new_AGEMA_signal_6833, SubBytesIns_Inst_Sbox_4_M53}), .b ({new_AGEMA_signal_6837, SubBytesIns_Inst_Sbox_4_L4}), .c ({new_AGEMA_signal_7029, SubBytesIns_Inst_Sbox_4_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L11_U1 ( .a ({new_AGEMA_signal_6380, SubBytesIns_Inst_Sbox_4_M60}), .b ({new_AGEMA_signal_6835, SubBytesIns_Inst_Sbox_4_L2}), .c ({new_AGEMA_signal_7030, SubBytesIns_Inst_Sbox_4_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L12_U1 ( .a ({new_AGEMA_signal_6374, SubBytesIns_Inst_Sbox_4_M48}), .b ({new_AGEMA_signal_6376, SubBytesIns_Inst_Sbox_4_M51}), .c ({new_AGEMA_signal_6620, SubBytesIns_Inst_Sbox_4_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L13_U1 ( .a ({new_AGEMA_signal_6375, SubBytesIns_Inst_Sbox_4_M50}), .b ({new_AGEMA_signal_7025, SubBytesIns_Inst_Sbox_4_L0}), .c ({new_AGEMA_signal_7221, SubBytesIns_Inst_Sbox_4_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L14_U1 ( .a ({new_AGEMA_signal_6612, SubBytesIns_Inst_Sbox_4_M52}), .b ({new_AGEMA_signal_6616, SubBytesIns_Inst_Sbox_4_M61}), .c ({new_AGEMA_signal_6839, SubBytesIns_Inst_Sbox_4_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L15_U1 ( .a ({new_AGEMA_signal_6614, SubBytesIns_Inst_Sbox_4_M55}), .b ({new_AGEMA_signal_6618, SubBytesIns_Inst_Sbox_4_L1}), .c ({new_AGEMA_signal_6840, SubBytesIns_Inst_Sbox_4_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L16_U1 ( .a ({new_AGEMA_signal_6377, SubBytesIns_Inst_Sbox_4_M56}), .b ({new_AGEMA_signal_7025, SubBytesIns_Inst_Sbox_4_L0}), .c ({new_AGEMA_signal_7222, SubBytesIns_Inst_Sbox_4_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L17_U1 ( .a ({new_AGEMA_signal_6378, SubBytesIns_Inst_Sbox_4_M57}), .b ({new_AGEMA_signal_6618, SubBytesIns_Inst_Sbox_4_L1}), .c ({new_AGEMA_signal_6841, SubBytesIns_Inst_Sbox_4_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L18_U1 ( .a ({new_AGEMA_signal_6615, SubBytesIns_Inst_Sbox_4_M58}), .b ({new_AGEMA_signal_6619, SubBytesIns_Inst_Sbox_4_L8}), .c ({new_AGEMA_signal_6842, SubBytesIns_Inst_Sbox_4_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L19_U1 ( .a ({new_AGEMA_signal_6617, SubBytesIns_Inst_Sbox_4_M63}), .b ({new_AGEMA_signal_6837, SubBytesIns_Inst_Sbox_4_L4}), .c ({new_AGEMA_signal_7031, SubBytesIns_Inst_Sbox_4_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L20_U1 ( .a ({new_AGEMA_signal_7025, SubBytesIns_Inst_Sbox_4_L0}), .b ({new_AGEMA_signal_6618, SubBytesIns_Inst_Sbox_4_L1}), .c ({new_AGEMA_signal_7223, SubBytesIns_Inst_Sbox_4_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L21_U1 ( .a ({new_AGEMA_signal_6618, SubBytesIns_Inst_Sbox_4_L1}), .b ({new_AGEMA_signal_7027, SubBytesIns_Inst_Sbox_4_L7}), .c ({new_AGEMA_signal_7224, SubBytesIns_Inst_Sbox_4_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L22_U1 ( .a ({new_AGEMA_signal_6836, SubBytesIns_Inst_Sbox_4_L3}), .b ({new_AGEMA_signal_6620, SubBytesIns_Inst_Sbox_4_L12}), .c ({new_AGEMA_signal_7032, SubBytesIns_Inst_Sbox_4_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L23_U1 ( .a ({new_AGEMA_signal_6842, SubBytesIns_Inst_Sbox_4_L18}), .b ({new_AGEMA_signal_6835, SubBytesIns_Inst_Sbox_4_L2}), .c ({new_AGEMA_signal_7033, SubBytesIns_Inst_Sbox_4_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L24_U1 ( .a ({new_AGEMA_signal_6840, SubBytesIns_Inst_Sbox_4_L15}), .b ({new_AGEMA_signal_7028, SubBytesIns_Inst_Sbox_4_L9}), .c ({new_AGEMA_signal_7225, SubBytesIns_Inst_Sbox_4_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L25_U1 ( .a ({new_AGEMA_signal_7026, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_7029, SubBytesIns_Inst_Sbox_4_L10}), .c ({new_AGEMA_signal_7226, SubBytesIns_Inst_Sbox_4_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L26_U1 ( .a ({new_AGEMA_signal_7027, SubBytesIns_Inst_Sbox_4_L7}), .b ({new_AGEMA_signal_7028, SubBytesIns_Inst_Sbox_4_L9}), .c ({new_AGEMA_signal_7227, SubBytesIns_Inst_Sbox_4_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L27_U1 ( .a ({new_AGEMA_signal_6619, SubBytesIns_Inst_Sbox_4_L8}), .b ({new_AGEMA_signal_7029, SubBytesIns_Inst_Sbox_4_L10}), .c ({new_AGEMA_signal_7228, SubBytesIns_Inst_Sbox_4_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L28_U1 ( .a ({new_AGEMA_signal_7030, SubBytesIns_Inst_Sbox_4_L11}), .b ({new_AGEMA_signal_6839, SubBytesIns_Inst_Sbox_4_L14}), .c ({new_AGEMA_signal_7229, SubBytesIns_Inst_Sbox_4_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L29_U1 ( .a ({new_AGEMA_signal_7030, SubBytesIns_Inst_Sbox_4_L11}), .b ({new_AGEMA_signal_6841, SubBytesIns_Inst_Sbox_4_L17}), .c ({new_AGEMA_signal_7230, SubBytesIns_Inst_Sbox_4_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S0_U1 ( .a ({new_AGEMA_signal_7026, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_7225, SubBytesIns_Inst_Sbox_4_L24}), .c ({new_AGEMA_signal_7413, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S1_U1 ( .a ({new_AGEMA_signal_7222, SubBytesIns_Inst_Sbox_4_L16}), .b ({new_AGEMA_signal_7227, SubBytesIns_Inst_Sbox_4_L26}), .c ({new_AGEMA_signal_7414, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S2_U1 ( .a ({new_AGEMA_signal_7031, SubBytesIns_Inst_Sbox_4_L19}), .b ({new_AGEMA_signal_7229, SubBytesIns_Inst_Sbox_4_L28}), .c ({new_AGEMA_signal_7415, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S3_U1 ( .a ({new_AGEMA_signal_7026, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_7224, SubBytesIns_Inst_Sbox_4_L21}), .c ({new_AGEMA_signal_7416, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S4_U1 ( .a ({new_AGEMA_signal_7223, SubBytesIns_Inst_Sbox_4_L20}), .b ({new_AGEMA_signal_7032, SubBytesIns_Inst_Sbox_4_L22}), .c ({new_AGEMA_signal_7417, MixColumnsInput[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S5_U1 ( .a ({new_AGEMA_signal_7226, SubBytesIns_Inst_Sbox_4_L25}), .b ({new_AGEMA_signal_7230, SubBytesIns_Inst_Sbox_4_L29}), .c ({new_AGEMA_signal_7418, MixColumnsInput[2]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S6_U1 ( .a ({new_AGEMA_signal_7221, SubBytesIns_Inst_Sbox_4_L13}), .b ({new_AGEMA_signal_7228, SubBytesIns_Inst_Sbox_4_L27}), .c ({new_AGEMA_signal_7419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S7_U1 ( .a ({new_AGEMA_signal_7026, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_7033, SubBytesIns_Inst_Sbox_4_L23}), .c ({new_AGEMA_signal_7231, MixColumnsInput[0]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M46_U1 ( .a ({new_AGEMA_signal_6384, SubBytesIns_Inst_Sbox_5_M44}), .b ({new_AGEMA_signal_5205, SubBytesIns_Inst_Sbox_5_T6}), .clk (clk), .r (Fresh[410]), .c ({new_AGEMA_signal_6622, SubBytesIns_Inst_Sbox_5_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M47_U1 ( .a ({new_AGEMA_signal_6232, SubBytesIns_Inst_Sbox_5_M40}), .b ({new_AGEMA_signal_5410, SubBytesIns_Inst_Sbox_5_T8}), .clk (clk), .r (Fresh[411]), .c ({new_AGEMA_signal_6385, SubBytesIns_Inst_Sbox_5_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M48_U1 ( .a ({new_AGEMA_signal_6231, SubBytesIns_Inst_Sbox_5_M39}), .b ({ciphertext_s1[40], ciphertext_s0[40]}), .clk (clk), .r (Fresh[412]), .c ({new_AGEMA_signal_6386, SubBytesIns_Inst_Sbox_5_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M49_U1 ( .a ({new_AGEMA_signal_6383, SubBytesIns_Inst_Sbox_5_M43}), .b ({new_AGEMA_signal_5209, SubBytesIns_Inst_Sbox_5_T16}), .clk (clk), .r (Fresh[413]), .c ({new_AGEMA_signal_6623, SubBytesIns_Inst_Sbox_5_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M50_U1 ( .a ({new_AGEMA_signal_6230, SubBytesIns_Inst_Sbox_5_M38}), .b ({new_AGEMA_signal_5206, SubBytesIns_Inst_Sbox_5_T9}), .clk (clk), .r (Fresh[414]), .c ({new_AGEMA_signal_6387, SubBytesIns_Inst_Sbox_5_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M51_U1 ( .a ({new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_5413, SubBytesIns_Inst_Sbox_5_T17}), .clk (clk), .r (Fresh[415]), .c ({new_AGEMA_signal_6388, SubBytesIns_Inst_Sbox_5_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M52_U1 ( .a ({new_AGEMA_signal_6382, SubBytesIns_Inst_Sbox_5_M42}), .b ({new_AGEMA_signal_5208, SubBytesIns_Inst_Sbox_5_T15}), .clk (clk), .r (Fresh[416]), .c ({new_AGEMA_signal_6624, SubBytesIns_Inst_Sbox_5_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M53_U1 ( .a ({new_AGEMA_signal_6621, SubBytesIns_Inst_Sbox_5_M45}), .b ({new_AGEMA_signal_5212, SubBytesIns_Inst_Sbox_5_T27}), .clk (clk), .r (Fresh[417]), .c ({new_AGEMA_signal_6843, SubBytesIns_Inst_Sbox_5_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M54_U1 ( .a ({new_AGEMA_signal_6381, SubBytesIns_Inst_Sbox_5_M41}), .b ({new_AGEMA_signal_5411, SubBytesIns_Inst_Sbox_5_T10}), .clk (clk), .r (Fresh[418]), .c ({new_AGEMA_signal_6625, SubBytesIns_Inst_Sbox_5_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M55_U1 ( .a ({new_AGEMA_signal_6384, SubBytesIns_Inst_Sbox_5_M44}), .b ({new_AGEMA_signal_5207, SubBytesIns_Inst_Sbox_5_T13}), .clk (clk), .r (Fresh[419]), .c ({new_AGEMA_signal_6626, SubBytesIns_Inst_Sbox_5_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M56_U1 ( .a ({new_AGEMA_signal_6232, SubBytesIns_Inst_Sbox_5_M40}), .b ({new_AGEMA_signal_5415, SubBytesIns_Inst_Sbox_5_T23}), .clk (clk), .r (Fresh[420]), .c ({new_AGEMA_signal_6389, SubBytesIns_Inst_Sbox_5_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M57_U1 ( .a ({new_AGEMA_signal_6231, SubBytesIns_Inst_Sbox_5_M39}), .b ({new_AGEMA_signal_5210, SubBytesIns_Inst_Sbox_5_T19}), .clk (clk), .r (Fresh[421]), .c ({new_AGEMA_signal_6390, SubBytesIns_Inst_Sbox_5_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M58_U1 ( .a ({new_AGEMA_signal_6383, SubBytesIns_Inst_Sbox_5_M43}), .b ({new_AGEMA_signal_5025, SubBytesIns_Inst_Sbox_5_T3}), .clk (clk), .r (Fresh[422]), .c ({new_AGEMA_signal_6627, SubBytesIns_Inst_Sbox_5_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M59_U1 ( .a ({new_AGEMA_signal_6230, SubBytesIns_Inst_Sbox_5_M38}), .b ({new_AGEMA_signal_5211, SubBytesIns_Inst_Sbox_5_T22}), .clk (clk), .r (Fresh[423]), .c ({new_AGEMA_signal_6391, SubBytesIns_Inst_Sbox_5_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M60_U1 ( .a ({new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_5414, SubBytesIns_Inst_Sbox_5_T20}), .clk (clk), .r (Fresh[424]), .c ({new_AGEMA_signal_6392, SubBytesIns_Inst_Sbox_5_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M61_U1 ( .a ({new_AGEMA_signal_6382, SubBytesIns_Inst_Sbox_5_M42}), .b ({new_AGEMA_signal_5023, SubBytesIns_Inst_Sbox_5_T1}), .clk (clk), .r (Fresh[425]), .c ({new_AGEMA_signal_6628, SubBytesIns_Inst_Sbox_5_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M62_U1 ( .a ({new_AGEMA_signal_6621, SubBytesIns_Inst_Sbox_5_M45}), .b ({new_AGEMA_signal_5026, SubBytesIns_Inst_Sbox_5_T4}), .clk (clk), .r (Fresh[426]), .c ({new_AGEMA_signal_6844, SubBytesIns_Inst_Sbox_5_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M63_U1 ( .a ({new_AGEMA_signal_6381, SubBytesIns_Inst_Sbox_5_M41}), .b ({new_AGEMA_signal_5024, SubBytesIns_Inst_Sbox_5_T2}), .clk (clk), .r (Fresh[427]), .c ({new_AGEMA_signal_6629, SubBytesIns_Inst_Sbox_5_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L0_U1 ( .a ({new_AGEMA_signal_6628, SubBytesIns_Inst_Sbox_5_M61}), .b ({new_AGEMA_signal_6844, SubBytesIns_Inst_Sbox_5_M62}), .c ({new_AGEMA_signal_7034, SubBytesIns_Inst_Sbox_5_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L1_U1 ( .a ({new_AGEMA_signal_6387, SubBytesIns_Inst_Sbox_5_M50}), .b ({new_AGEMA_signal_6389, SubBytesIns_Inst_Sbox_5_M56}), .c ({new_AGEMA_signal_6630, SubBytesIns_Inst_Sbox_5_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L2_U1 ( .a ({new_AGEMA_signal_6622, SubBytesIns_Inst_Sbox_5_M46}), .b ({new_AGEMA_signal_6386, SubBytesIns_Inst_Sbox_5_M48}), .c ({new_AGEMA_signal_6845, SubBytesIns_Inst_Sbox_5_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L3_U1 ( .a ({new_AGEMA_signal_6385, SubBytesIns_Inst_Sbox_5_M47}), .b ({new_AGEMA_signal_6626, SubBytesIns_Inst_Sbox_5_M55}), .c ({new_AGEMA_signal_6846, SubBytesIns_Inst_Sbox_5_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L4_U1 ( .a ({new_AGEMA_signal_6625, SubBytesIns_Inst_Sbox_5_M54}), .b ({new_AGEMA_signal_6627, SubBytesIns_Inst_Sbox_5_M58}), .c ({new_AGEMA_signal_6847, SubBytesIns_Inst_Sbox_5_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L5_U1 ( .a ({new_AGEMA_signal_6623, SubBytesIns_Inst_Sbox_5_M49}), .b ({new_AGEMA_signal_6628, SubBytesIns_Inst_Sbox_5_M61}), .c ({new_AGEMA_signal_6848, SubBytesIns_Inst_Sbox_5_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L6_U1 ( .a ({new_AGEMA_signal_6844, SubBytesIns_Inst_Sbox_5_M62}), .b ({new_AGEMA_signal_6848, SubBytesIns_Inst_Sbox_5_L5}), .c ({new_AGEMA_signal_7035, SubBytesIns_Inst_Sbox_5_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L7_U1 ( .a ({new_AGEMA_signal_6622, SubBytesIns_Inst_Sbox_5_M46}), .b ({new_AGEMA_signal_6846, SubBytesIns_Inst_Sbox_5_L3}), .c ({new_AGEMA_signal_7036, SubBytesIns_Inst_Sbox_5_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L8_U1 ( .a ({new_AGEMA_signal_6388, SubBytesIns_Inst_Sbox_5_M51}), .b ({new_AGEMA_signal_6391, SubBytesIns_Inst_Sbox_5_M59}), .c ({new_AGEMA_signal_6631, SubBytesIns_Inst_Sbox_5_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L9_U1 ( .a ({new_AGEMA_signal_6624, SubBytesIns_Inst_Sbox_5_M52}), .b ({new_AGEMA_signal_6843, SubBytesIns_Inst_Sbox_5_M53}), .c ({new_AGEMA_signal_7037, SubBytesIns_Inst_Sbox_5_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L10_U1 ( .a ({new_AGEMA_signal_6843, SubBytesIns_Inst_Sbox_5_M53}), .b ({new_AGEMA_signal_6847, SubBytesIns_Inst_Sbox_5_L4}), .c ({new_AGEMA_signal_7038, SubBytesIns_Inst_Sbox_5_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L11_U1 ( .a ({new_AGEMA_signal_6392, SubBytesIns_Inst_Sbox_5_M60}), .b ({new_AGEMA_signal_6845, SubBytesIns_Inst_Sbox_5_L2}), .c ({new_AGEMA_signal_7039, SubBytesIns_Inst_Sbox_5_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L12_U1 ( .a ({new_AGEMA_signal_6386, SubBytesIns_Inst_Sbox_5_M48}), .b ({new_AGEMA_signal_6388, SubBytesIns_Inst_Sbox_5_M51}), .c ({new_AGEMA_signal_6632, SubBytesIns_Inst_Sbox_5_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L13_U1 ( .a ({new_AGEMA_signal_6387, SubBytesIns_Inst_Sbox_5_M50}), .b ({new_AGEMA_signal_7034, SubBytesIns_Inst_Sbox_5_L0}), .c ({new_AGEMA_signal_7232, SubBytesIns_Inst_Sbox_5_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L14_U1 ( .a ({new_AGEMA_signal_6624, SubBytesIns_Inst_Sbox_5_M52}), .b ({new_AGEMA_signal_6628, SubBytesIns_Inst_Sbox_5_M61}), .c ({new_AGEMA_signal_6849, SubBytesIns_Inst_Sbox_5_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L15_U1 ( .a ({new_AGEMA_signal_6626, SubBytesIns_Inst_Sbox_5_M55}), .b ({new_AGEMA_signal_6630, SubBytesIns_Inst_Sbox_5_L1}), .c ({new_AGEMA_signal_6850, SubBytesIns_Inst_Sbox_5_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L16_U1 ( .a ({new_AGEMA_signal_6389, SubBytesIns_Inst_Sbox_5_M56}), .b ({new_AGEMA_signal_7034, SubBytesIns_Inst_Sbox_5_L0}), .c ({new_AGEMA_signal_7233, SubBytesIns_Inst_Sbox_5_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L17_U1 ( .a ({new_AGEMA_signal_6390, SubBytesIns_Inst_Sbox_5_M57}), .b ({new_AGEMA_signal_6630, SubBytesIns_Inst_Sbox_5_L1}), .c ({new_AGEMA_signal_6851, SubBytesIns_Inst_Sbox_5_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L18_U1 ( .a ({new_AGEMA_signal_6627, SubBytesIns_Inst_Sbox_5_M58}), .b ({new_AGEMA_signal_6631, SubBytesIns_Inst_Sbox_5_L8}), .c ({new_AGEMA_signal_6852, SubBytesIns_Inst_Sbox_5_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L19_U1 ( .a ({new_AGEMA_signal_6629, SubBytesIns_Inst_Sbox_5_M63}), .b ({new_AGEMA_signal_6847, SubBytesIns_Inst_Sbox_5_L4}), .c ({new_AGEMA_signal_7040, SubBytesIns_Inst_Sbox_5_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L20_U1 ( .a ({new_AGEMA_signal_7034, SubBytesIns_Inst_Sbox_5_L0}), .b ({new_AGEMA_signal_6630, SubBytesIns_Inst_Sbox_5_L1}), .c ({new_AGEMA_signal_7234, SubBytesIns_Inst_Sbox_5_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L21_U1 ( .a ({new_AGEMA_signal_6630, SubBytesIns_Inst_Sbox_5_L1}), .b ({new_AGEMA_signal_7036, SubBytesIns_Inst_Sbox_5_L7}), .c ({new_AGEMA_signal_7235, SubBytesIns_Inst_Sbox_5_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L22_U1 ( .a ({new_AGEMA_signal_6846, SubBytesIns_Inst_Sbox_5_L3}), .b ({new_AGEMA_signal_6632, SubBytesIns_Inst_Sbox_5_L12}), .c ({new_AGEMA_signal_7041, SubBytesIns_Inst_Sbox_5_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L23_U1 ( .a ({new_AGEMA_signal_6852, SubBytesIns_Inst_Sbox_5_L18}), .b ({new_AGEMA_signal_6845, SubBytesIns_Inst_Sbox_5_L2}), .c ({new_AGEMA_signal_7042, SubBytesIns_Inst_Sbox_5_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L24_U1 ( .a ({new_AGEMA_signal_6850, SubBytesIns_Inst_Sbox_5_L15}), .b ({new_AGEMA_signal_7037, SubBytesIns_Inst_Sbox_5_L9}), .c ({new_AGEMA_signal_7236, SubBytesIns_Inst_Sbox_5_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L25_U1 ( .a ({new_AGEMA_signal_7035, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_7038, SubBytesIns_Inst_Sbox_5_L10}), .c ({new_AGEMA_signal_7237, SubBytesIns_Inst_Sbox_5_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L26_U1 ( .a ({new_AGEMA_signal_7036, SubBytesIns_Inst_Sbox_5_L7}), .b ({new_AGEMA_signal_7037, SubBytesIns_Inst_Sbox_5_L9}), .c ({new_AGEMA_signal_7238, SubBytesIns_Inst_Sbox_5_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L27_U1 ( .a ({new_AGEMA_signal_6631, SubBytesIns_Inst_Sbox_5_L8}), .b ({new_AGEMA_signal_7038, SubBytesIns_Inst_Sbox_5_L10}), .c ({new_AGEMA_signal_7239, SubBytesIns_Inst_Sbox_5_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L28_U1 ( .a ({new_AGEMA_signal_7039, SubBytesIns_Inst_Sbox_5_L11}), .b ({new_AGEMA_signal_6849, SubBytesIns_Inst_Sbox_5_L14}), .c ({new_AGEMA_signal_7240, SubBytesIns_Inst_Sbox_5_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L29_U1 ( .a ({new_AGEMA_signal_7039, SubBytesIns_Inst_Sbox_5_L11}), .b ({new_AGEMA_signal_6851, SubBytesIns_Inst_Sbox_5_L17}), .c ({new_AGEMA_signal_7241, SubBytesIns_Inst_Sbox_5_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S0_U1 ( .a ({new_AGEMA_signal_7035, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_7236, SubBytesIns_Inst_Sbox_5_L24}), .c ({new_AGEMA_signal_7420, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S1_U1 ( .a ({new_AGEMA_signal_7233, SubBytesIns_Inst_Sbox_5_L16}), .b ({new_AGEMA_signal_7238, SubBytesIns_Inst_Sbox_5_L26}), .c ({new_AGEMA_signal_7421, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S2_U1 ( .a ({new_AGEMA_signal_7040, SubBytesIns_Inst_Sbox_5_L19}), .b ({new_AGEMA_signal_7240, SubBytesIns_Inst_Sbox_5_L28}), .c ({new_AGEMA_signal_7422, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S3_U1 ( .a ({new_AGEMA_signal_7035, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_7235, SubBytesIns_Inst_Sbox_5_L21}), .c ({new_AGEMA_signal_7423, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S4_U1 ( .a ({new_AGEMA_signal_7234, SubBytesIns_Inst_Sbox_5_L20}), .b ({new_AGEMA_signal_7041, SubBytesIns_Inst_Sbox_5_L22}), .c ({new_AGEMA_signal_7424, MixColumnsInput[107]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S5_U1 ( .a ({new_AGEMA_signal_7237, SubBytesIns_Inst_Sbox_5_L25}), .b ({new_AGEMA_signal_7241, SubBytesIns_Inst_Sbox_5_L29}), .c ({new_AGEMA_signal_7425, MixColumnsInput[106]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S6_U1 ( .a ({new_AGEMA_signal_7232, SubBytesIns_Inst_Sbox_5_L13}), .b ({new_AGEMA_signal_7239, SubBytesIns_Inst_Sbox_5_L27}), .c ({new_AGEMA_signal_7426, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S7_U1 ( .a ({new_AGEMA_signal_7035, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_7042, SubBytesIns_Inst_Sbox_5_L23}), .c ({new_AGEMA_signal_7242, MixColumnsInput[104]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M46_U1 ( .a ({new_AGEMA_signal_6396, SubBytesIns_Inst_Sbox_6_M44}), .b ({new_AGEMA_signal_5213, SubBytesIns_Inst_Sbox_6_T6}), .clk (clk), .r (Fresh[428]), .c ({new_AGEMA_signal_6634, SubBytesIns_Inst_Sbox_6_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M47_U1 ( .a ({new_AGEMA_signal_6236, SubBytesIns_Inst_Sbox_6_M40}), .b ({new_AGEMA_signal_5423, SubBytesIns_Inst_Sbox_6_T8}), .clk (clk), .r (Fresh[429]), .c ({new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_6_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M48_U1 ( .a ({new_AGEMA_signal_6235, SubBytesIns_Inst_Sbox_6_M39}), .b ({ciphertext_s1[48], ciphertext_s0[48]}), .clk (clk), .r (Fresh[430]), .c ({new_AGEMA_signal_6398, SubBytesIns_Inst_Sbox_6_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M49_U1 ( .a ({new_AGEMA_signal_6395, SubBytesIns_Inst_Sbox_6_M43}), .b ({new_AGEMA_signal_5217, SubBytesIns_Inst_Sbox_6_T16}), .clk (clk), .r (Fresh[431]), .c ({new_AGEMA_signal_6635, SubBytesIns_Inst_Sbox_6_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M50_U1 ( .a ({new_AGEMA_signal_6234, SubBytesIns_Inst_Sbox_6_M38}), .b ({new_AGEMA_signal_5214, SubBytesIns_Inst_Sbox_6_T9}), .clk (clk), .r (Fresh[432]), .c ({new_AGEMA_signal_6399, SubBytesIns_Inst_Sbox_6_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M51_U1 ( .a ({new_AGEMA_signal_6233, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_5426, SubBytesIns_Inst_Sbox_6_T17}), .clk (clk), .r (Fresh[433]), .c ({new_AGEMA_signal_6400, SubBytesIns_Inst_Sbox_6_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M52_U1 ( .a ({new_AGEMA_signal_6394, SubBytesIns_Inst_Sbox_6_M42}), .b ({new_AGEMA_signal_5216, SubBytesIns_Inst_Sbox_6_T15}), .clk (clk), .r (Fresh[434]), .c ({new_AGEMA_signal_6636, SubBytesIns_Inst_Sbox_6_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M53_U1 ( .a ({new_AGEMA_signal_6633, SubBytesIns_Inst_Sbox_6_M45}), .b ({new_AGEMA_signal_5220, SubBytesIns_Inst_Sbox_6_T27}), .clk (clk), .r (Fresh[435]), .c ({new_AGEMA_signal_6853, SubBytesIns_Inst_Sbox_6_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M54_U1 ( .a ({new_AGEMA_signal_6393, SubBytesIns_Inst_Sbox_6_M41}), .b ({new_AGEMA_signal_5424, SubBytesIns_Inst_Sbox_6_T10}), .clk (clk), .r (Fresh[436]), .c ({new_AGEMA_signal_6637, SubBytesIns_Inst_Sbox_6_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M55_U1 ( .a ({new_AGEMA_signal_6396, SubBytesIns_Inst_Sbox_6_M44}), .b ({new_AGEMA_signal_5215, SubBytesIns_Inst_Sbox_6_T13}), .clk (clk), .r (Fresh[437]), .c ({new_AGEMA_signal_6638, SubBytesIns_Inst_Sbox_6_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M56_U1 ( .a ({new_AGEMA_signal_6236, SubBytesIns_Inst_Sbox_6_M40}), .b ({new_AGEMA_signal_5428, SubBytesIns_Inst_Sbox_6_T23}), .clk (clk), .r (Fresh[438]), .c ({new_AGEMA_signal_6401, SubBytesIns_Inst_Sbox_6_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M57_U1 ( .a ({new_AGEMA_signal_6235, SubBytesIns_Inst_Sbox_6_M39}), .b ({new_AGEMA_signal_5218, SubBytesIns_Inst_Sbox_6_T19}), .clk (clk), .r (Fresh[439]), .c ({new_AGEMA_signal_6402, SubBytesIns_Inst_Sbox_6_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M58_U1 ( .a ({new_AGEMA_signal_6395, SubBytesIns_Inst_Sbox_6_M43}), .b ({new_AGEMA_signal_5035, SubBytesIns_Inst_Sbox_6_T3}), .clk (clk), .r (Fresh[440]), .c ({new_AGEMA_signal_6639, SubBytesIns_Inst_Sbox_6_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M59_U1 ( .a ({new_AGEMA_signal_6234, SubBytesIns_Inst_Sbox_6_M38}), .b ({new_AGEMA_signal_5219, SubBytesIns_Inst_Sbox_6_T22}), .clk (clk), .r (Fresh[441]), .c ({new_AGEMA_signal_6403, SubBytesIns_Inst_Sbox_6_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M60_U1 ( .a ({new_AGEMA_signal_6233, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_5427, SubBytesIns_Inst_Sbox_6_T20}), .clk (clk), .r (Fresh[442]), .c ({new_AGEMA_signal_6404, SubBytesIns_Inst_Sbox_6_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M61_U1 ( .a ({new_AGEMA_signal_6394, SubBytesIns_Inst_Sbox_6_M42}), .b ({new_AGEMA_signal_5033, SubBytesIns_Inst_Sbox_6_T1}), .clk (clk), .r (Fresh[443]), .c ({new_AGEMA_signal_6640, SubBytesIns_Inst_Sbox_6_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M62_U1 ( .a ({new_AGEMA_signal_6633, SubBytesIns_Inst_Sbox_6_M45}), .b ({new_AGEMA_signal_5036, SubBytesIns_Inst_Sbox_6_T4}), .clk (clk), .r (Fresh[444]), .c ({new_AGEMA_signal_6854, SubBytesIns_Inst_Sbox_6_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M63_U1 ( .a ({new_AGEMA_signal_6393, SubBytesIns_Inst_Sbox_6_M41}), .b ({new_AGEMA_signal_5034, SubBytesIns_Inst_Sbox_6_T2}), .clk (clk), .r (Fresh[445]), .c ({new_AGEMA_signal_6641, SubBytesIns_Inst_Sbox_6_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L0_U1 ( .a ({new_AGEMA_signal_6640, SubBytesIns_Inst_Sbox_6_M61}), .b ({new_AGEMA_signal_6854, SubBytesIns_Inst_Sbox_6_M62}), .c ({new_AGEMA_signal_7043, SubBytesIns_Inst_Sbox_6_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L1_U1 ( .a ({new_AGEMA_signal_6399, SubBytesIns_Inst_Sbox_6_M50}), .b ({new_AGEMA_signal_6401, SubBytesIns_Inst_Sbox_6_M56}), .c ({new_AGEMA_signal_6642, SubBytesIns_Inst_Sbox_6_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L2_U1 ( .a ({new_AGEMA_signal_6634, SubBytesIns_Inst_Sbox_6_M46}), .b ({new_AGEMA_signal_6398, SubBytesIns_Inst_Sbox_6_M48}), .c ({new_AGEMA_signal_6855, SubBytesIns_Inst_Sbox_6_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L3_U1 ( .a ({new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_6_M47}), .b ({new_AGEMA_signal_6638, SubBytesIns_Inst_Sbox_6_M55}), .c ({new_AGEMA_signal_6856, SubBytesIns_Inst_Sbox_6_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L4_U1 ( .a ({new_AGEMA_signal_6637, SubBytesIns_Inst_Sbox_6_M54}), .b ({new_AGEMA_signal_6639, SubBytesIns_Inst_Sbox_6_M58}), .c ({new_AGEMA_signal_6857, SubBytesIns_Inst_Sbox_6_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L5_U1 ( .a ({new_AGEMA_signal_6635, SubBytesIns_Inst_Sbox_6_M49}), .b ({new_AGEMA_signal_6640, SubBytesIns_Inst_Sbox_6_M61}), .c ({new_AGEMA_signal_6858, SubBytesIns_Inst_Sbox_6_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L6_U1 ( .a ({new_AGEMA_signal_6854, SubBytesIns_Inst_Sbox_6_M62}), .b ({new_AGEMA_signal_6858, SubBytesIns_Inst_Sbox_6_L5}), .c ({new_AGEMA_signal_7044, SubBytesIns_Inst_Sbox_6_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L7_U1 ( .a ({new_AGEMA_signal_6634, SubBytesIns_Inst_Sbox_6_M46}), .b ({new_AGEMA_signal_6856, SubBytesIns_Inst_Sbox_6_L3}), .c ({new_AGEMA_signal_7045, SubBytesIns_Inst_Sbox_6_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L8_U1 ( .a ({new_AGEMA_signal_6400, SubBytesIns_Inst_Sbox_6_M51}), .b ({new_AGEMA_signal_6403, SubBytesIns_Inst_Sbox_6_M59}), .c ({new_AGEMA_signal_6643, SubBytesIns_Inst_Sbox_6_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L9_U1 ( .a ({new_AGEMA_signal_6636, SubBytesIns_Inst_Sbox_6_M52}), .b ({new_AGEMA_signal_6853, SubBytesIns_Inst_Sbox_6_M53}), .c ({new_AGEMA_signal_7046, SubBytesIns_Inst_Sbox_6_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L10_U1 ( .a ({new_AGEMA_signal_6853, SubBytesIns_Inst_Sbox_6_M53}), .b ({new_AGEMA_signal_6857, SubBytesIns_Inst_Sbox_6_L4}), .c ({new_AGEMA_signal_7047, SubBytesIns_Inst_Sbox_6_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L11_U1 ( .a ({new_AGEMA_signal_6404, SubBytesIns_Inst_Sbox_6_M60}), .b ({new_AGEMA_signal_6855, SubBytesIns_Inst_Sbox_6_L2}), .c ({new_AGEMA_signal_7048, SubBytesIns_Inst_Sbox_6_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L12_U1 ( .a ({new_AGEMA_signal_6398, SubBytesIns_Inst_Sbox_6_M48}), .b ({new_AGEMA_signal_6400, SubBytesIns_Inst_Sbox_6_M51}), .c ({new_AGEMA_signal_6644, SubBytesIns_Inst_Sbox_6_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L13_U1 ( .a ({new_AGEMA_signal_6399, SubBytesIns_Inst_Sbox_6_M50}), .b ({new_AGEMA_signal_7043, SubBytesIns_Inst_Sbox_6_L0}), .c ({new_AGEMA_signal_7243, SubBytesIns_Inst_Sbox_6_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L14_U1 ( .a ({new_AGEMA_signal_6636, SubBytesIns_Inst_Sbox_6_M52}), .b ({new_AGEMA_signal_6640, SubBytesIns_Inst_Sbox_6_M61}), .c ({new_AGEMA_signal_6859, SubBytesIns_Inst_Sbox_6_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L15_U1 ( .a ({new_AGEMA_signal_6638, SubBytesIns_Inst_Sbox_6_M55}), .b ({new_AGEMA_signal_6642, SubBytesIns_Inst_Sbox_6_L1}), .c ({new_AGEMA_signal_6860, SubBytesIns_Inst_Sbox_6_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L16_U1 ( .a ({new_AGEMA_signal_6401, SubBytesIns_Inst_Sbox_6_M56}), .b ({new_AGEMA_signal_7043, SubBytesIns_Inst_Sbox_6_L0}), .c ({new_AGEMA_signal_7244, SubBytesIns_Inst_Sbox_6_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L17_U1 ( .a ({new_AGEMA_signal_6402, SubBytesIns_Inst_Sbox_6_M57}), .b ({new_AGEMA_signal_6642, SubBytesIns_Inst_Sbox_6_L1}), .c ({new_AGEMA_signal_6861, SubBytesIns_Inst_Sbox_6_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L18_U1 ( .a ({new_AGEMA_signal_6639, SubBytesIns_Inst_Sbox_6_M58}), .b ({new_AGEMA_signal_6643, SubBytesIns_Inst_Sbox_6_L8}), .c ({new_AGEMA_signal_6862, SubBytesIns_Inst_Sbox_6_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L19_U1 ( .a ({new_AGEMA_signal_6641, SubBytesIns_Inst_Sbox_6_M63}), .b ({new_AGEMA_signal_6857, SubBytesIns_Inst_Sbox_6_L4}), .c ({new_AGEMA_signal_7049, SubBytesIns_Inst_Sbox_6_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L20_U1 ( .a ({new_AGEMA_signal_7043, SubBytesIns_Inst_Sbox_6_L0}), .b ({new_AGEMA_signal_6642, SubBytesIns_Inst_Sbox_6_L1}), .c ({new_AGEMA_signal_7245, SubBytesIns_Inst_Sbox_6_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L21_U1 ( .a ({new_AGEMA_signal_6642, SubBytesIns_Inst_Sbox_6_L1}), .b ({new_AGEMA_signal_7045, SubBytesIns_Inst_Sbox_6_L7}), .c ({new_AGEMA_signal_7246, SubBytesIns_Inst_Sbox_6_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L22_U1 ( .a ({new_AGEMA_signal_6856, SubBytesIns_Inst_Sbox_6_L3}), .b ({new_AGEMA_signal_6644, SubBytesIns_Inst_Sbox_6_L12}), .c ({new_AGEMA_signal_7050, SubBytesIns_Inst_Sbox_6_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L23_U1 ( .a ({new_AGEMA_signal_6862, SubBytesIns_Inst_Sbox_6_L18}), .b ({new_AGEMA_signal_6855, SubBytesIns_Inst_Sbox_6_L2}), .c ({new_AGEMA_signal_7051, SubBytesIns_Inst_Sbox_6_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L24_U1 ( .a ({new_AGEMA_signal_6860, SubBytesIns_Inst_Sbox_6_L15}), .b ({new_AGEMA_signal_7046, SubBytesIns_Inst_Sbox_6_L9}), .c ({new_AGEMA_signal_7247, SubBytesIns_Inst_Sbox_6_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L25_U1 ( .a ({new_AGEMA_signal_7044, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_7047, SubBytesIns_Inst_Sbox_6_L10}), .c ({new_AGEMA_signal_7248, SubBytesIns_Inst_Sbox_6_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L26_U1 ( .a ({new_AGEMA_signal_7045, SubBytesIns_Inst_Sbox_6_L7}), .b ({new_AGEMA_signal_7046, SubBytesIns_Inst_Sbox_6_L9}), .c ({new_AGEMA_signal_7249, SubBytesIns_Inst_Sbox_6_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L27_U1 ( .a ({new_AGEMA_signal_6643, SubBytesIns_Inst_Sbox_6_L8}), .b ({new_AGEMA_signal_7047, SubBytesIns_Inst_Sbox_6_L10}), .c ({new_AGEMA_signal_7250, SubBytesIns_Inst_Sbox_6_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L28_U1 ( .a ({new_AGEMA_signal_7048, SubBytesIns_Inst_Sbox_6_L11}), .b ({new_AGEMA_signal_6859, SubBytesIns_Inst_Sbox_6_L14}), .c ({new_AGEMA_signal_7251, SubBytesIns_Inst_Sbox_6_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L29_U1 ( .a ({new_AGEMA_signal_7048, SubBytesIns_Inst_Sbox_6_L11}), .b ({new_AGEMA_signal_6861, SubBytesIns_Inst_Sbox_6_L17}), .c ({new_AGEMA_signal_7252, SubBytesIns_Inst_Sbox_6_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S0_U1 ( .a ({new_AGEMA_signal_7044, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_7247, SubBytesIns_Inst_Sbox_6_L24}), .c ({new_AGEMA_signal_7427, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S1_U1 ( .a ({new_AGEMA_signal_7244, SubBytesIns_Inst_Sbox_6_L16}), .b ({new_AGEMA_signal_7249, SubBytesIns_Inst_Sbox_6_L26}), .c ({new_AGEMA_signal_7428, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S2_U1 ( .a ({new_AGEMA_signal_7049, SubBytesIns_Inst_Sbox_6_L19}), .b ({new_AGEMA_signal_7251, SubBytesIns_Inst_Sbox_6_L28}), .c ({new_AGEMA_signal_7429, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S3_U1 ( .a ({new_AGEMA_signal_7044, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_7246, SubBytesIns_Inst_Sbox_6_L21}), .c ({new_AGEMA_signal_7430, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S4_U1 ( .a ({new_AGEMA_signal_7245, SubBytesIns_Inst_Sbox_6_L20}), .b ({new_AGEMA_signal_7050, SubBytesIns_Inst_Sbox_6_L22}), .c ({new_AGEMA_signal_7431, MixColumnsInput[83]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S5_U1 ( .a ({new_AGEMA_signal_7248, SubBytesIns_Inst_Sbox_6_L25}), .b ({new_AGEMA_signal_7252, SubBytesIns_Inst_Sbox_6_L29}), .c ({new_AGEMA_signal_7432, MixColumnsInput[82]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S6_U1 ( .a ({new_AGEMA_signal_7243, SubBytesIns_Inst_Sbox_6_L13}), .b ({new_AGEMA_signal_7250, SubBytesIns_Inst_Sbox_6_L27}), .c ({new_AGEMA_signal_7433, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S7_U1 ( .a ({new_AGEMA_signal_7044, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_7051, SubBytesIns_Inst_Sbox_6_L23}), .c ({new_AGEMA_signal_7253, MixColumnsInput[80]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M46_U1 ( .a ({new_AGEMA_signal_6408, SubBytesIns_Inst_Sbox_7_M44}), .b ({new_AGEMA_signal_5221, SubBytesIns_Inst_Sbox_7_T6}), .clk (clk), .r (Fresh[446]), .c ({new_AGEMA_signal_6646, SubBytesIns_Inst_Sbox_7_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M47_U1 ( .a ({new_AGEMA_signal_6240, SubBytesIns_Inst_Sbox_7_M40}), .b ({new_AGEMA_signal_5436, SubBytesIns_Inst_Sbox_7_T8}), .clk (clk), .r (Fresh[447]), .c ({new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_7_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M48_U1 ( .a ({new_AGEMA_signal_6239, SubBytesIns_Inst_Sbox_7_M39}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .clk (clk), .r (Fresh[448]), .c ({new_AGEMA_signal_6410, SubBytesIns_Inst_Sbox_7_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M49_U1 ( .a ({new_AGEMA_signal_6407, SubBytesIns_Inst_Sbox_7_M43}), .b ({new_AGEMA_signal_5225, SubBytesIns_Inst_Sbox_7_T16}), .clk (clk), .r (Fresh[449]), .c ({new_AGEMA_signal_6647, SubBytesIns_Inst_Sbox_7_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M50_U1 ( .a ({new_AGEMA_signal_6238, SubBytesIns_Inst_Sbox_7_M38}), .b ({new_AGEMA_signal_5222, SubBytesIns_Inst_Sbox_7_T9}), .clk (clk), .r (Fresh[450]), .c ({new_AGEMA_signal_6411, SubBytesIns_Inst_Sbox_7_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M51_U1 ( .a ({new_AGEMA_signal_6237, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_5439, SubBytesIns_Inst_Sbox_7_T17}), .clk (clk), .r (Fresh[451]), .c ({new_AGEMA_signal_6412, SubBytesIns_Inst_Sbox_7_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M52_U1 ( .a ({new_AGEMA_signal_6406, SubBytesIns_Inst_Sbox_7_M42}), .b ({new_AGEMA_signal_5224, SubBytesIns_Inst_Sbox_7_T15}), .clk (clk), .r (Fresh[452]), .c ({new_AGEMA_signal_6648, SubBytesIns_Inst_Sbox_7_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M53_U1 ( .a ({new_AGEMA_signal_6645, SubBytesIns_Inst_Sbox_7_M45}), .b ({new_AGEMA_signal_5228, SubBytesIns_Inst_Sbox_7_T27}), .clk (clk), .r (Fresh[453]), .c ({new_AGEMA_signal_6863, SubBytesIns_Inst_Sbox_7_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M54_U1 ( .a ({new_AGEMA_signal_6405, SubBytesIns_Inst_Sbox_7_M41}), .b ({new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_7_T10}), .clk (clk), .r (Fresh[454]), .c ({new_AGEMA_signal_6649, SubBytesIns_Inst_Sbox_7_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M55_U1 ( .a ({new_AGEMA_signal_6408, SubBytesIns_Inst_Sbox_7_M44}), .b ({new_AGEMA_signal_5223, SubBytesIns_Inst_Sbox_7_T13}), .clk (clk), .r (Fresh[455]), .c ({new_AGEMA_signal_6650, SubBytesIns_Inst_Sbox_7_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M56_U1 ( .a ({new_AGEMA_signal_6240, SubBytesIns_Inst_Sbox_7_M40}), .b ({new_AGEMA_signal_5441, SubBytesIns_Inst_Sbox_7_T23}), .clk (clk), .r (Fresh[456]), .c ({new_AGEMA_signal_6413, SubBytesIns_Inst_Sbox_7_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M57_U1 ( .a ({new_AGEMA_signal_6239, SubBytesIns_Inst_Sbox_7_M39}), .b ({new_AGEMA_signal_5226, SubBytesIns_Inst_Sbox_7_T19}), .clk (clk), .r (Fresh[457]), .c ({new_AGEMA_signal_6414, SubBytesIns_Inst_Sbox_7_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M58_U1 ( .a ({new_AGEMA_signal_6407, SubBytesIns_Inst_Sbox_7_M43}), .b ({new_AGEMA_signal_5045, SubBytesIns_Inst_Sbox_7_T3}), .clk (clk), .r (Fresh[458]), .c ({new_AGEMA_signal_6651, SubBytesIns_Inst_Sbox_7_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M59_U1 ( .a ({new_AGEMA_signal_6238, SubBytesIns_Inst_Sbox_7_M38}), .b ({new_AGEMA_signal_5227, SubBytesIns_Inst_Sbox_7_T22}), .clk (clk), .r (Fresh[459]), .c ({new_AGEMA_signal_6415, SubBytesIns_Inst_Sbox_7_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M60_U1 ( .a ({new_AGEMA_signal_6237, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_5440, SubBytesIns_Inst_Sbox_7_T20}), .clk (clk), .r (Fresh[460]), .c ({new_AGEMA_signal_6416, SubBytesIns_Inst_Sbox_7_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M61_U1 ( .a ({new_AGEMA_signal_6406, SubBytesIns_Inst_Sbox_7_M42}), .b ({new_AGEMA_signal_5043, SubBytesIns_Inst_Sbox_7_T1}), .clk (clk), .r (Fresh[461]), .c ({new_AGEMA_signal_6652, SubBytesIns_Inst_Sbox_7_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M62_U1 ( .a ({new_AGEMA_signal_6645, SubBytesIns_Inst_Sbox_7_M45}), .b ({new_AGEMA_signal_5046, SubBytesIns_Inst_Sbox_7_T4}), .clk (clk), .r (Fresh[462]), .c ({new_AGEMA_signal_6864, SubBytesIns_Inst_Sbox_7_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M63_U1 ( .a ({new_AGEMA_signal_6405, SubBytesIns_Inst_Sbox_7_M41}), .b ({new_AGEMA_signal_5044, SubBytesIns_Inst_Sbox_7_T2}), .clk (clk), .r (Fresh[463]), .c ({new_AGEMA_signal_6653, SubBytesIns_Inst_Sbox_7_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L0_U1 ( .a ({new_AGEMA_signal_6652, SubBytesIns_Inst_Sbox_7_M61}), .b ({new_AGEMA_signal_6864, SubBytesIns_Inst_Sbox_7_M62}), .c ({new_AGEMA_signal_7052, SubBytesIns_Inst_Sbox_7_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L1_U1 ( .a ({new_AGEMA_signal_6411, SubBytesIns_Inst_Sbox_7_M50}), .b ({new_AGEMA_signal_6413, SubBytesIns_Inst_Sbox_7_M56}), .c ({new_AGEMA_signal_6654, SubBytesIns_Inst_Sbox_7_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L2_U1 ( .a ({new_AGEMA_signal_6646, SubBytesIns_Inst_Sbox_7_M46}), .b ({new_AGEMA_signal_6410, SubBytesIns_Inst_Sbox_7_M48}), .c ({new_AGEMA_signal_6865, SubBytesIns_Inst_Sbox_7_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L3_U1 ( .a ({new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_7_M47}), .b ({new_AGEMA_signal_6650, SubBytesIns_Inst_Sbox_7_M55}), .c ({new_AGEMA_signal_6866, SubBytesIns_Inst_Sbox_7_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L4_U1 ( .a ({new_AGEMA_signal_6649, SubBytesIns_Inst_Sbox_7_M54}), .b ({new_AGEMA_signal_6651, SubBytesIns_Inst_Sbox_7_M58}), .c ({new_AGEMA_signal_6867, SubBytesIns_Inst_Sbox_7_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L5_U1 ( .a ({new_AGEMA_signal_6647, SubBytesIns_Inst_Sbox_7_M49}), .b ({new_AGEMA_signal_6652, SubBytesIns_Inst_Sbox_7_M61}), .c ({new_AGEMA_signal_6868, SubBytesIns_Inst_Sbox_7_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L6_U1 ( .a ({new_AGEMA_signal_6864, SubBytesIns_Inst_Sbox_7_M62}), .b ({new_AGEMA_signal_6868, SubBytesIns_Inst_Sbox_7_L5}), .c ({new_AGEMA_signal_7053, SubBytesIns_Inst_Sbox_7_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L7_U1 ( .a ({new_AGEMA_signal_6646, SubBytesIns_Inst_Sbox_7_M46}), .b ({new_AGEMA_signal_6866, SubBytesIns_Inst_Sbox_7_L3}), .c ({new_AGEMA_signal_7054, SubBytesIns_Inst_Sbox_7_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L8_U1 ( .a ({new_AGEMA_signal_6412, SubBytesIns_Inst_Sbox_7_M51}), .b ({new_AGEMA_signal_6415, SubBytesIns_Inst_Sbox_7_M59}), .c ({new_AGEMA_signal_6655, SubBytesIns_Inst_Sbox_7_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L9_U1 ( .a ({new_AGEMA_signal_6648, SubBytesIns_Inst_Sbox_7_M52}), .b ({new_AGEMA_signal_6863, SubBytesIns_Inst_Sbox_7_M53}), .c ({new_AGEMA_signal_7055, SubBytesIns_Inst_Sbox_7_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L10_U1 ( .a ({new_AGEMA_signal_6863, SubBytesIns_Inst_Sbox_7_M53}), .b ({new_AGEMA_signal_6867, SubBytesIns_Inst_Sbox_7_L4}), .c ({new_AGEMA_signal_7056, SubBytesIns_Inst_Sbox_7_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L11_U1 ( .a ({new_AGEMA_signal_6416, SubBytesIns_Inst_Sbox_7_M60}), .b ({new_AGEMA_signal_6865, SubBytesIns_Inst_Sbox_7_L2}), .c ({new_AGEMA_signal_7057, SubBytesIns_Inst_Sbox_7_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L12_U1 ( .a ({new_AGEMA_signal_6410, SubBytesIns_Inst_Sbox_7_M48}), .b ({new_AGEMA_signal_6412, SubBytesIns_Inst_Sbox_7_M51}), .c ({new_AGEMA_signal_6656, SubBytesIns_Inst_Sbox_7_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L13_U1 ( .a ({new_AGEMA_signal_6411, SubBytesIns_Inst_Sbox_7_M50}), .b ({new_AGEMA_signal_7052, SubBytesIns_Inst_Sbox_7_L0}), .c ({new_AGEMA_signal_7254, SubBytesIns_Inst_Sbox_7_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L14_U1 ( .a ({new_AGEMA_signal_6648, SubBytesIns_Inst_Sbox_7_M52}), .b ({new_AGEMA_signal_6652, SubBytesIns_Inst_Sbox_7_M61}), .c ({new_AGEMA_signal_6869, SubBytesIns_Inst_Sbox_7_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L15_U1 ( .a ({new_AGEMA_signal_6650, SubBytesIns_Inst_Sbox_7_M55}), .b ({new_AGEMA_signal_6654, SubBytesIns_Inst_Sbox_7_L1}), .c ({new_AGEMA_signal_6870, SubBytesIns_Inst_Sbox_7_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L16_U1 ( .a ({new_AGEMA_signal_6413, SubBytesIns_Inst_Sbox_7_M56}), .b ({new_AGEMA_signal_7052, SubBytesIns_Inst_Sbox_7_L0}), .c ({new_AGEMA_signal_7255, SubBytesIns_Inst_Sbox_7_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L17_U1 ( .a ({new_AGEMA_signal_6414, SubBytesIns_Inst_Sbox_7_M57}), .b ({new_AGEMA_signal_6654, SubBytesIns_Inst_Sbox_7_L1}), .c ({new_AGEMA_signal_6871, SubBytesIns_Inst_Sbox_7_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L18_U1 ( .a ({new_AGEMA_signal_6651, SubBytesIns_Inst_Sbox_7_M58}), .b ({new_AGEMA_signal_6655, SubBytesIns_Inst_Sbox_7_L8}), .c ({new_AGEMA_signal_6872, SubBytesIns_Inst_Sbox_7_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L19_U1 ( .a ({new_AGEMA_signal_6653, SubBytesIns_Inst_Sbox_7_M63}), .b ({new_AGEMA_signal_6867, SubBytesIns_Inst_Sbox_7_L4}), .c ({new_AGEMA_signal_7058, SubBytesIns_Inst_Sbox_7_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L20_U1 ( .a ({new_AGEMA_signal_7052, SubBytesIns_Inst_Sbox_7_L0}), .b ({new_AGEMA_signal_6654, SubBytesIns_Inst_Sbox_7_L1}), .c ({new_AGEMA_signal_7256, SubBytesIns_Inst_Sbox_7_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L21_U1 ( .a ({new_AGEMA_signal_6654, SubBytesIns_Inst_Sbox_7_L1}), .b ({new_AGEMA_signal_7054, SubBytesIns_Inst_Sbox_7_L7}), .c ({new_AGEMA_signal_7257, SubBytesIns_Inst_Sbox_7_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L22_U1 ( .a ({new_AGEMA_signal_6866, SubBytesIns_Inst_Sbox_7_L3}), .b ({new_AGEMA_signal_6656, SubBytesIns_Inst_Sbox_7_L12}), .c ({new_AGEMA_signal_7059, SubBytesIns_Inst_Sbox_7_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L23_U1 ( .a ({new_AGEMA_signal_6872, SubBytesIns_Inst_Sbox_7_L18}), .b ({new_AGEMA_signal_6865, SubBytesIns_Inst_Sbox_7_L2}), .c ({new_AGEMA_signal_7060, SubBytesIns_Inst_Sbox_7_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L24_U1 ( .a ({new_AGEMA_signal_6870, SubBytesIns_Inst_Sbox_7_L15}), .b ({new_AGEMA_signal_7055, SubBytesIns_Inst_Sbox_7_L9}), .c ({new_AGEMA_signal_7258, SubBytesIns_Inst_Sbox_7_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L25_U1 ( .a ({new_AGEMA_signal_7053, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_7056, SubBytesIns_Inst_Sbox_7_L10}), .c ({new_AGEMA_signal_7259, SubBytesIns_Inst_Sbox_7_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L26_U1 ( .a ({new_AGEMA_signal_7054, SubBytesIns_Inst_Sbox_7_L7}), .b ({new_AGEMA_signal_7055, SubBytesIns_Inst_Sbox_7_L9}), .c ({new_AGEMA_signal_7260, SubBytesIns_Inst_Sbox_7_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L27_U1 ( .a ({new_AGEMA_signal_6655, SubBytesIns_Inst_Sbox_7_L8}), .b ({new_AGEMA_signal_7056, SubBytesIns_Inst_Sbox_7_L10}), .c ({new_AGEMA_signal_7261, SubBytesIns_Inst_Sbox_7_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L28_U1 ( .a ({new_AGEMA_signal_7057, SubBytesIns_Inst_Sbox_7_L11}), .b ({new_AGEMA_signal_6869, SubBytesIns_Inst_Sbox_7_L14}), .c ({new_AGEMA_signal_7262, SubBytesIns_Inst_Sbox_7_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L29_U1 ( .a ({new_AGEMA_signal_7057, SubBytesIns_Inst_Sbox_7_L11}), .b ({new_AGEMA_signal_6871, SubBytesIns_Inst_Sbox_7_L17}), .c ({new_AGEMA_signal_7263, SubBytesIns_Inst_Sbox_7_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S0_U1 ( .a ({new_AGEMA_signal_7053, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_7258, SubBytesIns_Inst_Sbox_7_L24}), .c ({new_AGEMA_signal_7434, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S1_U1 ( .a ({new_AGEMA_signal_7255, SubBytesIns_Inst_Sbox_7_L16}), .b ({new_AGEMA_signal_7260, SubBytesIns_Inst_Sbox_7_L26}), .c ({new_AGEMA_signal_7435, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S2_U1 ( .a ({new_AGEMA_signal_7058, SubBytesIns_Inst_Sbox_7_L19}), .b ({new_AGEMA_signal_7262, SubBytesIns_Inst_Sbox_7_L28}), .c ({new_AGEMA_signal_7436, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S3_U1 ( .a ({new_AGEMA_signal_7053, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_7257, SubBytesIns_Inst_Sbox_7_L21}), .c ({new_AGEMA_signal_7437, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S4_U1 ( .a ({new_AGEMA_signal_7256, SubBytesIns_Inst_Sbox_7_L20}), .b ({new_AGEMA_signal_7059, SubBytesIns_Inst_Sbox_7_L22}), .c ({new_AGEMA_signal_7438, MixColumnsInput[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S5_U1 ( .a ({new_AGEMA_signal_7259, SubBytesIns_Inst_Sbox_7_L25}), .b ({new_AGEMA_signal_7263, SubBytesIns_Inst_Sbox_7_L29}), .c ({new_AGEMA_signal_7439, MixColumnsInput[58]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S6_U1 ( .a ({new_AGEMA_signal_7254, SubBytesIns_Inst_Sbox_7_L13}), .b ({new_AGEMA_signal_7261, SubBytesIns_Inst_Sbox_7_L27}), .c ({new_AGEMA_signal_7440, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S7_U1 ( .a ({new_AGEMA_signal_7053, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_7060, SubBytesIns_Inst_Sbox_7_L23}), .c ({new_AGEMA_signal_7264, MixColumnsInput[56]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M46_U1 ( .a ({new_AGEMA_signal_6420, SubBytesIns_Inst_Sbox_8_M44}), .b ({new_AGEMA_signal_5229, SubBytesIns_Inst_Sbox_8_T6}), .clk (clk), .r (Fresh[464]), .c ({new_AGEMA_signal_6658, SubBytesIns_Inst_Sbox_8_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M47_U1 ( .a ({new_AGEMA_signal_6244, SubBytesIns_Inst_Sbox_8_M40}), .b ({new_AGEMA_signal_5449, SubBytesIns_Inst_Sbox_8_T8}), .clk (clk), .r (Fresh[465]), .c ({new_AGEMA_signal_6421, SubBytesIns_Inst_Sbox_8_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M48_U1 ( .a ({new_AGEMA_signal_6243, SubBytesIns_Inst_Sbox_8_M39}), .b ({ciphertext_s1[64], ciphertext_s0[64]}), .clk (clk), .r (Fresh[466]), .c ({new_AGEMA_signal_6422, SubBytesIns_Inst_Sbox_8_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M49_U1 ( .a ({new_AGEMA_signal_6419, SubBytesIns_Inst_Sbox_8_M43}), .b ({new_AGEMA_signal_5233, SubBytesIns_Inst_Sbox_8_T16}), .clk (clk), .r (Fresh[467]), .c ({new_AGEMA_signal_6659, SubBytesIns_Inst_Sbox_8_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M50_U1 ( .a ({new_AGEMA_signal_6242, SubBytesIns_Inst_Sbox_8_M38}), .b ({new_AGEMA_signal_5230, SubBytesIns_Inst_Sbox_8_T9}), .clk (clk), .r (Fresh[468]), .c ({new_AGEMA_signal_6423, SubBytesIns_Inst_Sbox_8_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M51_U1 ( .a ({new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_5452, SubBytesIns_Inst_Sbox_8_T17}), .clk (clk), .r (Fresh[469]), .c ({new_AGEMA_signal_6424, SubBytesIns_Inst_Sbox_8_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M52_U1 ( .a ({new_AGEMA_signal_6418, SubBytesIns_Inst_Sbox_8_M42}), .b ({new_AGEMA_signal_5232, SubBytesIns_Inst_Sbox_8_T15}), .clk (clk), .r (Fresh[470]), .c ({new_AGEMA_signal_6660, SubBytesIns_Inst_Sbox_8_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M53_U1 ( .a ({new_AGEMA_signal_6657, SubBytesIns_Inst_Sbox_8_M45}), .b ({new_AGEMA_signal_5236, SubBytesIns_Inst_Sbox_8_T27}), .clk (clk), .r (Fresh[471]), .c ({new_AGEMA_signal_6873, SubBytesIns_Inst_Sbox_8_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M54_U1 ( .a ({new_AGEMA_signal_6417, SubBytesIns_Inst_Sbox_8_M41}), .b ({new_AGEMA_signal_5450, SubBytesIns_Inst_Sbox_8_T10}), .clk (clk), .r (Fresh[472]), .c ({new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_8_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M55_U1 ( .a ({new_AGEMA_signal_6420, SubBytesIns_Inst_Sbox_8_M44}), .b ({new_AGEMA_signal_5231, SubBytesIns_Inst_Sbox_8_T13}), .clk (clk), .r (Fresh[473]), .c ({new_AGEMA_signal_6662, SubBytesIns_Inst_Sbox_8_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M56_U1 ( .a ({new_AGEMA_signal_6244, SubBytesIns_Inst_Sbox_8_M40}), .b ({new_AGEMA_signal_5454, SubBytesIns_Inst_Sbox_8_T23}), .clk (clk), .r (Fresh[474]), .c ({new_AGEMA_signal_6425, SubBytesIns_Inst_Sbox_8_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M57_U1 ( .a ({new_AGEMA_signal_6243, SubBytesIns_Inst_Sbox_8_M39}), .b ({new_AGEMA_signal_5234, SubBytesIns_Inst_Sbox_8_T19}), .clk (clk), .r (Fresh[475]), .c ({new_AGEMA_signal_6426, SubBytesIns_Inst_Sbox_8_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M58_U1 ( .a ({new_AGEMA_signal_6419, SubBytesIns_Inst_Sbox_8_M43}), .b ({new_AGEMA_signal_5055, SubBytesIns_Inst_Sbox_8_T3}), .clk (clk), .r (Fresh[476]), .c ({new_AGEMA_signal_6663, SubBytesIns_Inst_Sbox_8_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M59_U1 ( .a ({new_AGEMA_signal_6242, SubBytesIns_Inst_Sbox_8_M38}), .b ({new_AGEMA_signal_5235, SubBytesIns_Inst_Sbox_8_T22}), .clk (clk), .r (Fresh[477]), .c ({new_AGEMA_signal_6427, SubBytesIns_Inst_Sbox_8_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M60_U1 ( .a ({new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_5453, SubBytesIns_Inst_Sbox_8_T20}), .clk (clk), .r (Fresh[478]), .c ({new_AGEMA_signal_6428, SubBytesIns_Inst_Sbox_8_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M61_U1 ( .a ({new_AGEMA_signal_6418, SubBytesIns_Inst_Sbox_8_M42}), .b ({new_AGEMA_signal_5053, SubBytesIns_Inst_Sbox_8_T1}), .clk (clk), .r (Fresh[479]), .c ({new_AGEMA_signal_6664, SubBytesIns_Inst_Sbox_8_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M62_U1 ( .a ({new_AGEMA_signal_6657, SubBytesIns_Inst_Sbox_8_M45}), .b ({new_AGEMA_signal_5056, SubBytesIns_Inst_Sbox_8_T4}), .clk (clk), .r (Fresh[480]), .c ({new_AGEMA_signal_6874, SubBytesIns_Inst_Sbox_8_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M63_U1 ( .a ({new_AGEMA_signal_6417, SubBytesIns_Inst_Sbox_8_M41}), .b ({new_AGEMA_signal_5054, SubBytesIns_Inst_Sbox_8_T2}), .clk (clk), .r (Fresh[481]), .c ({new_AGEMA_signal_6665, SubBytesIns_Inst_Sbox_8_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L0_U1 ( .a ({new_AGEMA_signal_6664, SubBytesIns_Inst_Sbox_8_M61}), .b ({new_AGEMA_signal_6874, SubBytesIns_Inst_Sbox_8_M62}), .c ({new_AGEMA_signal_7061, SubBytesIns_Inst_Sbox_8_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L1_U1 ( .a ({new_AGEMA_signal_6423, SubBytesIns_Inst_Sbox_8_M50}), .b ({new_AGEMA_signal_6425, SubBytesIns_Inst_Sbox_8_M56}), .c ({new_AGEMA_signal_6666, SubBytesIns_Inst_Sbox_8_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L2_U1 ( .a ({new_AGEMA_signal_6658, SubBytesIns_Inst_Sbox_8_M46}), .b ({new_AGEMA_signal_6422, SubBytesIns_Inst_Sbox_8_M48}), .c ({new_AGEMA_signal_6875, SubBytesIns_Inst_Sbox_8_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L3_U1 ( .a ({new_AGEMA_signal_6421, SubBytesIns_Inst_Sbox_8_M47}), .b ({new_AGEMA_signal_6662, SubBytesIns_Inst_Sbox_8_M55}), .c ({new_AGEMA_signal_6876, SubBytesIns_Inst_Sbox_8_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L4_U1 ( .a ({new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_8_M54}), .b ({new_AGEMA_signal_6663, SubBytesIns_Inst_Sbox_8_M58}), .c ({new_AGEMA_signal_6877, SubBytesIns_Inst_Sbox_8_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L5_U1 ( .a ({new_AGEMA_signal_6659, SubBytesIns_Inst_Sbox_8_M49}), .b ({new_AGEMA_signal_6664, SubBytesIns_Inst_Sbox_8_M61}), .c ({new_AGEMA_signal_6878, SubBytesIns_Inst_Sbox_8_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L6_U1 ( .a ({new_AGEMA_signal_6874, SubBytesIns_Inst_Sbox_8_M62}), .b ({new_AGEMA_signal_6878, SubBytesIns_Inst_Sbox_8_L5}), .c ({new_AGEMA_signal_7062, SubBytesIns_Inst_Sbox_8_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L7_U1 ( .a ({new_AGEMA_signal_6658, SubBytesIns_Inst_Sbox_8_M46}), .b ({new_AGEMA_signal_6876, SubBytesIns_Inst_Sbox_8_L3}), .c ({new_AGEMA_signal_7063, SubBytesIns_Inst_Sbox_8_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L8_U1 ( .a ({new_AGEMA_signal_6424, SubBytesIns_Inst_Sbox_8_M51}), .b ({new_AGEMA_signal_6427, SubBytesIns_Inst_Sbox_8_M59}), .c ({new_AGEMA_signal_6667, SubBytesIns_Inst_Sbox_8_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L9_U1 ( .a ({new_AGEMA_signal_6660, SubBytesIns_Inst_Sbox_8_M52}), .b ({new_AGEMA_signal_6873, SubBytesIns_Inst_Sbox_8_M53}), .c ({new_AGEMA_signal_7064, SubBytesIns_Inst_Sbox_8_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L10_U1 ( .a ({new_AGEMA_signal_6873, SubBytesIns_Inst_Sbox_8_M53}), .b ({new_AGEMA_signal_6877, SubBytesIns_Inst_Sbox_8_L4}), .c ({new_AGEMA_signal_7065, SubBytesIns_Inst_Sbox_8_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L11_U1 ( .a ({new_AGEMA_signal_6428, SubBytesIns_Inst_Sbox_8_M60}), .b ({new_AGEMA_signal_6875, SubBytesIns_Inst_Sbox_8_L2}), .c ({new_AGEMA_signal_7066, SubBytesIns_Inst_Sbox_8_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L12_U1 ( .a ({new_AGEMA_signal_6422, SubBytesIns_Inst_Sbox_8_M48}), .b ({new_AGEMA_signal_6424, SubBytesIns_Inst_Sbox_8_M51}), .c ({new_AGEMA_signal_6668, SubBytesIns_Inst_Sbox_8_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L13_U1 ( .a ({new_AGEMA_signal_6423, SubBytesIns_Inst_Sbox_8_M50}), .b ({new_AGEMA_signal_7061, SubBytesIns_Inst_Sbox_8_L0}), .c ({new_AGEMA_signal_7265, SubBytesIns_Inst_Sbox_8_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L14_U1 ( .a ({new_AGEMA_signal_6660, SubBytesIns_Inst_Sbox_8_M52}), .b ({new_AGEMA_signal_6664, SubBytesIns_Inst_Sbox_8_M61}), .c ({new_AGEMA_signal_6879, SubBytesIns_Inst_Sbox_8_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L15_U1 ( .a ({new_AGEMA_signal_6662, SubBytesIns_Inst_Sbox_8_M55}), .b ({new_AGEMA_signal_6666, SubBytesIns_Inst_Sbox_8_L1}), .c ({new_AGEMA_signal_6880, SubBytesIns_Inst_Sbox_8_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L16_U1 ( .a ({new_AGEMA_signal_6425, SubBytesIns_Inst_Sbox_8_M56}), .b ({new_AGEMA_signal_7061, SubBytesIns_Inst_Sbox_8_L0}), .c ({new_AGEMA_signal_7266, SubBytesIns_Inst_Sbox_8_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L17_U1 ( .a ({new_AGEMA_signal_6426, SubBytesIns_Inst_Sbox_8_M57}), .b ({new_AGEMA_signal_6666, SubBytesIns_Inst_Sbox_8_L1}), .c ({new_AGEMA_signal_6881, SubBytesIns_Inst_Sbox_8_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L18_U1 ( .a ({new_AGEMA_signal_6663, SubBytesIns_Inst_Sbox_8_M58}), .b ({new_AGEMA_signal_6667, SubBytesIns_Inst_Sbox_8_L8}), .c ({new_AGEMA_signal_6882, SubBytesIns_Inst_Sbox_8_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L19_U1 ( .a ({new_AGEMA_signal_6665, SubBytesIns_Inst_Sbox_8_M63}), .b ({new_AGEMA_signal_6877, SubBytesIns_Inst_Sbox_8_L4}), .c ({new_AGEMA_signal_7067, SubBytesIns_Inst_Sbox_8_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L20_U1 ( .a ({new_AGEMA_signal_7061, SubBytesIns_Inst_Sbox_8_L0}), .b ({new_AGEMA_signal_6666, SubBytesIns_Inst_Sbox_8_L1}), .c ({new_AGEMA_signal_7267, SubBytesIns_Inst_Sbox_8_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L21_U1 ( .a ({new_AGEMA_signal_6666, SubBytesIns_Inst_Sbox_8_L1}), .b ({new_AGEMA_signal_7063, SubBytesIns_Inst_Sbox_8_L7}), .c ({new_AGEMA_signal_7268, SubBytesIns_Inst_Sbox_8_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L22_U1 ( .a ({new_AGEMA_signal_6876, SubBytesIns_Inst_Sbox_8_L3}), .b ({new_AGEMA_signal_6668, SubBytesIns_Inst_Sbox_8_L12}), .c ({new_AGEMA_signal_7068, SubBytesIns_Inst_Sbox_8_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L23_U1 ( .a ({new_AGEMA_signal_6882, SubBytesIns_Inst_Sbox_8_L18}), .b ({new_AGEMA_signal_6875, SubBytesIns_Inst_Sbox_8_L2}), .c ({new_AGEMA_signal_7069, SubBytesIns_Inst_Sbox_8_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L24_U1 ( .a ({new_AGEMA_signal_6880, SubBytesIns_Inst_Sbox_8_L15}), .b ({new_AGEMA_signal_7064, SubBytesIns_Inst_Sbox_8_L9}), .c ({new_AGEMA_signal_7269, SubBytesIns_Inst_Sbox_8_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L25_U1 ( .a ({new_AGEMA_signal_7062, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_7065, SubBytesIns_Inst_Sbox_8_L10}), .c ({new_AGEMA_signal_7270, SubBytesIns_Inst_Sbox_8_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L26_U1 ( .a ({new_AGEMA_signal_7063, SubBytesIns_Inst_Sbox_8_L7}), .b ({new_AGEMA_signal_7064, SubBytesIns_Inst_Sbox_8_L9}), .c ({new_AGEMA_signal_7271, SubBytesIns_Inst_Sbox_8_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L27_U1 ( .a ({new_AGEMA_signal_6667, SubBytesIns_Inst_Sbox_8_L8}), .b ({new_AGEMA_signal_7065, SubBytesIns_Inst_Sbox_8_L10}), .c ({new_AGEMA_signal_7272, SubBytesIns_Inst_Sbox_8_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L28_U1 ( .a ({new_AGEMA_signal_7066, SubBytesIns_Inst_Sbox_8_L11}), .b ({new_AGEMA_signal_6879, SubBytesIns_Inst_Sbox_8_L14}), .c ({new_AGEMA_signal_7273, SubBytesIns_Inst_Sbox_8_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L29_U1 ( .a ({new_AGEMA_signal_7066, SubBytesIns_Inst_Sbox_8_L11}), .b ({new_AGEMA_signal_6881, SubBytesIns_Inst_Sbox_8_L17}), .c ({new_AGEMA_signal_7274, SubBytesIns_Inst_Sbox_8_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S0_U1 ( .a ({new_AGEMA_signal_7062, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_7269, SubBytesIns_Inst_Sbox_8_L24}), .c ({new_AGEMA_signal_7441, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S1_U1 ( .a ({new_AGEMA_signal_7266, SubBytesIns_Inst_Sbox_8_L16}), .b ({new_AGEMA_signal_7271, SubBytesIns_Inst_Sbox_8_L26}), .c ({new_AGEMA_signal_7442, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S2_U1 ( .a ({new_AGEMA_signal_7067, SubBytesIns_Inst_Sbox_8_L19}), .b ({new_AGEMA_signal_7273, SubBytesIns_Inst_Sbox_8_L28}), .c ({new_AGEMA_signal_7443, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S3_U1 ( .a ({new_AGEMA_signal_7062, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_7268, SubBytesIns_Inst_Sbox_8_L21}), .c ({new_AGEMA_signal_7444, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S4_U1 ( .a ({new_AGEMA_signal_7267, SubBytesIns_Inst_Sbox_8_L20}), .b ({new_AGEMA_signal_7068, SubBytesIns_Inst_Sbox_8_L22}), .c ({new_AGEMA_signal_7445, MixColumnsInput[35]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S5_U1 ( .a ({new_AGEMA_signal_7270, SubBytesIns_Inst_Sbox_8_L25}), .b ({new_AGEMA_signal_7274, SubBytesIns_Inst_Sbox_8_L29}), .c ({new_AGEMA_signal_7446, MixColumnsInput[34]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S6_U1 ( .a ({new_AGEMA_signal_7265, SubBytesIns_Inst_Sbox_8_L13}), .b ({new_AGEMA_signal_7272, SubBytesIns_Inst_Sbox_8_L27}), .c ({new_AGEMA_signal_7447, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S7_U1 ( .a ({new_AGEMA_signal_7062, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_7069, SubBytesIns_Inst_Sbox_8_L23}), .c ({new_AGEMA_signal_7275, MixColumnsInput[32]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M46_U1 ( .a ({new_AGEMA_signal_6432, SubBytesIns_Inst_Sbox_9_M44}), .b ({new_AGEMA_signal_5237, SubBytesIns_Inst_Sbox_9_T6}), .clk (clk), .r (Fresh[482]), .c ({new_AGEMA_signal_6670, SubBytesIns_Inst_Sbox_9_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M47_U1 ( .a ({new_AGEMA_signal_6248, SubBytesIns_Inst_Sbox_9_M40}), .b ({new_AGEMA_signal_5462, SubBytesIns_Inst_Sbox_9_T8}), .clk (clk), .r (Fresh[483]), .c ({new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_9_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M48_U1 ( .a ({new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_9_M39}), .b ({ciphertext_s1[72], ciphertext_s0[72]}), .clk (clk), .r (Fresh[484]), .c ({new_AGEMA_signal_6434, SubBytesIns_Inst_Sbox_9_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M49_U1 ( .a ({new_AGEMA_signal_6431, SubBytesIns_Inst_Sbox_9_M43}), .b ({new_AGEMA_signal_5241, SubBytesIns_Inst_Sbox_9_T16}), .clk (clk), .r (Fresh[485]), .c ({new_AGEMA_signal_6671, SubBytesIns_Inst_Sbox_9_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M50_U1 ( .a ({new_AGEMA_signal_6246, SubBytesIns_Inst_Sbox_9_M38}), .b ({new_AGEMA_signal_5238, SubBytesIns_Inst_Sbox_9_T9}), .clk (clk), .r (Fresh[486]), .c ({new_AGEMA_signal_6435, SubBytesIns_Inst_Sbox_9_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M51_U1 ( .a ({new_AGEMA_signal_6245, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_5465, SubBytesIns_Inst_Sbox_9_T17}), .clk (clk), .r (Fresh[487]), .c ({new_AGEMA_signal_6436, SubBytesIns_Inst_Sbox_9_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M52_U1 ( .a ({new_AGEMA_signal_6430, SubBytesIns_Inst_Sbox_9_M42}), .b ({new_AGEMA_signal_5240, SubBytesIns_Inst_Sbox_9_T15}), .clk (clk), .r (Fresh[488]), .c ({new_AGEMA_signal_6672, SubBytesIns_Inst_Sbox_9_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M53_U1 ( .a ({new_AGEMA_signal_6669, SubBytesIns_Inst_Sbox_9_M45}), .b ({new_AGEMA_signal_5244, SubBytesIns_Inst_Sbox_9_T27}), .clk (clk), .r (Fresh[489]), .c ({new_AGEMA_signal_6883, SubBytesIns_Inst_Sbox_9_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M54_U1 ( .a ({new_AGEMA_signal_6429, SubBytesIns_Inst_Sbox_9_M41}), .b ({new_AGEMA_signal_5463, SubBytesIns_Inst_Sbox_9_T10}), .clk (clk), .r (Fresh[490]), .c ({new_AGEMA_signal_6673, SubBytesIns_Inst_Sbox_9_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M55_U1 ( .a ({new_AGEMA_signal_6432, SubBytesIns_Inst_Sbox_9_M44}), .b ({new_AGEMA_signal_5239, SubBytesIns_Inst_Sbox_9_T13}), .clk (clk), .r (Fresh[491]), .c ({new_AGEMA_signal_6674, SubBytesIns_Inst_Sbox_9_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M56_U1 ( .a ({new_AGEMA_signal_6248, SubBytesIns_Inst_Sbox_9_M40}), .b ({new_AGEMA_signal_5467, SubBytesIns_Inst_Sbox_9_T23}), .clk (clk), .r (Fresh[492]), .c ({new_AGEMA_signal_6437, SubBytesIns_Inst_Sbox_9_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M57_U1 ( .a ({new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_9_M39}), .b ({new_AGEMA_signal_5242, SubBytesIns_Inst_Sbox_9_T19}), .clk (clk), .r (Fresh[493]), .c ({new_AGEMA_signal_6438, SubBytesIns_Inst_Sbox_9_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M58_U1 ( .a ({new_AGEMA_signal_6431, SubBytesIns_Inst_Sbox_9_M43}), .b ({new_AGEMA_signal_5065, SubBytesIns_Inst_Sbox_9_T3}), .clk (clk), .r (Fresh[494]), .c ({new_AGEMA_signal_6675, SubBytesIns_Inst_Sbox_9_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M59_U1 ( .a ({new_AGEMA_signal_6246, SubBytesIns_Inst_Sbox_9_M38}), .b ({new_AGEMA_signal_5243, SubBytesIns_Inst_Sbox_9_T22}), .clk (clk), .r (Fresh[495]), .c ({new_AGEMA_signal_6439, SubBytesIns_Inst_Sbox_9_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M60_U1 ( .a ({new_AGEMA_signal_6245, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_5466, SubBytesIns_Inst_Sbox_9_T20}), .clk (clk), .r (Fresh[496]), .c ({new_AGEMA_signal_6440, SubBytesIns_Inst_Sbox_9_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M61_U1 ( .a ({new_AGEMA_signal_6430, SubBytesIns_Inst_Sbox_9_M42}), .b ({new_AGEMA_signal_5063, SubBytesIns_Inst_Sbox_9_T1}), .clk (clk), .r (Fresh[497]), .c ({new_AGEMA_signal_6676, SubBytesIns_Inst_Sbox_9_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M62_U1 ( .a ({new_AGEMA_signal_6669, SubBytesIns_Inst_Sbox_9_M45}), .b ({new_AGEMA_signal_5066, SubBytesIns_Inst_Sbox_9_T4}), .clk (clk), .r (Fresh[498]), .c ({new_AGEMA_signal_6884, SubBytesIns_Inst_Sbox_9_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M63_U1 ( .a ({new_AGEMA_signal_6429, SubBytesIns_Inst_Sbox_9_M41}), .b ({new_AGEMA_signal_5064, SubBytesIns_Inst_Sbox_9_T2}), .clk (clk), .r (Fresh[499]), .c ({new_AGEMA_signal_6677, SubBytesIns_Inst_Sbox_9_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L0_U1 ( .a ({new_AGEMA_signal_6676, SubBytesIns_Inst_Sbox_9_M61}), .b ({new_AGEMA_signal_6884, SubBytesIns_Inst_Sbox_9_M62}), .c ({new_AGEMA_signal_7070, SubBytesIns_Inst_Sbox_9_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L1_U1 ( .a ({new_AGEMA_signal_6435, SubBytesIns_Inst_Sbox_9_M50}), .b ({new_AGEMA_signal_6437, SubBytesIns_Inst_Sbox_9_M56}), .c ({new_AGEMA_signal_6678, SubBytesIns_Inst_Sbox_9_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L2_U1 ( .a ({new_AGEMA_signal_6670, SubBytesIns_Inst_Sbox_9_M46}), .b ({new_AGEMA_signal_6434, SubBytesIns_Inst_Sbox_9_M48}), .c ({new_AGEMA_signal_6885, SubBytesIns_Inst_Sbox_9_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L3_U1 ( .a ({new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_9_M47}), .b ({new_AGEMA_signal_6674, SubBytesIns_Inst_Sbox_9_M55}), .c ({new_AGEMA_signal_6886, SubBytesIns_Inst_Sbox_9_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L4_U1 ( .a ({new_AGEMA_signal_6673, SubBytesIns_Inst_Sbox_9_M54}), .b ({new_AGEMA_signal_6675, SubBytesIns_Inst_Sbox_9_M58}), .c ({new_AGEMA_signal_6887, SubBytesIns_Inst_Sbox_9_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L5_U1 ( .a ({new_AGEMA_signal_6671, SubBytesIns_Inst_Sbox_9_M49}), .b ({new_AGEMA_signal_6676, SubBytesIns_Inst_Sbox_9_M61}), .c ({new_AGEMA_signal_6888, SubBytesIns_Inst_Sbox_9_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L6_U1 ( .a ({new_AGEMA_signal_6884, SubBytesIns_Inst_Sbox_9_M62}), .b ({new_AGEMA_signal_6888, SubBytesIns_Inst_Sbox_9_L5}), .c ({new_AGEMA_signal_7071, SubBytesIns_Inst_Sbox_9_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L7_U1 ( .a ({new_AGEMA_signal_6670, SubBytesIns_Inst_Sbox_9_M46}), .b ({new_AGEMA_signal_6886, SubBytesIns_Inst_Sbox_9_L3}), .c ({new_AGEMA_signal_7072, SubBytesIns_Inst_Sbox_9_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L8_U1 ( .a ({new_AGEMA_signal_6436, SubBytesIns_Inst_Sbox_9_M51}), .b ({new_AGEMA_signal_6439, SubBytesIns_Inst_Sbox_9_M59}), .c ({new_AGEMA_signal_6679, SubBytesIns_Inst_Sbox_9_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L9_U1 ( .a ({new_AGEMA_signal_6672, SubBytesIns_Inst_Sbox_9_M52}), .b ({new_AGEMA_signal_6883, SubBytesIns_Inst_Sbox_9_M53}), .c ({new_AGEMA_signal_7073, SubBytesIns_Inst_Sbox_9_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L10_U1 ( .a ({new_AGEMA_signal_6883, SubBytesIns_Inst_Sbox_9_M53}), .b ({new_AGEMA_signal_6887, SubBytesIns_Inst_Sbox_9_L4}), .c ({new_AGEMA_signal_7074, SubBytesIns_Inst_Sbox_9_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L11_U1 ( .a ({new_AGEMA_signal_6440, SubBytesIns_Inst_Sbox_9_M60}), .b ({new_AGEMA_signal_6885, SubBytesIns_Inst_Sbox_9_L2}), .c ({new_AGEMA_signal_7075, SubBytesIns_Inst_Sbox_9_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L12_U1 ( .a ({new_AGEMA_signal_6434, SubBytesIns_Inst_Sbox_9_M48}), .b ({new_AGEMA_signal_6436, SubBytesIns_Inst_Sbox_9_M51}), .c ({new_AGEMA_signal_6680, SubBytesIns_Inst_Sbox_9_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L13_U1 ( .a ({new_AGEMA_signal_6435, SubBytesIns_Inst_Sbox_9_M50}), .b ({new_AGEMA_signal_7070, SubBytesIns_Inst_Sbox_9_L0}), .c ({new_AGEMA_signal_7276, SubBytesIns_Inst_Sbox_9_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L14_U1 ( .a ({new_AGEMA_signal_6672, SubBytesIns_Inst_Sbox_9_M52}), .b ({new_AGEMA_signal_6676, SubBytesIns_Inst_Sbox_9_M61}), .c ({new_AGEMA_signal_6889, SubBytesIns_Inst_Sbox_9_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L15_U1 ( .a ({new_AGEMA_signal_6674, SubBytesIns_Inst_Sbox_9_M55}), .b ({new_AGEMA_signal_6678, SubBytesIns_Inst_Sbox_9_L1}), .c ({new_AGEMA_signal_6890, SubBytesIns_Inst_Sbox_9_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L16_U1 ( .a ({new_AGEMA_signal_6437, SubBytesIns_Inst_Sbox_9_M56}), .b ({new_AGEMA_signal_7070, SubBytesIns_Inst_Sbox_9_L0}), .c ({new_AGEMA_signal_7277, SubBytesIns_Inst_Sbox_9_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L17_U1 ( .a ({new_AGEMA_signal_6438, SubBytesIns_Inst_Sbox_9_M57}), .b ({new_AGEMA_signal_6678, SubBytesIns_Inst_Sbox_9_L1}), .c ({new_AGEMA_signal_6891, SubBytesIns_Inst_Sbox_9_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L18_U1 ( .a ({new_AGEMA_signal_6675, SubBytesIns_Inst_Sbox_9_M58}), .b ({new_AGEMA_signal_6679, SubBytesIns_Inst_Sbox_9_L8}), .c ({new_AGEMA_signal_6892, SubBytesIns_Inst_Sbox_9_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L19_U1 ( .a ({new_AGEMA_signal_6677, SubBytesIns_Inst_Sbox_9_M63}), .b ({new_AGEMA_signal_6887, SubBytesIns_Inst_Sbox_9_L4}), .c ({new_AGEMA_signal_7076, SubBytesIns_Inst_Sbox_9_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L20_U1 ( .a ({new_AGEMA_signal_7070, SubBytesIns_Inst_Sbox_9_L0}), .b ({new_AGEMA_signal_6678, SubBytesIns_Inst_Sbox_9_L1}), .c ({new_AGEMA_signal_7278, SubBytesIns_Inst_Sbox_9_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L21_U1 ( .a ({new_AGEMA_signal_6678, SubBytesIns_Inst_Sbox_9_L1}), .b ({new_AGEMA_signal_7072, SubBytesIns_Inst_Sbox_9_L7}), .c ({new_AGEMA_signal_7279, SubBytesIns_Inst_Sbox_9_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L22_U1 ( .a ({new_AGEMA_signal_6886, SubBytesIns_Inst_Sbox_9_L3}), .b ({new_AGEMA_signal_6680, SubBytesIns_Inst_Sbox_9_L12}), .c ({new_AGEMA_signal_7077, SubBytesIns_Inst_Sbox_9_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L23_U1 ( .a ({new_AGEMA_signal_6892, SubBytesIns_Inst_Sbox_9_L18}), .b ({new_AGEMA_signal_6885, SubBytesIns_Inst_Sbox_9_L2}), .c ({new_AGEMA_signal_7078, SubBytesIns_Inst_Sbox_9_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L24_U1 ( .a ({new_AGEMA_signal_6890, SubBytesIns_Inst_Sbox_9_L15}), .b ({new_AGEMA_signal_7073, SubBytesIns_Inst_Sbox_9_L9}), .c ({new_AGEMA_signal_7280, SubBytesIns_Inst_Sbox_9_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L25_U1 ( .a ({new_AGEMA_signal_7071, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_7074, SubBytesIns_Inst_Sbox_9_L10}), .c ({new_AGEMA_signal_7281, SubBytesIns_Inst_Sbox_9_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L26_U1 ( .a ({new_AGEMA_signal_7072, SubBytesIns_Inst_Sbox_9_L7}), .b ({new_AGEMA_signal_7073, SubBytesIns_Inst_Sbox_9_L9}), .c ({new_AGEMA_signal_7282, SubBytesIns_Inst_Sbox_9_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L27_U1 ( .a ({new_AGEMA_signal_6679, SubBytesIns_Inst_Sbox_9_L8}), .b ({new_AGEMA_signal_7074, SubBytesIns_Inst_Sbox_9_L10}), .c ({new_AGEMA_signal_7283, SubBytesIns_Inst_Sbox_9_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L28_U1 ( .a ({new_AGEMA_signal_7075, SubBytesIns_Inst_Sbox_9_L11}), .b ({new_AGEMA_signal_6889, SubBytesIns_Inst_Sbox_9_L14}), .c ({new_AGEMA_signal_7284, SubBytesIns_Inst_Sbox_9_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L29_U1 ( .a ({new_AGEMA_signal_7075, SubBytesIns_Inst_Sbox_9_L11}), .b ({new_AGEMA_signal_6891, SubBytesIns_Inst_Sbox_9_L17}), .c ({new_AGEMA_signal_7285, SubBytesIns_Inst_Sbox_9_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S0_U1 ( .a ({new_AGEMA_signal_7071, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_7280, SubBytesIns_Inst_Sbox_9_L24}), .c ({new_AGEMA_signal_7448, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S1_U1 ( .a ({new_AGEMA_signal_7277, SubBytesIns_Inst_Sbox_9_L16}), .b ({new_AGEMA_signal_7282, SubBytesIns_Inst_Sbox_9_L26}), .c ({new_AGEMA_signal_7449, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S2_U1 ( .a ({new_AGEMA_signal_7076, SubBytesIns_Inst_Sbox_9_L19}), .b ({new_AGEMA_signal_7284, SubBytesIns_Inst_Sbox_9_L28}), .c ({new_AGEMA_signal_7450, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S3_U1 ( .a ({new_AGEMA_signal_7071, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_7279, SubBytesIns_Inst_Sbox_9_L21}), .c ({new_AGEMA_signal_7451, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S4_U1 ( .a ({new_AGEMA_signal_7278, SubBytesIns_Inst_Sbox_9_L20}), .b ({new_AGEMA_signal_7077, SubBytesIns_Inst_Sbox_9_L22}), .c ({new_AGEMA_signal_7452, MixColumnsInput[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S5_U1 ( .a ({new_AGEMA_signal_7281, SubBytesIns_Inst_Sbox_9_L25}), .b ({new_AGEMA_signal_7285, SubBytesIns_Inst_Sbox_9_L29}), .c ({new_AGEMA_signal_7453, MixColumnsInput[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S6_U1 ( .a ({new_AGEMA_signal_7276, SubBytesIns_Inst_Sbox_9_L13}), .b ({new_AGEMA_signal_7283, SubBytesIns_Inst_Sbox_9_L27}), .c ({new_AGEMA_signal_7454, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S7_U1 ( .a ({new_AGEMA_signal_7071, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_7078, SubBytesIns_Inst_Sbox_9_L23}), .c ({new_AGEMA_signal_7286, MixColumnsInput[8]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M46_U1 ( .a ({new_AGEMA_signal_6444, SubBytesIns_Inst_Sbox_10_M44}), .b ({new_AGEMA_signal_5245, SubBytesIns_Inst_Sbox_10_T6}), .clk (clk), .r (Fresh[500]), .c ({new_AGEMA_signal_6682, SubBytesIns_Inst_Sbox_10_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M47_U1 ( .a ({new_AGEMA_signal_6252, SubBytesIns_Inst_Sbox_10_M40}), .b ({new_AGEMA_signal_5475, SubBytesIns_Inst_Sbox_10_T8}), .clk (clk), .r (Fresh[501]), .c ({new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_10_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M48_U1 ( .a ({new_AGEMA_signal_6251, SubBytesIns_Inst_Sbox_10_M39}), .b ({ciphertext_s1[80], ciphertext_s0[80]}), .clk (clk), .r (Fresh[502]), .c ({new_AGEMA_signal_6446, SubBytesIns_Inst_Sbox_10_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M49_U1 ( .a ({new_AGEMA_signal_6443, SubBytesIns_Inst_Sbox_10_M43}), .b ({new_AGEMA_signal_5249, SubBytesIns_Inst_Sbox_10_T16}), .clk (clk), .r (Fresh[503]), .c ({new_AGEMA_signal_6683, SubBytesIns_Inst_Sbox_10_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M50_U1 ( .a ({new_AGEMA_signal_6250, SubBytesIns_Inst_Sbox_10_M38}), .b ({new_AGEMA_signal_5246, SubBytesIns_Inst_Sbox_10_T9}), .clk (clk), .r (Fresh[504]), .c ({new_AGEMA_signal_6447, SubBytesIns_Inst_Sbox_10_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M51_U1 ( .a ({new_AGEMA_signal_6249, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_5478, SubBytesIns_Inst_Sbox_10_T17}), .clk (clk), .r (Fresh[505]), .c ({new_AGEMA_signal_6448, SubBytesIns_Inst_Sbox_10_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M52_U1 ( .a ({new_AGEMA_signal_6442, SubBytesIns_Inst_Sbox_10_M42}), .b ({new_AGEMA_signal_5248, SubBytesIns_Inst_Sbox_10_T15}), .clk (clk), .r (Fresh[506]), .c ({new_AGEMA_signal_6684, SubBytesIns_Inst_Sbox_10_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M53_U1 ( .a ({new_AGEMA_signal_6681, SubBytesIns_Inst_Sbox_10_M45}), .b ({new_AGEMA_signal_5252, SubBytesIns_Inst_Sbox_10_T27}), .clk (clk), .r (Fresh[507]), .c ({new_AGEMA_signal_6893, SubBytesIns_Inst_Sbox_10_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M54_U1 ( .a ({new_AGEMA_signal_6441, SubBytesIns_Inst_Sbox_10_M41}), .b ({new_AGEMA_signal_5476, SubBytesIns_Inst_Sbox_10_T10}), .clk (clk), .r (Fresh[508]), .c ({new_AGEMA_signal_6685, SubBytesIns_Inst_Sbox_10_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M55_U1 ( .a ({new_AGEMA_signal_6444, SubBytesIns_Inst_Sbox_10_M44}), .b ({new_AGEMA_signal_5247, SubBytesIns_Inst_Sbox_10_T13}), .clk (clk), .r (Fresh[509]), .c ({new_AGEMA_signal_6686, SubBytesIns_Inst_Sbox_10_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M56_U1 ( .a ({new_AGEMA_signal_6252, SubBytesIns_Inst_Sbox_10_M40}), .b ({new_AGEMA_signal_5480, SubBytesIns_Inst_Sbox_10_T23}), .clk (clk), .r (Fresh[510]), .c ({new_AGEMA_signal_6449, SubBytesIns_Inst_Sbox_10_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M57_U1 ( .a ({new_AGEMA_signal_6251, SubBytesIns_Inst_Sbox_10_M39}), .b ({new_AGEMA_signal_5250, SubBytesIns_Inst_Sbox_10_T19}), .clk (clk), .r (Fresh[511]), .c ({new_AGEMA_signal_6450, SubBytesIns_Inst_Sbox_10_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M58_U1 ( .a ({new_AGEMA_signal_6443, SubBytesIns_Inst_Sbox_10_M43}), .b ({new_AGEMA_signal_5075, SubBytesIns_Inst_Sbox_10_T3}), .clk (clk), .r (Fresh[512]), .c ({new_AGEMA_signal_6687, SubBytesIns_Inst_Sbox_10_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M59_U1 ( .a ({new_AGEMA_signal_6250, SubBytesIns_Inst_Sbox_10_M38}), .b ({new_AGEMA_signal_5251, SubBytesIns_Inst_Sbox_10_T22}), .clk (clk), .r (Fresh[513]), .c ({new_AGEMA_signal_6451, SubBytesIns_Inst_Sbox_10_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M60_U1 ( .a ({new_AGEMA_signal_6249, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_5479, SubBytesIns_Inst_Sbox_10_T20}), .clk (clk), .r (Fresh[514]), .c ({new_AGEMA_signal_6452, SubBytesIns_Inst_Sbox_10_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M61_U1 ( .a ({new_AGEMA_signal_6442, SubBytesIns_Inst_Sbox_10_M42}), .b ({new_AGEMA_signal_5073, SubBytesIns_Inst_Sbox_10_T1}), .clk (clk), .r (Fresh[515]), .c ({new_AGEMA_signal_6688, SubBytesIns_Inst_Sbox_10_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M62_U1 ( .a ({new_AGEMA_signal_6681, SubBytesIns_Inst_Sbox_10_M45}), .b ({new_AGEMA_signal_5076, SubBytesIns_Inst_Sbox_10_T4}), .clk (clk), .r (Fresh[516]), .c ({new_AGEMA_signal_6894, SubBytesIns_Inst_Sbox_10_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M63_U1 ( .a ({new_AGEMA_signal_6441, SubBytesIns_Inst_Sbox_10_M41}), .b ({new_AGEMA_signal_5074, SubBytesIns_Inst_Sbox_10_T2}), .clk (clk), .r (Fresh[517]), .c ({new_AGEMA_signal_6689, SubBytesIns_Inst_Sbox_10_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L0_U1 ( .a ({new_AGEMA_signal_6688, SubBytesIns_Inst_Sbox_10_M61}), .b ({new_AGEMA_signal_6894, SubBytesIns_Inst_Sbox_10_M62}), .c ({new_AGEMA_signal_7079, SubBytesIns_Inst_Sbox_10_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L1_U1 ( .a ({new_AGEMA_signal_6447, SubBytesIns_Inst_Sbox_10_M50}), .b ({new_AGEMA_signal_6449, SubBytesIns_Inst_Sbox_10_M56}), .c ({new_AGEMA_signal_6690, SubBytesIns_Inst_Sbox_10_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L2_U1 ( .a ({new_AGEMA_signal_6682, SubBytesIns_Inst_Sbox_10_M46}), .b ({new_AGEMA_signal_6446, SubBytesIns_Inst_Sbox_10_M48}), .c ({new_AGEMA_signal_6895, SubBytesIns_Inst_Sbox_10_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L3_U1 ( .a ({new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_10_M47}), .b ({new_AGEMA_signal_6686, SubBytesIns_Inst_Sbox_10_M55}), .c ({new_AGEMA_signal_6896, SubBytesIns_Inst_Sbox_10_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L4_U1 ( .a ({new_AGEMA_signal_6685, SubBytesIns_Inst_Sbox_10_M54}), .b ({new_AGEMA_signal_6687, SubBytesIns_Inst_Sbox_10_M58}), .c ({new_AGEMA_signal_6897, SubBytesIns_Inst_Sbox_10_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L5_U1 ( .a ({new_AGEMA_signal_6683, SubBytesIns_Inst_Sbox_10_M49}), .b ({new_AGEMA_signal_6688, SubBytesIns_Inst_Sbox_10_M61}), .c ({new_AGEMA_signal_6898, SubBytesIns_Inst_Sbox_10_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L6_U1 ( .a ({new_AGEMA_signal_6894, SubBytesIns_Inst_Sbox_10_M62}), .b ({new_AGEMA_signal_6898, SubBytesIns_Inst_Sbox_10_L5}), .c ({new_AGEMA_signal_7080, SubBytesIns_Inst_Sbox_10_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L7_U1 ( .a ({new_AGEMA_signal_6682, SubBytesIns_Inst_Sbox_10_M46}), .b ({new_AGEMA_signal_6896, SubBytesIns_Inst_Sbox_10_L3}), .c ({new_AGEMA_signal_7081, SubBytesIns_Inst_Sbox_10_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L8_U1 ( .a ({new_AGEMA_signal_6448, SubBytesIns_Inst_Sbox_10_M51}), .b ({new_AGEMA_signal_6451, SubBytesIns_Inst_Sbox_10_M59}), .c ({new_AGEMA_signal_6691, SubBytesIns_Inst_Sbox_10_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L9_U1 ( .a ({new_AGEMA_signal_6684, SubBytesIns_Inst_Sbox_10_M52}), .b ({new_AGEMA_signal_6893, SubBytesIns_Inst_Sbox_10_M53}), .c ({new_AGEMA_signal_7082, SubBytesIns_Inst_Sbox_10_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L10_U1 ( .a ({new_AGEMA_signal_6893, SubBytesIns_Inst_Sbox_10_M53}), .b ({new_AGEMA_signal_6897, SubBytesIns_Inst_Sbox_10_L4}), .c ({new_AGEMA_signal_7083, SubBytesIns_Inst_Sbox_10_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L11_U1 ( .a ({new_AGEMA_signal_6452, SubBytesIns_Inst_Sbox_10_M60}), .b ({new_AGEMA_signal_6895, SubBytesIns_Inst_Sbox_10_L2}), .c ({new_AGEMA_signal_7084, SubBytesIns_Inst_Sbox_10_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L12_U1 ( .a ({new_AGEMA_signal_6446, SubBytesIns_Inst_Sbox_10_M48}), .b ({new_AGEMA_signal_6448, SubBytesIns_Inst_Sbox_10_M51}), .c ({new_AGEMA_signal_6692, SubBytesIns_Inst_Sbox_10_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L13_U1 ( .a ({new_AGEMA_signal_6447, SubBytesIns_Inst_Sbox_10_M50}), .b ({new_AGEMA_signal_7079, SubBytesIns_Inst_Sbox_10_L0}), .c ({new_AGEMA_signal_7287, SubBytesIns_Inst_Sbox_10_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L14_U1 ( .a ({new_AGEMA_signal_6684, SubBytesIns_Inst_Sbox_10_M52}), .b ({new_AGEMA_signal_6688, SubBytesIns_Inst_Sbox_10_M61}), .c ({new_AGEMA_signal_6899, SubBytesIns_Inst_Sbox_10_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L15_U1 ( .a ({new_AGEMA_signal_6686, SubBytesIns_Inst_Sbox_10_M55}), .b ({new_AGEMA_signal_6690, SubBytesIns_Inst_Sbox_10_L1}), .c ({new_AGEMA_signal_6900, SubBytesIns_Inst_Sbox_10_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L16_U1 ( .a ({new_AGEMA_signal_6449, SubBytesIns_Inst_Sbox_10_M56}), .b ({new_AGEMA_signal_7079, SubBytesIns_Inst_Sbox_10_L0}), .c ({new_AGEMA_signal_7288, SubBytesIns_Inst_Sbox_10_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L17_U1 ( .a ({new_AGEMA_signal_6450, SubBytesIns_Inst_Sbox_10_M57}), .b ({new_AGEMA_signal_6690, SubBytesIns_Inst_Sbox_10_L1}), .c ({new_AGEMA_signal_6901, SubBytesIns_Inst_Sbox_10_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L18_U1 ( .a ({new_AGEMA_signal_6687, SubBytesIns_Inst_Sbox_10_M58}), .b ({new_AGEMA_signal_6691, SubBytesIns_Inst_Sbox_10_L8}), .c ({new_AGEMA_signal_6902, SubBytesIns_Inst_Sbox_10_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L19_U1 ( .a ({new_AGEMA_signal_6689, SubBytesIns_Inst_Sbox_10_M63}), .b ({new_AGEMA_signal_6897, SubBytesIns_Inst_Sbox_10_L4}), .c ({new_AGEMA_signal_7085, SubBytesIns_Inst_Sbox_10_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L20_U1 ( .a ({new_AGEMA_signal_7079, SubBytesIns_Inst_Sbox_10_L0}), .b ({new_AGEMA_signal_6690, SubBytesIns_Inst_Sbox_10_L1}), .c ({new_AGEMA_signal_7289, SubBytesIns_Inst_Sbox_10_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L21_U1 ( .a ({new_AGEMA_signal_6690, SubBytesIns_Inst_Sbox_10_L1}), .b ({new_AGEMA_signal_7081, SubBytesIns_Inst_Sbox_10_L7}), .c ({new_AGEMA_signal_7290, SubBytesIns_Inst_Sbox_10_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L22_U1 ( .a ({new_AGEMA_signal_6896, SubBytesIns_Inst_Sbox_10_L3}), .b ({new_AGEMA_signal_6692, SubBytesIns_Inst_Sbox_10_L12}), .c ({new_AGEMA_signal_7086, SubBytesIns_Inst_Sbox_10_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L23_U1 ( .a ({new_AGEMA_signal_6902, SubBytesIns_Inst_Sbox_10_L18}), .b ({new_AGEMA_signal_6895, SubBytesIns_Inst_Sbox_10_L2}), .c ({new_AGEMA_signal_7087, SubBytesIns_Inst_Sbox_10_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L24_U1 ( .a ({new_AGEMA_signal_6900, SubBytesIns_Inst_Sbox_10_L15}), .b ({new_AGEMA_signal_7082, SubBytesIns_Inst_Sbox_10_L9}), .c ({new_AGEMA_signal_7291, SubBytesIns_Inst_Sbox_10_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L25_U1 ( .a ({new_AGEMA_signal_7080, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_7083, SubBytesIns_Inst_Sbox_10_L10}), .c ({new_AGEMA_signal_7292, SubBytesIns_Inst_Sbox_10_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L26_U1 ( .a ({new_AGEMA_signal_7081, SubBytesIns_Inst_Sbox_10_L7}), .b ({new_AGEMA_signal_7082, SubBytesIns_Inst_Sbox_10_L9}), .c ({new_AGEMA_signal_7293, SubBytesIns_Inst_Sbox_10_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L27_U1 ( .a ({new_AGEMA_signal_6691, SubBytesIns_Inst_Sbox_10_L8}), .b ({new_AGEMA_signal_7083, SubBytesIns_Inst_Sbox_10_L10}), .c ({new_AGEMA_signal_7294, SubBytesIns_Inst_Sbox_10_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L28_U1 ( .a ({new_AGEMA_signal_7084, SubBytesIns_Inst_Sbox_10_L11}), .b ({new_AGEMA_signal_6899, SubBytesIns_Inst_Sbox_10_L14}), .c ({new_AGEMA_signal_7295, SubBytesIns_Inst_Sbox_10_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L29_U1 ( .a ({new_AGEMA_signal_7084, SubBytesIns_Inst_Sbox_10_L11}), .b ({new_AGEMA_signal_6901, SubBytesIns_Inst_Sbox_10_L17}), .c ({new_AGEMA_signal_7296, SubBytesIns_Inst_Sbox_10_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S0_U1 ( .a ({new_AGEMA_signal_7080, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_7291, SubBytesIns_Inst_Sbox_10_L24}), .c ({new_AGEMA_signal_7455, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S1_U1 ( .a ({new_AGEMA_signal_7288, SubBytesIns_Inst_Sbox_10_L16}), .b ({new_AGEMA_signal_7293, SubBytesIns_Inst_Sbox_10_L26}), .c ({new_AGEMA_signal_7456, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S2_U1 ( .a ({new_AGEMA_signal_7085, SubBytesIns_Inst_Sbox_10_L19}), .b ({new_AGEMA_signal_7295, SubBytesIns_Inst_Sbox_10_L28}), .c ({new_AGEMA_signal_7457, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S3_U1 ( .a ({new_AGEMA_signal_7080, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_7290, SubBytesIns_Inst_Sbox_10_L21}), .c ({new_AGEMA_signal_7458, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S4_U1 ( .a ({new_AGEMA_signal_7289, SubBytesIns_Inst_Sbox_10_L20}), .b ({new_AGEMA_signal_7086, SubBytesIns_Inst_Sbox_10_L22}), .c ({new_AGEMA_signal_7459, MixColumnsInput[115]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S5_U1 ( .a ({new_AGEMA_signal_7292, SubBytesIns_Inst_Sbox_10_L25}), .b ({new_AGEMA_signal_7296, SubBytesIns_Inst_Sbox_10_L29}), .c ({new_AGEMA_signal_7460, MixColumnsInput[114]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S6_U1 ( .a ({new_AGEMA_signal_7287, SubBytesIns_Inst_Sbox_10_L13}), .b ({new_AGEMA_signal_7294, SubBytesIns_Inst_Sbox_10_L27}), .c ({new_AGEMA_signal_7461, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S7_U1 ( .a ({new_AGEMA_signal_7080, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_7087, SubBytesIns_Inst_Sbox_10_L23}), .c ({new_AGEMA_signal_7297, MixColumnsInput[112]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M46_U1 ( .a ({new_AGEMA_signal_6456, SubBytesIns_Inst_Sbox_11_M44}), .b ({new_AGEMA_signal_5253, SubBytesIns_Inst_Sbox_11_T6}), .clk (clk), .r (Fresh[518]), .c ({new_AGEMA_signal_6694, SubBytesIns_Inst_Sbox_11_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M47_U1 ( .a ({new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_11_M40}), .b ({new_AGEMA_signal_5488, SubBytesIns_Inst_Sbox_11_T8}), .clk (clk), .r (Fresh[519]), .c ({new_AGEMA_signal_6457, SubBytesIns_Inst_Sbox_11_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M48_U1 ( .a ({new_AGEMA_signal_6255, SubBytesIns_Inst_Sbox_11_M39}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .clk (clk), .r (Fresh[520]), .c ({new_AGEMA_signal_6458, SubBytesIns_Inst_Sbox_11_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M49_U1 ( .a ({new_AGEMA_signal_6455, SubBytesIns_Inst_Sbox_11_M43}), .b ({new_AGEMA_signal_5257, SubBytesIns_Inst_Sbox_11_T16}), .clk (clk), .r (Fresh[521]), .c ({new_AGEMA_signal_6695, SubBytesIns_Inst_Sbox_11_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M50_U1 ( .a ({new_AGEMA_signal_6254, SubBytesIns_Inst_Sbox_11_M38}), .b ({new_AGEMA_signal_5254, SubBytesIns_Inst_Sbox_11_T9}), .clk (clk), .r (Fresh[522]), .c ({new_AGEMA_signal_6459, SubBytesIns_Inst_Sbox_11_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M51_U1 ( .a ({new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_5491, SubBytesIns_Inst_Sbox_11_T17}), .clk (clk), .r (Fresh[523]), .c ({new_AGEMA_signal_6460, SubBytesIns_Inst_Sbox_11_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M52_U1 ( .a ({new_AGEMA_signal_6454, SubBytesIns_Inst_Sbox_11_M42}), .b ({new_AGEMA_signal_5256, SubBytesIns_Inst_Sbox_11_T15}), .clk (clk), .r (Fresh[524]), .c ({new_AGEMA_signal_6696, SubBytesIns_Inst_Sbox_11_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M53_U1 ( .a ({new_AGEMA_signal_6693, SubBytesIns_Inst_Sbox_11_M45}), .b ({new_AGEMA_signal_5260, SubBytesIns_Inst_Sbox_11_T27}), .clk (clk), .r (Fresh[525]), .c ({new_AGEMA_signal_6903, SubBytesIns_Inst_Sbox_11_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M54_U1 ( .a ({new_AGEMA_signal_6453, SubBytesIns_Inst_Sbox_11_M41}), .b ({new_AGEMA_signal_5489, SubBytesIns_Inst_Sbox_11_T10}), .clk (clk), .r (Fresh[526]), .c ({new_AGEMA_signal_6697, SubBytesIns_Inst_Sbox_11_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M55_U1 ( .a ({new_AGEMA_signal_6456, SubBytesIns_Inst_Sbox_11_M44}), .b ({new_AGEMA_signal_5255, SubBytesIns_Inst_Sbox_11_T13}), .clk (clk), .r (Fresh[527]), .c ({new_AGEMA_signal_6698, SubBytesIns_Inst_Sbox_11_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M56_U1 ( .a ({new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_11_M40}), .b ({new_AGEMA_signal_5493, SubBytesIns_Inst_Sbox_11_T23}), .clk (clk), .r (Fresh[528]), .c ({new_AGEMA_signal_6461, SubBytesIns_Inst_Sbox_11_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M57_U1 ( .a ({new_AGEMA_signal_6255, SubBytesIns_Inst_Sbox_11_M39}), .b ({new_AGEMA_signal_5258, SubBytesIns_Inst_Sbox_11_T19}), .clk (clk), .r (Fresh[529]), .c ({new_AGEMA_signal_6462, SubBytesIns_Inst_Sbox_11_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M58_U1 ( .a ({new_AGEMA_signal_6455, SubBytesIns_Inst_Sbox_11_M43}), .b ({new_AGEMA_signal_5085, SubBytesIns_Inst_Sbox_11_T3}), .clk (clk), .r (Fresh[530]), .c ({new_AGEMA_signal_6699, SubBytesIns_Inst_Sbox_11_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M59_U1 ( .a ({new_AGEMA_signal_6254, SubBytesIns_Inst_Sbox_11_M38}), .b ({new_AGEMA_signal_5259, SubBytesIns_Inst_Sbox_11_T22}), .clk (clk), .r (Fresh[531]), .c ({new_AGEMA_signal_6463, SubBytesIns_Inst_Sbox_11_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M60_U1 ( .a ({new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_5492, SubBytesIns_Inst_Sbox_11_T20}), .clk (clk), .r (Fresh[532]), .c ({new_AGEMA_signal_6464, SubBytesIns_Inst_Sbox_11_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M61_U1 ( .a ({new_AGEMA_signal_6454, SubBytesIns_Inst_Sbox_11_M42}), .b ({new_AGEMA_signal_5083, SubBytesIns_Inst_Sbox_11_T1}), .clk (clk), .r (Fresh[533]), .c ({new_AGEMA_signal_6700, SubBytesIns_Inst_Sbox_11_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M62_U1 ( .a ({new_AGEMA_signal_6693, SubBytesIns_Inst_Sbox_11_M45}), .b ({new_AGEMA_signal_5086, SubBytesIns_Inst_Sbox_11_T4}), .clk (clk), .r (Fresh[534]), .c ({new_AGEMA_signal_6904, SubBytesIns_Inst_Sbox_11_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M63_U1 ( .a ({new_AGEMA_signal_6453, SubBytesIns_Inst_Sbox_11_M41}), .b ({new_AGEMA_signal_5084, SubBytesIns_Inst_Sbox_11_T2}), .clk (clk), .r (Fresh[535]), .c ({new_AGEMA_signal_6701, SubBytesIns_Inst_Sbox_11_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L0_U1 ( .a ({new_AGEMA_signal_6700, SubBytesIns_Inst_Sbox_11_M61}), .b ({new_AGEMA_signal_6904, SubBytesIns_Inst_Sbox_11_M62}), .c ({new_AGEMA_signal_7088, SubBytesIns_Inst_Sbox_11_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L1_U1 ( .a ({new_AGEMA_signal_6459, SubBytesIns_Inst_Sbox_11_M50}), .b ({new_AGEMA_signal_6461, SubBytesIns_Inst_Sbox_11_M56}), .c ({new_AGEMA_signal_6702, SubBytesIns_Inst_Sbox_11_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L2_U1 ( .a ({new_AGEMA_signal_6694, SubBytesIns_Inst_Sbox_11_M46}), .b ({new_AGEMA_signal_6458, SubBytesIns_Inst_Sbox_11_M48}), .c ({new_AGEMA_signal_6905, SubBytesIns_Inst_Sbox_11_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L3_U1 ( .a ({new_AGEMA_signal_6457, SubBytesIns_Inst_Sbox_11_M47}), .b ({new_AGEMA_signal_6698, SubBytesIns_Inst_Sbox_11_M55}), .c ({new_AGEMA_signal_6906, SubBytesIns_Inst_Sbox_11_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L4_U1 ( .a ({new_AGEMA_signal_6697, SubBytesIns_Inst_Sbox_11_M54}), .b ({new_AGEMA_signal_6699, SubBytesIns_Inst_Sbox_11_M58}), .c ({new_AGEMA_signal_6907, SubBytesIns_Inst_Sbox_11_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L5_U1 ( .a ({new_AGEMA_signal_6695, SubBytesIns_Inst_Sbox_11_M49}), .b ({new_AGEMA_signal_6700, SubBytesIns_Inst_Sbox_11_M61}), .c ({new_AGEMA_signal_6908, SubBytesIns_Inst_Sbox_11_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L6_U1 ( .a ({new_AGEMA_signal_6904, SubBytesIns_Inst_Sbox_11_M62}), .b ({new_AGEMA_signal_6908, SubBytesIns_Inst_Sbox_11_L5}), .c ({new_AGEMA_signal_7089, SubBytesIns_Inst_Sbox_11_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L7_U1 ( .a ({new_AGEMA_signal_6694, SubBytesIns_Inst_Sbox_11_M46}), .b ({new_AGEMA_signal_6906, SubBytesIns_Inst_Sbox_11_L3}), .c ({new_AGEMA_signal_7090, SubBytesIns_Inst_Sbox_11_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L8_U1 ( .a ({new_AGEMA_signal_6460, SubBytesIns_Inst_Sbox_11_M51}), .b ({new_AGEMA_signal_6463, SubBytesIns_Inst_Sbox_11_M59}), .c ({new_AGEMA_signal_6703, SubBytesIns_Inst_Sbox_11_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L9_U1 ( .a ({new_AGEMA_signal_6696, SubBytesIns_Inst_Sbox_11_M52}), .b ({new_AGEMA_signal_6903, SubBytesIns_Inst_Sbox_11_M53}), .c ({new_AGEMA_signal_7091, SubBytesIns_Inst_Sbox_11_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L10_U1 ( .a ({new_AGEMA_signal_6903, SubBytesIns_Inst_Sbox_11_M53}), .b ({new_AGEMA_signal_6907, SubBytesIns_Inst_Sbox_11_L4}), .c ({new_AGEMA_signal_7092, SubBytesIns_Inst_Sbox_11_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L11_U1 ( .a ({new_AGEMA_signal_6464, SubBytesIns_Inst_Sbox_11_M60}), .b ({new_AGEMA_signal_6905, SubBytesIns_Inst_Sbox_11_L2}), .c ({new_AGEMA_signal_7093, SubBytesIns_Inst_Sbox_11_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L12_U1 ( .a ({new_AGEMA_signal_6458, SubBytesIns_Inst_Sbox_11_M48}), .b ({new_AGEMA_signal_6460, SubBytesIns_Inst_Sbox_11_M51}), .c ({new_AGEMA_signal_6704, SubBytesIns_Inst_Sbox_11_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L13_U1 ( .a ({new_AGEMA_signal_6459, SubBytesIns_Inst_Sbox_11_M50}), .b ({new_AGEMA_signal_7088, SubBytesIns_Inst_Sbox_11_L0}), .c ({new_AGEMA_signal_7298, SubBytesIns_Inst_Sbox_11_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L14_U1 ( .a ({new_AGEMA_signal_6696, SubBytesIns_Inst_Sbox_11_M52}), .b ({new_AGEMA_signal_6700, SubBytesIns_Inst_Sbox_11_M61}), .c ({new_AGEMA_signal_6909, SubBytesIns_Inst_Sbox_11_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L15_U1 ( .a ({new_AGEMA_signal_6698, SubBytesIns_Inst_Sbox_11_M55}), .b ({new_AGEMA_signal_6702, SubBytesIns_Inst_Sbox_11_L1}), .c ({new_AGEMA_signal_6910, SubBytesIns_Inst_Sbox_11_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L16_U1 ( .a ({new_AGEMA_signal_6461, SubBytesIns_Inst_Sbox_11_M56}), .b ({new_AGEMA_signal_7088, SubBytesIns_Inst_Sbox_11_L0}), .c ({new_AGEMA_signal_7299, SubBytesIns_Inst_Sbox_11_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L17_U1 ( .a ({new_AGEMA_signal_6462, SubBytesIns_Inst_Sbox_11_M57}), .b ({new_AGEMA_signal_6702, SubBytesIns_Inst_Sbox_11_L1}), .c ({new_AGEMA_signal_6911, SubBytesIns_Inst_Sbox_11_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L18_U1 ( .a ({new_AGEMA_signal_6699, SubBytesIns_Inst_Sbox_11_M58}), .b ({new_AGEMA_signal_6703, SubBytesIns_Inst_Sbox_11_L8}), .c ({new_AGEMA_signal_6912, SubBytesIns_Inst_Sbox_11_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L19_U1 ( .a ({new_AGEMA_signal_6701, SubBytesIns_Inst_Sbox_11_M63}), .b ({new_AGEMA_signal_6907, SubBytesIns_Inst_Sbox_11_L4}), .c ({new_AGEMA_signal_7094, SubBytesIns_Inst_Sbox_11_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L20_U1 ( .a ({new_AGEMA_signal_7088, SubBytesIns_Inst_Sbox_11_L0}), .b ({new_AGEMA_signal_6702, SubBytesIns_Inst_Sbox_11_L1}), .c ({new_AGEMA_signal_7300, SubBytesIns_Inst_Sbox_11_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L21_U1 ( .a ({new_AGEMA_signal_6702, SubBytesIns_Inst_Sbox_11_L1}), .b ({new_AGEMA_signal_7090, SubBytesIns_Inst_Sbox_11_L7}), .c ({new_AGEMA_signal_7301, SubBytesIns_Inst_Sbox_11_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L22_U1 ( .a ({new_AGEMA_signal_6906, SubBytesIns_Inst_Sbox_11_L3}), .b ({new_AGEMA_signal_6704, SubBytesIns_Inst_Sbox_11_L12}), .c ({new_AGEMA_signal_7095, SubBytesIns_Inst_Sbox_11_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L23_U1 ( .a ({new_AGEMA_signal_6912, SubBytesIns_Inst_Sbox_11_L18}), .b ({new_AGEMA_signal_6905, SubBytesIns_Inst_Sbox_11_L2}), .c ({new_AGEMA_signal_7096, SubBytesIns_Inst_Sbox_11_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L24_U1 ( .a ({new_AGEMA_signal_6910, SubBytesIns_Inst_Sbox_11_L15}), .b ({new_AGEMA_signal_7091, SubBytesIns_Inst_Sbox_11_L9}), .c ({new_AGEMA_signal_7302, SubBytesIns_Inst_Sbox_11_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L25_U1 ( .a ({new_AGEMA_signal_7089, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_7092, SubBytesIns_Inst_Sbox_11_L10}), .c ({new_AGEMA_signal_7303, SubBytesIns_Inst_Sbox_11_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L26_U1 ( .a ({new_AGEMA_signal_7090, SubBytesIns_Inst_Sbox_11_L7}), .b ({new_AGEMA_signal_7091, SubBytesIns_Inst_Sbox_11_L9}), .c ({new_AGEMA_signal_7304, SubBytesIns_Inst_Sbox_11_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L27_U1 ( .a ({new_AGEMA_signal_6703, SubBytesIns_Inst_Sbox_11_L8}), .b ({new_AGEMA_signal_7092, SubBytesIns_Inst_Sbox_11_L10}), .c ({new_AGEMA_signal_7305, SubBytesIns_Inst_Sbox_11_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L28_U1 ( .a ({new_AGEMA_signal_7093, SubBytesIns_Inst_Sbox_11_L11}), .b ({new_AGEMA_signal_6909, SubBytesIns_Inst_Sbox_11_L14}), .c ({new_AGEMA_signal_7306, SubBytesIns_Inst_Sbox_11_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L29_U1 ( .a ({new_AGEMA_signal_7093, SubBytesIns_Inst_Sbox_11_L11}), .b ({new_AGEMA_signal_6911, SubBytesIns_Inst_Sbox_11_L17}), .c ({new_AGEMA_signal_7307, SubBytesIns_Inst_Sbox_11_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S0_U1 ( .a ({new_AGEMA_signal_7089, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_7302, SubBytesIns_Inst_Sbox_11_L24}), .c ({new_AGEMA_signal_7462, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S1_U1 ( .a ({new_AGEMA_signal_7299, SubBytesIns_Inst_Sbox_11_L16}), .b ({new_AGEMA_signal_7304, SubBytesIns_Inst_Sbox_11_L26}), .c ({new_AGEMA_signal_7463, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S2_U1 ( .a ({new_AGEMA_signal_7094, SubBytesIns_Inst_Sbox_11_L19}), .b ({new_AGEMA_signal_7306, SubBytesIns_Inst_Sbox_11_L28}), .c ({new_AGEMA_signal_7464, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S3_U1 ( .a ({new_AGEMA_signal_7089, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_7301, SubBytesIns_Inst_Sbox_11_L21}), .c ({new_AGEMA_signal_7465, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S4_U1 ( .a ({new_AGEMA_signal_7300, SubBytesIns_Inst_Sbox_11_L20}), .b ({new_AGEMA_signal_7095, SubBytesIns_Inst_Sbox_11_L22}), .c ({new_AGEMA_signal_7466, MixColumnsInput[91]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S5_U1 ( .a ({new_AGEMA_signal_7303, SubBytesIns_Inst_Sbox_11_L25}), .b ({new_AGEMA_signal_7307, SubBytesIns_Inst_Sbox_11_L29}), .c ({new_AGEMA_signal_7467, MixColumnsInput[90]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S6_U1 ( .a ({new_AGEMA_signal_7298, SubBytesIns_Inst_Sbox_11_L13}), .b ({new_AGEMA_signal_7305, SubBytesIns_Inst_Sbox_11_L27}), .c ({new_AGEMA_signal_7468, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S7_U1 ( .a ({new_AGEMA_signal_7089, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_7096, SubBytesIns_Inst_Sbox_11_L23}), .c ({new_AGEMA_signal_7308, MixColumnsInput[88]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M46_U1 ( .a ({new_AGEMA_signal_6468, SubBytesIns_Inst_Sbox_12_M44}), .b ({new_AGEMA_signal_5261, SubBytesIns_Inst_Sbox_12_T6}), .clk (clk), .r (Fresh[536]), .c ({new_AGEMA_signal_6706, SubBytesIns_Inst_Sbox_12_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M47_U1 ( .a ({new_AGEMA_signal_6260, SubBytesIns_Inst_Sbox_12_M40}), .b ({new_AGEMA_signal_5501, SubBytesIns_Inst_Sbox_12_T8}), .clk (clk), .r (Fresh[537]), .c ({new_AGEMA_signal_6469, SubBytesIns_Inst_Sbox_12_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M48_U1 ( .a ({new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_12_M39}), .b ({ciphertext_s1[96], ciphertext_s0[96]}), .clk (clk), .r (Fresh[538]), .c ({new_AGEMA_signal_6470, SubBytesIns_Inst_Sbox_12_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M49_U1 ( .a ({new_AGEMA_signal_6467, SubBytesIns_Inst_Sbox_12_M43}), .b ({new_AGEMA_signal_5265, SubBytesIns_Inst_Sbox_12_T16}), .clk (clk), .r (Fresh[539]), .c ({new_AGEMA_signal_6707, SubBytesIns_Inst_Sbox_12_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M50_U1 ( .a ({new_AGEMA_signal_6258, SubBytesIns_Inst_Sbox_12_M38}), .b ({new_AGEMA_signal_5262, SubBytesIns_Inst_Sbox_12_T9}), .clk (clk), .r (Fresh[540]), .c ({new_AGEMA_signal_6471, SubBytesIns_Inst_Sbox_12_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M51_U1 ( .a ({new_AGEMA_signal_6257, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_5504, SubBytesIns_Inst_Sbox_12_T17}), .clk (clk), .r (Fresh[541]), .c ({new_AGEMA_signal_6472, SubBytesIns_Inst_Sbox_12_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M52_U1 ( .a ({new_AGEMA_signal_6466, SubBytesIns_Inst_Sbox_12_M42}), .b ({new_AGEMA_signal_5264, SubBytesIns_Inst_Sbox_12_T15}), .clk (clk), .r (Fresh[542]), .c ({new_AGEMA_signal_6708, SubBytesIns_Inst_Sbox_12_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M53_U1 ( .a ({new_AGEMA_signal_6705, SubBytesIns_Inst_Sbox_12_M45}), .b ({new_AGEMA_signal_5268, SubBytesIns_Inst_Sbox_12_T27}), .clk (clk), .r (Fresh[543]), .c ({new_AGEMA_signal_6913, SubBytesIns_Inst_Sbox_12_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M54_U1 ( .a ({new_AGEMA_signal_6465, SubBytesIns_Inst_Sbox_12_M41}), .b ({new_AGEMA_signal_5502, SubBytesIns_Inst_Sbox_12_T10}), .clk (clk), .r (Fresh[544]), .c ({new_AGEMA_signal_6709, SubBytesIns_Inst_Sbox_12_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M55_U1 ( .a ({new_AGEMA_signal_6468, SubBytesIns_Inst_Sbox_12_M44}), .b ({new_AGEMA_signal_5263, SubBytesIns_Inst_Sbox_12_T13}), .clk (clk), .r (Fresh[545]), .c ({new_AGEMA_signal_6710, SubBytesIns_Inst_Sbox_12_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M56_U1 ( .a ({new_AGEMA_signal_6260, SubBytesIns_Inst_Sbox_12_M40}), .b ({new_AGEMA_signal_5506, SubBytesIns_Inst_Sbox_12_T23}), .clk (clk), .r (Fresh[546]), .c ({new_AGEMA_signal_6473, SubBytesIns_Inst_Sbox_12_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M57_U1 ( .a ({new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_12_M39}), .b ({new_AGEMA_signal_5266, SubBytesIns_Inst_Sbox_12_T19}), .clk (clk), .r (Fresh[547]), .c ({new_AGEMA_signal_6474, SubBytesIns_Inst_Sbox_12_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M58_U1 ( .a ({new_AGEMA_signal_6467, SubBytesIns_Inst_Sbox_12_M43}), .b ({new_AGEMA_signal_5095, SubBytesIns_Inst_Sbox_12_T3}), .clk (clk), .r (Fresh[548]), .c ({new_AGEMA_signal_6711, SubBytesIns_Inst_Sbox_12_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M59_U1 ( .a ({new_AGEMA_signal_6258, SubBytesIns_Inst_Sbox_12_M38}), .b ({new_AGEMA_signal_5267, SubBytesIns_Inst_Sbox_12_T22}), .clk (clk), .r (Fresh[549]), .c ({new_AGEMA_signal_6475, SubBytesIns_Inst_Sbox_12_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M60_U1 ( .a ({new_AGEMA_signal_6257, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_5505, SubBytesIns_Inst_Sbox_12_T20}), .clk (clk), .r (Fresh[550]), .c ({new_AGEMA_signal_6476, SubBytesIns_Inst_Sbox_12_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M61_U1 ( .a ({new_AGEMA_signal_6466, SubBytesIns_Inst_Sbox_12_M42}), .b ({new_AGEMA_signal_5093, SubBytesIns_Inst_Sbox_12_T1}), .clk (clk), .r (Fresh[551]), .c ({new_AGEMA_signal_6712, SubBytesIns_Inst_Sbox_12_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M62_U1 ( .a ({new_AGEMA_signal_6705, SubBytesIns_Inst_Sbox_12_M45}), .b ({new_AGEMA_signal_5096, SubBytesIns_Inst_Sbox_12_T4}), .clk (clk), .r (Fresh[552]), .c ({new_AGEMA_signal_6914, SubBytesIns_Inst_Sbox_12_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M63_U1 ( .a ({new_AGEMA_signal_6465, SubBytesIns_Inst_Sbox_12_M41}), .b ({new_AGEMA_signal_5094, SubBytesIns_Inst_Sbox_12_T2}), .clk (clk), .r (Fresh[553]), .c ({new_AGEMA_signal_6713, SubBytesIns_Inst_Sbox_12_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L0_U1 ( .a ({new_AGEMA_signal_6712, SubBytesIns_Inst_Sbox_12_M61}), .b ({new_AGEMA_signal_6914, SubBytesIns_Inst_Sbox_12_M62}), .c ({new_AGEMA_signal_7097, SubBytesIns_Inst_Sbox_12_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L1_U1 ( .a ({new_AGEMA_signal_6471, SubBytesIns_Inst_Sbox_12_M50}), .b ({new_AGEMA_signal_6473, SubBytesIns_Inst_Sbox_12_M56}), .c ({new_AGEMA_signal_6714, SubBytesIns_Inst_Sbox_12_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L2_U1 ( .a ({new_AGEMA_signal_6706, SubBytesIns_Inst_Sbox_12_M46}), .b ({new_AGEMA_signal_6470, SubBytesIns_Inst_Sbox_12_M48}), .c ({new_AGEMA_signal_6915, SubBytesIns_Inst_Sbox_12_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L3_U1 ( .a ({new_AGEMA_signal_6469, SubBytesIns_Inst_Sbox_12_M47}), .b ({new_AGEMA_signal_6710, SubBytesIns_Inst_Sbox_12_M55}), .c ({new_AGEMA_signal_6916, SubBytesIns_Inst_Sbox_12_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L4_U1 ( .a ({new_AGEMA_signal_6709, SubBytesIns_Inst_Sbox_12_M54}), .b ({new_AGEMA_signal_6711, SubBytesIns_Inst_Sbox_12_M58}), .c ({new_AGEMA_signal_6917, SubBytesIns_Inst_Sbox_12_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L5_U1 ( .a ({new_AGEMA_signal_6707, SubBytesIns_Inst_Sbox_12_M49}), .b ({new_AGEMA_signal_6712, SubBytesIns_Inst_Sbox_12_M61}), .c ({new_AGEMA_signal_6918, SubBytesIns_Inst_Sbox_12_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L6_U1 ( .a ({new_AGEMA_signal_6914, SubBytesIns_Inst_Sbox_12_M62}), .b ({new_AGEMA_signal_6918, SubBytesIns_Inst_Sbox_12_L5}), .c ({new_AGEMA_signal_7098, SubBytesIns_Inst_Sbox_12_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L7_U1 ( .a ({new_AGEMA_signal_6706, SubBytesIns_Inst_Sbox_12_M46}), .b ({new_AGEMA_signal_6916, SubBytesIns_Inst_Sbox_12_L3}), .c ({new_AGEMA_signal_7099, SubBytesIns_Inst_Sbox_12_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L8_U1 ( .a ({new_AGEMA_signal_6472, SubBytesIns_Inst_Sbox_12_M51}), .b ({new_AGEMA_signal_6475, SubBytesIns_Inst_Sbox_12_M59}), .c ({new_AGEMA_signal_6715, SubBytesIns_Inst_Sbox_12_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L9_U1 ( .a ({new_AGEMA_signal_6708, SubBytesIns_Inst_Sbox_12_M52}), .b ({new_AGEMA_signal_6913, SubBytesIns_Inst_Sbox_12_M53}), .c ({new_AGEMA_signal_7100, SubBytesIns_Inst_Sbox_12_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L10_U1 ( .a ({new_AGEMA_signal_6913, SubBytesIns_Inst_Sbox_12_M53}), .b ({new_AGEMA_signal_6917, SubBytesIns_Inst_Sbox_12_L4}), .c ({new_AGEMA_signal_7101, SubBytesIns_Inst_Sbox_12_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L11_U1 ( .a ({new_AGEMA_signal_6476, SubBytesIns_Inst_Sbox_12_M60}), .b ({new_AGEMA_signal_6915, SubBytesIns_Inst_Sbox_12_L2}), .c ({new_AGEMA_signal_7102, SubBytesIns_Inst_Sbox_12_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L12_U1 ( .a ({new_AGEMA_signal_6470, SubBytesIns_Inst_Sbox_12_M48}), .b ({new_AGEMA_signal_6472, SubBytesIns_Inst_Sbox_12_M51}), .c ({new_AGEMA_signal_6716, SubBytesIns_Inst_Sbox_12_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L13_U1 ( .a ({new_AGEMA_signal_6471, SubBytesIns_Inst_Sbox_12_M50}), .b ({new_AGEMA_signal_7097, SubBytesIns_Inst_Sbox_12_L0}), .c ({new_AGEMA_signal_7309, SubBytesIns_Inst_Sbox_12_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L14_U1 ( .a ({new_AGEMA_signal_6708, SubBytesIns_Inst_Sbox_12_M52}), .b ({new_AGEMA_signal_6712, SubBytesIns_Inst_Sbox_12_M61}), .c ({new_AGEMA_signal_6919, SubBytesIns_Inst_Sbox_12_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L15_U1 ( .a ({new_AGEMA_signal_6710, SubBytesIns_Inst_Sbox_12_M55}), .b ({new_AGEMA_signal_6714, SubBytesIns_Inst_Sbox_12_L1}), .c ({new_AGEMA_signal_6920, SubBytesIns_Inst_Sbox_12_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L16_U1 ( .a ({new_AGEMA_signal_6473, SubBytesIns_Inst_Sbox_12_M56}), .b ({new_AGEMA_signal_7097, SubBytesIns_Inst_Sbox_12_L0}), .c ({new_AGEMA_signal_7310, SubBytesIns_Inst_Sbox_12_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L17_U1 ( .a ({new_AGEMA_signal_6474, SubBytesIns_Inst_Sbox_12_M57}), .b ({new_AGEMA_signal_6714, SubBytesIns_Inst_Sbox_12_L1}), .c ({new_AGEMA_signal_6921, SubBytesIns_Inst_Sbox_12_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L18_U1 ( .a ({new_AGEMA_signal_6711, SubBytesIns_Inst_Sbox_12_M58}), .b ({new_AGEMA_signal_6715, SubBytesIns_Inst_Sbox_12_L8}), .c ({new_AGEMA_signal_6922, SubBytesIns_Inst_Sbox_12_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L19_U1 ( .a ({new_AGEMA_signal_6713, SubBytesIns_Inst_Sbox_12_M63}), .b ({new_AGEMA_signal_6917, SubBytesIns_Inst_Sbox_12_L4}), .c ({new_AGEMA_signal_7103, SubBytesIns_Inst_Sbox_12_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L20_U1 ( .a ({new_AGEMA_signal_7097, SubBytesIns_Inst_Sbox_12_L0}), .b ({new_AGEMA_signal_6714, SubBytesIns_Inst_Sbox_12_L1}), .c ({new_AGEMA_signal_7311, SubBytesIns_Inst_Sbox_12_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L21_U1 ( .a ({new_AGEMA_signal_6714, SubBytesIns_Inst_Sbox_12_L1}), .b ({new_AGEMA_signal_7099, SubBytesIns_Inst_Sbox_12_L7}), .c ({new_AGEMA_signal_7312, SubBytesIns_Inst_Sbox_12_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L22_U1 ( .a ({new_AGEMA_signal_6916, SubBytesIns_Inst_Sbox_12_L3}), .b ({new_AGEMA_signal_6716, SubBytesIns_Inst_Sbox_12_L12}), .c ({new_AGEMA_signal_7104, SubBytesIns_Inst_Sbox_12_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L23_U1 ( .a ({new_AGEMA_signal_6922, SubBytesIns_Inst_Sbox_12_L18}), .b ({new_AGEMA_signal_6915, SubBytesIns_Inst_Sbox_12_L2}), .c ({new_AGEMA_signal_7105, SubBytesIns_Inst_Sbox_12_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L24_U1 ( .a ({new_AGEMA_signal_6920, SubBytesIns_Inst_Sbox_12_L15}), .b ({new_AGEMA_signal_7100, SubBytesIns_Inst_Sbox_12_L9}), .c ({new_AGEMA_signal_7313, SubBytesIns_Inst_Sbox_12_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L25_U1 ( .a ({new_AGEMA_signal_7098, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_7101, SubBytesIns_Inst_Sbox_12_L10}), .c ({new_AGEMA_signal_7314, SubBytesIns_Inst_Sbox_12_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L26_U1 ( .a ({new_AGEMA_signal_7099, SubBytesIns_Inst_Sbox_12_L7}), .b ({new_AGEMA_signal_7100, SubBytesIns_Inst_Sbox_12_L9}), .c ({new_AGEMA_signal_7315, SubBytesIns_Inst_Sbox_12_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L27_U1 ( .a ({new_AGEMA_signal_6715, SubBytesIns_Inst_Sbox_12_L8}), .b ({new_AGEMA_signal_7101, SubBytesIns_Inst_Sbox_12_L10}), .c ({new_AGEMA_signal_7316, SubBytesIns_Inst_Sbox_12_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L28_U1 ( .a ({new_AGEMA_signal_7102, SubBytesIns_Inst_Sbox_12_L11}), .b ({new_AGEMA_signal_6919, SubBytesIns_Inst_Sbox_12_L14}), .c ({new_AGEMA_signal_7317, SubBytesIns_Inst_Sbox_12_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L29_U1 ( .a ({new_AGEMA_signal_7102, SubBytesIns_Inst_Sbox_12_L11}), .b ({new_AGEMA_signal_6921, SubBytesIns_Inst_Sbox_12_L17}), .c ({new_AGEMA_signal_7318, SubBytesIns_Inst_Sbox_12_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S0_U1 ( .a ({new_AGEMA_signal_7098, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_7313, SubBytesIns_Inst_Sbox_12_L24}), .c ({new_AGEMA_signal_7469, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S1_U1 ( .a ({new_AGEMA_signal_7310, SubBytesIns_Inst_Sbox_12_L16}), .b ({new_AGEMA_signal_7315, SubBytesIns_Inst_Sbox_12_L26}), .c ({new_AGEMA_signal_7470, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S2_U1 ( .a ({new_AGEMA_signal_7103, SubBytesIns_Inst_Sbox_12_L19}), .b ({new_AGEMA_signal_7317, SubBytesIns_Inst_Sbox_12_L28}), .c ({new_AGEMA_signal_7471, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S3_U1 ( .a ({new_AGEMA_signal_7098, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_7312, SubBytesIns_Inst_Sbox_12_L21}), .c ({new_AGEMA_signal_7472, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S4_U1 ( .a ({new_AGEMA_signal_7311, SubBytesIns_Inst_Sbox_12_L20}), .b ({new_AGEMA_signal_7104, SubBytesIns_Inst_Sbox_12_L22}), .c ({new_AGEMA_signal_7473, MixColumnsInput[67]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S5_U1 ( .a ({new_AGEMA_signal_7314, SubBytesIns_Inst_Sbox_12_L25}), .b ({new_AGEMA_signal_7318, SubBytesIns_Inst_Sbox_12_L29}), .c ({new_AGEMA_signal_7474, MixColumnsInput[66]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S6_U1 ( .a ({new_AGEMA_signal_7309, SubBytesIns_Inst_Sbox_12_L13}), .b ({new_AGEMA_signal_7316, SubBytesIns_Inst_Sbox_12_L27}), .c ({new_AGEMA_signal_7475, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S7_U1 ( .a ({new_AGEMA_signal_7098, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_7105, SubBytesIns_Inst_Sbox_12_L23}), .c ({new_AGEMA_signal_7319, MixColumnsInput[64]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M46_U1 ( .a ({new_AGEMA_signal_6480, SubBytesIns_Inst_Sbox_13_M44}), .b ({new_AGEMA_signal_5269, SubBytesIns_Inst_Sbox_13_T6}), .clk (clk), .r (Fresh[554]), .c ({new_AGEMA_signal_6718, SubBytesIns_Inst_Sbox_13_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M47_U1 ( .a ({new_AGEMA_signal_6264, SubBytesIns_Inst_Sbox_13_M40}), .b ({new_AGEMA_signal_5514, SubBytesIns_Inst_Sbox_13_T8}), .clk (clk), .r (Fresh[555]), .c ({new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_13_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M48_U1 ( .a ({new_AGEMA_signal_6263, SubBytesIns_Inst_Sbox_13_M39}), .b ({ciphertext_s1[104], ciphertext_s0[104]}), .clk (clk), .r (Fresh[556]), .c ({new_AGEMA_signal_6482, SubBytesIns_Inst_Sbox_13_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M49_U1 ( .a ({new_AGEMA_signal_6479, SubBytesIns_Inst_Sbox_13_M43}), .b ({new_AGEMA_signal_5273, SubBytesIns_Inst_Sbox_13_T16}), .clk (clk), .r (Fresh[557]), .c ({new_AGEMA_signal_6719, SubBytesIns_Inst_Sbox_13_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M50_U1 ( .a ({new_AGEMA_signal_6262, SubBytesIns_Inst_Sbox_13_M38}), .b ({new_AGEMA_signal_5270, SubBytesIns_Inst_Sbox_13_T9}), .clk (clk), .r (Fresh[558]), .c ({new_AGEMA_signal_6483, SubBytesIns_Inst_Sbox_13_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M51_U1 ( .a ({new_AGEMA_signal_6261, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_5517, SubBytesIns_Inst_Sbox_13_T17}), .clk (clk), .r (Fresh[559]), .c ({new_AGEMA_signal_6484, SubBytesIns_Inst_Sbox_13_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M52_U1 ( .a ({new_AGEMA_signal_6478, SubBytesIns_Inst_Sbox_13_M42}), .b ({new_AGEMA_signal_5272, SubBytesIns_Inst_Sbox_13_T15}), .clk (clk), .r (Fresh[560]), .c ({new_AGEMA_signal_6720, SubBytesIns_Inst_Sbox_13_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M53_U1 ( .a ({new_AGEMA_signal_6717, SubBytesIns_Inst_Sbox_13_M45}), .b ({new_AGEMA_signal_5276, SubBytesIns_Inst_Sbox_13_T27}), .clk (clk), .r (Fresh[561]), .c ({new_AGEMA_signal_6923, SubBytesIns_Inst_Sbox_13_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M54_U1 ( .a ({new_AGEMA_signal_6477, SubBytesIns_Inst_Sbox_13_M41}), .b ({new_AGEMA_signal_5515, SubBytesIns_Inst_Sbox_13_T10}), .clk (clk), .r (Fresh[562]), .c ({new_AGEMA_signal_6721, SubBytesIns_Inst_Sbox_13_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M55_U1 ( .a ({new_AGEMA_signal_6480, SubBytesIns_Inst_Sbox_13_M44}), .b ({new_AGEMA_signal_5271, SubBytesIns_Inst_Sbox_13_T13}), .clk (clk), .r (Fresh[563]), .c ({new_AGEMA_signal_6722, SubBytesIns_Inst_Sbox_13_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M56_U1 ( .a ({new_AGEMA_signal_6264, SubBytesIns_Inst_Sbox_13_M40}), .b ({new_AGEMA_signal_5519, SubBytesIns_Inst_Sbox_13_T23}), .clk (clk), .r (Fresh[564]), .c ({new_AGEMA_signal_6485, SubBytesIns_Inst_Sbox_13_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M57_U1 ( .a ({new_AGEMA_signal_6263, SubBytesIns_Inst_Sbox_13_M39}), .b ({new_AGEMA_signal_5274, SubBytesIns_Inst_Sbox_13_T19}), .clk (clk), .r (Fresh[565]), .c ({new_AGEMA_signal_6486, SubBytesIns_Inst_Sbox_13_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M58_U1 ( .a ({new_AGEMA_signal_6479, SubBytesIns_Inst_Sbox_13_M43}), .b ({new_AGEMA_signal_5105, SubBytesIns_Inst_Sbox_13_T3}), .clk (clk), .r (Fresh[566]), .c ({new_AGEMA_signal_6723, SubBytesIns_Inst_Sbox_13_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M59_U1 ( .a ({new_AGEMA_signal_6262, SubBytesIns_Inst_Sbox_13_M38}), .b ({new_AGEMA_signal_5275, SubBytesIns_Inst_Sbox_13_T22}), .clk (clk), .r (Fresh[567]), .c ({new_AGEMA_signal_6487, SubBytesIns_Inst_Sbox_13_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M60_U1 ( .a ({new_AGEMA_signal_6261, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_5518, SubBytesIns_Inst_Sbox_13_T20}), .clk (clk), .r (Fresh[568]), .c ({new_AGEMA_signal_6488, SubBytesIns_Inst_Sbox_13_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M61_U1 ( .a ({new_AGEMA_signal_6478, SubBytesIns_Inst_Sbox_13_M42}), .b ({new_AGEMA_signal_5103, SubBytesIns_Inst_Sbox_13_T1}), .clk (clk), .r (Fresh[569]), .c ({new_AGEMA_signal_6724, SubBytesIns_Inst_Sbox_13_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M62_U1 ( .a ({new_AGEMA_signal_6717, SubBytesIns_Inst_Sbox_13_M45}), .b ({new_AGEMA_signal_5106, SubBytesIns_Inst_Sbox_13_T4}), .clk (clk), .r (Fresh[570]), .c ({new_AGEMA_signal_6924, SubBytesIns_Inst_Sbox_13_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M63_U1 ( .a ({new_AGEMA_signal_6477, SubBytesIns_Inst_Sbox_13_M41}), .b ({new_AGEMA_signal_5104, SubBytesIns_Inst_Sbox_13_T2}), .clk (clk), .r (Fresh[571]), .c ({new_AGEMA_signal_6725, SubBytesIns_Inst_Sbox_13_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L0_U1 ( .a ({new_AGEMA_signal_6724, SubBytesIns_Inst_Sbox_13_M61}), .b ({new_AGEMA_signal_6924, SubBytesIns_Inst_Sbox_13_M62}), .c ({new_AGEMA_signal_7106, SubBytesIns_Inst_Sbox_13_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L1_U1 ( .a ({new_AGEMA_signal_6483, SubBytesIns_Inst_Sbox_13_M50}), .b ({new_AGEMA_signal_6485, SubBytesIns_Inst_Sbox_13_M56}), .c ({new_AGEMA_signal_6726, SubBytesIns_Inst_Sbox_13_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L2_U1 ( .a ({new_AGEMA_signal_6718, SubBytesIns_Inst_Sbox_13_M46}), .b ({new_AGEMA_signal_6482, SubBytesIns_Inst_Sbox_13_M48}), .c ({new_AGEMA_signal_6925, SubBytesIns_Inst_Sbox_13_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L3_U1 ( .a ({new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_13_M47}), .b ({new_AGEMA_signal_6722, SubBytesIns_Inst_Sbox_13_M55}), .c ({new_AGEMA_signal_6926, SubBytesIns_Inst_Sbox_13_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L4_U1 ( .a ({new_AGEMA_signal_6721, SubBytesIns_Inst_Sbox_13_M54}), .b ({new_AGEMA_signal_6723, SubBytesIns_Inst_Sbox_13_M58}), .c ({new_AGEMA_signal_6927, SubBytesIns_Inst_Sbox_13_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L5_U1 ( .a ({new_AGEMA_signal_6719, SubBytesIns_Inst_Sbox_13_M49}), .b ({new_AGEMA_signal_6724, SubBytesIns_Inst_Sbox_13_M61}), .c ({new_AGEMA_signal_6928, SubBytesIns_Inst_Sbox_13_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L6_U1 ( .a ({new_AGEMA_signal_6924, SubBytesIns_Inst_Sbox_13_M62}), .b ({new_AGEMA_signal_6928, SubBytesIns_Inst_Sbox_13_L5}), .c ({new_AGEMA_signal_7107, SubBytesIns_Inst_Sbox_13_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L7_U1 ( .a ({new_AGEMA_signal_6718, SubBytesIns_Inst_Sbox_13_M46}), .b ({new_AGEMA_signal_6926, SubBytesIns_Inst_Sbox_13_L3}), .c ({new_AGEMA_signal_7108, SubBytesIns_Inst_Sbox_13_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L8_U1 ( .a ({new_AGEMA_signal_6484, SubBytesIns_Inst_Sbox_13_M51}), .b ({new_AGEMA_signal_6487, SubBytesIns_Inst_Sbox_13_M59}), .c ({new_AGEMA_signal_6727, SubBytesIns_Inst_Sbox_13_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L9_U1 ( .a ({new_AGEMA_signal_6720, SubBytesIns_Inst_Sbox_13_M52}), .b ({new_AGEMA_signal_6923, SubBytesIns_Inst_Sbox_13_M53}), .c ({new_AGEMA_signal_7109, SubBytesIns_Inst_Sbox_13_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L10_U1 ( .a ({new_AGEMA_signal_6923, SubBytesIns_Inst_Sbox_13_M53}), .b ({new_AGEMA_signal_6927, SubBytesIns_Inst_Sbox_13_L4}), .c ({new_AGEMA_signal_7110, SubBytesIns_Inst_Sbox_13_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L11_U1 ( .a ({new_AGEMA_signal_6488, SubBytesIns_Inst_Sbox_13_M60}), .b ({new_AGEMA_signal_6925, SubBytesIns_Inst_Sbox_13_L2}), .c ({new_AGEMA_signal_7111, SubBytesIns_Inst_Sbox_13_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L12_U1 ( .a ({new_AGEMA_signal_6482, SubBytesIns_Inst_Sbox_13_M48}), .b ({new_AGEMA_signal_6484, SubBytesIns_Inst_Sbox_13_M51}), .c ({new_AGEMA_signal_6728, SubBytesIns_Inst_Sbox_13_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L13_U1 ( .a ({new_AGEMA_signal_6483, SubBytesIns_Inst_Sbox_13_M50}), .b ({new_AGEMA_signal_7106, SubBytesIns_Inst_Sbox_13_L0}), .c ({new_AGEMA_signal_7320, SubBytesIns_Inst_Sbox_13_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L14_U1 ( .a ({new_AGEMA_signal_6720, SubBytesIns_Inst_Sbox_13_M52}), .b ({new_AGEMA_signal_6724, SubBytesIns_Inst_Sbox_13_M61}), .c ({new_AGEMA_signal_6929, SubBytesIns_Inst_Sbox_13_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L15_U1 ( .a ({new_AGEMA_signal_6722, SubBytesIns_Inst_Sbox_13_M55}), .b ({new_AGEMA_signal_6726, SubBytesIns_Inst_Sbox_13_L1}), .c ({new_AGEMA_signal_6930, SubBytesIns_Inst_Sbox_13_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L16_U1 ( .a ({new_AGEMA_signal_6485, SubBytesIns_Inst_Sbox_13_M56}), .b ({new_AGEMA_signal_7106, SubBytesIns_Inst_Sbox_13_L0}), .c ({new_AGEMA_signal_7321, SubBytesIns_Inst_Sbox_13_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L17_U1 ( .a ({new_AGEMA_signal_6486, SubBytesIns_Inst_Sbox_13_M57}), .b ({new_AGEMA_signal_6726, SubBytesIns_Inst_Sbox_13_L1}), .c ({new_AGEMA_signal_6931, SubBytesIns_Inst_Sbox_13_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L18_U1 ( .a ({new_AGEMA_signal_6723, SubBytesIns_Inst_Sbox_13_M58}), .b ({new_AGEMA_signal_6727, SubBytesIns_Inst_Sbox_13_L8}), .c ({new_AGEMA_signal_6932, SubBytesIns_Inst_Sbox_13_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L19_U1 ( .a ({new_AGEMA_signal_6725, SubBytesIns_Inst_Sbox_13_M63}), .b ({new_AGEMA_signal_6927, SubBytesIns_Inst_Sbox_13_L4}), .c ({new_AGEMA_signal_7112, SubBytesIns_Inst_Sbox_13_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L20_U1 ( .a ({new_AGEMA_signal_7106, SubBytesIns_Inst_Sbox_13_L0}), .b ({new_AGEMA_signal_6726, SubBytesIns_Inst_Sbox_13_L1}), .c ({new_AGEMA_signal_7322, SubBytesIns_Inst_Sbox_13_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L21_U1 ( .a ({new_AGEMA_signal_6726, SubBytesIns_Inst_Sbox_13_L1}), .b ({new_AGEMA_signal_7108, SubBytesIns_Inst_Sbox_13_L7}), .c ({new_AGEMA_signal_7323, SubBytesIns_Inst_Sbox_13_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L22_U1 ( .a ({new_AGEMA_signal_6926, SubBytesIns_Inst_Sbox_13_L3}), .b ({new_AGEMA_signal_6728, SubBytesIns_Inst_Sbox_13_L12}), .c ({new_AGEMA_signal_7113, SubBytesIns_Inst_Sbox_13_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L23_U1 ( .a ({new_AGEMA_signal_6932, SubBytesIns_Inst_Sbox_13_L18}), .b ({new_AGEMA_signal_6925, SubBytesIns_Inst_Sbox_13_L2}), .c ({new_AGEMA_signal_7114, SubBytesIns_Inst_Sbox_13_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L24_U1 ( .a ({new_AGEMA_signal_6930, SubBytesIns_Inst_Sbox_13_L15}), .b ({new_AGEMA_signal_7109, SubBytesIns_Inst_Sbox_13_L9}), .c ({new_AGEMA_signal_7324, SubBytesIns_Inst_Sbox_13_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L25_U1 ( .a ({new_AGEMA_signal_7107, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_7110, SubBytesIns_Inst_Sbox_13_L10}), .c ({new_AGEMA_signal_7325, SubBytesIns_Inst_Sbox_13_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L26_U1 ( .a ({new_AGEMA_signal_7108, SubBytesIns_Inst_Sbox_13_L7}), .b ({new_AGEMA_signal_7109, SubBytesIns_Inst_Sbox_13_L9}), .c ({new_AGEMA_signal_7326, SubBytesIns_Inst_Sbox_13_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L27_U1 ( .a ({new_AGEMA_signal_6727, SubBytesIns_Inst_Sbox_13_L8}), .b ({new_AGEMA_signal_7110, SubBytesIns_Inst_Sbox_13_L10}), .c ({new_AGEMA_signal_7327, SubBytesIns_Inst_Sbox_13_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L28_U1 ( .a ({new_AGEMA_signal_7111, SubBytesIns_Inst_Sbox_13_L11}), .b ({new_AGEMA_signal_6929, SubBytesIns_Inst_Sbox_13_L14}), .c ({new_AGEMA_signal_7328, SubBytesIns_Inst_Sbox_13_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L29_U1 ( .a ({new_AGEMA_signal_7111, SubBytesIns_Inst_Sbox_13_L11}), .b ({new_AGEMA_signal_6931, SubBytesIns_Inst_Sbox_13_L17}), .c ({new_AGEMA_signal_7329, SubBytesIns_Inst_Sbox_13_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S0_U1 ( .a ({new_AGEMA_signal_7107, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_7324, SubBytesIns_Inst_Sbox_13_L24}), .c ({new_AGEMA_signal_7476, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S1_U1 ( .a ({new_AGEMA_signal_7321, SubBytesIns_Inst_Sbox_13_L16}), .b ({new_AGEMA_signal_7326, SubBytesIns_Inst_Sbox_13_L26}), .c ({new_AGEMA_signal_7477, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S2_U1 ( .a ({new_AGEMA_signal_7112, SubBytesIns_Inst_Sbox_13_L19}), .b ({new_AGEMA_signal_7328, SubBytesIns_Inst_Sbox_13_L28}), .c ({new_AGEMA_signal_7478, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S3_U1 ( .a ({new_AGEMA_signal_7107, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_7323, SubBytesIns_Inst_Sbox_13_L21}), .c ({new_AGEMA_signal_7479, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S4_U1 ( .a ({new_AGEMA_signal_7322, SubBytesIns_Inst_Sbox_13_L20}), .b ({new_AGEMA_signal_7113, SubBytesIns_Inst_Sbox_13_L22}), .c ({new_AGEMA_signal_7480, MixColumnsInput[43]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S5_U1 ( .a ({new_AGEMA_signal_7325, SubBytesIns_Inst_Sbox_13_L25}), .b ({new_AGEMA_signal_7329, SubBytesIns_Inst_Sbox_13_L29}), .c ({new_AGEMA_signal_7481, MixColumnsInput[42]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S6_U1 ( .a ({new_AGEMA_signal_7320, SubBytesIns_Inst_Sbox_13_L13}), .b ({new_AGEMA_signal_7327, SubBytesIns_Inst_Sbox_13_L27}), .c ({new_AGEMA_signal_7482, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S7_U1 ( .a ({new_AGEMA_signal_7107, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_7114, SubBytesIns_Inst_Sbox_13_L23}), .c ({new_AGEMA_signal_7330, MixColumnsInput[40]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M46_U1 ( .a ({new_AGEMA_signal_6492, SubBytesIns_Inst_Sbox_14_M44}), .b ({new_AGEMA_signal_5277, SubBytesIns_Inst_Sbox_14_T6}), .clk (clk), .r (Fresh[572]), .c ({new_AGEMA_signal_6730, SubBytesIns_Inst_Sbox_14_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M47_U1 ( .a ({new_AGEMA_signal_6268, SubBytesIns_Inst_Sbox_14_M40}), .b ({new_AGEMA_signal_5527, SubBytesIns_Inst_Sbox_14_T8}), .clk (clk), .r (Fresh[573]), .c ({new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_14_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M48_U1 ( .a ({new_AGEMA_signal_6267, SubBytesIns_Inst_Sbox_14_M39}), .b ({ciphertext_s1[112], ciphertext_s0[112]}), .clk (clk), .r (Fresh[574]), .c ({new_AGEMA_signal_6494, SubBytesIns_Inst_Sbox_14_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M49_U1 ( .a ({new_AGEMA_signal_6491, SubBytesIns_Inst_Sbox_14_M43}), .b ({new_AGEMA_signal_5281, SubBytesIns_Inst_Sbox_14_T16}), .clk (clk), .r (Fresh[575]), .c ({new_AGEMA_signal_6731, SubBytesIns_Inst_Sbox_14_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M50_U1 ( .a ({new_AGEMA_signal_6266, SubBytesIns_Inst_Sbox_14_M38}), .b ({new_AGEMA_signal_5278, SubBytesIns_Inst_Sbox_14_T9}), .clk (clk), .r (Fresh[576]), .c ({new_AGEMA_signal_6495, SubBytesIns_Inst_Sbox_14_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M51_U1 ( .a ({new_AGEMA_signal_6265, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_5530, SubBytesIns_Inst_Sbox_14_T17}), .clk (clk), .r (Fresh[577]), .c ({new_AGEMA_signal_6496, SubBytesIns_Inst_Sbox_14_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M52_U1 ( .a ({new_AGEMA_signal_6490, SubBytesIns_Inst_Sbox_14_M42}), .b ({new_AGEMA_signal_5280, SubBytesIns_Inst_Sbox_14_T15}), .clk (clk), .r (Fresh[578]), .c ({new_AGEMA_signal_6732, SubBytesIns_Inst_Sbox_14_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M53_U1 ( .a ({new_AGEMA_signal_6729, SubBytesIns_Inst_Sbox_14_M45}), .b ({new_AGEMA_signal_5284, SubBytesIns_Inst_Sbox_14_T27}), .clk (clk), .r (Fresh[579]), .c ({new_AGEMA_signal_6933, SubBytesIns_Inst_Sbox_14_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M54_U1 ( .a ({new_AGEMA_signal_6489, SubBytesIns_Inst_Sbox_14_M41}), .b ({new_AGEMA_signal_5528, SubBytesIns_Inst_Sbox_14_T10}), .clk (clk), .r (Fresh[580]), .c ({new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_14_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M55_U1 ( .a ({new_AGEMA_signal_6492, SubBytesIns_Inst_Sbox_14_M44}), .b ({new_AGEMA_signal_5279, SubBytesIns_Inst_Sbox_14_T13}), .clk (clk), .r (Fresh[581]), .c ({new_AGEMA_signal_6734, SubBytesIns_Inst_Sbox_14_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M56_U1 ( .a ({new_AGEMA_signal_6268, SubBytesIns_Inst_Sbox_14_M40}), .b ({new_AGEMA_signal_5532, SubBytesIns_Inst_Sbox_14_T23}), .clk (clk), .r (Fresh[582]), .c ({new_AGEMA_signal_6497, SubBytesIns_Inst_Sbox_14_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M57_U1 ( .a ({new_AGEMA_signal_6267, SubBytesIns_Inst_Sbox_14_M39}), .b ({new_AGEMA_signal_5282, SubBytesIns_Inst_Sbox_14_T19}), .clk (clk), .r (Fresh[583]), .c ({new_AGEMA_signal_6498, SubBytesIns_Inst_Sbox_14_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M58_U1 ( .a ({new_AGEMA_signal_6491, SubBytesIns_Inst_Sbox_14_M43}), .b ({new_AGEMA_signal_5115, SubBytesIns_Inst_Sbox_14_T3}), .clk (clk), .r (Fresh[584]), .c ({new_AGEMA_signal_6735, SubBytesIns_Inst_Sbox_14_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M59_U1 ( .a ({new_AGEMA_signal_6266, SubBytesIns_Inst_Sbox_14_M38}), .b ({new_AGEMA_signal_5283, SubBytesIns_Inst_Sbox_14_T22}), .clk (clk), .r (Fresh[585]), .c ({new_AGEMA_signal_6499, SubBytesIns_Inst_Sbox_14_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M60_U1 ( .a ({new_AGEMA_signal_6265, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_5531, SubBytesIns_Inst_Sbox_14_T20}), .clk (clk), .r (Fresh[586]), .c ({new_AGEMA_signal_6500, SubBytesIns_Inst_Sbox_14_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M61_U1 ( .a ({new_AGEMA_signal_6490, SubBytesIns_Inst_Sbox_14_M42}), .b ({new_AGEMA_signal_5113, SubBytesIns_Inst_Sbox_14_T1}), .clk (clk), .r (Fresh[587]), .c ({new_AGEMA_signal_6736, SubBytesIns_Inst_Sbox_14_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M62_U1 ( .a ({new_AGEMA_signal_6729, SubBytesIns_Inst_Sbox_14_M45}), .b ({new_AGEMA_signal_5116, SubBytesIns_Inst_Sbox_14_T4}), .clk (clk), .r (Fresh[588]), .c ({new_AGEMA_signal_6934, SubBytesIns_Inst_Sbox_14_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M63_U1 ( .a ({new_AGEMA_signal_6489, SubBytesIns_Inst_Sbox_14_M41}), .b ({new_AGEMA_signal_5114, SubBytesIns_Inst_Sbox_14_T2}), .clk (clk), .r (Fresh[589]), .c ({new_AGEMA_signal_6737, SubBytesIns_Inst_Sbox_14_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L0_U1 ( .a ({new_AGEMA_signal_6736, SubBytesIns_Inst_Sbox_14_M61}), .b ({new_AGEMA_signal_6934, SubBytesIns_Inst_Sbox_14_M62}), .c ({new_AGEMA_signal_7115, SubBytesIns_Inst_Sbox_14_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L1_U1 ( .a ({new_AGEMA_signal_6495, SubBytesIns_Inst_Sbox_14_M50}), .b ({new_AGEMA_signal_6497, SubBytesIns_Inst_Sbox_14_M56}), .c ({new_AGEMA_signal_6738, SubBytesIns_Inst_Sbox_14_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L2_U1 ( .a ({new_AGEMA_signal_6730, SubBytesIns_Inst_Sbox_14_M46}), .b ({new_AGEMA_signal_6494, SubBytesIns_Inst_Sbox_14_M48}), .c ({new_AGEMA_signal_6935, SubBytesIns_Inst_Sbox_14_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L3_U1 ( .a ({new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_14_M47}), .b ({new_AGEMA_signal_6734, SubBytesIns_Inst_Sbox_14_M55}), .c ({new_AGEMA_signal_6936, SubBytesIns_Inst_Sbox_14_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L4_U1 ( .a ({new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_14_M54}), .b ({new_AGEMA_signal_6735, SubBytesIns_Inst_Sbox_14_M58}), .c ({new_AGEMA_signal_6937, SubBytesIns_Inst_Sbox_14_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L5_U1 ( .a ({new_AGEMA_signal_6731, SubBytesIns_Inst_Sbox_14_M49}), .b ({new_AGEMA_signal_6736, SubBytesIns_Inst_Sbox_14_M61}), .c ({new_AGEMA_signal_6938, SubBytesIns_Inst_Sbox_14_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L6_U1 ( .a ({new_AGEMA_signal_6934, SubBytesIns_Inst_Sbox_14_M62}), .b ({new_AGEMA_signal_6938, SubBytesIns_Inst_Sbox_14_L5}), .c ({new_AGEMA_signal_7116, SubBytesIns_Inst_Sbox_14_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L7_U1 ( .a ({new_AGEMA_signal_6730, SubBytesIns_Inst_Sbox_14_M46}), .b ({new_AGEMA_signal_6936, SubBytesIns_Inst_Sbox_14_L3}), .c ({new_AGEMA_signal_7117, SubBytesIns_Inst_Sbox_14_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L8_U1 ( .a ({new_AGEMA_signal_6496, SubBytesIns_Inst_Sbox_14_M51}), .b ({new_AGEMA_signal_6499, SubBytesIns_Inst_Sbox_14_M59}), .c ({new_AGEMA_signal_6739, SubBytesIns_Inst_Sbox_14_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L9_U1 ( .a ({new_AGEMA_signal_6732, SubBytesIns_Inst_Sbox_14_M52}), .b ({new_AGEMA_signal_6933, SubBytesIns_Inst_Sbox_14_M53}), .c ({new_AGEMA_signal_7118, SubBytesIns_Inst_Sbox_14_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L10_U1 ( .a ({new_AGEMA_signal_6933, SubBytesIns_Inst_Sbox_14_M53}), .b ({new_AGEMA_signal_6937, SubBytesIns_Inst_Sbox_14_L4}), .c ({new_AGEMA_signal_7119, SubBytesIns_Inst_Sbox_14_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L11_U1 ( .a ({new_AGEMA_signal_6500, SubBytesIns_Inst_Sbox_14_M60}), .b ({new_AGEMA_signal_6935, SubBytesIns_Inst_Sbox_14_L2}), .c ({new_AGEMA_signal_7120, SubBytesIns_Inst_Sbox_14_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L12_U1 ( .a ({new_AGEMA_signal_6494, SubBytesIns_Inst_Sbox_14_M48}), .b ({new_AGEMA_signal_6496, SubBytesIns_Inst_Sbox_14_M51}), .c ({new_AGEMA_signal_6740, SubBytesIns_Inst_Sbox_14_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L13_U1 ( .a ({new_AGEMA_signal_6495, SubBytesIns_Inst_Sbox_14_M50}), .b ({new_AGEMA_signal_7115, SubBytesIns_Inst_Sbox_14_L0}), .c ({new_AGEMA_signal_7331, SubBytesIns_Inst_Sbox_14_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L14_U1 ( .a ({new_AGEMA_signal_6732, SubBytesIns_Inst_Sbox_14_M52}), .b ({new_AGEMA_signal_6736, SubBytesIns_Inst_Sbox_14_M61}), .c ({new_AGEMA_signal_6939, SubBytesIns_Inst_Sbox_14_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L15_U1 ( .a ({new_AGEMA_signal_6734, SubBytesIns_Inst_Sbox_14_M55}), .b ({new_AGEMA_signal_6738, SubBytesIns_Inst_Sbox_14_L1}), .c ({new_AGEMA_signal_6940, SubBytesIns_Inst_Sbox_14_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L16_U1 ( .a ({new_AGEMA_signal_6497, SubBytesIns_Inst_Sbox_14_M56}), .b ({new_AGEMA_signal_7115, SubBytesIns_Inst_Sbox_14_L0}), .c ({new_AGEMA_signal_7332, SubBytesIns_Inst_Sbox_14_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L17_U1 ( .a ({new_AGEMA_signal_6498, SubBytesIns_Inst_Sbox_14_M57}), .b ({new_AGEMA_signal_6738, SubBytesIns_Inst_Sbox_14_L1}), .c ({new_AGEMA_signal_6941, SubBytesIns_Inst_Sbox_14_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L18_U1 ( .a ({new_AGEMA_signal_6735, SubBytesIns_Inst_Sbox_14_M58}), .b ({new_AGEMA_signal_6739, SubBytesIns_Inst_Sbox_14_L8}), .c ({new_AGEMA_signal_6942, SubBytesIns_Inst_Sbox_14_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L19_U1 ( .a ({new_AGEMA_signal_6737, SubBytesIns_Inst_Sbox_14_M63}), .b ({new_AGEMA_signal_6937, SubBytesIns_Inst_Sbox_14_L4}), .c ({new_AGEMA_signal_7121, SubBytesIns_Inst_Sbox_14_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L20_U1 ( .a ({new_AGEMA_signal_7115, SubBytesIns_Inst_Sbox_14_L0}), .b ({new_AGEMA_signal_6738, SubBytesIns_Inst_Sbox_14_L1}), .c ({new_AGEMA_signal_7333, SubBytesIns_Inst_Sbox_14_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L21_U1 ( .a ({new_AGEMA_signal_6738, SubBytesIns_Inst_Sbox_14_L1}), .b ({new_AGEMA_signal_7117, SubBytesIns_Inst_Sbox_14_L7}), .c ({new_AGEMA_signal_7334, SubBytesIns_Inst_Sbox_14_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L22_U1 ( .a ({new_AGEMA_signal_6936, SubBytesIns_Inst_Sbox_14_L3}), .b ({new_AGEMA_signal_6740, SubBytesIns_Inst_Sbox_14_L12}), .c ({new_AGEMA_signal_7122, SubBytesIns_Inst_Sbox_14_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L23_U1 ( .a ({new_AGEMA_signal_6942, SubBytesIns_Inst_Sbox_14_L18}), .b ({new_AGEMA_signal_6935, SubBytesIns_Inst_Sbox_14_L2}), .c ({new_AGEMA_signal_7123, SubBytesIns_Inst_Sbox_14_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L24_U1 ( .a ({new_AGEMA_signal_6940, SubBytesIns_Inst_Sbox_14_L15}), .b ({new_AGEMA_signal_7118, SubBytesIns_Inst_Sbox_14_L9}), .c ({new_AGEMA_signal_7335, SubBytesIns_Inst_Sbox_14_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L25_U1 ( .a ({new_AGEMA_signal_7116, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_7119, SubBytesIns_Inst_Sbox_14_L10}), .c ({new_AGEMA_signal_7336, SubBytesIns_Inst_Sbox_14_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L26_U1 ( .a ({new_AGEMA_signal_7117, SubBytesIns_Inst_Sbox_14_L7}), .b ({new_AGEMA_signal_7118, SubBytesIns_Inst_Sbox_14_L9}), .c ({new_AGEMA_signal_7337, SubBytesIns_Inst_Sbox_14_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L27_U1 ( .a ({new_AGEMA_signal_6739, SubBytesIns_Inst_Sbox_14_L8}), .b ({new_AGEMA_signal_7119, SubBytesIns_Inst_Sbox_14_L10}), .c ({new_AGEMA_signal_7338, SubBytesIns_Inst_Sbox_14_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L28_U1 ( .a ({new_AGEMA_signal_7120, SubBytesIns_Inst_Sbox_14_L11}), .b ({new_AGEMA_signal_6939, SubBytesIns_Inst_Sbox_14_L14}), .c ({new_AGEMA_signal_7339, SubBytesIns_Inst_Sbox_14_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L29_U1 ( .a ({new_AGEMA_signal_7120, SubBytesIns_Inst_Sbox_14_L11}), .b ({new_AGEMA_signal_6941, SubBytesIns_Inst_Sbox_14_L17}), .c ({new_AGEMA_signal_7340, SubBytesIns_Inst_Sbox_14_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S0_U1 ( .a ({new_AGEMA_signal_7116, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_7335, SubBytesIns_Inst_Sbox_14_L24}), .c ({new_AGEMA_signal_7483, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S1_U1 ( .a ({new_AGEMA_signal_7332, SubBytesIns_Inst_Sbox_14_L16}), .b ({new_AGEMA_signal_7337, SubBytesIns_Inst_Sbox_14_L26}), .c ({new_AGEMA_signal_7484, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S2_U1 ( .a ({new_AGEMA_signal_7121, SubBytesIns_Inst_Sbox_14_L19}), .b ({new_AGEMA_signal_7339, SubBytesIns_Inst_Sbox_14_L28}), .c ({new_AGEMA_signal_7485, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S3_U1 ( .a ({new_AGEMA_signal_7116, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_7334, SubBytesIns_Inst_Sbox_14_L21}), .c ({new_AGEMA_signal_7486, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S4_U1 ( .a ({new_AGEMA_signal_7333, SubBytesIns_Inst_Sbox_14_L20}), .b ({new_AGEMA_signal_7122, SubBytesIns_Inst_Sbox_14_L22}), .c ({new_AGEMA_signal_7487, MixColumnsInput[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S5_U1 ( .a ({new_AGEMA_signal_7336, SubBytesIns_Inst_Sbox_14_L25}), .b ({new_AGEMA_signal_7340, SubBytesIns_Inst_Sbox_14_L29}), .c ({new_AGEMA_signal_7488, MixColumnsInput[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S6_U1 ( .a ({new_AGEMA_signal_7331, SubBytesIns_Inst_Sbox_14_L13}), .b ({new_AGEMA_signal_7338, SubBytesIns_Inst_Sbox_14_L27}), .c ({new_AGEMA_signal_7489, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S7_U1 ( .a ({new_AGEMA_signal_7116, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_7123, SubBytesIns_Inst_Sbox_14_L23}), .c ({new_AGEMA_signal_7341, MixColumnsInput[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M46_U1 ( .a ({new_AGEMA_signal_6504, SubBytesIns_Inst_Sbox_15_M44}), .b ({new_AGEMA_signal_5285, SubBytesIns_Inst_Sbox_15_T6}), .clk (clk), .r (Fresh[590]), .c ({new_AGEMA_signal_6742, SubBytesIns_Inst_Sbox_15_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M47_U1 ( .a ({new_AGEMA_signal_6272, SubBytesIns_Inst_Sbox_15_M40}), .b ({new_AGEMA_signal_5540, SubBytesIns_Inst_Sbox_15_T8}), .clk (clk), .r (Fresh[591]), .c ({new_AGEMA_signal_6505, SubBytesIns_Inst_Sbox_15_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M48_U1 ( .a ({new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_M39}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .clk (clk), .r (Fresh[592]), .c ({new_AGEMA_signal_6506, SubBytesIns_Inst_Sbox_15_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M49_U1 ( .a ({new_AGEMA_signal_6503, SubBytesIns_Inst_Sbox_15_M43}), .b ({new_AGEMA_signal_5289, SubBytesIns_Inst_Sbox_15_T16}), .clk (clk), .r (Fresh[593]), .c ({new_AGEMA_signal_6743, SubBytesIns_Inst_Sbox_15_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M50_U1 ( .a ({new_AGEMA_signal_6270, SubBytesIns_Inst_Sbox_15_M38}), .b ({new_AGEMA_signal_5286, SubBytesIns_Inst_Sbox_15_T9}), .clk (clk), .r (Fresh[594]), .c ({new_AGEMA_signal_6507, SubBytesIns_Inst_Sbox_15_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M51_U1 ( .a ({new_AGEMA_signal_6269, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_5543, SubBytesIns_Inst_Sbox_15_T17}), .clk (clk), .r (Fresh[595]), .c ({new_AGEMA_signal_6508, SubBytesIns_Inst_Sbox_15_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M52_U1 ( .a ({new_AGEMA_signal_6502, SubBytesIns_Inst_Sbox_15_M42}), .b ({new_AGEMA_signal_5288, SubBytesIns_Inst_Sbox_15_T15}), .clk (clk), .r (Fresh[596]), .c ({new_AGEMA_signal_6744, SubBytesIns_Inst_Sbox_15_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M53_U1 ( .a ({new_AGEMA_signal_6741, SubBytesIns_Inst_Sbox_15_M45}), .b ({new_AGEMA_signal_5292, SubBytesIns_Inst_Sbox_15_T27}), .clk (clk), .r (Fresh[597]), .c ({new_AGEMA_signal_6943, SubBytesIns_Inst_Sbox_15_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M54_U1 ( .a ({new_AGEMA_signal_6501, SubBytesIns_Inst_Sbox_15_M41}), .b ({new_AGEMA_signal_5541, SubBytesIns_Inst_Sbox_15_T10}), .clk (clk), .r (Fresh[598]), .c ({new_AGEMA_signal_6745, SubBytesIns_Inst_Sbox_15_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M55_U1 ( .a ({new_AGEMA_signal_6504, SubBytesIns_Inst_Sbox_15_M44}), .b ({new_AGEMA_signal_5287, SubBytesIns_Inst_Sbox_15_T13}), .clk (clk), .r (Fresh[599]), .c ({new_AGEMA_signal_6746, SubBytesIns_Inst_Sbox_15_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M56_U1 ( .a ({new_AGEMA_signal_6272, SubBytesIns_Inst_Sbox_15_M40}), .b ({new_AGEMA_signal_5545, SubBytesIns_Inst_Sbox_15_T23}), .clk (clk), .r (Fresh[600]), .c ({new_AGEMA_signal_6509, SubBytesIns_Inst_Sbox_15_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M57_U1 ( .a ({new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_M39}), .b ({new_AGEMA_signal_5290, SubBytesIns_Inst_Sbox_15_T19}), .clk (clk), .r (Fresh[601]), .c ({new_AGEMA_signal_6510, SubBytesIns_Inst_Sbox_15_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M58_U1 ( .a ({new_AGEMA_signal_6503, SubBytesIns_Inst_Sbox_15_M43}), .b ({new_AGEMA_signal_5125, SubBytesIns_Inst_Sbox_15_T3}), .clk (clk), .r (Fresh[602]), .c ({new_AGEMA_signal_6747, SubBytesIns_Inst_Sbox_15_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M59_U1 ( .a ({new_AGEMA_signal_6270, SubBytesIns_Inst_Sbox_15_M38}), .b ({new_AGEMA_signal_5291, SubBytesIns_Inst_Sbox_15_T22}), .clk (clk), .r (Fresh[603]), .c ({new_AGEMA_signal_6511, SubBytesIns_Inst_Sbox_15_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M60_U1 ( .a ({new_AGEMA_signal_6269, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_5544, SubBytesIns_Inst_Sbox_15_T20}), .clk (clk), .r (Fresh[604]), .c ({new_AGEMA_signal_6512, SubBytesIns_Inst_Sbox_15_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M61_U1 ( .a ({new_AGEMA_signal_6502, SubBytesIns_Inst_Sbox_15_M42}), .b ({new_AGEMA_signal_5123, SubBytesIns_Inst_Sbox_15_T1}), .clk (clk), .r (Fresh[605]), .c ({new_AGEMA_signal_6748, SubBytesIns_Inst_Sbox_15_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M62_U1 ( .a ({new_AGEMA_signal_6741, SubBytesIns_Inst_Sbox_15_M45}), .b ({new_AGEMA_signal_5126, SubBytesIns_Inst_Sbox_15_T4}), .clk (clk), .r (Fresh[606]), .c ({new_AGEMA_signal_6944, SubBytesIns_Inst_Sbox_15_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M63_U1 ( .a ({new_AGEMA_signal_6501, SubBytesIns_Inst_Sbox_15_M41}), .b ({new_AGEMA_signal_5124, SubBytesIns_Inst_Sbox_15_T2}), .clk (clk), .r (Fresh[607]), .c ({new_AGEMA_signal_6749, SubBytesIns_Inst_Sbox_15_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L0_U1 ( .a ({new_AGEMA_signal_6748, SubBytesIns_Inst_Sbox_15_M61}), .b ({new_AGEMA_signal_6944, SubBytesIns_Inst_Sbox_15_M62}), .c ({new_AGEMA_signal_7124, SubBytesIns_Inst_Sbox_15_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L1_U1 ( .a ({new_AGEMA_signal_6507, SubBytesIns_Inst_Sbox_15_M50}), .b ({new_AGEMA_signal_6509, SubBytesIns_Inst_Sbox_15_M56}), .c ({new_AGEMA_signal_6750, SubBytesIns_Inst_Sbox_15_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L2_U1 ( .a ({new_AGEMA_signal_6742, SubBytesIns_Inst_Sbox_15_M46}), .b ({new_AGEMA_signal_6506, SubBytesIns_Inst_Sbox_15_M48}), .c ({new_AGEMA_signal_6945, SubBytesIns_Inst_Sbox_15_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L3_U1 ( .a ({new_AGEMA_signal_6505, SubBytesIns_Inst_Sbox_15_M47}), .b ({new_AGEMA_signal_6746, SubBytesIns_Inst_Sbox_15_M55}), .c ({new_AGEMA_signal_6946, SubBytesIns_Inst_Sbox_15_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L4_U1 ( .a ({new_AGEMA_signal_6745, SubBytesIns_Inst_Sbox_15_M54}), .b ({new_AGEMA_signal_6747, SubBytesIns_Inst_Sbox_15_M58}), .c ({new_AGEMA_signal_6947, SubBytesIns_Inst_Sbox_15_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L5_U1 ( .a ({new_AGEMA_signal_6743, SubBytesIns_Inst_Sbox_15_M49}), .b ({new_AGEMA_signal_6748, SubBytesIns_Inst_Sbox_15_M61}), .c ({new_AGEMA_signal_6948, SubBytesIns_Inst_Sbox_15_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L6_U1 ( .a ({new_AGEMA_signal_6944, SubBytesIns_Inst_Sbox_15_M62}), .b ({new_AGEMA_signal_6948, SubBytesIns_Inst_Sbox_15_L5}), .c ({new_AGEMA_signal_7125, SubBytesIns_Inst_Sbox_15_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L7_U1 ( .a ({new_AGEMA_signal_6742, SubBytesIns_Inst_Sbox_15_M46}), .b ({new_AGEMA_signal_6946, SubBytesIns_Inst_Sbox_15_L3}), .c ({new_AGEMA_signal_7126, SubBytesIns_Inst_Sbox_15_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L8_U1 ( .a ({new_AGEMA_signal_6508, SubBytesIns_Inst_Sbox_15_M51}), .b ({new_AGEMA_signal_6511, SubBytesIns_Inst_Sbox_15_M59}), .c ({new_AGEMA_signal_6751, SubBytesIns_Inst_Sbox_15_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L9_U1 ( .a ({new_AGEMA_signal_6744, SubBytesIns_Inst_Sbox_15_M52}), .b ({new_AGEMA_signal_6943, SubBytesIns_Inst_Sbox_15_M53}), .c ({new_AGEMA_signal_7127, SubBytesIns_Inst_Sbox_15_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L10_U1 ( .a ({new_AGEMA_signal_6943, SubBytesIns_Inst_Sbox_15_M53}), .b ({new_AGEMA_signal_6947, SubBytesIns_Inst_Sbox_15_L4}), .c ({new_AGEMA_signal_7128, SubBytesIns_Inst_Sbox_15_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L11_U1 ( .a ({new_AGEMA_signal_6512, SubBytesIns_Inst_Sbox_15_M60}), .b ({new_AGEMA_signal_6945, SubBytesIns_Inst_Sbox_15_L2}), .c ({new_AGEMA_signal_7129, SubBytesIns_Inst_Sbox_15_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L12_U1 ( .a ({new_AGEMA_signal_6506, SubBytesIns_Inst_Sbox_15_M48}), .b ({new_AGEMA_signal_6508, SubBytesIns_Inst_Sbox_15_M51}), .c ({new_AGEMA_signal_6752, SubBytesIns_Inst_Sbox_15_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L13_U1 ( .a ({new_AGEMA_signal_6507, SubBytesIns_Inst_Sbox_15_M50}), .b ({new_AGEMA_signal_7124, SubBytesIns_Inst_Sbox_15_L0}), .c ({new_AGEMA_signal_7342, SubBytesIns_Inst_Sbox_15_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L14_U1 ( .a ({new_AGEMA_signal_6744, SubBytesIns_Inst_Sbox_15_M52}), .b ({new_AGEMA_signal_6748, SubBytesIns_Inst_Sbox_15_M61}), .c ({new_AGEMA_signal_6949, SubBytesIns_Inst_Sbox_15_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L15_U1 ( .a ({new_AGEMA_signal_6746, SubBytesIns_Inst_Sbox_15_M55}), .b ({new_AGEMA_signal_6750, SubBytesIns_Inst_Sbox_15_L1}), .c ({new_AGEMA_signal_6950, SubBytesIns_Inst_Sbox_15_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L16_U1 ( .a ({new_AGEMA_signal_6509, SubBytesIns_Inst_Sbox_15_M56}), .b ({new_AGEMA_signal_7124, SubBytesIns_Inst_Sbox_15_L0}), .c ({new_AGEMA_signal_7343, SubBytesIns_Inst_Sbox_15_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L17_U1 ( .a ({new_AGEMA_signal_6510, SubBytesIns_Inst_Sbox_15_M57}), .b ({new_AGEMA_signal_6750, SubBytesIns_Inst_Sbox_15_L1}), .c ({new_AGEMA_signal_6951, SubBytesIns_Inst_Sbox_15_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L18_U1 ( .a ({new_AGEMA_signal_6747, SubBytesIns_Inst_Sbox_15_M58}), .b ({new_AGEMA_signal_6751, SubBytesIns_Inst_Sbox_15_L8}), .c ({new_AGEMA_signal_6952, SubBytesIns_Inst_Sbox_15_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L19_U1 ( .a ({new_AGEMA_signal_6749, SubBytesIns_Inst_Sbox_15_M63}), .b ({new_AGEMA_signal_6947, SubBytesIns_Inst_Sbox_15_L4}), .c ({new_AGEMA_signal_7130, SubBytesIns_Inst_Sbox_15_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L20_U1 ( .a ({new_AGEMA_signal_7124, SubBytesIns_Inst_Sbox_15_L0}), .b ({new_AGEMA_signal_6750, SubBytesIns_Inst_Sbox_15_L1}), .c ({new_AGEMA_signal_7344, SubBytesIns_Inst_Sbox_15_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L21_U1 ( .a ({new_AGEMA_signal_6750, SubBytesIns_Inst_Sbox_15_L1}), .b ({new_AGEMA_signal_7126, SubBytesIns_Inst_Sbox_15_L7}), .c ({new_AGEMA_signal_7345, SubBytesIns_Inst_Sbox_15_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L22_U1 ( .a ({new_AGEMA_signal_6946, SubBytesIns_Inst_Sbox_15_L3}), .b ({new_AGEMA_signal_6752, SubBytesIns_Inst_Sbox_15_L12}), .c ({new_AGEMA_signal_7131, SubBytesIns_Inst_Sbox_15_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L23_U1 ( .a ({new_AGEMA_signal_6952, SubBytesIns_Inst_Sbox_15_L18}), .b ({new_AGEMA_signal_6945, SubBytesIns_Inst_Sbox_15_L2}), .c ({new_AGEMA_signal_7132, SubBytesIns_Inst_Sbox_15_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L24_U1 ( .a ({new_AGEMA_signal_6950, SubBytesIns_Inst_Sbox_15_L15}), .b ({new_AGEMA_signal_7127, SubBytesIns_Inst_Sbox_15_L9}), .c ({new_AGEMA_signal_7346, SubBytesIns_Inst_Sbox_15_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L25_U1 ( .a ({new_AGEMA_signal_7125, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_7128, SubBytesIns_Inst_Sbox_15_L10}), .c ({new_AGEMA_signal_7347, SubBytesIns_Inst_Sbox_15_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L26_U1 ( .a ({new_AGEMA_signal_7126, SubBytesIns_Inst_Sbox_15_L7}), .b ({new_AGEMA_signal_7127, SubBytesIns_Inst_Sbox_15_L9}), .c ({new_AGEMA_signal_7348, SubBytesIns_Inst_Sbox_15_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L27_U1 ( .a ({new_AGEMA_signal_6751, SubBytesIns_Inst_Sbox_15_L8}), .b ({new_AGEMA_signal_7128, SubBytesIns_Inst_Sbox_15_L10}), .c ({new_AGEMA_signal_7349, SubBytesIns_Inst_Sbox_15_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L28_U1 ( .a ({new_AGEMA_signal_7129, SubBytesIns_Inst_Sbox_15_L11}), .b ({new_AGEMA_signal_6949, SubBytesIns_Inst_Sbox_15_L14}), .c ({new_AGEMA_signal_7350, SubBytesIns_Inst_Sbox_15_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L29_U1 ( .a ({new_AGEMA_signal_7129, SubBytesIns_Inst_Sbox_15_L11}), .b ({new_AGEMA_signal_6951, SubBytesIns_Inst_Sbox_15_L17}), .c ({new_AGEMA_signal_7351, SubBytesIns_Inst_Sbox_15_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S0_U1 ( .a ({new_AGEMA_signal_7125, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_7346, SubBytesIns_Inst_Sbox_15_L24}), .c ({new_AGEMA_signal_7490, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S1_U1 ( .a ({new_AGEMA_signal_7343, SubBytesIns_Inst_Sbox_15_L16}), .b ({new_AGEMA_signal_7348, SubBytesIns_Inst_Sbox_15_L26}), .c ({new_AGEMA_signal_7491, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S2_U1 ( .a ({new_AGEMA_signal_7130, SubBytesIns_Inst_Sbox_15_L19}), .b ({new_AGEMA_signal_7350, SubBytesIns_Inst_Sbox_15_L28}), .c ({new_AGEMA_signal_7492, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S3_U1 ( .a ({new_AGEMA_signal_7125, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_7345, SubBytesIns_Inst_Sbox_15_L21}), .c ({new_AGEMA_signal_7493, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S4_U1 ( .a ({new_AGEMA_signal_7344, SubBytesIns_Inst_Sbox_15_L20}), .b ({new_AGEMA_signal_7131, SubBytesIns_Inst_Sbox_15_L22}), .c ({new_AGEMA_signal_7494, MixColumnsInput[123]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S5_U1 ( .a ({new_AGEMA_signal_7347, SubBytesIns_Inst_Sbox_15_L25}), .b ({new_AGEMA_signal_7351, SubBytesIns_Inst_Sbox_15_L29}), .c ({new_AGEMA_signal_7495, MixColumnsInput[122]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S6_U1 ( .a ({new_AGEMA_signal_7342, SubBytesIns_Inst_Sbox_15_L13}), .b ({new_AGEMA_signal_7349, SubBytesIns_Inst_Sbox_15_L27}), .c ({new_AGEMA_signal_7496, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S7_U1 ( .a ({new_AGEMA_signal_7125, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_7132, SubBytesIns_Inst_Sbox_15_L23}), .c ({new_AGEMA_signal_7352, MixColumnsInput[120]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U96 ( .a ({new_AGEMA_signal_7969, MixColumnsIns_MixOneColumnInst_0_n64}), .b ({new_AGEMA_signal_7461, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .c ({new_AGEMA_signal_8270, MixColumnsOutput[105]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U95 ( .a ({new_AGEMA_signal_7766, MixColumnsIns_MixOneColumnInst_0_n63}), .b ({new_AGEMA_signal_7762, MixColumnsIns_MixOneColumnInst_0_n62}), .c ({new_AGEMA_signal_7969, MixColumnsIns_MixOneColumnInst_0_n64}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U94 ( .a ({new_AGEMA_signal_7745, MixColumnsIns_MixOneColumnInst_0_n61}), .b ({new_AGEMA_signal_7544, MixColumnsIns_MixOneColumnInst_0_n60}), .c ({new_AGEMA_signal_7970, MixColumnsOutput[104]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U93 ( .a ({new_AGEMA_signal_7554, MixColumnsIns_MixOneColumnInst_0_n59}), .b ({new_AGEMA_signal_7297, MixColumnsInput[112]}), .c ({new_AGEMA_signal_7745, MixColumnsIns_MixOneColumnInst_0_n61}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U92 ( .a ({new_AGEMA_signal_7746, MixColumnsIns_MixOneColumnInst_0_n58}), .b ({new_AGEMA_signal_7535, MixColumnsIns_MixOneColumnInst_0_n57}), .c ({new_AGEMA_signal_7971, MixColumnsOutput[103]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U91 ( .a ({new_AGEMA_signal_7546, MixColumnsIns_MixOneColumnInst_0_n56}), .b ({new_AGEMA_signal_7420, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .c ({new_AGEMA_signal_7746, MixColumnsIns_MixOneColumnInst_0_n58}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U90 ( .a ({new_AGEMA_signal_7747, MixColumnsIns_MixOneColumnInst_0_n55}), .b ({new_AGEMA_signal_7536, MixColumnsIns_MixOneColumnInst_0_n54}), .c ({new_AGEMA_signal_7972, MixColumnsOutput[102]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U89 ( .a ({new_AGEMA_signal_7548, MixColumnsIns_MixOneColumnInst_0_n53}), .b ({new_AGEMA_signal_7421, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .c ({new_AGEMA_signal_7747, MixColumnsIns_MixOneColumnInst_0_n55}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U88 ( .a ({new_AGEMA_signal_7748, MixColumnsIns_MixOneColumnInst_0_n52}), .b ({new_AGEMA_signal_7537, MixColumnsIns_MixOneColumnInst_0_n51}), .c ({new_AGEMA_signal_7973, MixColumnsOutput[101]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U87 ( .a ({new_AGEMA_signal_7550, MixColumnsIns_MixOneColumnInst_0_n50}), .b ({new_AGEMA_signal_7422, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .c ({new_AGEMA_signal_7748, MixColumnsIns_MixOneColumnInst_0_n52}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U86 ( .a ({new_AGEMA_signal_7974, MixColumnsIns_MixOneColumnInst_0_n49}), .b ({new_AGEMA_signal_7753, MixColumnsIns_MixOneColumnInst_0_n48}), .c ({new_AGEMA_signal_8271, MixColumnsOutput[100]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U85 ( .a ({new_AGEMA_signal_7772, MixColumnsIns_MixOneColumnInst_0_n47}), .b ({new_AGEMA_signal_7423, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .c ({new_AGEMA_signal_7974, MixColumnsIns_MixOneColumnInst_0_n49}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U84 ( .a ({new_AGEMA_signal_7975, MixColumnsIns_MixOneColumnInst_0_n46}), .b ({new_AGEMA_signal_7754, MixColumnsIns_MixOneColumnInst_0_n45}), .c ({new_AGEMA_signal_8272, MixColumnsOutput[99]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U83 ( .a ({new_AGEMA_signal_7774, MixColumnsIns_MixOneColumnInst_0_n44}), .b ({new_AGEMA_signal_7424, MixColumnsInput[107]}), .c ({new_AGEMA_signal_7975, MixColumnsIns_MixOneColumnInst_0_n46}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U82 ( .a ({new_AGEMA_signal_7749, MixColumnsIns_MixOneColumnInst_0_n43}), .b ({new_AGEMA_signal_7535, MixColumnsIns_MixOneColumnInst_0_n57}), .c ({new_AGEMA_signal_7976, MixColumnsOutput[127]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U81 ( .a ({new_AGEMA_signal_7455, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_7491, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .c ({new_AGEMA_signal_7535, MixColumnsIns_MixOneColumnInst_0_n57}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U80 ( .a ({new_AGEMA_signal_7385, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_7539, MixColumnsIns_MixOneColumnInst_0_n42}), .c ({new_AGEMA_signal_7749, MixColumnsIns_MixOneColumnInst_0_n43}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U79 ( .a ({new_AGEMA_signal_7750, MixColumnsIns_MixOneColumnInst_0_n41}), .b ({new_AGEMA_signal_7536, MixColumnsIns_MixOneColumnInst_0_n54}), .c ({new_AGEMA_signal_7977, MixColumnsOutput[126]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U78 ( .a ({new_AGEMA_signal_7456, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .b ({new_AGEMA_signal_7492, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .c ({new_AGEMA_signal_7536, MixColumnsIns_MixOneColumnInst_0_n54}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U77 ( .a ({new_AGEMA_signal_7386, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .b ({new_AGEMA_signal_7540, MixColumnsIns_MixOneColumnInst_0_n40}), .c ({new_AGEMA_signal_7750, MixColumnsIns_MixOneColumnInst_0_n41}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U76 ( .a ({new_AGEMA_signal_7751, MixColumnsIns_MixOneColumnInst_0_n39}), .b ({new_AGEMA_signal_7538, MixColumnsIns_MixOneColumnInst_0_n38}), .c ({new_AGEMA_signal_7978, MixColumnsOutput[98]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U75 ( .a ({new_AGEMA_signal_7552, MixColumnsIns_MixOneColumnInst_0_n37}), .b ({new_AGEMA_signal_7425, MixColumnsInput[106]}), .c ({new_AGEMA_signal_7751, MixColumnsIns_MixOneColumnInst_0_n39}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U74 ( .a ({new_AGEMA_signal_7752, MixColumnsIns_MixOneColumnInst_0_n36}), .b ({new_AGEMA_signal_7537, MixColumnsIns_MixOneColumnInst_0_n51}), .c ({new_AGEMA_signal_7979, MixColumnsOutput[125]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U73 ( .a ({new_AGEMA_signal_7457, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .b ({new_AGEMA_signal_7493, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .c ({new_AGEMA_signal_7537, MixColumnsIns_MixOneColumnInst_0_n51}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U72 ( .a ({new_AGEMA_signal_7387, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .b ({new_AGEMA_signal_7541, MixColumnsIns_MixOneColumnInst_0_n35}), .c ({new_AGEMA_signal_7752, MixColumnsIns_MixOneColumnInst_0_n36}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U71 ( .a ({new_AGEMA_signal_7980, MixColumnsIns_MixOneColumnInst_0_n34}), .b ({new_AGEMA_signal_7753, MixColumnsIns_MixOneColumnInst_0_n48}), .c ({new_AGEMA_signal_8273, MixColumnsOutput[124]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U70 ( .a ({new_AGEMA_signal_7458, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .b ({new_AGEMA_signal_7555, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]}), .c ({new_AGEMA_signal_7753, MixColumnsIns_MixOneColumnInst_0_n48}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U69 ( .a ({new_AGEMA_signal_7388, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .b ({new_AGEMA_signal_7760, MixColumnsIns_MixOneColumnInst_0_n33}), .c ({new_AGEMA_signal_7980, MixColumnsIns_MixOneColumnInst_0_n34}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U68 ( .a ({new_AGEMA_signal_7981, MixColumnsIns_MixOneColumnInst_0_n32}), .b ({new_AGEMA_signal_7754, MixColumnsIns_MixOneColumnInst_0_n45}), .c ({new_AGEMA_signal_8274, MixColumnsOutput[123]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U67 ( .a ({new_AGEMA_signal_7459, MixColumnsInput[115]}), .b ({new_AGEMA_signal_7556, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]}), .c ({new_AGEMA_signal_7754, MixColumnsIns_MixOneColumnInst_0_n45}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U66 ( .a ({new_AGEMA_signal_7389, MixColumnsInput[99]}), .b ({new_AGEMA_signal_7763, MixColumnsIns_MixOneColumnInst_0_n31}), .c ({new_AGEMA_signal_7981, MixColumnsIns_MixOneColumnInst_0_n32}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U65 ( .a ({new_AGEMA_signal_7755, MixColumnsIns_MixOneColumnInst_0_n30}), .b ({new_AGEMA_signal_7538, MixColumnsIns_MixOneColumnInst_0_n38}), .c ({new_AGEMA_signal_7982, MixColumnsOutput[122]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U64 ( .a ({new_AGEMA_signal_7460, MixColumnsInput[114]}), .b ({new_AGEMA_signal_7496, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .c ({new_AGEMA_signal_7538, MixColumnsIns_MixOneColumnInst_0_n38}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U63 ( .a ({new_AGEMA_signal_7390, MixColumnsInput[98]}), .b ({new_AGEMA_signal_7542, MixColumnsIns_MixOneColumnInst_0_n29}), .c ({new_AGEMA_signal_7755, MixColumnsIns_MixOneColumnInst_0_n30}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U62 ( .a ({new_AGEMA_signal_7983, MixColumnsIns_MixOneColumnInst_0_n28}), .b ({new_AGEMA_signal_7761, MixColumnsIns_MixOneColumnInst_0_n27}), .c ({new_AGEMA_signal_8275, MixColumnsOutput[121]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U61 ( .a ({new_AGEMA_signal_7391, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .b ({new_AGEMA_signal_7765, MixColumnsIns_MixOneColumnInst_0_n26}), .c ({new_AGEMA_signal_7983, MixColumnsIns_MixOneColumnInst_0_n28}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U60 ( .a ({new_AGEMA_signal_7756, MixColumnsIns_MixOneColumnInst_0_n25}), .b ({new_AGEMA_signal_7543, MixColumnsIns_MixOneColumnInst_0_n24}), .c ({new_AGEMA_signal_7984, MixColumnsOutput[120]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U59 ( .a ({new_AGEMA_signal_7553, MixColumnsIns_MixOneColumnInst_0_n23}), .b ({new_AGEMA_signal_7187, MixColumnsInput[96]}), .c ({new_AGEMA_signal_7756, MixColumnsIns_MixOneColumnInst_0_n25}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U58 ( .a ({new_AGEMA_signal_7757, MixColumnsIns_MixOneColumnInst_0_n22}), .b ({new_AGEMA_signal_7539, MixColumnsIns_MixOneColumnInst_0_n42}), .c ({new_AGEMA_signal_7985, MixColumnsOutput[119]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U57 ( .a ({new_AGEMA_signal_7420, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_7456, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .c ({new_AGEMA_signal_7539, MixColumnsIns_MixOneColumnInst_0_n42}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U56 ( .a ({new_AGEMA_signal_7490, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_7545, MixColumnsIns_MixOneColumnInst_0_n21}), .c ({new_AGEMA_signal_7757, MixColumnsIns_MixOneColumnInst_0_n22}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U55 ( .a ({new_AGEMA_signal_7758, MixColumnsIns_MixOneColumnInst_0_n20}), .b ({new_AGEMA_signal_7540, MixColumnsIns_MixOneColumnInst_0_n40}), .c ({new_AGEMA_signal_7986, MixColumnsOutput[118]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U54 ( .a ({new_AGEMA_signal_7421, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .b ({new_AGEMA_signal_7457, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .c ({new_AGEMA_signal_7540, MixColumnsIns_MixOneColumnInst_0_n40}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U53 ( .a ({new_AGEMA_signal_7491, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .b ({new_AGEMA_signal_7547, MixColumnsIns_MixOneColumnInst_0_n19}), .c ({new_AGEMA_signal_7758, MixColumnsIns_MixOneColumnInst_0_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U52 ( .a ({new_AGEMA_signal_7759, MixColumnsIns_MixOneColumnInst_0_n18}), .b ({new_AGEMA_signal_7541, MixColumnsIns_MixOneColumnInst_0_n35}), .c ({new_AGEMA_signal_7987, MixColumnsOutput[117]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U51 ( .a ({new_AGEMA_signal_7422, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .b ({new_AGEMA_signal_7458, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .c ({new_AGEMA_signal_7541, MixColumnsIns_MixOneColumnInst_0_n35}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U50 ( .a ({new_AGEMA_signal_7492, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .b ({new_AGEMA_signal_7549, MixColumnsIns_MixOneColumnInst_0_n17}), .c ({new_AGEMA_signal_7759, MixColumnsIns_MixOneColumnInst_0_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U49 ( .a ({new_AGEMA_signal_7988, MixColumnsIns_MixOneColumnInst_0_n16}), .b ({new_AGEMA_signal_7760, MixColumnsIns_MixOneColumnInst_0_n33}), .c ({new_AGEMA_signal_8276, MixColumnsOutput[116]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U48 ( .a ({new_AGEMA_signal_7423, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .b ({new_AGEMA_signal_7558, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]}), .c ({new_AGEMA_signal_7760, MixColumnsIns_MixOneColumnInst_0_n33}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U47 ( .a ({new_AGEMA_signal_7493, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .b ({new_AGEMA_signal_7771, MixColumnsIns_MixOneColumnInst_0_n15}), .c ({new_AGEMA_signal_7988, MixColumnsIns_MixOneColumnInst_0_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U46 ( .a ({new_AGEMA_signal_7989, MixColumnsIns_MixOneColumnInst_0_n14}), .b ({new_AGEMA_signal_7761, MixColumnsIns_MixOneColumnInst_0_n27}), .c ({new_AGEMA_signal_8277, MixColumnsOutput[97]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U45 ( .a ({new_AGEMA_signal_7461, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .b ({new_AGEMA_signal_7557, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]}), .c ({new_AGEMA_signal_7761, MixColumnsIns_MixOneColumnInst_0_n27}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U44 ( .a ({new_AGEMA_signal_7426, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .b ({new_AGEMA_signal_7762, MixColumnsIns_MixOneColumnInst_0_n62}), .c ({new_AGEMA_signal_7989, MixColumnsIns_MixOneColumnInst_0_n14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U43 ( .a ({new_AGEMA_signal_7496, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .b ({new_AGEMA_signal_7566, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]}), .c ({new_AGEMA_signal_7762, MixColumnsIns_MixOneColumnInst_0_n62}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U42 ( .a ({new_AGEMA_signal_7990, MixColumnsIns_MixOneColumnInst_0_n13}), .b ({new_AGEMA_signal_7763, MixColumnsIns_MixOneColumnInst_0_n31}), .c ({new_AGEMA_signal_8278, MixColumnsOutput[115]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U41 ( .a ({new_AGEMA_signal_7424, MixColumnsInput[107]}), .b ({new_AGEMA_signal_7559, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]}), .c ({new_AGEMA_signal_7763, MixColumnsIns_MixOneColumnInst_0_n31}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U40 ( .a ({new_AGEMA_signal_7494, MixColumnsInput[123]}), .b ({new_AGEMA_signal_7773, MixColumnsIns_MixOneColumnInst_0_n12}), .c ({new_AGEMA_signal_7990, MixColumnsIns_MixOneColumnInst_0_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U39 ( .a ({new_AGEMA_signal_7764, MixColumnsIns_MixOneColumnInst_0_n11}), .b ({new_AGEMA_signal_7542, MixColumnsIns_MixOneColumnInst_0_n29}), .c ({new_AGEMA_signal_7991, MixColumnsOutput[114]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U38 ( .a ({new_AGEMA_signal_7425, MixColumnsInput[106]}), .b ({new_AGEMA_signal_7461, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .c ({new_AGEMA_signal_7542, MixColumnsIns_MixOneColumnInst_0_n29}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U37 ( .a ({new_AGEMA_signal_7495, MixColumnsInput[122]}), .b ({new_AGEMA_signal_7551, MixColumnsIns_MixOneColumnInst_0_n10}), .c ({new_AGEMA_signal_7764, MixColumnsIns_MixOneColumnInst_0_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U36 ( .a ({new_AGEMA_signal_7992, MixColumnsIns_MixOneColumnInst_0_n9}), .b ({new_AGEMA_signal_7765, MixColumnsIns_MixOneColumnInst_0_n26}), .c ({new_AGEMA_signal_8279, MixColumnsOutput[113]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U35 ( .a ({new_AGEMA_signal_7560, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]}), .b ({new_AGEMA_signal_7426, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .c ({new_AGEMA_signal_7765, MixColumnsIns_MixOneColumnInst_0_n26}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U34 ( .a ({new_AGEMA_signal_7766, MixColumnsIns_MixOneColumnInst_0_n63}), .b ({new_AGEMA_signal_7496, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .c ({new_AGEMA_signal_7992, MixColumnsIns_MixOneColumnInst_0_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U33 ( .a ({new_AGEMA_signal_7563, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]}), .b ({new_AGEMA_signal_7391, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .c ({new_AGEMA_signal_7766, MixColumnsIns_MixOneColumnInst_0_n63}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U32 ( .a ({new_AGEMA_signal_7767, MixColumnsIns_MixOneColumnInst_0_n8}), .b ({new_AGEMA_signal_7543, MixColumnsIns_MixOneColumnInst_0_n24}), .c ({new_AGEMA_signal_7993, MixColumnsOutput[112]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U31 ( .a ({new_AGEMA_signal_7242, MixColumnsInput[104]}), .b ({new_AGEMA_signal_7455, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .c ({new_AGEMA_signal_7543, MixColumnsIns_MixOneColumnInst_0_n24}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U30 ( .a ({new_AGEMA_signal_7352, MixColumnsInput[120]}), .b ({new_AGEMA_signal_7544, MixColumnsIns_MixOneColumnInst_0_n60}), .c ({new_AGEMA_signal_7767, MixColumnsIns_MixOneColumnInst_0_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U29 ( .a ({new_AGEMA_signal_7420, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_7187, MixColumnsInput[96]}), .c ({new_AGEMA_signal_7544, MixColumnsIns_MixOneColumnInst_0_n60}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U28 ( .a ({new_AGEMA_signal_7768, MixColumnsIns_MixOneColumnInst_0_n7}), .b ({new_AGEMA_signal_7545, MixColumnsIns_MixOneColumnInst_0_n21}), .c ({new_AGEMA_signal_7994, MixColumnsOutput[111]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U27 ( .a ({new_AGEMA_signal_7385, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_7421, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .c ({new_AGEMA_signal_7545, MixColumnsIns_MixOneColumnInst_0_n21}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U26 ( .a ({new_AGEMA_signal_7546, MixColumnsIns_MixOneColumnInst_0_n56}), .b ({new_AGEMA_signal_7455, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .c ({new_AGEMA_signal_7768, MixColumnsIns_MixOneColumnInst_0_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U25 ( .a ({new_AGEMA_signal_7386, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .b ({new_AGEMA_signal_7490, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .c ({new_AGEMA_signal_7546, MixColumnsIns_MixOneColumnInst_0_n56}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U24 ( .a ({new_AGEMA_signal_7769, MixColumnsIns_MixOneColumnInst_0_n6}), .b ({new_AGEMA_signal_7547, MixColumnsIns_MixOneColumnInst_0_n19}), .c ({new_AGEMA_signal_7995, MixColumnsOutput[110]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U23 ( .a ({new_AGEMA_signal_7386, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .b ({new_AGEMA_signal_7422, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .c ({new_AGEMA_signal_7547, MixColumnsIns_MixOneColumnInst_0_n19}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U22 ( .a ({new_AGEMA_signal_7548, MixColumnsIns_MixOneColumnInst_0_n53}), .b ({new_AGEMA_signal_7456, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .c ({new_AGEMA_signal_7769, MixColumnsIns_MixOneColumnInst_0_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U21 ( .a ({new_AGEMA_signal_7387, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .b ({new_AGEMA_signal_7491, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .c ({new_AGEMA_signal_7548, MixColumnsIns_MixOneColumnInst_0_n53}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U20 ( .a ({new_AGEMA_signal_7770, MixColumnsIns_MixOneColumnInst_0_n5}), .b ({new_AGEMA_signal_7549, MixColumnsIns_MixOneColumnInst_0_n17}), .c ({new_AGEMA_signal_7996, MixColumnsOutput[109]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U19 ( .a ({new_AGEMA_signal_7387, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .b ({new_AGEMA_signal_7423, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .c ({new_AGEMA_signal_7549, MixColumnsIns_MixOneColumnInst_0_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U18 ( .a ({new_AGEMA_signal_7550, MixColumnsIns_MixOneColumnInst_0_n50}), .b ({new_AGEMA_signal_7457, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .c ({new_AGEMA_signal_7770, MixColumnsIns_MixOneColumnInst_0_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U17 ( .a ({new_AGEMA_signal_7388, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .b ({new_AGEMA_signal_7492, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .c ({new_AGEMA_signal_7550, MixColumnsIns_MixOneColumnInst_0_n50}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U16 ( .a ({new_AGEMA_signal_7997, MixColumnsIns_MixOneColumnInst_0_n4}), .b ({new_AGEMA_signal_7771, MixColumnsIns_MixOneColumnInst_0_n15}), .c ({new_AGEMA_signal_8280, MixColumnsOutput[108]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U15 ( .a ({new_AGEMA_signal_7388, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .b ({new_AGEMA_signal_7561, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]}), .c ({new_AGEMA_signal_7771, MixColumnsIns_MixOneColumnInst_0_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U14 ( .a ({new_AGEMA_signal_7772, MixColumnsIns_MixOneColumnInst_0_n47}), .b ({new_AGEMA_signal_7458, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .c ({new_AGEMA_signal_7997, MixColumnsIns_MixOneColumnInst_0_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U13 ( .a ({new_AGEMA_signal_7564, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]}), .b ({new_AGEMA_signal_7493, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .c ({new_AGEMA_signal_7772, MixColumnsIns_MixOneColumnInst_0_n47}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U12 ( .a ({new_AGEMA_signal_7998, MixColumnsIns_MixOneColumnInst_0_n3}), .b ({new_AGEMA_signal_7773, MixColumnsIns_MixOneColumnInst_0_n12}), .c ({new_AGEMA_signal_8281, MixColumnsOutput[107]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U11 ( .a ({new_AGEMA_signal_7389, MixColumnsInput[99]}), .b ({new_AGEMA_signal_7562, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]}), .c ({new_AGEMA_signal_7773, MixColumnsIns_MixOneColumnInst_0_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U10 ( .a ({new_AGEMA_signal_7774, MixColumnsIns_MixOneColumnInst_0_n44}), .b ({new_AGEMA_signal_7459, MixColumnsInput[115]}), .c ({new_AGEMA_signal_7998, MixColumnsIns_MixOneColumnInst_0_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U9 ( .a ({new_AGEMA_signal_7565, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]}), .b ({new_AGEMA_signal_7494, MixColumnsInput[123]}), .c ({new_AGEMA_signal_7774, MixColumnsIns_MixOneColumnInst_0_n44}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U8 ( .a ({new_AGEMA_signal_7775, MixColumnsIns_MixOneColumnInst_0_n2}), .b ({new_AGEMA_signal_7551, MixColumnsIns_MixOneColumnInst_0_n10}), .c ({new_AGEMA_signal_7999, MixColumnsOutput[106]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U7 ( .a ({new_AGEMA_signal_7390, MixColumnsInput[98]}), .b ({new_AGEMA_signal_7426, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .c ({new_AGEMA_signal_7551, MixColumnsIns_MixOneColumnInst_0_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U6 ( .a ({new_AGEMA_signal_7552, MixColumnsIns_MixOneColumnInst_0_n37}), .b ({new_AGEMA_signal_7460, MixColumnsInput[114]}), .c ({new_AGEMA_signal_7775, MixColumnsIns_MixOneColumnInst_0_n2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U5 ( .a ({new_AGEMA_signal_7391, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .b ({new_AGEMA_signal_7495, MixColumnsInput[122]}), .c ({new_AGEMA_signal_7552, MixColumnsIns_MixOneColumnInst_0_n37}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U4 ( .a ({new_AGEMA_signal_7776, MixColumnsIns_MixOneColumnInst_0_n1}), .b ({new_AGEMA_signal_7242, MixColumnsInput[104]}), .c ({new_AGEMA_signal_8000, MixColumnsOutput[96]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U3 ( .a ({new_AGEMA_signal_7554, MixColumnsIns_MixOneColumnInst_0_n59}), .b ({new_AGEMA_signal_7553, MixColumnsIns_MixOneColumnInst_0_n23}), .c ({new_AGEMA_signal_7776, MixColumnsIns_MixOneColumnInst_0_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U2 ( .a ({new_AGEMA_signal_7297, MixColumnsInput[112]}), .b ({new_AGEMA_signal_7490, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .c ({new_AGEMA_signal_7553, MixColumnsIns_MixOneColumnInst_0_n23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U1 ( .a ({new_AGEMA_signal_7385, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_7352, MixColumnsInput[120]}), .c ({new_AGEMA_signal_7554, MixColumnsIns_MixOneColumnInst_0_n59}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_7490, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_7494, MixColumnsInput[123]}), .c ({new_AGEMA_signal_7555, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_7490, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_7495, MixColumnsInput[122]}), .c ({new_AGEMA_signal_7556, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_7490, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_7352, MixColumnsInput[120]}), .c ({new_AGEMA_signal_7557, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_7455, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_7459, MixColumnsInput[115]}), .c ({new_AGEMA_signal_7558, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_7455, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_7460, MixColumnsInput[114]}), .c ({new_AGEMA_signal_7559, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_7455, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_7297, MixColumnsInput[112]}), .c ({new_AGEMA_signal_7560, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_7420, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_7424, MixColumnsInput[107]}), .c ({new_AGEMA_signal_7561, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_7420, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_7425, MixColumnsInput[106]}), .c ({new_AGEMA_signal_7562, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_7420, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_7242, MixColumnsInput[104]}), .c ({new_AGEMA_signal_7563, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_7385, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_7389, MixColumnsInput[99]}), .c ({new_AGEMA_signal_7564, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_7385, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_7390, MixColumnsInput[98]}), .c ({new_AGEMA_signal_7565, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_7385, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_7187, MixColumnsInput[96]}), .c ({new_AGEMA_signal_7566, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U96 ( .a ({new_AGEMA_signal_8001, MixColumnsIns_MixOneColumnInst_1_n64}), .b ({new_AGEMA_signal_7433, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .c ({new_AGEMA_signal_8282, MixColumnsOutput[73]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U95 ( .a ({new_AGEMA_signal_7798, MixColumnsIns_MixOneColumnInst_1_n63}), .b ({new_AGEMA_signal_7794, MixColumnsIns_MixOneColumnInst_1_n62}), .c ({new_AGEMA_signal_8001, MixColumnsIns_MixOneColumnInst_1_n64}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U94 ( .a ({new_AGEMA_signal_7777, MixColumnsIns_MixOneColumnInst_1_n61}), .b ({new_AGEMA_signal_7576, MixColumnsIns_MixOneColumnInst_1_n60}), .c ({new_AGEMA_signal_8002, MixColumnsOutput[72]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U93 ( .a ({new_AGEMA_signal_7586, MixColumnsIns_MixOneColumnInst_1_n59}), .b ({new_AGEMA_signal_7253, MixColumnsInput[80]}), .c ({new_AGEMA_signal_7777, MixColumnsIns_MixOneColumnInst_1_n61}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U92 ( .a ({new_AGEMA_signal_7778, MixColumnsIns_MixOneColumnInst_1_n58}), .b ({new_AGEMA_signal_7567, MixColumnsIns_MixOneColumnInst_1_n57}), .c ({new_AGEMA_signal_8003, MixColumnsOutput[71]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U91 ( .a ({new_AGEMA_signal_7578, MixColumnsIns_MixOneColumnInst_1_n56}), .b ({new_AGEMA_signal_7392, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .c ({new_AGEMA_signal_7778, MixColumnsIns_MixOneColumnInst_1_n58}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U90 ( .a ({new_AGEMA_signal_7779, MixColumnsIns_MixOneColumnInst_1_n55}), .b ({new_AGEMA_signal_7568, MixColumnsIns_MixOneColumnInst_1_n54}), .c ({new_AGEMA_signal_8004, MixColumnsOutput[70]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U89 ( .a ({new_AGEMA_signal_7580, MixColumnsIns_MixOneColumnInst_1_n53}), .b ({new_AGEMA_signal_7393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .c ({new_AGEMA_signal_7779, MixColumnsIns_MixOneColumnInst_1_n55}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U88 ( .a ({new_AGEMA_signal_7780, MixColumnsIns_MixOneColumnInst_1_n52}), .b ({new_AGEMA_signal_7569, MixColumnsIns_MixOneColumnInst_1_n51}), .c ({new_AGEMA_signal_8005, MixColumnsOutput[69]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U87 ( .a ({new_AGEMA_signal_7582, MixColumnsIns_MixOneColumnInst_1_n50}), .b ({new_AGEMA_signal_7394, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .c ({new_AGEMA_signal_7780, MixColumnsIns_MixOneColumnInst_1_n52}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U86 ( .a ({new_AGEMA_signal_8006, MixColumnsIns_MixOneColumnInst_1_n49}), .b ({new_AGEMA_signal_7785, MixColumnsIns_MixOneColumnInst_1_n48}), .c ({new_AGEMA_signal_8283, MixColumnsOutput[68]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U85 ( .a ({new_AGEMA_signal_7804, MixColumnsIns_MixOneColumnInst_1_n47}), .b ({new_AGEMA_signal_7395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .c ({new_AGEMA_signal_8006, MixColumnsIns_MixOneColumnInst_1_n49}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U84 ( .a ({new_AGEMA_signal_8007, MixColumnsIns_MixOneColumnInst_1_n46}), .b ({new_AGEMA_signal_7786, MixColumnsIns_MixOneColumnInst_1_n45}), .c ({new_AGEMA_signal_8284, MixColumnsOutput[67]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U83 ( .a ({new_AGEMA_signal_7806, MixColumnsIns_MixOneColumnInst_1_n44}), .b ({new_AGEMA_signal_7396, MixColumnsInput[75]}), .c ({new_AGEMA_signal_8007, MixColumnsIns_MixOneColumnInst_1_n46}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U82 ( .a ({new_AGEMA_signal_7781, MixColumnsIns_MixOneColumnInst_1_n43}), .b ({new_AGEMA_signal_7567, MixColumnsIns_MixOneColumnInst_1_n57}), .c ({new_AGEMA_signal_8008, MixColumnsOutput[95]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U81 ( .a ({new_AGEMA_signal_7427, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_7463, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .c ({new_AGEMA_signal_7567, MixColumnsIns_MixOneColumnInst_1_n57}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U80 ( .a ({new_AGEMA_signal_7469, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_7571, MixColumnsIns_MixOneColumnInst_1_n42}), .c ({new_AGEMA_signal_7781, MixColumnsIns_MixOneColumnInst_1_n43}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U79 ( .a ({new_AGEMA_signal_7782, MixColumnsIns_MixOneColumnInst_1_n41}), .b ({new_AGEMA_signal_7568, MixColumnsIns_MixOneColumnInst_1_n54}), .c ({new_AGEMA_signal_8009, MixColumnsOutput[94]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U78 ( .a ({new_AGEMA_signal_7428, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .b ({new_AGEMA_signal_7464, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .c ({new_AGEMA_signal_7568, MixColumnsIns_MixOneColumnInst_1_n54}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U77 ( .a ({new_AGEMA_signal_7470, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .b ({new_AGEMA_signal_7572, MixColumnsIns_MixOneColumnInst_1_n40}), .c ({new_AGEMA_signal_7782, MixColumnsIns_MixOneColumnInst_1_n41}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U76 ( .a ({new_AGEMA_signal_7783, MixColumnsIns_MixOneColumnInst_1_n39}), .b ({new_AGEMA_signal_7570, MixColumnsIns_MixOneColumnInst_1_n38}), .c ({new_AGEMA_signal_8010, MixColumnsOutput[66]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U75 ( .a ({new_AGEMA_signal_7584, MixColumnsIns_MixOneColumnInst_1_n37}), .b ({new_AGEMA_signal_7397, MixColumnsInput[74]}), .c ({new_AGEMA_signal_7783, MixColumnsIns_MixOneColumnInst_1_n39}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U74 ( .a ({new_AGEMA_signal_7784, MixColumnsIns_MixOneColumnInst_1_n36}), .b ({new_AGEMA_signal_7569, MixColumnsIns_MixOneColumnInst_1_n51}), .c ({new_AGEMA_signal_8011, MixColumnsOutput[93]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U73 ( .a ({new_AGEMA_signal_7429, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .b ({new_AGEMA_signal_7465, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .c ({new_AGEMA_signal_7569, MixColumnsIns_MixOneColumnInst_1_n51}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U72 ( .a ({new_AGEMA_signal_7471, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .b ({new_AGEMA_signal_7573, MixColumnsIns_MixOneColumnInst_1_n35}), .c ({new_AGEMA_signal_7784, MixColumnsIns_MixOneColumnInst_1_n36}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U71 ( .a ({new_AGEMA_signal_8012, MixColumnsIns_MixOneColumnInst_1_n34}), .b ({new_AGEMA_signal_7785, MixColumnsIns_MixOneColumnInst_1_n48}), .c ({new_AGEMA_signal_8285, MixColumnsOutput[92]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U70 ( .a ({new_AGEMA_signal_7430, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .b ({new_AGEMA_signal_7587, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]}), .c ({new_AGEMA_signal_7785, MixColumnsIns_MixOneColumnInst_1_n48}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U69 ( .a ({new_AGEMA_signal_7472, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .b ({new_AGEMA_signal_7792, MixColumnsIns_MixOneColumnInst_1_n33}), .c ({new_AGEMA_signal_8012, MixColumnsIns_MixOneColumnInst_1_n34}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U68 ( .a ({new_AGEMA_signal_8013, MixColumnsIns_MixOneColumnInst_1_n32}), .b ({new_AGEMA_signal_7786, MixColumnsIns_MixOneColumnInst_1_n45}), .c ({new_AGEMA_signal_8286, MixColumnsOutput[91]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U67 ( .a ({new_AGEMA_signal_7431, MixColumnsInput[83]}), .b ({new_AGEMA_signal_7588, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]}), .c ({new_AGEMA_signal_7786, MixColumnsIns_MixOneColumnInst_1_n45}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U66 ( .a ({new_AGEMA_signal_7473, MixColumnsInput[67]}), .b ({new_AGEMA_signal_7795, MixColumnsIns_MixOneColumnInst_1_n31}), .c ({new_AGEMA_signal_8013, MixColumnsIns_MixOneColumnInst_1_n32}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U65 ( .a ({new_AGEMA_signal_7787, MixColumnsIns_MixOneColumnInst_1_n30}), .b ({new_AGEMA_signal_7570, MixColumnsIns_MixOneColumnInst_1_n38}), .c ({new_AGEMA_signal_8014, MixColumnsOutput[90]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U64 ( .a ({new_AGEMA_signal_7432, MixColumnsInput[82]}), .b ({new_AGEMA_signal_7468, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .c ({new_AGEMA_signal_7570, MixColumnsIns_MixOneColumnInst_1_n38}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U63 ( .a ({new_AGEMA_signal_7474, MixColumnsInput[66]}), .b ({new_AGEMA_signal_7574, MixColumnsIns_MixOneColumnInst_1_n29}), .c ({new_AGEMA_signal_7787, MixColumnsIns_MixOneColumnInst_1_n30}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U62 ( .a ({new_AGEMA_signal_8015, MixColumnsIns_MixOneColumnInst_1_n28}), .b ({new_AGEMA_signal_7793, MixColumnsIns_MixOneColumnInst_1_n27}), .c ({new_AGEMA_signal_8287, MixColumnsOutput[89]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U61 ( .a ({new_AGEMA_signal_7475, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .b ({new_AGEMA_signal_7797, MixColumnsIns_MixOneColumnInst_1_n26}), .c ({new_AGEMA_signal_8015, MixColumnsIns_MixOneColumnInst_1_n28}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U60 ( .a ({new_AGEMA_signal_7788, MixColumnsIns_MixOneColumnInst_1_n25}), .b ({new_AGEMA_signal_7575, MixColumnsIns_MixOneColumnInst_1_n24}), .c ({new_AGEMA_signal_8016, MixColumnsOutput[88]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U59 ( .a ({new_AGEMA_signal_7585, MixColumnsIns_MixOneColumnInst_1_n23}), .b ({new_AGEMA_signal_7319, MixColumnsInput[64]}), .c ({new_AGEMA_signal_7788, MixColumnsIns_MixOneColumnInst_1_n25}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U58 ( .a ({new_AGEMA_signal_7789, MixColumnsIns_MixOneColumnInst_1_n22}), .b ({new_AGEMA_signal_7571, MixColumnsIns_MixOneColumnInst_1_n42}), .c ({new_AGEMA_signal_8017, MixColumnsOutput[87]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U57 ( .a ({new_AGEMA_signal_7392, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_7428, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .c ({new_AGEMA_signal_7571, MixColumnsIns_MixOneColumnInst_1_n42}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U56 ( .a ({new_AGEMA_signal_7462, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_7577, MixColumnsIns_MixOneColumnInst_1_n21}), .c ({new_AGEMA_signal_7789, MixColumnsIns_MixOneColumnInst_1_n22}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U55 ( .a ({new_AGEMA_signal_7790, MixColumnsIns_MixOneColumnInst_1_n20}), .b ({new_AGEMA_signal_7572, MixColumnsIns_MixOneColumnInst_1_n40}), .c ({new_AGEMA_signal_8018, MixColumnsOutput[86]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U54 ( .a ({new_AGEMA_signal_7393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .b ({new_AGEMA_signal_7429, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .c ({new_AGEMA_signal_7572, MixColumnsIns_MixOneColumnInst_1_n40}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U53 ( .a ({new_AGEMA_signal_7463, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .b ({new_AGEMA_signal_7579, MixColumnsIns_MixOneColumnInst_1_n19}), .c ({new_AGEMA_signal_7790, MixColumnsIns_MixOneColumnInst_1_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U52 ( .a ({new_AGEMA_signal_7791, MixColumnsIns_MixOneColumnInst_1_n18}), .b ({new_AGEMA_signal_7573, MixColumnsIns_MixOneColumnInst_1_n35}), .c ({new_AGEMA_signal_8019, MixColumnsOutput[85]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U51 ( .a ({new_AGEMA_signal_7394, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .b ({new_AGEMA_signal_7430, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .c ({new_AGEMA_signal_7573, MixColumnsIns_MixOneColumnInst_1_n35}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U50 ( .a ({new_AGEMA_signal_7464, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .b ({new_AGEMA_signal_7581, MixColumnsIns_MixOneColumnInst_1_n17}), .c ({new_AGEMA_signal_7791, MixColumnsIns_MixOneColumnInst_1_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U49 ( .a ({new_AGEMA_signal_8020, MixColumnsIns_MixOneColumnInst_1_n16}), .b ({new_AGEMA_signal_7792, MixColumnsIns_MixOneColumnInst_1_n33}), .c ({new_AGEMA_signal_8288, MixColumnsOutput[84]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U48 ( .a ({new_AGEMA_signal_7395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .b ({new_AGEMA_signal_7590, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]}), .c ({new_AGEMA_signal_7792, MixColumnsIns_MixOneColumnInst_1_n33}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U47 ( .a ({new_AGEMA_signal_7465, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .b ({new_AGEMA_signal_7803, MixColumnsIns_MixOneColumnInst_1_n15}), .c ({new_AGEMA_signal_8020, MixColumnsIns_MixOneColumnInst_1_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U46 ( .a ({new_AGEMA_signal_8021, MixColumnsIns_MixOneColumnInst_1_n14}), .b ({new_AGEMA_signal_7793, MixColumnsIns_MixOneColumnInst_1_n27}), .c ({new_AGEMA_signal_8289, MixColumnsOutput[65]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U45 ( .a ({new_AGEMA_signal_7433, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .b ({new_AGEMA_signal_7589, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]}), .c ({new_AGEMA_signal_7793, MixColumnsIns_MixOneColumnInst_1_n27}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U44 ( .a ({new_AGEMA_signal_7398, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .b ({new_AGEMA_signal_7794, MixColumnsIns_MixOneColumnInst_1_n62}), .c ({new_AGEMA_signal_8021, MixColumnsIns_MixOneColumnInst_1_n14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U43 ( .a ({new_AGEMA_signal_7468, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .b ({new_AGEMA_signal_7598, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]}), .c ({new_AGEMA_signal_7794, MixColumnsIns_MixOneColumnInst_1_n62}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U42 ( .a ({new_AGEMA_signal_8022, MixColumnsIns_MixOneColumnInst_1_n13}), .b ({new_AGEMA_signal_7795, MixColumnsIns_MixOneColumnInst_1_n31}), .c ({new_AGEMA_signal_8290, MixColumnsOutput[83]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U41 ( .a ({new_AGEMA_signal_7396, MixColumnsInput[75]}), .b ({new_AGEMA_signal_7591, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]}), .c ({new_AGEMA_signal_7795, MixColumnsIns_MixOneColumnInst_1_n31}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U40 ( .a ({new_AGEMA_signal_7466, MixColumnsInput[91]}), .b ({new_AGEMA_signal_7805, MixColumnsIns_MixOneColumnInst_1_n12}), .c ({new_AGEMA_signal_8022, MixColumnsIns_MixOneColumnInst_1_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U39 ( .a ({new_AGEMA_signal_7796, MixColumnsIns_MixOneColumnInst_1_n11}), .b ({new_AGEMA_signal_7574, MixColumnsIns_MixOneColumnInst_1_n29}), .c ({new_AGEMA_signal_8023, MixColumnsOutput[82]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U38 ( .a ({new_AGEMA_signal_7397, MixColumnsInput[74]}), .b ({new_AGEMA_signal_7433, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .c ({new_AGEMA_signal_7574, MixColumnsIns_MixOneColumnInst_1_n29}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U37 ( .a ({new_AGEMA_signal_7467, MixColumnsInput[90]}), .b ({new_AGEMA_signal_7583, MixColumnsIns_MixOneColumnInst_1_n10}), .c ({new_AGEMA_signal_7796, MixColumnsIns_MixOneColumnInst_1_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U36 ( .a ({new_AGEMA_signal_8024, MixColumnsIns_MixOneColumnInst_1_n9}), .b ({new_AGEMA_signal_7797, MixColumnsIns_MixOneColumnInst_1_n26}), .c ({new_AGEMA_signal_8291, MixColumnsOutput[81]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U35 ( .a ({new_AGEMA_signal_7592, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]}), .b ({new_AGEMA_signal_7398, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .c ({new_AGEMA_signal_7797, MixColumnsIns_MixOneColumnInst_1_n26}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U34 ( .a ({new_AGEMA_signal_7798, MixColumnsIns_MixOneColumnInst_1_n63}), .b ({new_AGEMA_signal_7468, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .c ({new_AGEMA_signal_8024, MixColumnsIns_MixOneColumnInst_1_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U33 ( .a ({new_AGEMA_signal_7595, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]}), .b ({new_AGEMA_signal_7475, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .c ({new_AGEMA_signal_7798, MixColumnsIns_MixOneColumnInst_1_n63}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U32 ( .a ({new_AGEMA_signal_7799, MixColumnsIns_MixOneColumnInst_1_n8}), .b ({new_AGEMA_signal_7575, MixColumnsIns_MixOneColumnInst_1_n24}), .c ({new_AGEMA_signal_8025, MixColumnsOutput[80]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U31 ( .a ({new_AGEMA_signal_7198, MixColumnsInput[72]}), .b ({new_AGEMA_signal_7427, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .c ({new_AGEMA_signal_7575, MixColumnsIns_MixOneColumnInst_1_n24}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U30 ( .a ({new_AGEMA_signal_7308, MixColumnsInput[88]}), .b ({new_AGEMA_signal_7576, MixColumnsIns_MixOneColumnInst_1_n60}), .c ({new_AGEMA_signal_7799, MixColumnsIns_MixOneColumnInst_1_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U29 ( .a ({new_AGEMA_signal_7392, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_7319, MixColumnsInput[64]}), .c ({new_AGEMA_signal_7576, MixColumnsIns_MixOneColumnInst_1_n60}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U28 ( .a ({new_AGEMA_signal_7800, MixColumnsIns_MixOneColumnInst_1_n7}), .b ({new_AGEMA_signal_7577, MixColumnsIns_MixOneColumnInst_1_n21}), .c ({new_AGEMA_signal_8026, MixColumnsOutput[79]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U27 ( .a ({new_AGEMA_signal_7469, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_7393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .c ({new_AGEMA_signal_7577, MixColumnsIns_MixOneColumnInst_1_n21}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U26 ( .a ({new_AGEMA_signal_7578, MixColumnsIns_MixOneColumnInst_1_n56}), .b ({new_AGEMA_signal_7427, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .c ({new_AGEMA_signal_7800, MixColumnsIns_MixOneColumnInst_1_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U25 ( .a ({new_AGEMA_signal_7470, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .b ({new_AGEMA_signal_7462, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .c ({new_AGEMA_signal_7578, MixColumnsIns_MixOneColumnInst_1_n56}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U24 ( .a ({new_AGEMA_signal_7801, MixColumnsIns_MixOneColumnInst_1_n6}), .b ({new_AGEMA_signal_7579, MixColumnsIns_MixOneColumnInst_1_n19}), .c ({new_AGEMA_signal_8027, MixColumnsOutput[78]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U23 ( .a ({new_AGEMA_signal_7470, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .b ({new_AGEMA_signal_7394, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .c ({new_AGEMA_signal_7579, MixColumnsIns_MixOneColumnInst_1_n19}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U22 ( .a ({new_AGEMA_signal_7580, MixColumnsIns_MixOneColumnInst_1_n53}), .b ({new_AGEMA_signal_7428, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .c ({new_AGEMA_signal_7801, MixColumnsIns_MixOneColumnInst_1_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U21 ( .a ({new_AGEMA_signal_7471, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .b ({new_AGEMA_signal_7463, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .c ({new_AGEMA_signal_7580, MixColumnsIns_MixOneColumnInst_1_n53}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U20 ( .a ({new_AGEMA_signal_7802, MixColumnsIns_MixOneColumnInst_1_n5}), .b ({new_AGEMA_signal_7581, MixColumnsIns_MixOneColumnInst_1_n17}), .c ({new_AGEMA_signal_8028, MixColumnsOutput[77]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U19 ( .a ({new_AGEMA_signal_7471, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .b ({new_AGEMA_signal_7395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .c ({new_AGEMA_signal_7581, MixColumnsIns_MixOneColumnInst_1_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U18 ( .a ({new_AGEMA_signal_7582, MixColumnsIns_MixOneColumnInst_1_n50}), .b ({new_AGEMA_signal_7429, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .c ({new_AGEMA_signal_7802, MixColumnsIns_MixOneColumnInst_1_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U17 ( .a ({new_AGEMA_signal_7472, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .b ({new_AGEMA_signal_7464, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .c ({new_AGEMA_signal_7582, MixColumnsIns_MixOneColumnInst_1_n50}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U16 ( .a ({new_AGEMA_signal_8029, MixColumnsIns_MixOneColumnInst_1_n4}), .b ({new_AGEMA_signal_7803, MixColumnsIns_MixOneColumnInst_1_n15}), .c ({new_AGEMA_signal_8292, MixColumnsOutput[76]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U15 ( .a ({new_AGEMA_signal_7472, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .b ({new_AGEMA_signal_7593, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]}), .c ({new_AGEMA_signal_7803, MixColumnsIns_MixOneColumnInst_1_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U14 ( .a ({new_AGEMA_signal_7804, MixColumnsIns_MixOneColumnInst_1_n47}), .b ({new_AGEMA_signal_7430, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .c ({new_AGEMA_signal_8029, MixColumnsIns_MixOneColumnInst_1_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U13 ( .a ({new_AGEMA_signal_7596, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]}), .b ({new_AGEMA_signal_7465, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .c ({new_AGEMA_signal_7804, MixColumnsIns_MixOneColumnInst_1_n47}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U12 ( .a ({new_AGEMA_signal_8030, MixColumnsIns_MixOneColumnInst_1_n3}), .b ({new_AGEMA_signal_7805, MixColumnsIns_MixOneColumnInst_1_n12}), .c ({new_AGEMA_signal_8293, MixColumnsOutput[75]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U11 ( .a ({new_AGEMA_signal_7473, MixColumnsInput[67]}), .b ({new_AGEMA_signal_7594, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]}), .c ({new_AGEMA_signal_7805, MixColumnsIns_MixOneColumnInst_1_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U10 ( .a ({new_AGEMA_signal_7806, MixColumnsIns_MixOneColumnInst_1_n44}), .b ({new_AGEMA_signal_7431, MixColumnsInput[83]}), .c ({new_AGEMA_signal_8030, MixColumnsIns_MixOneColumnInst_1_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U9 ( .a ({new_AGEMA_signal_7597, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]}), .b ({new_AGEMA_signal_7466, MixColumnsInput[91]}), .c ({new_AGEMA_signal_7806, MixColumnsIns_MixOneColumnInst_1_n44}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U8 ( .a ({new_AGEMA_signal_7807, MixColumnsIns_MixOneColumnInst_1_n2}), .b ({new_AGEMA_signal_7583, MixColumnsIns_MixOneColumnInst_1_n10}), .c ({new_AGEMA_signal_8031, MixColumnsOutput[74]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U7 ( .a ({new_AGEMA_signal_7474, MixColumnsInput[66]}), .b ({new_AGEMA_signal_7398, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .c ({new_AGEMA_signal_7583, MixColumnsIns_MixOneColumnInst_1_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U6 ( .a ({new_AGEMA_signal_7584, MixColumnsIns_MixOneColumnInst_1_n37}), .b ({new_AGEMA_signal_7432, MixColumnsInput[82]}), .c ({new_AGEMA_signal_7807, MixColumnsIns_MixOneColumnInst_1_n2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U5 ( .a ({new_AGEMA_signal_7475, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .b ({new_AGEMA_signal_7467, MixColumnsInput[90]}), .c ({new_AGEMA_signal_7584, MixColumnsIns_MixOneColumnInst_1_n37}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U4 ( .a ({new_AGEMA_signal_7808, MixColumnsIns_MixOneColumnInst_1_n1}), .b ({new_AGEMA_signal_7198, MixColumnsInput[72]}), .c ({new_AGEMA_signal_8032, MixColumnsOutput[64]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U3 ( .a ({new_AGEMA_signal_7586, MixColumnsIns_MixOneColumnInst_1_n59}), .b ({new_AGEMA_signal_7585, MixColumnsIns_MixOneColumnInst_1_n23}), .c ({new_AGEMA_signal_7808, MixColumnsIns_MixOneColumnInst_1_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U2 ( .a ({new_AGEMA_signal_7253, MixColumnsInput[80]}), .b ({new_AGEMA_signal_7462, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .c ({new_AGEMA_signal_7585, MixColumnsIns_MixOneColumnInst_1_n23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U1 ( .a ({new_AGEMA_signal_7469, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_7308, MixColumnsInput[88]}), .c ({new_AGEMA_signal_7586, MixColumnsIns_MixOneColumnInst_1_n59}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_7462, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_7466, MixColumnsInput[91]}), .c ({new_AGEMA_signal_7587, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_7462, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_7467, MixColumnsInput[90]}), .c ({new_AGEMA_signal_7588, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_7462, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_7308, MixColumnsInput[88]}), .c ({new_AGEMA_signal_7589, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_7427, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_7431, MixColumnsInput[83]}), .c ({new_AGEMA_signal_7590, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_7427, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_7432, MixColumnsInput[82]}), .c ({new_AGEMA_signal_7591, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_7427, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_7253, MixColumnsInput[80]}), .c ({new_AGEMA_signal_7592, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_7392, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_7396, MixColumnsInput[75]}), .c ({new_AGEMA_signal_7593, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_7392, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_7397, MixColumnsInput[74]}), .c ({new_AGEMA_signal_7594, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_7392, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_7198, MixColumnsInput[72]}), .c ({new_AGEMA_signal_7595, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_7469, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_7473, MixColumnsInput[67]}), .c ({new_AGEMA_signal_7596, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_7469, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_7474, MixColumnsInput[66]}), .c ({new_AGEMA_signal_7597, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_7469, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_7319, MixColumnsInput[64]}), .c ({new_AGEMA_signal_7598, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U96 ( .a ({new_AGEMA_signal_8033, MixColumnsIns_MixOneColumnInst_2_n64}), .b ({new_AGEMA_signal_7405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .c ({new_AGEMA_signal_8294, MixColumnsOutput[41]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U95 ( .a ({new_AGEMA_signal_7830, MixColumnsIns_MixOneColumnInst_2_n63}), .b ({new_AGEMA_signal_7826, MixColumnsIns_MixOneColumnInst_2_n62}), .c ({new_AGEMA_signal_8033, MixColumnsIns_MixOneColumnInst_2_n64}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U94 ( .a ({new_AGEMA_signal_7809, MixColumnsIns_MixOneColumnInst_2_n61}), .b ({new_AGEMA_signal_7608, MixColumnsIns_MixOneColumnInst_2_n60}), .c ({new_AGEMA_signal_8034, MixColumnsOutput[40]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U93 ( .a ({new_AGEMA_signal_7618, MixColumnsIns_MixOneColumnInst_2_n59}), .b ({new_AGEMA_signal_7209, MixColumnsInput[48]}), .c ({new_AGEMA_signal_7809, MixColumnsIns_MixOneColumnInst_2_n61}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U92 ( .a ({new_AGEMA_signal_7810, MixColumnsIns_MixOneColumnInst_2_n58}), .b ({new_AGEMA_signal_7599, MixColumnsIns_MixOneColumnInst_2_n57}), .c ({new_AGEMA_signal_8035, MixColumnsOutput[39]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U91 ( .a ({new_AGEMA_signal_7610, MixColumnsIns_MixOneColumnInst_2_n56}), .b ({new_AGEMA_signal_7476, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .c ({new_AGEMA_signal_7810, MixColumnsIns_MixOneColumnInst_2_n58}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U90 ( .a ({new_AGEMA_signal_7811, MixColumnsIns_MixOneColumnInst_2_n55}), .b ({new_AGEMA_signal_7600, MixColumnsIns_MixOneColumnInst_2_n54}), .c ({new_AGEMA_signal_8036, MixColumnsOutput[38]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U89 ( .a ({new_AGEMA_signal_7612, MixColumnsIns_MixOneColumnInst_2_n53}), .b ({new_AGEMA_signal_7477, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .c ({new_AGEMA_signal_7811, MixColumnsIns_MixOneColumnInst_2_n55}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U88 ( .a ({new_AGEMA_signal_7812, MixColumnsIns_MixOneColumnInst_2_n52}), .b ({new_AGEMA_signal_7601, MixColumnsIns_MixOneColumnInst_2_n51}), .c ({new_AGEMA_signal_8037, MixColumnsOutput[37]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U87 ( .a ({new_AGEMA_signal_7614, MixColumnsIns_MixOneColumnInst_2_n50}), .b ({new_AGEMA_signal_7478, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .c ({new_AGEMA_signal_7812, MixColumnsIns_MixOneColumnInst_2_n52}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U86 ( .a ({new_AGEMA_signal_8038, MixColumnsIns_MixOneColumnInst_2_n49}), .b ({new_AGEMA_signal_7817, MixColumnsIns_MixOneColumnInst_2_n48}), .c ({new_AGEMA_signal_8295, MixColumnsOutput[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U85 ( .a ({new_AGEMA_signal_7836, MixColumnsIns_MixOneColumnInst_2_n47}), .b ({new_AGEMA_signal_7479, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .c ({new_AGEMA_signal_8038, MixColumnsIns_MixOneColumnInst_2_n49}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U84 ( .a ({new_AGEMA_signal_8039, MixColumnsIns_MixOneColumnInst_2_n46}), .b ({new_AGEMA_signal_7818, MixColumnsIns_MixOneColumnInst_2_n45}), .c ({new_AGEMA_signal_8296, MixColumnsOutput[35]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U83 ( .a ({new_AGEMA_signal_7838, MixColumnsIns_MixOneColumnInst_2_n44}), .b ({new_AGEMA_signal_7480, MixColumnsInput[43]}), .c ({new_AGEMA_signal_8039, MixColumnsIns_MixOneColumnInst_2_n46}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U82 ( .a ({new_AGEMA_signal_7813, MixColumnsIns_MixOneColumnInst_2_n43}), .b ({new_AGEMA_signal_7599, MixColumnsIns_MixOneColumnInst_2_n57}), .c ({new_AGEMA_signal_8040, MixColumnsOutput[63]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U81 ( .a ({new_AGEMA_signal_7399, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_7435, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .c ({new_AGEMA_signal_7599, MixColumnsIns_MixOneColumnInst_2_n57}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U80 ( .a ({new_AGEMA_signal_7441, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_7603, MixColumnsIns_MixOneColumnInst_2_n42}), .c ({new_AGEMA_signal_7813, MixColumnsIns_MixOneColumnInst_2_n43}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U79 ( .a ({new_AGEMA_signal_7814, MixColumnsIns_MixOneColumnInst_2_n41}), .b ({new_AGEMA_signal_7600, MixColumnsIns_MixOneColumnInst_2_n54}), .c ({new_AGEMA_signal_8041, MixColumnsOutput[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U78 ( .a ({new_AGEMA_signal_7400, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .b ({new_AGEMA_signal_7436, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .c ({new_AGEMA_signal_7600, MixColumnsIns_MixOneColumnInst_2_n54}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U77 ( .a ({new_AGEMA_signal_7442, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .b ({new_AGEMA_signal_7604, MixColumnsIns_MixOneColumnInst_2_n40}), .c ({new_AGEMA_signal_7814, MixColumnsIns_MixOneColumnInst_2_n41}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U76 ( .a ({new_AGEMA_signal_7815, MixColumnsIns_MixOneColumnInst_2_n39}), .b ({new_AGEMA_signal_7602, MixColumnsIns_MixOneColumnInst_2_n38}), .c ({new_AGEMA_signal_8042, MixColumnsOutput[34]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U75 ( .a ({new_AGEMA_signal_7616, MixColumnsIns_MixOneColumnInst_2_n37}), .b ({new_AGEMA_signal_7481, MixColumnsInput[42]}), .c ({new_AGEMA_signal_7815, MixColumnsIns_MixOneColumnInst_2_n39}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U74 ( .a ({new_AGEMA_signal_7816, MixColumnsIns_MixOneColumnInst_2_n36}), .b ({new_AGEMA_signal_7601, MixColumnsIns_MixOneColumnInst_2_n51}), .c ({new_AGEMA_signal_8043, MixColumnsOutput[61]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U73 ( .a ({new_AGEMA_signal_7401, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .b ({new_AGEMA_signal_7437, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .c ({new_AGEMA_signal_7601, MixColumnsIns_MixOneColumnInst_2_n51}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U72 ( .a ({new_AGEMA_signal_7443, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .b ({new_AGEMA_signal_7605, MixColumnsIns_MixOneColumnInst_2_n35}), .c ({new_AGEMA_signal_7816, MixColumnsIns_MixOneColumnInst_2_n36}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U71 ( .a ({new_AGEMA_signal_8044, MixColumnsIns_MixOneColumnInst_2_n34}), .b ({new_AGEMA_signal_7817, MixColumnsIns_MixOneColumnInst_2_n48}), .c ({new_AGEMA_signal_8297, MixColumnsOutput[60]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U70 ( .a ({new_AGEMA_signal_7402, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .b ({new_AGEMA_signal_7619, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]}), .c ({new_AGEMA_signal_7817, MixColumnsIns_MixOneColumnInst_2_n48}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U69 ( .a ({new_AGEMA_signal_7444, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .b ({new_AGEMA_signal_7824, MixColumnsIns_MixOneColumnInst_2_n33}), .c ({new_AGEMA_signal_8044, MixColumnsIns_MixOneColumnInst_2_n34}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U68 ( .a ({new_AGEMA_signal_8045, MixColumnsIns_MixOneColumnInst_2_n32}), .b ({new_AGEMA_signal_7818, MixColumnsIns_MixOneColumnInst_2_n45}), .c ({new_AGEMA_signal_8298, MixColumnsOutput[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U67 ( .a ({new_AGEMA_signal_7403, MixColumnsInput[51]}), .b ({new_AGEMA_signal_7620, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]}), .c ({new_AGEMA_signal_7818, MixColumnsIns_MixOneColumnInst_2_n45}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U66 ( .a ({new_AGEMA_signal_7445, MixColumnsInput[35]}), .b ({new_AGEMA_signal_7827, MixColumnsIns_MixOneColumnInst_2_n31}), .c ({new_AGEMA_signal_8045, MixColumnsIns_MixOneColumnInst_2_n32}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U65 ( .a ({new_AGEMA_signal_7819, MixColumnsIns_MixOneColumnInst_2_n30}), .b ({new_AGEMA_signal_7602, MixColumnsIns_MixOneColumnInst_2_n38}), .c ({new_AGEMA_signal_8046, MixColumnsOutput[58]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U64 ( .a ({new_AGEMA_signal_7404, MixColumnsInput[50]}), .b ({new_AGEMA_signal_7440, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .c ({new_AGEMA_signal_7602, MixColumnsIns_MixOneColumnInst_2_n38}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U63 ( .a ({new_AGEMA_signal_7446, MixColumnsInput[34]}), .b ({new_AGEMA_signal_7606, MixColumnsIns_MixOneColumnInst_2_n29}), .c ({new_AGEMA_signal_7819, MixColumnsIns_MixOneColumnInst_2_n30}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U62 ( .a ({new_AGEMA_signal_8047, MixColumnsIns_MixOneColumnInst_2_n28}), .b ({new_AGEMA_signal_7825, MixColumnsIns_MixOneColumnInst_2_n27}), .c ({new_AGEMA_signal_8299, MixColumnsOutput[57]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U61 ( .a ({new_AGEMA_signal_7447, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .b ({new_AGEMA_signal_7829, MixColumnsIns_MixOneColumnInst_2_n26}), .c ({new_AGEMA_signal_8047, MixColumnsIns_MixOneColumnInst_2_n28}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U60 ( .a ({new_AGEMA_signal_7820, MixColumnsIns_MixOneColumnInst_2_n25}), .b ({new_AGEMA_signal_7607, MixColumnsIns_MixOneColumnInst_2_n24}), .c ({new_AGEMA_signal_8048, MixColumnsOutput[56]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U59 ( .a ({new_AGEMA_signal_7617, MixColumnsIns_MixOneColumnInst_2_n23}), .b ({new_AGEMA_signal_7275, MixColumnsInput[32]}), .c ({new_AGEMA_signal_7820, MixColumnsIns_MixOneColumnInst_2_n25}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U58 ( .a ({new_AGEMA_signal_7821, MixColumnsIns_MixOneColumnInst_2_n22}), .b ({new_AGEMA_signal_7603, MixColumnsIns_MixOneColumnInst_2_n42}), .c ({new_AGEMA_signal_8049, MixColumnsOutput[55]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U57 ( .a ({new_AGEMA_signal_7476, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_7400, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .c ({new_AGEMA_signal_7603, MixColumnsIns_MixOneColumnInst_2_n42}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U56 ( .a ({new_AGEMA_signal_7434, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_7609, MixColumnsIns_MixOneColumnInst_2_n21}), .c ({new_AGEMA_signal_7821, MixColumnsIns_MixOneColumnInst_2_n22}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U55 ( .a ({new_AGEMA_signal_7822, MixColumnsIns_MixOneColumnInst_2_n20}), .b ({new_AGEMA_signal_7604, MixColumnsIns_MixOneColumnInst_2_n40}), .c ({new_AGEMA_signal_8050, MixColumnsOutput[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U54 ( .a ({new_AGEMA_signal_7477, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .b ({new_AGEMA_signal_7401, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .c ({new_AGEMA_signal_7604, MixColumnsIns_MixOneColumnInst_2_n40}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U53 ( .a ({new_AGEMA_signal_7435, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .b ({new_AGEMA_signal_7611, MixColumnsIns_MixOneColumnInst_2_n19}), .c ({new_AGEMA_signal_7822, MixColumnsIns_MixOneColumnInst_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U52 ( .a ({new_AGEMA_signal_7823, MixColumnsIns_MixOneColumnInst_2_n18}), .b ({new_AGEMA_signal_7605, MixColumnsIns_MixOneColumnInst_2_n35}), .c ({new_AGEMA_signal_8051, MixColumnsOutput[53]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U51 ( .a ({new_AGEMA_signal_7478, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .b ({new_AGEMA_signal_7402, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .c ({new_AGEMA_signal_7605, MixColumnsIns_MixOneColumnInst_2_n35}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U50 ( .a ({new_AGEMA_signal_7436, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .b ({new_AGEMA_signal_7613, MixColumnsIns_MixOneColumnInst_2_n17}), .c ({new_AGEMA_signal_7823, MixColumnsIns_MixOneColumnInst_2_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U49 ( .a ({new_AGEMA_signal_8052, MixColumnsIns_MixOneColumnInst_2_n16}), .b ({new_AGEMA_signal_7824, MixColumnsIns_MixOneColumnInst_2_n33}), .c ({new_AGEMA_signal_8300, MixColumnsOutput[52]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U48 ( .a ({new_AGEMA_signal_7479, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .b ({new_AGEMA_signal_7622, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]}), .c ({new_AGEMA_signal_7824, MixColumnsIns_MixOneColumnInst_2_n33}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U47 ( .a ({new_AGEMA_signal_7437, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .b ({new_AGEMA_signal_7835, MixColumnsIns_MixOneColumnInst_2_n15}), .c ({new_AGEMA_signal_8052, MixColumnsIns_MixOneColumnInst_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U46 ( .a ({new_AGEMA_signal_8053, MixColumnsIns_MixOneColumnInst_2_n14}), .b ({new_AGEMA_signal_7825, MixColumnsIns_MixOneColumnInst_2_n27}), .c ({new_AGEMA_signal_8301, MixColumnsOutput[33]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U45 ( .a ({new_AGEMA_signal_7405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .b ({new_AGEMA_signal_7621, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]}), .c ({new_AGEMA_signal_7825, MixColumnsIns_MixOneColumnInst_2_n27}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U44 ( .a ({new_AGEMA_signal_7482, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .b ({new_AGEMA_signal_7826, MixColumnsIns_MixOneColumnInst_2_n62}), .c ({new_AGEMA_signal_8053, MixColumnsIns_MixOneColumnInst_2_n14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U43 ( .a ({new_AGEMA_signal_7440, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .b ({new_AGEMA_signal_7630, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]}), .c ({new_AGEMA_signal_7826, MixColumnsIns_MixOneColumnInst_2_n62}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U42 ( .a ({new_AGEMA_signal_8054, MixColumnsIns_MixOneColumnInst_2_n13}), .b ({new_AGEMA_signal_7827, MixColumnsIns_MixOneColumnInst_2_n31}), .c ({new_AGEMA_signal_8302, MixColumnsOutput[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U41 ( .a ({new_AGEMA_signal_7480, MixColumnsInput[43]}), .b ({new_AGEMA_signal_7623, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]}), .c ({new_AGEMA_signal_7827, MixColumnsIns_MixOneColumnInst_2_n31}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U40 ( .a ({new_AGEMA_signal_7438, MixColumnsInput[59]}), .b ({new_AGEMA_signal_7837, MixColumnsIns_MixOneColumnInst_2_n12}), .c ({new_AGEMA_signal_8054, MixColumnsIns_MixOneColumnInst_2_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U39 ( .a ({new_AGEMA_signal_7828, MixColumnsIns_MixOneColumnInst_2_n11}), .b ({new_AGEMA_signal_7606, MixColumnsIns_MixOneColumnInst_2_n29}), .c ({new_AGEMA_signal_8055, MixColumnsOutput[50]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U38 ( .a ({new_AGEMA_signal_7481, MixColumnsInput[42]}), .b ({new_AGEMA_signal_7405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .c ({new_AGEMA_signal_7606, MixColumnsIns_MixOneColumnInst_2_n29}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U37 ( .a ({new_AGEMA_signal_7439, MixColumnsInput[58]}), .b ({new_AGEMA_signal_7615, MixColumnsIns_MixOneColumnInst_2_n10}), .c ({new_AGEMA_signal_7828, MixColumnsIns_MixOneColumnInst_2_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U36 ( .a ({new_AGEMA_signal_8056, MixColumnsIns_MixOneColumnInst_2_n9}), .b ({new_AGEMA_signal_7829, MixColumnsIns_MixOneColumnInst_2_n26}), .c ({new_AGEMA_signal_8303, MixColumnsOutput[49]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U35 ( .a ({new_AGEMA_signal_7624, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]}), .b ({new_AGEMA_signal_7482, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .c ({new_AGEMA_signal_7829, MixColumnsIns_MixOneColumnInst_2_n26}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U34 ( .a ({new_AGEMA_signal_7830, MixColumnsIns_MixOneColumnInst_2_n63}), .b ({new_AGEMA_signal_7440, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .c ({new_AGEMA_signal_8056, MixColumnsIns_MixOneColumnInst_2_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U33 ( .a ({new_AGEMA_signal_7627, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]}), .b ({new_AGEMA_signal_7447, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .c ({new_AGEMA_signal_7830, MixColumnsIns_MixOneColumnInst_2_n63}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U32 ( .a ({new_AGEMA_signal_7831, MixColumnsIns_MixOneColumnInst_2_n8}), .b ({new_AGEMA_signal_7607, MixColumnsIns_MixOneColumnInst_2_n24}), .c ({new_AGEMA_signal_8057, MixColumnsOutput[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U31 ( .a ({new_AGEMA_signal_7330, MixColumnsInput[40]}), .b ({new_AGEMA_signal_7399, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .c ({new_AGEMA_signal_7607, MixColumnsIns_MixOneColumnInst_2_n24}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U30 ( .a ({new_AGEMA_signal_7264, MixColumnsInput[56]}), .b ({new_AGEMA_signal_7608, MixColumnsIns_MixOneColumnInst_2_n60}), .c ({new_AGEMA_signal_7831, MixColumnsIns_MixOneColumnInst_2_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U29 ( .a ({new_AGEMA_signal_7476, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_7275, MixColumnsInput[32]}), .c ({new_AGEMA_signal_7608, MixColumnsIns_MixOneColumnInst_2_n60}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U28 ( .a ({new_AGEMA_signal_7832, MixColumnsIns_MixOneColumnInst_2_n7}), .b ({new_AGEMA_signal_7609, MixColumnsIns_MixOneColumnInst_2_n21}), .c ({new_AGEMA_signal_8058, MixColumnsOutput[47]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U27 ( .a ({new_AGEMA_signal_7441, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_7477, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .c ({new_AGEMA_signal_7609, MixColumnsIns_MixOneColumnInst_2_n21}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U26 ( .a ({new_AGEMA_signal_7610, MixColumnsIns_MixOneColumnInst_2_n56}), .b ({new_AGEMA_signal_7399, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .c ({new_AGEMA_signal_7832, MixColumnsIns_MixOneColumnInst_2_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U25 ( .a ({new_AGEMA_signal_7442, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .b ({new_AGEMA_signal_7434, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .c ({new_AGEMA_signal_7610, MixColumnsIns_MixOneColumnInst_2_n56}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U24 ( .a ({new_AGEMA_signal_7833, MixColumnsIns_MixOneColumnInst_2_n6}), .b ({new_AGEMA_signal_7611, MixColumnsIns_MixOneColumnInst_2_n19}), .c ({new_AGEMA_signal_8059, MixColumnsOutput[46]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U23 ( .a ({new_AGEMA_signal_7442, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .b ({new_AGEMA_signal_7478, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .c ({new_AGEMA_signal_7611, MixColumnsIns_MixOneColumnInst_2_n19}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U22 ( .a ({new_AGEMA_signal_7612, MixColumnsIns_MixOneColumnInst_2_n53}), .b ({new_AGEMA_signal_7400, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .c ({new_AGEMA_signal_7833, MixColumnsIns_MixOneColumnInst_2_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U21 ( .a ({new_AGEMA_signal_7443, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .b ({new_AGEMA_signal_7435, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .c ({new_AGEMA_signal_7612, MixColumnsIns_MixOneColumnInst_2_n53}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U20 ( .a ({new_AGEMA_signal_7834, MixColumnsIns_MixOneColumnInst_2_n5}), .b ({new_AGEMA_signal_7613, MixColumnsIns_MixOneColumnInst_2_n17}), .c ({new_AGEMA_signal_8060, MixColumnsOutput[45]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U19 ( .a ({new_AGEMA_signal_7443, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .b ({new_AGEMA_signal_7479, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .c ({new_AGEMA_signal_7613, MixColumnsIns_MixOneColumnInst_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U18 ( .a ({new_AGEMA_signal_7614, MixColumnsIns_MixOneColumnInst_2_n50}), .b ({new_AGEMA_signal_7401, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .c ({new_AGEMA_signal_7834, MixColumnsIns_MixOneColumnInst_2_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U17 ( .a ({new_AGEMA_signal_7444, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .b ({new_AGEMA_signal_7436, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .c ({new_AGEMA_signal_7614, MixColumnsIns_MixOneColumnInst_2_n50}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U16 ( .a ({new_AGEMA_signal_8061, MixColumnsIns_MixOneColumnInst_2_n4}), .b ({new_AGEMA_signal_7835, MixColumnsIns_MixOneColumnInst_2_n15}), .c ({new_AGEMA_signal_8304, MixColumnsOutput[44]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U15 ( .a ({new_AGEMA_signal_7444, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .b ({new_AGEMA_signal_7625, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]}), .c ({new_AGEMA_signal_7835, MixColumnsIns_MixOneColumnInst_2_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U14 ( .a ({new_AGEMA_signal_7836, MixColumnsIns_MixOneColumnInst_2_n47}), .b ({new_AGEMA_signal_7402, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .c ({new_AGEMA_signal_8061, MixColumnsIns_MixOneColumnInst_2_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U13 ( .a ({new_AGEMA_signal_7628, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]}), .b ({new_AGEMA_signal_7437, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .c ({new_AGEMA_signal_7836, MixColumnsIns_MixOneColumnInst_2_n47}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U12 ( .a ({new_AGEMA_signal_8062, MixColumnsIns_MixOneColumnInst_2_n3}), .b ({new_AGEMA_signal_7837, MixColumnsIns_MixOneColumnInst_2_n12}), .c ({new_AGEMA_signal_8305, MixColumnsOutput[43]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U11 ( .a ({new_AGEMA_signal_7445, MixColumnsInput[35]}), .b ({new_AGEMA_signal_7626, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]}), .c ({new_AGEMA_signal_7837, MixColumnsIns_MixOneColumnInst_2_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U10 ( .a ({new_AGEMA_signal_7838, MixColumnsIns_MixOneColumnInst_2_n44}), .b ({new_AGEMA_signal_7403, MixColumnsInput[51]}), .c ({new_AGEMA_signal_8062, MixColumnsIns_MixOneColumnInst_2_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U9 ( .a ({new_AGEMA_signal_7629, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]}), .b ({new_AGEMA_signal_7438, MixColumnsInput[59]}), .c ({new_AGEMA_signal_7838, MixColumnsIns_MixOneColumnInst_2_n44}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U8 ( .a ({new_AGEMA_signal_7839, MixColumnsIns_MixOneColumnInst_2_n2}), .b ({new_AGEMA_signal_7615, MixColumnsIns_MixOneColumnInst_2_n10}), .c ({new_AGEMA_signal_8063, MixColumnsOutput[42]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U7 ( .a ({new_AGEMA_signal_7446, MixColumnsInput[34]}), .b ({new_AGEMA_signal_7482, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .c ({new_AGEMA_signal_7615, MixColumnsIns_MixOneColumnInst_2_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U6 ( .a ({new_AGEMA_signal_7616, MixColumnsIns_MixOneColumnInst_2_n37}), .b ({new_AGEMA_signal_7404, MixColumnsInput[50]}), .c ({new_AGEMA_signal_7839, MixColumnsIns_MixOneColumnInst_2_n2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U5 ( .a ({new_AGEMA_signal_7447, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .b ({new_AGEMA_signal_7439, MixColumnsInput[58]}), .c ({new_AGEMA_signal_7616, MixColumnsIns_MixOneColumnInst_2_n37}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U4 ( .a ({new_AGEMA_signal_7840, MixColumnsIns_MixOneColumnInst_2_n1}), .b ({new_AGEMA_signal_7330, MixColumnsInput[40]}), .c ({new_AGEMA_signal_8064, MixColumnsOutput[32]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U3 ( .a ({new_AGEMA_signal_7618, MixColumnsIns_MixOneColumnInst_2_n59}), .b ({new_AGEMA_signal_7617, MixColumnsIns_MixOneColumnInst_2_n23}), .c ({new_AGEMA_signal_7840, MixColumnsIns_MixOneColumnInst_2_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U2 ( .a ({new_AGEMA_signal_7209, MixColumnsInput[48]}), .b ({new_AGEMA_signal_7434, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .c ({new_AGEMA_signal_7617, MixColumnsIns_MixOneColumnInst_2_n23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U1 ( .a ({new_AGEMA_signal_7441, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_7264, MixColumnsInput[56]}), .c ({new_AGEMA_signal_7618, MixColumnsIns_MixOneColumnInst_2_n59}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_7434, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_7438, MixColumnsInput[59]}), .c ({new_AGEMA_signal_7619, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_7434, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_7439, MixColumnsInput[58]}), .c ({new_AGEMA_signal_7620, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_7434, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_7264, MixColumnsInput[56]}), .c ({new_AGEMA_signal_7621, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_7399, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_7403, MixColumnsInput[51]}), .c ({new_AGEMA_signal_7622, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_7399, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_7404, MixColumnsInput[50]}), .c ({new_AGEMA_signal_7623, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_7399, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_7209, MixColumnsInput[48]}), .c ({new_AGEMA_signal_7624, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_7476, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_7480, MixColumnsInput[43]}), .c ({new_AGEMA_signal_7625, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_7476, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_7481, MixColumnsInput[42]}), .c ({new_AGEMA_signal_7626, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_7476, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_7330, MixColumnsInput[40]}), .c ({new_AGEMA_signal_7627, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_7441, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_7445, MixColumnsInput[35]}), .c ({new_AGEMA_signal_7628, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_7441, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_7446, MixColumnsInput[34]}), .c ({new_AGEMA_signal_7629, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_7441, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_7275, MixColumnsInput[32]}), .c ({new_AGEMA_signal_7630, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U96 ( .a ({new_AGEMA_signal_8065, MixColumnsIns_MixOneColumnInst_3_n64}), .b ({new_AGEMA_signal_7489, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .c ({new_AGEMA_signal_8306, MixColumnsOutput[9]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U95 ( .a ({new_AGEMA_signal_7862, MixColumnsIns_MixOneColumnInst_3_n63}), .b ({new_AGEMA_signal_7858, MixColumnsIns_MixOneColumnInst_3_n62}), .c ({new_AGEMA_signal_8065, MixColumnsIns_MixOneColumnInst_3_n64}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U94 ( .a ({new_AGEMA_signal_7841, MixColumnsIns_MixOneColumnInst_3_n61}), .b ({new_AGEMA_signal_7640, MixColumnsIns_MixOneColumnInst_3_n60}), .c ({new_AGEMA_signal_8066, MixColumnsOutput[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U93 ( .a ({new_AGEMA_signal_7650, MixColumnsIns_MixOneColumnInst_3_n59}), .b ({new_AGEMA_signal_7341, MixColumnsInput[16]}), .c ({new_AGEMA_signal_7841, MixColumnsIns_MixOneColumnInst_3_n61}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U92 ( .a ({new_AGEMA_signal_7842, MixColumnsIns_MixOneColumnInst_3_n58}), .b ({new_AGEMA_signal_7631, MixColumnsIns_MixOneColumnInst_3_n57}), .c ({new_AGEMA_signal_8067, MixColumnsOutput[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U91 ( .a ({new_AGEMA_signal_7642, MixColumnsIns_MixOneColumnInst_3_n56}), .b ({new_AGEMA_signal_7448, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .c ({new_AGEMA_signal_7842, MixColumnsIns_MixOneColumnInst_3_n58}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U90 ( .a ({new_AGEMA_signal_7843, MixColumnsIns_MixOneColumnInst_3_n55}), .b ({new_AGEMA_signal_7632, MixColumnsIns_MixOneColumnInst_3_n54}), .c ({new_AGEMA_signal_8068, MixColumnsOutput[6]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U89 ( .a ({new_AGEMA_signal_7644, MixColumnsIns_MixOneColumnInst_3_n53}), .b ({new_AGEMA_signal_7449, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .c ({new_AGEMA_signal_7843, MixColumnsIns_MixOneColumnInst_3_n55}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U88 ( .a ({new_AGEMA_signal_7844, MixColumnsIns_MixOneColumnInst_3_n52}), .b ({new_AGEMA_signal_7633, MixColumnsIns_MixOneColumnInst_3_n51}), .c ({new_AGEMA_signal_8069, MixColumnsOutput[5]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U87 ( .a ({new_AGEMA_signal_7646, MixColumnsIns_MixOneColumnInst_3_n50}), .b ({new_AGEMA_signal_7450, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .c ({new_AGEMA_signal_7844, MixColumnsIns_MixOneColumnInst_3_n52}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U86 ( .a ({new_AGEMA_signal_8070, MixColumnsIns_MixOneColumnInst_3_n49}), .b ({new_AGEMA_signal_7849, MixColumnsIns_MixOneColumnInst_3_n48}), .c ({new_AGEMA_signal_8307, MixColumnsOutput[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U85 ( .a ({new_AGEMA_signal_7868, MixColumnsIns_MixOneColumnInst_3_n47}), .b ({new_AGEMA_signal_7451, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .c ({new_AGEMA_signal_8070, MixColumnsIns_MixOneColumnInst_3_n49}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U84 ( .a ({new_AGEMA_signal_8071, MixColumnsIns_MixOneColumnInst_3_n46}), .b ({new_AGEMA_signal_7850, MixColumnsIns_MixOneColumnInst_3_n45}), .c ({new_AGEMA_signal_8308, MixColumnsOutput[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U83 ( .a ({new_AGEMA_signal_7870, MixColumnsIns_MixOneColumnInst_3_n44}), .b ({new_AGEMA_signal_7452, MixColumnsInput[11]}), .c ({new_AGEMA_signal_8071, MixColumnsIns_MixOneColumnInst_3_n46}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U82 ( .a ({new_AGEMA_signal_7845, MixColumnsIns_MixOneColumnInst_3_n43}), .b ({new_AGEMA_signal_7631, MixColumnsIns_MixOneColumnInst_3_n57}), .c ({new_AGEMA_signal_8072, MixColumnsOutput[31]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U81 ( .a ({new_AGEMA_signal_7483, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_7407, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .c ({new_AGEMA_signal_7631, MixColumnsIns_MixOneColumnInst_3_n57}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U80 ( .a ({new_AGEMA_signal_7413, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_7635, MixColumnsIns_MixOneColumnInst_3_n42}), .c ({new_AGEMA_signal_7845, MixColumnsIns_MixOneColumnInst_3_n43}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U79 ( .a ({new_AGEMA_signal_7846, MixColumnsIns_MixOneColumnInst_3_n41}), .b ({new_AGEMA_signal_7632, MixColumnsIns_MixOneColumnInst_3_n54}), .c ({new_AGEMA_signal_8073, MixColumnsOutput[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U78 ( .a ({new_AGEMA_signal_7484, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .b ({new_AGEMA_signal_7408, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .c ({new_AGEMA_signal_7632, MixColumnsIns_MixOneColumnInst_3_n54}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U77 ( .a ({new_AGEMA_signal_7414, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .b ({new_AGEMA_signal_7636, MixColumnsIns_MixOneColumnInst_3_n40}), .c ({new_AGEMA_signal_7846, MixColumnsIns_MixOneColumnInst_3_n41}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U76 ( .a ({new_AGEMA_signal_7847, MixColumnsIns_MixOneColumnInst_3_n39}), .b ({new_AGEMA_signal_7634, MixColumnsIns_MixOneColumnInst_3_n38}), .c ({new_AGEMA_signal_8074, MixColumnsOutput[2]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U75 ( .a ({new_AGEMA_signal_7648, MixColumnsIns_MixOneColumnInst_3_n37}), .b ({new_AGEMA_signal_7453, MixColumnsInput[10]}), .c ({new_AGEMA_signal_7847, MixColumnsIns_MixOneColumnInst_3_n39}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U74 ( .a ({new_AGEMA_signal_7848, MixColumnsIns_MixOneColumnInst_3_n36}), .b ({new_AGEMA_signal_7633, MixColumnsIns_MixOneColumnInst_3_n51}), .c ({new_AGEMA_signal_8075, MixColumnsOutput[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U73 ( .a ({new_AGEMA_signal_7485, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .b ({new_AGEMA_signal_7409, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .c ({new_AGEMA_signal_7633, MixColumnsIns_MixOneColumnInst_3_n51}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U72 ( .a ({new_AGEMA_signal_7415, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .b ({new_AGEMA_signal_7637, MixColumnsIns_MixOneColumnInst_3_n35}), .c ({new_AGEMA_signal_7848, MixColumnsIns_MixOneColumnInst_3_n36}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U71 ( .a ({new_AGEMA_signal_8076, MixColumnsIns_MixOneColumnInst_3_n34}), .b ({new_AGEMA_signal_7849, MixColumnsIns_MixOneColumnInst_3_n48}), .c ({new_AGEMA_signal_8309, MixColumnsOutput[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U70 ( .a ({new_AGEMA_signal_7486, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .b ({new_AGEMA_signal_7651, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]}), .c ({new_AGEMA_signal_7849, MixColumnsIns_MixOneColumnInst_3_n48}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U69 ( .a ({new_AGEMA_signal_7416, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .b ({new_AGEMA_signal_7856, MixColumnsIns_MixOneColumnInst_3_n33}), .c ({new_AGEMA_signal_8076, MixColumnsIns_MixOneColumnInst_3_n34}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U68 ( .a ({new_AGEMA_signal_8077, MixColumnsIns_MixOneColumnInst_3_n32}), .b ({new_AGEMA_signal_7850, MixColumnsIns_MixOneColumnInst_3_n45}), .c ({new_AGEMA_signal_8310, MixColumnsOutput[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U67 ( .a ({new_AGEMA_signal_7487, MixColumnsInput[19]}), .b ({new_AGEMA_signal_7652, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]}), .c ({new_AGEMA_signal_7850, MixColumnsIns_MixOneColumnInst_3_n45}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U66 ( .a ({new_AGEMA_signal_7417, MixColumnsInput[3]}), .b ({new_AGEMA_signal_7859, MixColumnsIns_MixOneColumnInst_3_n31}), .c ({new_AGEMA_signal_8077, MixColumnsIns_MixOneColumnInst_3_n32}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U65 ( .a ({new_AGEMA_signal_7851, MixColumnsIns_MixOneColumnInst_3_n30}), .b ({new_AGEMA_signal_7634, MixColumnsIns_MixOneColumnInst_3_n38}), .c ({new_AGEMA_signal_8078, MixColumnsOutput[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U64 ( .a ({new_AGEMA_signal_7488, MixColumnsInput[18]}), .b ({new_AGEMA_signal_7412, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .c ({new_AGEMA_signal_7634, MixColumnsIns_MixOneColumnInst_3_n38}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U63 ( .a ({new_AGEMA_signal_7418, MixColumnsInput[2]}), .b ({new_AGEMA_signal_7638, MixColumnsIns_MixOneColumnInst_3_n29}), .c ({new_AGEMA_signal_7851, MixColumnsIns_MixOneColumnInst_3_n30}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U62 ( .a ({new_AGEMA_signal_8079, MixColumnsIns_MixOneColumnInst_3_n28}), .b ({new_AGEMA_signal_7857, MixColumnsIns_MixOneColumnInst_3_n27}), .c ({new_AGEMA_signal_8311, MixColumnsOutput[25]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U61 ( .a ({new_AGEMA_signal_7419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .b ({new_AGEMA_signal_7861, MixColumnsIns_MixOneColumnInst_3_n26}), .c ({new_AGEMA_signal_8079, MixColumnsIns_MixOneColumnInst_3_n28}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U60 ( .a ({new_AGEMA_signal_7852, MixColumnsIns_MixOneColumnInst_3_n25}), .b ({new_AGEMA_signal_7639, MixColumnsIns_MixOneColumnInst_3_n24}), .c ({new_AGEMA_signal_8080, MixColumnsOutput[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U59 ( .a ({new_AGEMA_signal_7649, MixColumnsIns_MixOneColumnInst_3_n23}), .b ({new_AGEMA_signal_7231, MixColumnsInput[0]}), .c ({new_AGEMA_signal_7852, MixColumnsIns_MixOneColumnInst_3_n25}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U58 ( .a ({new_AGEMA_signal_7853, MixColumnsIns_MixOneColumnInst_3_n22}), .b ({new_AGEMA_signal_7635, MixColumnsIns_MixOneColumnInst_3_n42}), .c ({new_AGEMA_signal_8081, MixColumnsOutput[23]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U57 ( .a ({new_AGEMA_signal_7448, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_7484, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .c ({new_AGEMA_signal_7635, MixColumnsIns_MixOneColumnInst_3_n42}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U56 ( .a ({new_AGEMA_signal_7406, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_7641, MixColumnsIns_MixOneColumnInst_3_n21}), .c ({new_AGEMA_signal_7853, MixColumnsIns_MixOneColumnInst_3_n22}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U55 ( .a ({new_AGEMA_signal_7854, MixColumnsIns_MixOneColumnInst_3_n20}), .b ({new_AGEMA_signal_7636, MixColumnsIns_MixOneColumnInst_3_n40}), .c ({new_AGEMA_signal_8082, MixColumnsOutput[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U54 ( .a ({new_AGEMA_signal_7449, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .b ({new_AGEMA_signal_7485, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .c ({new_AGEMA_signal_7636, MixColumnsIns_MixOneColumnInst_3_n40}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U53 ( .a ({new_AGEMA_signal_7407, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .b ({new_AGEMA_signal_7643, MixColumnsIns_MixOneColumnInst_3_n19}), .c ({new_AGEMA_signal_7854, MixColumnsIns_MixOneColumnInst_3_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U52 ( .a ({new_AGEMA_signal_7855, MixColumnsIns_MixOneColumnInst_3_n18}), .b ({new_AGEMA_signal_7637, MixColumnsIns_MixOneColumnInst_3_n35}), .c ({new_AGEMA_signal_8083, MixColumnsOutput[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U51 ( .a ({new_AGEMA_signal_7450, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .b ({new_AGEMA_signal_7486, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .c ({new_AGEMA_signal_7637, MixColumnsIns_MixOneColumnInst_3_n35}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U50 ( .a ({new_AGEMA_signal_7408, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .b ({new_AGEMA_signal_7645, MixColumnsIns_MixOneColumnInst_3_n17}), .c ({new_AGEMA_signal_7855, MixColumnsIns_MixOneColumnInst_3_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U49 ( .a ({new_AGEMA_signal_8084, MixColumnsIns_MixOneColumnInst_3_n16}), .b ({new_AGEMA_signal_7856, MixColumnsIns_MixOneColumnInst_3_n33}), .c ({new_AGEMA_signal_8312, MixColumnsOutput[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U48 ( .a ({new_AGEMA_signal_7451, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .b ({new_AGEMA_signal_7654, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]}), .c ({new_AGEMA_signal_7856, MixColumnsIns_MixOneColumnInst_3_n33}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U47 ( .a ({new_AGEMA_signal_7409, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .b ({new_AGEMA_signal_7867, MixColumnsIns_MixOneColumnInst_3_n15}), .c ({new_AGEMA_signal_8084, MixColumnsIns_MixOneColumnInst_3_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U46 ( .a ({new_AGEMA_signal_8085, MixColumnsIns_MixOneColumnInst_3_n14}), .b ({new_AGEMA_signal_7857, MixColumnsIns_MixOneColumnInst_3_n27}), .c ({new_AGEMA_signal_8313, MixColumnsOutput[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U45 ( .a ({new_AGEMA_signal_7489, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .b ({new_AGEMA_signal_7653, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]}), .c ({new_AGEMA_signal_7857, MixColumnsIns_MixOneColumnInst_3_n27}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U44 ( .a ({new_AGEMA_signal_7454, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .b ({new_AGEMA_signal_7858, MixColumnsIns_MixOneColumnInst_3_n62}), .c ({new_AGEMA_signal_8085, MixColumnsIns_MixOneColumnInst_3_n14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U43 ( .a ({new_AGEMA_signal_7412, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .b ({new_AGEMA_signal_7662, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]}), .c ({new_AGEMA_signal_7858, MixColumnsIns_MixOneColumnInst_3_n62}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U42 ( .a ({new_AGEMA_signal_8086, MixColumnsIns_MixOneColumnInst_3_n13}), .b ({new_AGEMA_signal_7859, MixColumnsIns_MixOneColumnInst_3_n31}), .c ({new_AGEMA_signal_8314, MixColumnsOutput[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U41 ( .a ({new_AGEMA_signal_7452, MixColumnsInput[11]}), .b ({new_AGEMA_signal_7655, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]}), .c ({new_AGEMA_signal_7859, MixColumnsIns_MixOneColumnInst_3_n31}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U40 ( .a ({new_AGEMA_signal_7410, MixColumnsInput[27]}), .b ({new_AGEMA_signal_7869, MixColumnsIns_MixOneColumnInst_3_n12}), .c ({new_AGEMA_signal_8086, MixColumnsIns_MixOneColumnInst_3_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U39 ( .a ({new_AGEMA_signal_7860, MixColumnsIns_MixOneColumnInst_3_n11}), .b ({new_AGEMA_signal_7638, MixColumnsIns_MixOneColumnInst_3_n29}), .c ({new_AGEMA_signal_8087, MixColumnsOutput[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U38 ( .a ({new_AGEMA_signal_7453, MixColumnsInput[10]}), .b ({new_AGEMA_signal_7489, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .c ({new_AGEMA_signal_7638, MixColumnsIns_MixOneColumnInst_3_n29}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U37 ( .a ({new_AGEMA_signal_7411, MixColumnsInput[26]}), .b ({new_AGEMA_signal_7647, MixColumnsIns_MixOneColumnInst_3_n10}), .c ({new_AGEMA_signal_7860, MixColumnsIns_MixOneColumnInst_3_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U36 ( .a ({new_AGEMA_signal_8088, MixColumnsIns_MixOneColumnInst_3_n9}), .b ({new_AGEMA_signal_7861, MixColumnsIns_MixOneColumnInst_3_n26}), .c ({new_AGEMA_signal_8315, MixColumnsOutput[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U35 ( .a ({new_AGEMA_signal_7656, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]}), .b ({new_AGEMA_signal_7454, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .c ({new_AGEMA_signal_7861, MixColumnsIns_MixOneColumnInst_3_n26}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U34 ( .a ({new_AGEMA_signal_7862, MixColumnsIns_MixOneColumnInst_3_n63}), .b ({new_AGEMA_signal_7412, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .c ({new_AGEMA_signal_8088, MixColumnsIns_MixOneColumnInst_3_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U33 ( .a ({new_AGEMA_signal_7659, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]}), .b ({new_AGEMA_signal_7419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .c ({new_AGEMA_signal_7862, MixColumnsIns_MixOneColumnInst_3_n63}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U32 ( .a ({new_AGEMA_signal_7863, MixColumnsIns_MixOneColumnInst_3_n8}), .b ({new_AGEMA_signal_7639, MixColumnsIns_MixOneColumnInst_3_n24}), .c ({new_AGEMA_signal_8089, MixColumnsOutput[16]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U31 ( .a ({new_AGEMA_signal_7286, MixColumnsInput[8]}), .b ({new_AGEMA_signal_7483, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .c ({new_AGEMA_signal_7639, MixColumnsIns_MixOneColumnInst_3_n24}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U30 ( .a ({new_AGEMA_signal_7220, MixColumnsInput[24]}), .b ({new_AGEMA_signal_7640, MixColumnsIns_MixOneColumnInst_3_n60}), .c ({new_AGEMA_signal_7863, MixColumnsIns_MixOneColumnInst_3_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U29 ( .a ({new_AGEMA_signal_7448, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_7231, MixColumnsInput[0]}), .c ({new_AGEMA_signal_7640, MixColumnsIns_MixOneColumnInst_3_n60}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U28 ( .a ({new_AGEMA_signal_7864, MixColumnsIns_MixOneColumnInst_3_n7}), .b ({new_AGEMA_signal_7641, MixColumnsIns_MixOneColumnInst_3_n21}), .c ({new_AGEMA_signal_8090, MixColumnsOutput[15]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U27 ( .a ({new_AGEMA_signal_7413, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_7449, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .c ({new_AGEMA_signal_7641, MixColumnsIns_MixOneColumnInst_3_n21}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U26 ( .a ({new_AGEMA_signal_7642, MixColumnsIns_MixOneColumnInst_3_n56}), .b ({new_AGEMA_signal_7483, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .c ({new_AGEMA_signal_7864, MixColumnsIns_MixOneColumnInst_3_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U25 ( .a ({new_AGEMA_signal_7414, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .b ({new_AGEMA_signal_7406, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .c ({new_AGEMA_signal_7642, MixColumnsIns_MixOneColumnInst_3_n56}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U24 ( .a ({new_AGEMA_signal_7865, MixColumnsIns_MixOneColumnInst_3_n6}), .b ({new_AGEMA_signal_7643, MixColumnsIns_MixOneColumnInst_3_n19}), .c ({new_AGEMA_signal_8091, MixColumnsOutput[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U23 ( .a ({new_AGEMA_signal_7414, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .b ({new_AGEMA_signal_7450, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .c ({new_AGEMA_signal_7643, MixColumnsIns_MixOneColumnInst_3_n19}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U22 ( .a ({new_AGEMA_signal_7644, MixColumnsIns_MixOneColumnInst_3_n53}), .b ({new_AGEMA_signal_7484, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .c ({new_AGEMA_signal_7865, MixColumnsIns_MixOneColumnInst_3_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U21 ( .a ({new_AGEMA_signal_7415, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .b ({new_AGEMA_signal_7407, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .c ({new_AGEMA_signal_7644, MixColumnsIns_MixOneColumnInst_3_n53}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U20 ( .a ({new_AGEMA_signal_7866, MixColumnsIns_MixOneColumnInst_3_n5}), .b ({new_AGEMA_signal_7645, MixColumnsIns_MixOneColumnInst_3_n17}), .c ({new_AGEMA_signal_8092, MixColumnsOutput[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U19 ( .a ({new_AGEMA_signal_7415, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .b ({new_AGEMA_signal_7451, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .c ({new_AGEMA_signal_7645, MixColumnsIns_MixOneColumnInst_3_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U18 ( .a ({new_AGEMA_signal_7646, MixColumnsIns_MixOneColumnInst_3_n50}), .b ({new_AGEMA_signal_7485, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .c ({new_AGEMA_signal_7866, MixColumnsIns_MixOneColumnInst_3_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U17 ( .a ({new_AGEMA_signal_7416, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .b ({new_AGEMA_signal_7408, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .c ({new_AGEMA_signal_7646, MixColumnsIns_MixOneColumnInst_3_n50}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U16 ( .a ({new_AGEMA_signal_8093, MixColumnsIns_MixOneColumnInst_3_n4}), .b ({new_AGEMA_signal_7867, MixColumnsIns_MixOneColumnInst_3_n15}), .c ({new_AGEMA_signal_8316, MixColumnsOutput[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U15 ( .a ({new_AGEMA_signal_7416, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .b ({new_AGEMA_signal_7657, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]}), .c ({new_AGEMA_signal_7867, MixColumnsIns_MixOneColumnInst_3_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U14 ( .a ({new_AGEMA_signal_7868, MixColumnsIns_MixOneColumnInst_3_n47}), .b ({new_AGEMA_signal_7486, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .c ({new_AGEMA_signal_8093, MixColumnsIns_MixOneColumnInst_3_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U13 ( .a ({new_AGEMA_signal_7660, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]}), .b ({new_AGEMA_signal_7409, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .c ({new_AGEMA_signal_7868, MixColumnsIns_MixOneColumnInst_3_n47}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U12 ( .a ({new_AGEMA_signal_8094, MixColumnsIns_MixOneColumnInst_3_n3}), .b ({new_AGEMA_signal_7869, MixColumnsIns_MixOneColumnInst_3_n12}), .c ({new_AGEMA_signal_8317, MixColumnsOutput[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U11 ( .a ({new_AGEMA_signal_7417, MixColumnsInput[3]}), .b ({new_AGEMA_signal_7658, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]}), .c ({new_AGEMA_signal_7869, MixColumnsIns_MixOneColumnInst_3_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U10 ( .a ({new_AGEMA_signal_7870, MixColumnsIns_MixOneColumnInst_3_n44}), .b ({new_AGEMA_signal_7487, MixColumnsInput[19]}), .c ({new_AGEMA_signal_8094, MixColumnsIns_MixOneColumnInst_3_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U9 ( .a ({new_AGEMA_signal_7661, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]}), .b ({new_AGEMA_signal_7410, MixColumnsInput[27]}), .c ({new_AGEMA_signal_7870, MixColumnsIns_MixOneColumnInst_3_n44}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U8 ( .a ({new_AGEMA_signal_7871, MixColumnsIns_MixOneColumnInst_3_n2}), .b ({new_AGEMA_signal_7647, MixColumnsIns_MixOneColumnInst_3_n10}), .c ({new_AGEMA_signal_8095, MixColumnsOutput[10]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U7 ( .a ({new_AGEMA_signal_7418, MixColumnsInput[2]}), .b ({new_AGEMA_signal_7454, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .c ({new_AGEMA_signal_7647, MixColumnsIns_MixOneColumnInst_3_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U6 ( .a ({new_AGEMA_signal_7648, MixColumnsIns_MixOneColumnInst_3_n37}), .b ({new_AGEMA_signal_7488, MixColumnsInput[18]}), .c ({new_AGEMA_signal_7871, MixColumnsIns_MixOneColumnInst_3_n2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U5 ( .a ({new_AGEMA_signal_7419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .b ({new_AGEMA_signal_7411, MixColumnsInput[26]}), .c ({new_AGEMA_signal_7648, MixColumnsIns_MixOneColumnInst_3_n37}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U4 ( .a ({new_AGEMA_signal_7872, MixColumnsIns_MixOneColumnInst_3_n1}), .b ({new_AGEMA_signal_7286, MixColumnsInput[8]}), .c ({new_AGEMA_signal_8096, MixColumnsOutput[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U3 ( .a ({new_AGEMA_signal_7650, MixColumnsIns_MixOneColumnInst_3_n59}), .b ({new_AGEMA_signal_7649, MixColumnsIns_MixOneColumnInst_3_n23}), .c ({new_AGEMA_signal_7872, MixColumnsIns_MixOneColumnInst_3_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U2 ( .a ({new_AGEMA_signal_7341, MixColumnsInput[16]}), .b ({new_AGEMA_signal_7406, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .c ({new_AGEMA_signal_7649, MixColumnsIns_MixOneColumnInst_3_n23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U1 ( .a ({new_AGEMA_signal_7413, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_7220, MixColumnsInput[24]}), .c ({new_AGEMA_signal_7650, MixColumnsIns_MixOneColumnInst_3_n59}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_7406, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_7410, MixColumnsInput[27]}), .c ({new_AGEMA_signal_7651, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_7406, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_7411, MixColumnsInput[26]}), .c ({new_AGEMA_signal_7652, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_7406, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_7220, MixColumnsInput[24]}), .c ({new_AGEMA_signal_7653, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_7483, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_7487, MixColumnsInput[19]}), .c ({new_AGEMA_signal_7654, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_7483, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_7488, MixColumnsInput[18]}), .c ({new_AGEMA_signal_7655, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_7483, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_7341, MixColumnsInput[16]}), .c ({new_AGEMA_signal_7656, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_7448, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_7452, MixColumnsInput[11]}), .c ({new_AGEMA_signal_7657, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_7448, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_7453, MixColumnsInput[10]}), .c ({new_AGEMA_signal_7658, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_7448, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_7286, MixColumnsInput[8]}), .c ({new_AGEMA_signal_7659, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_7413, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_7417, MixColumnsInput[3]}), .c ({new_AGEMA_signal_7660, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_7413, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_7418, MixColumnsInput[2]}), .c ({new_AGEMA_signal_7661, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_7413, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_7231, MixColumnsInput[0]}), .c ({new_AGEMA_signal_7662, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7968, KeyExpansionOutput[0]}), .a ({key_s1[0], key_s0[0]}), .c ({new_AGEMA_signal_8098, KeyReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8180, KeyExpansionOutput[1]}), .a ({key_s1[1], key_s0[1]}), .c ({new_AGEMA_signal_8319, KeyReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8169, KeyExpansionOutput[2]}), .a ({key_s1[2], key_s0[2]}), .c ({new_AGEMA_signal_8321, KeyReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8166, KeyExpansionOutput[3]}), .a ({key_s1[3], key_s0[3]}), .c ({new_AGEMA_signal_8323, KeyReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8165, KeyExpansionOutput[4]}), .a ({key_s1[4], key_s0[4]}), .c ({new_AGEMA_signal_8325, KeyReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8164, KeyExpansionOutput[5]}), .a ({key_s1[5], key_s0[5]}), .c ({new_AGEMA_signal_8327, KeyReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8163, KeyExpansionOutput[6]}), .a ({key_s1[6], key_s0[6]}), .c ({new_AGEMA_signal_8329, KeyReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8162, KeyExpansionOutput[7]}), .a ({key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_8331, KeyReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7937, KeyExpansionOutput[8]}), .a ({key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_8100, KeyReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8161, KeyExpansionOutput[9]}), .a ({key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_8333, KeyReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8189, KeyExpansionOutput[10]}), .a ({key_s1[10], key_s0[10]}), .c ({new_AGEMA_signal_8335, KeyReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8188, KeyExpansionOutput[11]}), .a ({key_s1[11], key_s0[11]}), .c ({new_AGEMA_signal_8337, KeyReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8187, KeyExpansionOutput[12]}), .a ({key_s1[12], key_s0[12]}), .c ({new_AGEMA_signal_8339, KeyReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8186, KeyExpansionOutput[13]}), .a ({key_s1[13], key_s0[13]}), .c ({new_AGEMA_signal_8341, KeyReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8185, KeyExpansionOutput[14]}), .a ({key_s1[14], key_s0[14]}), .c ({new_AGEMA_signal_8343, KeyReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8184, KeyExpansionOutput[15]}), .a ({key_s1[15], key_s0[15]}), .c ({new_AGEMA_signal_8345, KeyReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7961, KeyExpansionOutput[16]}), .a ({key_s1[16], key_s0[16]}), .c ({new_AGEMA_signal_8102, KeyReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8183, KeyExpansionOutput[17]}), .a ({key_s1[17], key_s0[17]}), .c ({new_AGEMA_signal_8347, KeyReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8182, KeyExpansionOutput[18]}), .a ({key_s1[18], key_s0[18]}), .c ({new_AGEMA_signal_8349, KeyReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8181, KeyExpansionOutput[19]}), .a ({key_s1[19], key_s0[19]}), .c ({new_AGEMA_signal_8351, KeyReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8179, KeyExpansionOutput[20]}), .a ({key_s1[20], key_s0[20]}), .c ({new_AGEMA_signal_8353, KeyReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8178, KeyExpansionOutput[21]}), .a ({key_s1[21], key_s0[21]}), .c ({new_AGEMA_signal_8355, KeyReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8177, KeyExpansionOutput[22]}), .a ({key_s1[22], key_s0[22]}), .c ({new_AGEMA_signal_8357, KeyReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8176, KeyExpansionOutput[23]}), .a ({key_s1[23], key_s0[23]}), .c ({new_AGEMA_signal_8359, KeyReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8175, KeyExpansionOutput[24]}), .a ({key_s1[24], key_s0[24]}), .c ({new_AGEMA_signal_8361, KeyReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8382, KeyExpansionOutput[25]}), .a ({key_s1[25], key_s0[25]}), .c ({new_AGEMA_signal_8592, KeyReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8381, KeyExpansionOutput[26]}), .a ({key_s1[26], key_s0[26]}), .c ({new_AGEMA_signal_8594, KeyReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8380, KeyExpansionOutput[27]}), .a ({key_s1[27], key_s0[27]}), .c ({new_AGEMA_signal_8596, KeyReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8379, KeyExpansionOutput[28]}), .a ({key_s1[28], key_s0[28]}), .c ({new_AGEMA_signal_8598, KeyReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8378, KeyExpansionOutput[29]}), .a ({key_s1[29], key_s0[29]}), .c ({new_AGEMA_signal_8600, KeyReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8377, KeyExpansionOutput[30]}), .a ({key_s1[30], key_s0[30]}), .c ({new_AGEMA_signal_8602, KeyReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8376, KeyExpansionOutput[31]}), .a ({key_s1[31], key_s0[31]}), .c ({new_AGEMA_signal_8604, KeyReg_Inst_ff_SDE_31_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7744, KeyExpansionOutput[32]}), .a ({key_s1[32], key_s0[32]}), .c ({new_AGEMA_signal_7874, KeyReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7957, KeyExpansionOutput[33]}), .a ({key_s1[33], key_s0[33]}), .c ({new_AGEMA_signal_8104, KeyReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7946, KeyExpansionOutput[34]}), .a ({key_s1[34], key_s0[34]}), .c ({new_AGEMA_signal_8106, KeyReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7943, KeyExpansionOutput[35]}), .a ({key_s1[35], key_s0[35]}), .c ({new_AGEMA_signal_8108, KeyReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7942, KeyExpansionOutput[36]}), .a ({key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_8110, KeyReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7941, KeyExpansionOutput[37]}), .a ({key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_8112, KeyReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7940, KeyExpansionOutput[38]}), .a ({key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_8114, KeyReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7939, KeyExpansionOutput[39]}), .a ({key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_8116, KeyReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7714, KeyExpansionOutput[40]}), .a ({key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_7876, KeyReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7938, KeyExpansionOutput[41]}), .a ({key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_8118, KeyReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7967, KeyExpansionOutput[42]}), .a ({key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_8120, KeyReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7966, KeyExpansionOutput[43]}), .a ({key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_8122, KeyReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7965, KeyExpansionOutput[44]}), .a ({key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_8124, KeyReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7964, KeyExpansionOutput[45]}), .a ({key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_8126, KeyReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7963, KeyExpansionOutput[46]}), .a ({key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_8128, KeyReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7962, KeyExpansionOutput[47]}), .a ({key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_8130, KeyReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7730, KeyExpansionOutput[48]}), .a ({key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_7878, KeyReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7960, KeyExpansionOutput[49]}), .a ({key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_8132, KeyReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7959, KeyExpansionOutput[50]}), .a ({key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_8134, KeyReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7958, KeyExpansionOutput[51]}), .a ({key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_8136, KeyReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7956, KeyExpansionOutput[52]}), .a ({key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_8138, KeyReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7955, KeyExpansionOutput[53]}), .a ({key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_8140, KeyReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7954, KeyExpansionOutput[54]}), .a ({key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_8142, KeyReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7953, KeyExpansionOutput[55]}), .a ({key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_8144, KeyReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7952, KeyExpansionOutput[56]}), .a ({key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_8146, KeyReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8174, KeyExpansionOutput[57]}), .a ({key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_8363, KeyReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8173, KeyExpansionOutput[58]}), .a ({key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_8365, KeyReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8172, KeyExpansionOutput[59]}), .a ({key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_8367, KeyReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8171, KeyExpansionOutput[60]}), .a ({key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_8369, KeyReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8170, KeyExpansionOutput[61]}), .a ({key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_8371, KeyReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8168, KeyExpansionOutput[62]}), .a ({key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_8373, KeyReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_8167, KeyExpansionOutput[63]}), .a ({key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_8375, KeyReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7527, KeyExpansionOutput[64]}), .a ({key_s1[64], key_s0[64]}), .c ({new_AGEMA_signal_7664, KeyReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7726, KeyExpansionOutput[65]}), .a ({key_s1[65], key_s0[65]}), .c ({new_AGEMA_signal_7880, KeyReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7720, KeyExpansionOutput[66]}), .a ({key_s1[66], key_s0[66]}), .c ({new_AGEMA_signal_7882, KeyReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7719, KeyExpansionOutput[67]}), .a ({key_s1[67], key_s0[67]}), .c ({new_AGEMA_signal_7884, KeyReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7718, KeyExpansionOutput[68]}), .a ({key_s1[68], key_s0[68]}), .c ({new_AGEMA_signal_7886, KeyReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7717, KeyExpansionOutput[69]}), .a ({key_s1[69], key_s0[69]}), .c ({new_AGEMA_signal_7888, KeyReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7716, KeyExpansionOutput[70]}), .a ({key_s1[70], key_s0[70]}), .c ({new_AGEMA_signal_7890, KeyReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7715, KeyExpansionOutput[71]}), .a ({key_s1[71], key_s0[71]}), .c ({new_AGEMA_signal_7892, KeyReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7503, KeyExpansionOutput[72]}), .a ({key_s1[72], key_s0[72]}), .c ({new_AGEMA_signal_7666, KeyReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7713, KeyExpansionOutput[73]}), .a ({key_s1[73], key_s0[73]}), .c ({new_AGEMA_signal_7894, KeyReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7743, KeyExpansionOutput[74]}), .a ({key_s1[74], key_s0[74]}), .c ({new_AGEMA_signal_7896, KeyReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7742, KeyExpansionOutput[75]}), .a ({key_s1[75], key_s0[75]}), .c ({new_AGEMA_signal_7898, KeyReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7734, KeyExpansionOutput[76]}), .a ({key_s1[76], key_s0[76]}), .c ({new_AGEMA_signal_7900, KeyReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7733, KeyExpansionOutput[77]}), .a ({key_s1[77], key_s0[77]}), .c ({new_AGEMA_signal_7902, KeyReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7732, KeyExpansionOutput[78]}), .a ({key_s1[78], key_s0[78]}), .c ({new_AGEMA_signal_7904, KeyReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7731, KeyExpansionOutput[79]}), .a ({key_s1[79], key_s0[79]}), .c ({new_AGEMA_signal_7906, KeyReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7507, KeyExpansionOutput[80]}), .a ({key_s1[80], key_s0[80]}), .c ({new_AGEMA_signal_7668, KeyReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7729, KeyExpansionOutput[81]}), .a ({key_s1[81], key_s0[81]}), .c ({new_AGEMA_signal_7908, KeyReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7728, KeyExpansionOutput[82]}), .a ({key_s1[82], key_s0[82]}), .c ({new_AGEMA_signal_7910, KeyReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7727, KeyExpansionOutput[83]}), .a ({key_s1[83], key_s0[83]}), .c ({new_AGEMA_signal_7912, KeyReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7725, KeyExpansionOutput[84]}), .a ({key_s1[84], key_s0[84]}), .c ({new_AGEMA_signal_7914, KeyReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7724, KeyExpansionOutput[85]}), .a ({key_s1[85], key_s0[85]}), .c ({new_AGEMA_signal_7916, KeyReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7723, KeyExpansionOutput[86]}), .a ({key_s1[86], key_s0[86]}), .c ({new_AGEMA_signal_7918, KeyReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7722, KeyExpansionOutput[87]}), .a ({key_s1[87], key_s0[87]}), .c ({new_AGEMA_signal_7920, KeyReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7721, KeyExpansionOutput[88]}), .a ({key_s1[88], key_s0[88]}), .c ({new_AGEMA_signal_7922, KeyReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7951, KeyExpansionOutput[89]}), .a ({key_s1[89], key_s0[89]}), .c ({new_AGEMA_signal_8148, KeyReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7950, KeyExpansionOutput[90]}), .a ({key_s1[90], key_s0[90]}), .c ({new_AGEMA_signal_8150, KeyReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7949, KeyExpansionOutput[91]}), .a ({key_s1[91], key_s0[91]}), .c ({new_AGEMA_signal_8152, KeyReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7948, KeyExpansionOutput[92]}), .a ({key_s1[92], key_s0[92]}), .c ({new_AGEMA_signal_8154, KeyReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7947, KeyExpansionOutput[93]}), .a ({key_s1[93], key_s0[93]}), .c ({new_AGEMA_signal_8156, KeyReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7945, KeyExpansionOutput[94]}), .a ({key_s1[94], key_s0[94]}), .c ({new_AGEMA_signal_8158, KeyReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7944, KeyExpansionOutput[95]}), .a ({key_s1[95], key_s0[95]}), .c ({new_AGEMA_signal_8160, KeyReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7355, KeyExpansionOutput[96]}), .a ({key_s1[96], key_s0[96]}), .c ({new_AGEMA_signal_7498, KeyReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7506, KeyExpansionOutput[97]}), .a ({key_s1[97], key_s0[97]}), .c ({new_AGEMA_signal_7670, KeyReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7505, KeyExpansionOutput[98]}), .a ({key_s1[98], key_s0[98]}), .c ({new_AGEMA_signal_7672, KeyReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7504, KeyExpansionOutput[99]}), .a ({key_s1[99], key_s0[99]}), .c ({new_AGEMA_signal_7674, KeyReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7526, KeyExpansionOutput[100]}), .a ({key_s1[100], key_s0[100]}), .c ({new_AGEMA_signal_7676, KeyReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7525, KeyExpansionOutput[101]}), .a ({key_s1[101], key_s0[101]}), .c ({new_AGEMA_signal_7678, KeyReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7524, KeyExpansionOutput[102]}), .a ({key_s1[102], key_s0[102]}), .c ({new_AGEMA_signal_7680, KeyReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7523, KeyExpansionOutput[103]}), .a ({key_s1[103], key_s0[103]}), .c ({new_AGEMA_signal_7682, KeyReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7354, KeyExpansionOutput[104]}), .a ({key_s1[104], key_s0[104]}), .c ({new_AGEMA_signal_7500, KeyReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7522, KeyExpansionOutput[105]}), .a ({key_s1[105], key_s0[105]}), .c ({new_AGEMA_signal_7684, KeyReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7521, KeyExpansionOutput[106]}), .a ({key_s1[106], key_s0[106]}), .c ({new_AGEMA_signal_7686, KeyReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7520, KeyExpansionOutput[107]}), .a ({key_s1[107], key_s0[107]}), .c ({new_AGEMA_signal_7688, KeyReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7519, KeyExpansionOutput[108]}), .a ({key_s1[108], key_s0[108]}), .c ({new_AGEMA_signal_7690, KeyReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7518, KeyExpansionOutput[109]}), .a ({key_s1[109], key_s0[109]}), .c ({new_AGEMA_signal_7692, KeyReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7517, KeyExpansionOutput[110]}), .a ({key_s1[110], key_s0[110]}), .c ({new_AGEMA_signal_7694, KeyReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7516, KeyExpansionOutput[111]}), .a ({key_s1[111], key_s0[111]}), .c ({new_AGEMA_signal_7696, KeyReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7353, KeyExpansionOutput[112]}), .a ({key_s1[112], key_s0[112]}), .c ({new_AGEMA_signal_7502, KeyReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7515, KeyExpansionOutput[113]}), .a ({key_s1[113], key_s0[113]}), .c ({new_AGEMA_signal_7698, KeyReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7514, KeyExpansionOutput[114]}), .a ({key_s1[114], key_s0[114]}), .c ({new_AGEMA_signal_7700, KeyReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7513, KeyExpansionOutput[115]}), .a ({key_s1[115], key_s0[115]}), .c ({new_AGEMA_signal_7702, KeyReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7512, KeyExpansionOutput[116]}), .a ({key_s1[116], key_s0[116]}), .c ({new_AGEMA_signal_7704, KeyReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7511, KeyExpansionOutput[117]}), .a ({key_s1[117], key_s0[117]}), .c ({new_AGEMA_signal_7706, KeyReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7510, KeyExpansionOutput[118]}), .a ({key_s1[118], key_s0[118]}), .c ({new_AGEMA_signal_7708, KeyReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7509, KeyExpansionOutput[119]}), .a ({key_s1[119], key_s0[119]}), .c ({new_AGEMA_signal_7710, KeyReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7508, KeyExpansionOutput[120]}), .a ({key_s1[120], key_s0[120]}), .c ({new_AGEMA_signal_7712, KeyReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7741, KeyExpansionOutput[121]}), .a ({key_s1[121], key_s0[121]}), .c ({new_AGEMA_signal_7924, KeyReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7740, KeyExpansionOutput[122]}), .a ({key_s1[122], key_s0[122]}), .c ({new_AGEMA_signal_7926, KeyReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7739, KeyExpansionOutput[123]}), .a ({key_s1[123], key_s0[123]}), .c ({new_AGEMA_signal_7928, KeyReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7738, KeyExpansionOutput[124]}), .a ({key_s1[124], key_s0[124]}), .c ({new_AGEMA_signal_7930, KeyReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7737, KeyExpansionOutput[125]}), .a ({key_s1[125], key_s0[125]}), .c ({new_AGEMA_signal_7932, KeyReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7736, KeyExpansionOutput[126]}), .a ({key_s1[126], key_s0[126]}), .c ({new_AGEMA_signal_7934, KeyReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_7735, KeyExpansionOutput[127]}), .a ({key_s1[127], key_s0[127]}), .c ({new_AGEMA_signal_7936, KeyReg_Inst_ff_SDE_127_next_state}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U128 ( .a ({new_AGEMA_signal_4931, RoundKey[9]}), .b ({new_AGEMA_signal_7938, KeyExpansionOutput[41]}), .c ({new_AGEMA_signal_8161, KeyExpansionOutput[9]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U127 ( .a ({new_AGEMA_signal_4898, RoundKey[8]}), .b ({new_AGEMA_signal_7714, KeyExpansionOutput[40]}), .c ({new_AGEMA_signal_7937, KeyExpansionOutput[8]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U126 ( .a ({new_AGEMA_signal_4865, RoundKey[7]}), .b ({new_AGEMA_signal_7939, KeyExpansionOutput[39]}), .c ({new_AGEMA_signal_8162, KeyExpansionOutput[7]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U125 ( .a ({new_AGEMA_signal_4832, RoundKey[6]}), .b ({new_AGEMA_signal_7940, KeyExpansionOutput[38]}), .c ({new_AGEMA_signal_8163, KeyExpansionOutput[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U124 ( .a ({new_AGEMA_signal_4799, RoundKey[5]}), .b ({new_AGEMA_signal_7941, KeyExpansionOutput[37]}), .c ({new_AGEMA_signal_8164, KeyExpansionOutput[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U123 ( .a ({new_AGEMA_signal_4766, RoundKey[4]}), .b ({new_AGEMA_signal_7942, KeyExpansionOutput[36]}), .c ({new_AGEMA_signal_8165, KeyExpansionOutput[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U122 ( .a ({new_AGEMA_signal_4739, RoundKey[41]}), .b ({new_AGEMA_signal_7713, KeyExpansionOutput[73]}), .c ({new_AGEMA_signal_7938, KeyExpansionOutput[41]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U121 ( .a ({new_AGEMA_signal_4844, RoundKey[73]}), .b ({new_AGEMA_signal_7522, KeyExpansionOutput[105]}), .c ({new_AGEMA_signal_7713, KeyExpansionOutput[73]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U120 ( .a ({new_AGEMA_signal_4736, RoundKey[40]}), .b ({new_AGEMA_signal_7503, KeyExpansionOutput[72]}), .c ({new_AGEMA_signal_7714, KeyExpansionOutput[40]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U119 ( .a ({new_AGEMA_signal_4841, RoundKey[72]}), .b ({new_AGEMA_signal_7354, KeyExpansionOutput[104]}), .c ({new_AGEMA_signal_7503, KeyExpansionOutput[72]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U118 ( .a ({new_AGEMA_signal_4733, RoundKey[3]}), .b ({new_AGEMA_signal_7943, KeyExpansionOutput[35]}), .c ({new_AGEMA_signal_8166, KeyExpansionOutput[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U117 ( .a ({new_AGEMA_signal_4730, RoundKey[39]}), .b ({new_AGEMA_signal_7715, KeyExpansionOutput[71]}), .c ({new_AGEMA_signal_7939, KeyExpansionOutput[39]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U116 ( .a ({new_AGEMA_signal_4838, RoundKey[71]}), .b ({new_AGEMA_signal_7523, KeyExpansionOutput[103]}), .c ({new_AGEMA_signal_7715, KeyExpansionOutput[71]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U115 ( .a ({new_AGEMA_signal_4727, RoundKey[38]}), .b ({new_AGEMA_signal_7716, KeyExpansionOutput[70]}), .c ({new_AGEMA_signal_7940, KeyExpansionOutput[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U114 ( .a ({new_AGEMA_signal_4835, RoundKey[70]}), .b ({new_AGEMA_signal_7524, KeyExpansionOutput[102]}), .c ({new_AGEMA_signal_7716, KeyExpansionOutput[70]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U113 ( .a ({new_AGEMA_signal_4724, RoundKey[37]}), .b ({new_AGEMA_signal_7717, KeyExpansionOutput[69]}), .c ({new_AGEMA_signal_7941, KeyExpansionOutput[37]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U112 ( .a ({new_AGEMA_signal_4829, RoundKey[69]}), .b ({new_AGEMA_signal_7525, KeyExpansionOutput[101]}), .c ({new_AGEMA_signal_7717, KeyExpansionOutput[69]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U111 ( .a ({new_AGEMA_signal_4721, RoundKey[36]}), .b ({new_AGEMA_signal_7718, KeyExpansionOutput[68]}), .c ({new_AGEMA_signal_7942, KeyExpansionOutput[36]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U110 ( .a ({new_AGEMA_signal_4826, RoundKey[68]}), .b ({new_AGEMA_signal_7526, KeyExpansionOutput[100]}), .c ({new_AGEMA_signal_7718, KeyExpansionOutput[68]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U109 ( .a ({new_AGEMA_signal_4718, RoundKey[35]}), .b ({new_AGEMA_signal_7719, KeyExpansionOutput[67]}), .c ({new_AGEMA_signal_7943, KeyExpansionOutput[35]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U108 ( .a ({new_AGEMA_signal_4823, RoundKey[67]}), .b ({new_AGEMA_signal_7504, KeyExpansionOutput[99]}), .c ({new_AGEMA_signal_7719, KeyExpansionOutput[67]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U107 ( .a ({new_AGEMA_signal_4928, RoundKey[99]}), .b ({new_AGEMA_signal_7382, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_7504, KeyExpansionOutput[99]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U106 ( .a ({new_AGEMA_signal_4706, RoundKey[31]}), .b ({new_AGEMA_signal_8167, KeyExpansionOutput[63]}), .c ({new_AGEMA_signal_8376, KeyExpansionOutput[31]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U105 ( .a ({new_AGEMA_signal_4811, RoundKey[63]}), .b ({new_AGEMA_signal_7944, KeyExpansionOutput[95]}), .c ({new_AGEMA_signal_8167, KeyExpansionOutput[63]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U104 ( .a ({new_AGEMA_signal_4916, RoundKey[95]}), .b ({new_AGEMA_signal_7735, KeyExpansionOutput[127]}), .c ({new_AGEMA_signal_7944, KeyExpansionOutput[95]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U103 ( .a ({new_AGEMA_signal_4703, RoundKey[30]}), .b ({new_AGEMA_signal_8168, KeyExpansionOutput[62]}), .c ({new_AGEMA_signal_8377, KeyExpansionOutput[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U102 ( .a ({new_AGEMA_signal_4808, RoundKey[62]}), .b ({new_AGEMA_signal_7945, KeyExpansionOutput[94]}), .c ({new_AGEMA_signal_8168, KeyExpansionOutput[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U101 ( .a ({new_AGEMA_signal_4913, RoundKey[94]}), .b ({new_AGEMA_signal_7736, KeyExpansionOutput[126]}), .c ({new_AGEMA_signal_7945, KeyExpansionOutput[94]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U100 ( .a ({new_AGEMA_signal_4700, RoundKey[2]}), .b ({new_AGEMA_signal_7946, KeyExpansionOutput[34]}), .c ({new_AGEMA_signal_8169, KeyExpansionOutput[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U99 ( .a ({new_AGEMA_signal_4715, RoundKey[34]}), .b ({new_AGEMA_signal_7720, KeyExpansionOutput[66]}), .c ({new_AGEMA_signal_7946, KeyExpansionOutput[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U98 ( .a ({new_AGEMA_signal_4820, RoundKey[66]}), .b ({new_AGEMA_signal_7505, KeyExpansionOutput[98]}), .c ({new_AGEMA_signal_7720, KeyExpansionOutput[66]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U97 ( .a ({new_AGEMA_signal_4925, RoundKey[98]}), .b ({new_AGEMA_signal_7383, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_7505, KeyExpansionOutput[98]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U96 ( .a ({new_AGEMA_signal_4697, RoundKey[29]}), .b ({new_AGEMA_signal_8170, KeyExpansionOutput[61]}), .c ({new_AGEMA_signal_8378, KeyExpansionOutput[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U95 ( .a ({new_AGEMA_signal_4805, RoundKey[61]}), .b ({new_AGEMA_signal_7947, KeyExpansionOutput[93]}), .c ({new_AGEMA_signal_8170, KeyExpansionOutput[61]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U94 ( .a ({new_AGEMA_signal_4910, RoundKey[93]}), .b ({new_AGEMA_signal_7737, KeyExpansionOutput[125]}), .c ({new_AGEMA_signal_7947, KeyExpansionOutput[93]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U93 ( .a ({new_AGEMA_signal_4694, RoundKey[28]}), .b ({new_AGEMA_signal_8171, KeyExpansionOutput[60]}), .c ({new_AGEMA_signal_8379, KeyExpansionOutput[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U92 ( .a ({new_AGEMA_signal_4802, RoundKey[60]}), .b ({new_AGEMA_signal_7948, KeyExpansionOutput[92]}), .c ({new_AGEMA_signal_8171, KeyExpansionOutput[60]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U91 ( .a ({new_AGEMA_signal_4907, RoundKey[92]}), .b ({new_AGEMA_signal_7738, KeyExpansionOutput[124]}), .c ({new_AGEMA_signal_7948, KeyExpansionOutput[92]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U90 ( .a ({new_AGEMA_signal_4691, RoundKey[27]}), .b ({new_AGEMA_signal_8172, KeyExpansionOutput[59]}), .c ({new_AGEMA_signal_8380, KeyExpansionOutput[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U89 ( .a ({new_AGEMA_signal_4796, RoundKey[59]}), .b ({new_AGEMA_signal_7949, KeyExpansionOutput[91]}), .c ({new_AGEMA_signal_8172, KeyExpansionOutput[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U88 ( .a ({new_AGEMA_signal_4904, RoundKey[91]}), .b ({new_AGEMA_signal_7739, KeyExpansionOutput[123]}), .c ({new_AGEMA_signal_7949, KeyExpansionOutput[91]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U87 ( .a ({new_AGEMA_signal_4688, RoundKey[26]}), .b ({new_AGEMA_signal_8173, KeyExpansionOutput[58]}), .c ({new_AGEMA_signal_8381, KeyExpansionOutput[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U86 ( .a ({new_AGEMA_signal_4793, RoundKey[58]}), .b ({new_AGEMA_signal_7950, KeyExpansionOutput[90]}), .c ({new_AGEMA_signal_8173, KeyExpansionOutput[58]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U85 ( .a ({new_AGEMA_signal_4901, RoundKey[90]}), .b ({new_AGEMA_signal_7740, KeyExpansionOutput[122]}), .c ({new_AGEMA_signal_7950, KeyExpansionOutput[90]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U84 ( .a ({new_AGEMA_signal_4685, RoundKey[25]}), .b ({new_AGEMA_signal_8174, KeyExpansionOutput[57]}), .c ({new_AGEMA_signal_8382, KeyExpansionOutput[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U83 ( .a ({new_AGEMA_signal_4790, RoundKey[57]}), .b ({new_AGEMA_signal_7951, KeyExpansionOutput[89]}), .c ({new_AGEMA_signal_8174, KeyExpansionOutput[57]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U82 ( .a ({new_AGEMA_signal_4895, RoundKey[89]}), .b ({new_AGEMA_signal_7741, KeyExpansionOutput[121]}), .c ({new_AGEMA_signal_7951, KeyExpansionOutput[89]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U81 ( .a ({new_AGEMA_signal_4682, RoundKey[24]}), .b ({new_AGEMA_signal_7952, KeyExpansionOutput[56]}), .c ({new_AGEMA_signal_8175, KeyExpansionOutput[24]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U80 ( .a ({new_AGEMA_signal_4787, RoundKey[56]}), .b ({new_AGEMA_signal_7721, KeyExpansionOutput[88]}), .c ({new_AGEMA_signal_7952, KeyExpansionOutput[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U79 ( .a ({new_AGEMA_signal_4892, RoundKey[88]}), .b ({new_AGEMA_signal_7508, KeyExpansionOutput[120]}), .c ({new_AGEMA_signal_7721, KeyExpansionOutput[88]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U78 ( .a ({new_AGEMA_signal_4679, RoundKey[23]}), .b ({new_AGEMA_signal_7953, KeyExpansionOutput[55]}), .c ({new_AGEMA_signal_8176, KeyExpansionOutput[23]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U77 ( .a ({new_AGEMA_signal_4784, RoundKey[55]}), .b ({new_AGEMA_signal_7722, KeyExpansionOutput[87]}), .c ({new_AGEMA_signal_7953, KeyExpansionOutput[55]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U76 ( .a ({new_AGEMA_signal_4889, RoundKey[87]}), .b ({new_AGEMA_signal_7509, KeyExpansionOutput[119]}), .c ({new_AGEMA_signal_7722, KeyExpansionOutput[87]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U75 ( .a ({new_AGEMA_signal_4676, RoundKey[22]}), .b ({new_AGEMA_signal_7954, KeyExpansionOutput[54]}), .c ({new_AGEMA_signal_8177, KeyExpansionOutput[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U74 ( .a ({new_AGEMA_signal_4781, RoundKey[54]}), .b ({new_AGEMA_signal_7723, KeyExpansionOutput[86]}), .c ({new_AGEMA_signal_7954, KeyExpansionOutput[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U73 ( .a ({new_AGEMA_signal_4886, RoundKey[86]}), .b ({new_AGEMA_signal_7510, KeyExpansionOutput[118]}), .c ({new_AGEMA_signal_7723, KeyExpansionOutput[86]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U72 ( .a ({new_AGEMA_signal_4673, RoundKey[21]}), .b ({new_AGEMA_signal_7955, KeyExpansionOutput[53]}), .c ({new_AGEMA_signal_8178, KeyExpansionOutput[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U71 ( .a ({new_AGEMA_signal_4778, RoundKey[53]}), .b ({new_AGEMA_signal_7724, KeyExpansionOutput[85]}), .c ({new_AGEMA_signal_7955, KeyExpansionOutput[53]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U70 ( .a ({new_AGEMA_signal_4883, RoundKey[85]}), .b ({new_AGEMA_signal_7511, KeyExpansionOutput[117]}), .c ({new_AGEMA_signal_7724, KeyExpansionOutput[85]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U69 ( .a ({new_AGEMA_signal_4670, RoundKey[20]}), .b ({new_AGEMA_signal_7956, KeyExpansionOutput[52]}), .c ({new_AGEMA_signal_8179, KeyExpansionOutput[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U68 ( .a ({new_AGEMA_signal_4775, RoundKey[52]}), .b ({new_AGEMA_signal_7725, KeyExpansionOutput[84]}), .c ({new_AGEMA_signal_7956, KeyExpansionOutput[52]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U67 ( .a ({new_AGEMA_signal_4880, RoundKey[84]}), .b ({new_AGEMA_signal_7512, KeyExpansionOutput[116]}), .c ({new_AGEMA_signal_7725, KeyExpansionOutput[84]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U66 ( .a ({new_AGEMA_signal_4667, RoundKey[1]}), .b ({new_AGEMA_signal_7957, KeyExpansionOutput[33]}), .c ({new_AGEMA_signal_8180, KeyExpansionOutput[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U65 ( .a ({new_AGEMA_signal_4712, RoundKey[33]}), .b ({new_AGEMA_signal_7726, KeyExpansionOutput[65]}), .c ({new_AGEMA_signal_7957, KeyExpansionOutput[33]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U64 ( .a ({new_AGEMA_signal_4817, RoundKey[65]}), .b ({new_AGEMA_signal_7506, KeyExpansionOutput[97]}), .c ({new_AGEMA_signal_7726, KeyExpansionOutput[65]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U63 ( .a ({new_AGEMA_signal_4922, RoundKey[97]}), .b ({new_AGEMA_signal_7384, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_7506, KeyExpansionOutput[97]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U62 ( .a ({new_AGEMA_signal_4664, RoundKey[19]}), .b ({new_AGEMA_signal_7958, KeyExpansionOutput[51]}), .c ({new_AGEMA_signal_8181, KeyExpansionOutput[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U61 ( .a ({new_AGEMA_signal_4772, RoundKey[51]}), .b ({new_AGEMA_signal_7727, KeyExpansionOutput[83]}), .c ({new_AGEMA_signal_7958, KeyExpansionOutput[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U60 ( .a ({new_AGEMA_signal_4877, RoundKey[83]}), .b ({new_AGEMA_signal_7513, KeyExpansionOutput[115]}), .c ({new_AGEMA_signal_7727, KeyExpansionOutput[83]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U59 ( .a ({new_AGEMA_signal_4661, RoundKey[18]}), .b ({new_AGEMA_signal_7959, KeyExpansionOutput[50]}), .c ({new_AGEMA_signal_8182, KeyExpansionOutput[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U58 ( .a ({new_AGEMA_signal_4769, RoundKey[50]}), .b ({new_AGEMA_signal_7728, KeyExpansionOutput[82]}), .c ({new_AGEMA_signal_7959, KeyExpansionOutput[50]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U57 ( .a ({new_AGEMA_signal_4874, RoundKey[82]}), .b ({new_AGEMA_signal_7514, KeyExpansionOutput[114]}), .c ({new_AGEMA_signal_7728, KeyExpansionOutput[82]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U56 ( .a ({new_AGEMA_signal_4658, RoundKey[17]}), .b ({new_AGEMA_signal_7960, KeyExpansionOutput[49]}), .c ({new_AGEMA_signal_8183, KeyExpansionOutput[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U55 ( .a ({new_AGEMA_signal_4763, RoundKey[49]}), .b ({new_AGEMA_signal_7729, KeyExpansionOutput[81]}), .c ({new_AGEMA_signal_7960, KeyExpansionOutput[49]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U54 ( .a ({new_AGEMA_signal_4871, RoundKey[81]}), .b ({new_AGEMA_signal_7515, KeyExpansionOutput[113]}), .c ({new_AGEMA_signal_7729, KeyExpansionOutput[81]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U53 ( .a ({new_AGEMA_signal_4655, RoundKey[16]}), .b ({new_AGEMA_signal_7730, KeyExpansionOutput[48]}), .c ({new_AGEMA_signal_7961, KeyExpansionOutput[16]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U52 ( .a ({new_AGEMA_signal_4760, RoundKey[48]}), .b ({new_AGEMA_signal_7507, KeyExpansionOutput[80]}), .c ({new_AGEMA_signal_7730, KeyExpansionOutput[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U51 ( .a ({new_AGEMA_signal_4868, RoundKey[80]}), .b ({new_AGEMA_signal_7353, KeyExpansionOutput[112]}), .c ({new_AGEMA_signal_7507, KeyExpansionOutput[80]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U50 ( .a ({new_AGEMA_signal_4652, RoundKey[15]}), .b ({new_AGEMA_signal_7962, KeyExpansionOutput[47]}), .c ({new_AGEMA_signal_8184, KeyExpansionOutput[15]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U49 ( .a ({new_AGEMA_signal_4757, RoundKey[47]}), .b ({new_AGEMA_signal_7731, KeyExpansionOutput[79]}), .c ({new_AGEMA_signal_7962, KeyExpansionOutput[47]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U48 ( .a ({new_AGEMA_signal_4862, RoundKey[79]}), .b ({new_AGEMA_signal_7516, KeyExpansionOutput[111]}), .c ({new_AGEMA_signal_7731, KeyExpansionOutput[79]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U47 ( .a ({new_AGEMA_signal_4649, RoundKey[14]}), .b ({new_AGEMA_signal_7963, KeyExpansionOutput[46]}), .c ({new_AGEMA_signal_8185, KeyExpansionOutput[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U46 ( .a ({new_AGEMA_signal_4754, RoundKey[46]}), .b ({new_AGEMA_signal_7732, KeyExpansionOutput[78]}), .c ({new_AGEMA_signal_7963, KeyExpansionOutput[46]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U45 ( .a ({new_AGEMA_signal_4859, RoundKey[78]}), .b ({new_AGEMA_signal_7517, KeyExpansionOutput[110]}), .c ({new_AGEMA_signal_7732, KeyExpansionOutput[78]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U44 ( .a ({new_AGEMA_signal_4646, RoundKey[13]}), .b ({new_AGEMA_signal_7964, KeyExpansionOutput[45]}), .c ({new_AGEMA_signal_8186, KeyExpansionOutput[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U43 ( .a ({new_AGEMA_signal_4751, RoundKey[45]}), .b ({new_AGEMA_signal_7733, KeyExpansionOutput[77]}), .c ({new_AGEMA_signal_7964, KeyExpansionOutput[45]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U42 ( .a ({new_AGEMA_signal_4856, RoundKey[77]}), .b ({new_AGEMA_signal_7518, KeyExpansionOutput[109]}), .c ({new_AGEMA_signal_7733, KeyExpansionOutput[77]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U41 ( .a ({new_AGEMA_signal_4643, RoundKey[12]}), .b ({new_AGEMA_signal_7965, KeyExpansionOutput[44]}), .c ({new_AGEMA_signal_8187, KeyExpansionOutput[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U40 ( .a ({new_AGEMA_signal_4748, RoundKey[44]}), .b ({new_AGEMA_signal_7734, KeyExpansionOutput[76]}), .c ({new_AGEMA_signal_7965, KeyExpansionOutput[44]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U39 ( .a ({new_AGEMA_signal_4853, RoundKey[76]}), .b ({new_AGEMA_signal_7519, KeyExpansionOutput[108]}), .c ({new_AGEMA_signal_7734, KeyExpansionOutput[76]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U38 ( .a ({new_AGEMA_signal_4640, RoundKey[127]}), .b ({new_AGEMA_signal_7528, KeyExpansionIns_tmp[31]}), .c ({new_AGEMA_signal_7735, KeyExpansionOutput[127]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U37 ( .a ({new_AGEMA_signal_4637, RoundKey[126]}), .b ({new_AGEMA_signal_7529, KeyExpansionIns_tmp[30]}), .c ({new_AGEMA_signal_7736, KeyExpansionOutput[126]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U36 ( .a ({new_AGEMA_signal_4634, RoundKey[125]}), .b ({new_AGEMA_signal_7530, KeyExpansionIns_tmp[29]}), .c ({new_AGEMA_signal_7737, KeyExpansionOutput[125]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U35 ( .a ({new_AGEMA_signal_4631, RoundKey[124]}), .b ({new_AGEMA_signal_7531, KeyExpansionIns_tmp[28]}), .c ({new_AGEMA_signal_7738, KeyExpansionOutput[124]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U34 ( .a ({new_AGEMA_signal_4628, RoundKey[123]}), .b ({new_AGEMA_signal_7532, KeyExpansionIns_tmp[27]}), .c ({new_AGEMA_signal_7739, KeyExpansionOutput[123]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U33 ( .a ({new_AGEMA_signal_4625, RoundKey[122]}), .b ({new_AGEMA_signal_7533, KeyExpansionIns_tmp[26]}), .c ({new_AGEMA_signal_7740, KeyExpansionOutput[122]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U32 ( .a ({new_AGEMA_signal_4622, RoundKey[121]}), .b ({new_AGEMA_signal_7534, KeyExpansionIns_tmp[25]}), .c ({new_AGEMA_signal_7741, KeyExpansionOutput[121]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U31 ( .a ({new_AGEMA_signal_4619, RoundKey[120]}), .b ({new_AGEMA_signal_7356, KeyExpansionIns_tmp[24]}), .c ({new_AGEMA_signal_7508, KeyExpansionOutput[120]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U30 ( .a ({new_AGEMA_signal_4616, RoundKey[11]}), .b ({new_AGEMA_signal_7966, KeyExpansionOutput[43]}), .c ({new_AGEMA_signal_8188, KeyExpansionOutput[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U29 ( .a ({new_AGEMA_signal_4745, RoundKey[43]}), .b ({new_AGEMA_signal_7742, KeyExpansionOutput[75]}), .c ({new_AGEMA_signal_7966, KeyExpansionOutput[43]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U28 ( .a ({new_AGEMA_signal_4850, RoundKey[75]}), .b ({new_AGEMA_signal_7520, KeyExpansionOutput[107]}), .c ({new_AGEMA_signal_7742, KeyExpansionOutput[75]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U27 ( .a ({new_AGEMA_signal_4613, RoundKey[119]}), .b ({new_AGEMA_signal_7364, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_7509, KeyExpansionOutput[119]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U26 ( .a ({new_AGEMA_signal_4610, RoundKey[118]}), .b ({new_AGEMA_signal_7365, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_7510, KeyExpansionOutput[118]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U25 ( .a ({new_AGEMA_signal_4607, RoundKey[117]}), .b ({new_AGEMA_signal_7366, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_7511, KeyExpansionOutput[117]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U24 ( .a ({new_AGEMA_signal_4604, RoundKey[116]}), .b ({new_AGEMA_signal_7367, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_7512, KeyExpansionOutput[116]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U23 ( .a ({new_AGEMA_signal_4601, RoundKey[115]}), .b ({new_AGEMA_signal_7368, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_7513, KeyExpansionOutput[115]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U22 ( .a ({new_AGEMA_signal_4598, RoundKey[114]}), .b ({new_AGEMA_signal_7369, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_7514, KeyExpansionOutput[114]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U21 ( .a ({new_AGEMA_signal_4595, RoundKey[113]}), .b ({new_AGEMA_signal_7370, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_7515, KeyExpansionOutput[113]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U20 ( .a ({new_AGEMA_signal_4592, RoundKey[112]}), .b ({new_AGEMA_signal_7154, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_7353, KeyExpansionOutput[112]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U19 ( .a ({new_AGEMA_signal_4589, RoundKey[111]}), .b ({new_AGEMA_signal_7371, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_7516, KeyExpansionOutput[111]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U18 ( .a ({new_AGEMA_signal_4586, RoundKey[110]}), .b ({new_AGEMA_signal_7372, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_7517, KeyExpansionOutput[110]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U17 ( .a ({new_AGEMA_signal_4583, RoundKey[10]}), .b ({new_AGEMA_signal_7967, KeyExpansionOutput[42]}), .c ({new_AGEMA_signal_8189, KeyExpansionOutput[10]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U16 ( .a ({new_AGEMA_signal_4742, RoundKey[42]}), .b ({new_AGEMA_signal_7743, KeyExpansionOutput[74]}), .c ({new_AGEMA_signal_7967, KeyExpansionOutput[42]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U15 ( .a ({new_AGEMA_signal_4847, RoundKey[74]}), .b ({new_AGEMA_signal_7521, KeyExpansionOutput[106]}), .c ({new_AGEMA_signal_7743, KeyExpansionOutput[74]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U14 ( .a ({new_AGEMA_signal_4580, RoundKey[109]}), .b ({new_AGEMA_signal_7373, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_7518, KeyExpansionOutput[109]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U13 ( .a ({new_AGEMA_signal_4577, RoundKey[108]}), .b ({new_AGEMA_signal_7374, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_7519, KeyExpansionOutput[108]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U12 ( .a ({new_AGEMA_signal_4574, RoundKey[107]}), .b ({new_AGEMA_signal_7375, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_7520, KeyExpansionOutput[107]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U11 ( .a ({new_AGEMA_signal_4571, RoundKey[106]}), .b ({new_AGEMA_signal_7376, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_7521, KeyExpansionOutput[106]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U10 ( .a ({new_AGEMA_signal_4568, RoundKey[105]}), .b ({new_AGEMA_signal_7377, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_7522, KeyExpansionOutput[105]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U9 ( .a ({new_AGEMA_signal_4565, RoundKey[104]}), .b ({new_AGEMA_signal_7165, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_7354, KeyExpansionOutput[104]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U8 ( .a ({new_AGEMA_signal_4562, RoundKey[103]}), .b ({new_AGEMA_signal_7378, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_7523, KeyExpansionOutput[103]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U7 ( .a ({new_AGEMA_signal_4559, RoundKey[102]}), .b ({new_AGEMA_signal_7379, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_7524, KeyExpansionOutput[102]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U6 ( .a ({new_AGEMA_signal_4556, RoundKey[101]}), .b ({new_AGEMA_signal_7380, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_7525, KeyExpansionOutput[101]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U5 ( .a ({new_AGEMA_signal_4553, RoundKey[100]}), .b ({new_AGEMA_signal_7381, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_7526, KeyExpansionOutput[100]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U4 ( .a ({new_AGEMA_signal_4550, RoundKey[0]}), .b ({new_AGEMA_signal_7744, KeyExpansionOutput[32]}), .c ({new_AGEMA_signal_7968, KeyExpansionOutput[0]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U3 ( .a ({new_AGEMA_signal_4709, RoundKey[32]}), .b ({new_AGEMA_signal_7527, KeyExpansionOutput[64]}), .c ({new_AGEMA_signal_7744, KeyExpansionOutput[32]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U2 ( .a ({new_AGEMA_signal_4814, RoundKey[64]}), .b ({new_AGEMA_signal_7355, KeyExpansionOutput[96]}), .c ({new_AGEMA_signal_7527, KeyExpansionOutput[64]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_U1 ( .a ({new_AGEMA_signal_4919, RoundKey[96]}), .b ({new_AGEMA_signal_7176, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_7355, KeyExpansionOutput[96]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U8 ( .a ({new_AGEMA_signal_7357, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_}), .b ({1'b0, n283}), .c ({new_AGEMA_signal_7528, KeyExpansionIns_tmp[31]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U7 ( .a ({new_AGEMA_signal_7358, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_}), .b ({1'b0, n285}), .c ({new_AGEMA_signal_7529, KeyExpansionIns_tmp[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U6 ( .a ({new_AGEMA_signal_7359, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_}), .b ({1'b0, Rcon[5]}), .c ({new_AGEMA_signal_7530, KeyExpansionIns_tmp[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U5 ( .a ({new_AGEMA_signal_7360, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_}), .b ({1'b0, Rcon[4]}), .c ({new_AGEMA_signal_7531, KeyExpansionIns_tmp[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U4 ( .a ({new_AGEMA_signal_7361, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_}), .b ({1'b0, Rcon[3]}), .c ({new_AGEMA_signal_7532, KeyExpansionIns_tmp[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U3 ( .a ({new_AGEMA_signal_7362, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_}), .b ({1'b0, Rcon[2]}), .c ({new_AGEMA_signal_7533, KeyExpansionIns_tmp[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U2 ( .a ({new_AGEMA_signal_7363, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_}), .b ({1'b0, Rcon[1]}), .c ({new_AGEMA_signal_7534, KeyExpansionIns_tmp[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U1 ( .a ({new_AGEMA_signal_7143, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_}), .b ({1'b0, Rcon[0]}), .c ({new_AGEMA_signal_7356, KeyExpansionIns_tmp[24]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M46_U1 ( .a ({new_AGEMA_signal_6276, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_5133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .clk (clk), .r (Fresh[608]), .c ({new_AGEMA_signal_6514, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M47_U1 ( .a ({new_AGEMA_signal_6196, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_5293, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8}), .clk (clk), .r (Fresh[609]), .c ({new_AGEMA_signal_6277, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M48_U1 ( .a ({new_AGEMA_signal_6195, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_4655, RoundKey[16]}), .clk (clk), .r (Fresh[610]), .c ({new_AGEMA_signal_6278, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M49_U1 ( .a ({new_AGEMA_signal_6275, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_5137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .clk (clk), .r (Fresh[611]), .c ({new_AGEMA_signal_6515, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M50_U1 ( .a ({new_AGEMA_signal_6194, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_5134, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}), .clk (clk), .r (Fresh[612]), .c ({new_AGEMA_signal_6279, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M51_U1 ( .a ({new_AGEMA_signal_6193, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_5296, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}), .clk (clk), .r (Fresh[613]), .c ({new_AGEMA_signal_6280, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M52_U1 ( .a ({new_AGEMA_signal_6274, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_5136, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15}), .clk (clk), .r (Fresh[614]), .c ({new_AGEMA_signal_6516, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M53_U1 ( .a ({new_AGEMA_signal_6513, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_5140, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27}), .clk (clk), .r (Fresh[615]), .c ({new_AGEMA_signal_6753, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M54_U1 ( .a ({new_AGEMA_signal_6273, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_5294, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}), .clk (clk), .r (Fresh[616]), .c ({new_AGEMA_signal_6517, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M55_U1 ( .a ({new_AGEMA_signal_6276, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_5135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13}), .clk (clk), .r (Fresh[617]), .c ({new_AGEMA_signal_6518, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M56_U1 ( .a ({new_AGEMA_signal_6196, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_5298, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23}), .clk (clk), .r (Fresh[618]), .c ({new_AGEMA_signal_6281, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M57_U1 ( .a ({new_AGEMA_signal_6195, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_5138, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}), .clk (clk), .r (Fresh[619]), .c ({new_AGEMA_signal_6282, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M58_U1 ( .a ({new_AGEMA_signal_6275, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_4935, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .clk (clk), .r (Fresh[620]), .c ({new_AGEMA_signal_6519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M59_U1 ( .a ({new_AGEMA_signal_6194, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_5139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}), .clk (clk), .r (Fresh[621]), .c ({new_AGEMA_signal_6283, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M60_U1 ( .a ({new_AGEMA_signal_6193, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_5297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}), .clk (clk), .r (Fresh[622]), .c ({new_AGEMA_signal_6284, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M61_U1 ( .a ({new_AGEMA_signal_6274, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_4933, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .clk (clk), .r (Fresh[623]), .c ({new_AGEMA_signal_6520, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M62_U1 ( .a ({new_AGEMA_signal_6513, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_4936, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}), .clk (clk), .r (Fresh[624]), .c ({new_AGEMA_signal_6754, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M63_U1 ( .a ({new_AGEMA_signal_6273, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_4934, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .clk (clk), .r (Fresh[625]), .c ({new_AGEMA_signal_6521, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L0_U1 ( .a ({new_AGEMA_signal_6520, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}), .b ({new_AGEMA_signal_6754, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62}), .c ({new_AGEMA_signal_6953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L1_U1 ( .a ({new_AGEMA_signal_6279, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_6281, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56}), .c ({new_AGEMA_signal_6522, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L2_U1 ( .a ({new_AGEMA_signal_6514, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_6278, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48}), .c ({new_AGEMA_signal_6755, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L3_U1 ( .a ({new_AGEMA_signal_6277, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47}), .b ({new_AGEMA_signal_6518, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55}), .c ({new_AGEMA_signal_6756, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L4_U1 ( .a ({new_AGEMA_signal_6517, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54}), .b ({new_AGEMA_signal_6519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58}), .c ({new_AGEMA_signal_6757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L5_U1 ( .a ({new_AGEMA_signal_6515, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49}), .b ({new_AGEMA_signal_6520, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_6758, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L6_U1 ( .a ({new_AGEMA_signal_6754, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62}), .b ({new_AGEMA_signal_6758, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5}), .c ({new_AGEMA_signal_6954, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L7_U1 ( .a ({new_AGEMA_signal_6514, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_6756, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3}), .c ({new_AGEMA_signal_6955, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L8_U1 ( .a ({new_AGEMA_signal_6280, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51}), .b ({new_AGEMA_signal_6283, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59}), .c ({new_AGEMA_signal_6523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L9_U1 ( .a ({new_AGEMA_signal_6516, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_6753, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53}), .c ({new_AGEMA_signal_6956, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L10_U1 ( .a ({new_AGEMA_signal_6753, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53}), .b ({new_AGEMA_signal_6757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_6957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L11_U1 ( .a ({new_AGEMA_signal_6284, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60}), .b ({new_AGEMA_signal_6755, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_6958, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L12_U1 ( .a ({new_AGEMA_signal_6278, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48}), .b ({new_AGEMA_signal_6280, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51}), .c ({new_AGEMA_signal_6524, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L13_U1 ( .a ({new_AGEMA_signal_6279, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_6953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_7133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L14_U1 ( .a ({new_AGEMA_signal_6516, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_6520, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_6759, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L15_U1 ( .a ({new_AGEMA_signal_6518, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55}), .b ({new_AGEMA_signal_6522, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_6760, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L16_U1 ( .a ({new_AGEMA_signal_6281, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56}), .b ({new_AGEMA_signal_6953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_7134, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L17_U1 ( .a ({new_AGEMA_signal_6282, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57}), .b ({new_AGEMA_signal_6522, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_6761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L18_U1 ( .a ({new_AGEMA_signal_6519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58}), .b ({new_AGEMA_signal_6523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8}), .c ({new_AGEMA_signal_6762, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L19_U1 ( .a ({new_AGEMA_signal_6521, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63}), .b ({new_AGEMA_signal_6757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_6959, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L20_U1 ( .a ({new_AGEMA_signal_6953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}), .b ({new_AGEMA_signal_6522, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_7135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L21_U1 ( .a ({new_AGEMA_signal_6522, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .b ({new_AGEMA_signal_6955, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7}), .c ({new_AGEMA_signal_7136, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L22_U1 ( .a ({new_AGEMA_signal_6756, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3}), .b ({new_AGEMA_signal_6524, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12}), .c ({new_AGEMA_signal_6960, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L23_U1 ( .a ({new_AGEMA_signal_6762, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18}), .b ({new_AGEMA_signal_6755, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_6961, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L24_U1 ( .a ({new_AGEMA_signal_6760, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15}), .b ({new_AGEMA_signal_6956, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_7137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L25_U1 ( .a ({new_AGEMA_signal_6954, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_6957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_7138, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L26_U1 ( .a ({new_AGEMA_signal_6955, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7}), .b ({new_AGEMA_signal_6956, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_7139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L27_U1 ( .a ({new_AGEMA_signal_6523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8}), .b ({new_AGEMA_signal_6957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_7140, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L28_U1 ( .a ({new_AGEMA_signal_6958, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_6759, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14}), .c ({new_AGEMA_signal_7141, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L29_U1 ( .a ({new_AGEMA_signal_6958, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_6761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17}), .c ({new_AGEMA_signal_7142, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S0_U1 ( .a ({new_AGEMA_signal_6954, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_7137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24}), .c ({new_AGEMA_signal_7357, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S1_U1 ( .a ({new_AGEMA_signal_7134, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16}), .b ({new_AGEMA_signal_7139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26}), .c ({new_AGEMA_signal_7358, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S2_U1 ( .a ({new_AGEMA_signal_6959, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19}), .b ({new_AGEMA_signal_7141, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28}), .c ({new_AGEMA_signal_7359, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S3_U1 ( .a ({new_AGEMA_signal_6954, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_7136, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21}), .c ({new_AGEMA_signal_7360, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S4_U1 ( .a ({new_AGEMA_signal_7135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20}), .b ({new_AGEMA_signal_6960, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22}), .c ({new_AGEMA_signal_7361, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S5_U1 ( .a ({new_AGEMA_signal_7138, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25}), .b ({new_AGEMA_signal_7142, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29}), .c ({new_AGEMA_signal_7362, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S6_U1 ( .a ({new_AGEMA_signal_7133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13}), .b ({new_AGEMA_signal_7140, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27}), .c ({new_AGEMA_signal_7363, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S7_U1 ( .a ({new_AGEMA_signal_6954, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_6961, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23}), .c ({new_AGEMA_signal_7143, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M46_U1 ( .a ({new_AGEMA_signal_6288, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_5141, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .clk (clk), .r (Fresh[626]), .c ({new_AGEMA_signal_6526, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M47_U1 ( .a ({new_AGEMA_signal_6200, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_5306, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8}), .clk (clk), .r (Fresh[627]), .c ({new_AGEMA_signal_6289, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M48_U1 ( .a ({new_AGEMA_signal_6199, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_4898, RoundKey[8]}), .clk (clk), .r (Fresh[628]), .c ({new_AGEMA_signal_6290, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M49_U1 ( .a ({new_AGEMA_signal_6287, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_5145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .clk (clk), .r (Fresh[629]), .c ({new_AGEMA_signal_6527, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M50_U1 ( .a ({new_AGEMA_signal_6198, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_5142, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}), .clk (clk), .r (Fresh[630]), .c ({new_AGEMA_signal_6291, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M51_U1 ( .a ({new_AGEMA_signal_6197, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_5309, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}), .clk (clk), .r (Fresh[631]), .c ({new_AGEMA_signal_6292, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M52_U1 ( .a ({new_AGEMA_signal_6286, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_5144, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15}), .clk (clk), .r (Fresh[632]), .c ({new_AGEMA_signal_6528, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M53_U1 ( .a ({new_AGEMA_signal_6525, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_5148, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27}), .clk (clk), .r (Fresh[633]), .c ({new_AGEMA_signal_6763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M54_U1 ( .a ({new_AGEMA_signal_6285, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_5307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}), .clk (clk), .r (Fresh[634]), .c ({new_AGEMA_signal_6529, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M55_U1 ( .a ({new_AGEMA_signal_6288, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_5143, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13}), .clk (clk), .r (Fresh[635]), .c ({new_AGEMA_signal_6530, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M56_U1 ( .a ({new_AGEMA_signal_6200, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_5311, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23}), .clk (clk), .r (Fresh[636]), .c ({new_AGEMA_signal_6293, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M57_U1 ( .a ({new_AGEMA_signal_6199, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_5146, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}), .clk (clk), .r (Fresh[637]), .c ({new_AGEMA_signal_6294, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M58_U1 ( .a ({new_AGEMA_signal_6287, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_4945, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .clk (clk), .r (Fresh[638]), .c ({new_AGEMA_signal_6531, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M59_U1 ( .a ({new_AGEMA_signal_6198, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_5147, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}), .clk (clk), .r (Fresh[639]), .c ({new_AGEMA_signal_6295, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M60_U1 ( .a ({new_AGEMA_signal_6197, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_5310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}), .clk (clk), .r (Fresh[640]), .c ({new_AGEMA_signal_6296, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M61_U1 ( .a ({new_AGEMA_signal_6286, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_4943, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .clk (clk), .r (Fresh[641]), .c ({new_AGEMA_signal_6532, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M62_U1 ( .a ({new_AGEMA_signal_6525, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_4946, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}), .clk (clk), .r (Fresh[642]), .c ({new_AGEMA_signal_6764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M63_U1 ( .a ({new_AGEMA_signal_6285, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_4944, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .clk (clk), .r (Fresh[643]), .c ({new_AGEMA_signal_6533, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L0_U1 ( .a ({new_AGEMA_signal_6532, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}), .b ({new_AGEMA_signal_6764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62}), .c ({new_AGEMA_signal_6962, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L1_U1 ( .a ({new_AGEMA_signal_6291, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_6293, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56}), .c ({new_AGEMA_signal_6534, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L2_U1 ( .a ({new_AGEMA_signal_6526, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_6290, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48}), .c ({new_AGEMA_signal_6765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L3_U1 ( .a ({new_AGEMA_signal_6289, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47}), .b ({new_AGEMA_signal_6530, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55}), .c ({new_AGEMA_signal_6766, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L4_U1 ( .a ({new_AGEMA_signal_6529, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54}), .b ({new_AGEMA_signal_6531, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58}), .c ({new_AGEMA_signal_6767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L5_U1 ( .a ({new_AGEMA_signal_6527, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49}), .b ({new_AGEMA_signal_6532, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_6768, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L6_U1 ( .a ({new_AGEMA_signal_6764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62}), .b ({new_AGEMA_signal_6768, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5}), .c ({new_AGEMA_signal_6963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L7_U1 ( .a ({new_AGEMA_signal_6526, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_6766, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3}), .c ({new_AGEMA_signal_6964, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L8_U1 ( .a ({new_AGEMA_signal_6292, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51}), .b ({new_AGEMA_signal_6295, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59}), .c ({new_AGEMA_signal_6535, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L9_U1 ( .a ({new_AGEMA_signal_6528, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_6763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53}), .c ({new_AGEMA_signal_6965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L10_U1 ( .a ({new_AGEMA_signal_6763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53}), .b ({new_AGEMA_signal_6767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_6966, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L11_U1 ( .a ({new_AGEMA_signal_6296, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60}), .b ({new_AGEMA_signal_6765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_6967, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L12_U1 ( .a ({new_AGEMA_signal_6290, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48}), .b ({new_AGEMA_signal_6292, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51}), .c ({new_AGEMA_signal_6536, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L13_U1 ( .a ({new_AGEMA_signal_6291, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_6962, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_7144, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L14_U1 ( .a ({new_AGEMA_signal_6528, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_6532, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_6769, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L15_U1 ( .a ({new_AGEMA_signal_6530, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55}), .b ({new_AGEMA_signal_6534, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_6770, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L16_U1 ( .a ({new_AGEMA_signal_6293, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56}), .b ({new_AGEMA_signal_6962, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_7145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L17_U1 ( .a ({new_AGEMA_signal_6294, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57}), .b ({new_AGEMA_signal_6534, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_6771, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L18_U1 ( .a ({new_AGEMA_signal_6531, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58}), .b ({new_AGEMA_signal_6535, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8}), .c ({new_AGEMA_signal_6772, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L19_U1 ( .a ({new_AGEMA_signal_6533, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63}), .b ({new_AGEMA_signal_6767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_6968, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L20_U1 ( .a ({new_AGEMA_signal_6962, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}), .b ({new_AGEMA_signal_6534, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_7146, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L21_U1 ( .a ({new_AGEMA_signal_6534, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .b ({new_AGEMA_signal_6964, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7}), .c ({new_AGEMA_signal_7147, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L22_U1 ( .a ({new_AGEMA_signal_6766, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3}), .b ({new_AGEMA_signal_6536, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12}), .c ({new_AGEMA_signal_6969, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L23_U1 ( .a ({new_AGEMA_signal_6772, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18}), .b ({new_AGEMA_signal_6765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_6970, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L24_U1 ( .a ({new_AGEMA_signal_6770, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15}), .b ({new_AGEMA_signal_6965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_7148, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L25_U1 ( .a ({new_AGEMA_signal_6963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_6966, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_7149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L26_U1 ( .a ({new_AGEMA_signal_6964, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7}), .b ({new_AGEMA_signal_6965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_7150, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L27_U1 ( .a ({new_AGEMA_signal_6535, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8}), .b ({new_AGEMA_signal_6966, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_7151, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L28_U1 ( .a ({new_AGEMA_signal_6967, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_6769, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14}), .c ({new_AGEMA_signal_7152, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L29_U1 ( .a ({new_AGEMA_signal_6967, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_6771, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17}), .c ({new_AGEMA_signal_7153, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S0_U1 ( .a ({new_AGEMA_signal_6963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_7148, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24}), .c ({new_AGEMA_signal_7364, KeyExpansionIns_tmp[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S1_U1 ( .a ({new_AGEMA_signal_7145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16}), .b ({new_AGEMA_signal_7150, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26}), .c ({new_AGEMA_signal_7365, KeyExpansionIns_tmp[22]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S2_U1 ( .a ({new_AGEMA_signal_6968, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19}), .b ({new_AGEMA_signal_7152, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28}), .c ({new_AGEMA_signal_7366, KeyExpansionIns_tmp[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S3_U1 ( .a ({new_AGEMA_signal_6963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_7147, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21}), .c ({new_AGEMA_signal_7367, KeyExpansionIns_tmp[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S4_U1 ( .a ({new_AGEMA_signal_7146, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20}), .b ({new_AGEMA_signal_6969, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22}), .c ({new_AGEMA_signal_7368, KeyExpansionIns_tmp[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S5_U1 ( .a ({new_AGEMA_signal_7149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25}), .b ({new_AGEMA_signal_7153, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29}), .c ({new_AGEMA_signal_7369, KeyExpansionIns_tmp[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S6_U1 ( .a ({new_AGEMA_signal_7144, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13}), .b ({new_AGEMA_signal_7151, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27}), .c ({new_AGEMA_signal_7370, KeyExpansionIns_tmp[17]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S7_U1 ( .a ({new_AGEMA_signal_6963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_6970, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23}), .c ({new_AGEMA_signal_7154, KeyExpansionIns_tmp[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M46_U1 ( .a ({new_AGEMA_signal_6300, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_5149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .clk (clk), .r (Fresh[644]), .c ({new_AGEMA_signal_6538, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M47_U1 ( .a ({new_AGEMA_signal_6204, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_5319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8}), .clk (clk), .r (Fresh[645]), .c ({new_AGEMA_signal_6301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M48_U1 ( .a ({new_AGEMA_signal_6203, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_4550, RoundKey[0]}), .clk (clk), .r (Fresh[646]), .c ({new_AGEMA_signal_6302, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M49_U1 ( .a ({new_AGEMA_signal_6299, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_5153, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .clk (clk), .r (Fresh[647]), .c ({new_AGEMA_signal_6539, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M50_U1 ( .a ({new_AGEMA_signal_6202, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_5150, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}), .clk (clk), .r (Fresh[648]), .c ({new_AGEMA_signal_6303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M51_U1 ( .a ({new_AGEMA_signal_6201, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_5322, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}), .clk (clk), .r (Fresh[649]), .c ({new_AGEMA_signal_6304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M52_U1 ( .a ({new_AGEMA_signal_6298, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_5152, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15}), .clk (clk), .r (Fresh[650]), .c ({new_AGEMA_signal_6540, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M53_U1 ( .a ({new_AGEMA_signal_6537, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_5156, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27}), .clk (clk), .r (Fresh[651]), .c ({new_AGEMA_signal_6773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M54_U1 ( .a ({new_AGEMA_signal_6297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_5320, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}), .clk (clk), .r (Fresh[652]), .c ({new_AGEMA_signal_6541, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M55_U1 ( .a ({new_AGEMA_signal_6300, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_5151, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13}), .clk (clk), .r (Fresh[653]), .c ({new_AGEMA_signal_6542, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M56_U1 ( .a ({new_AGEMA_signal_6204, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_5324, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23}), .clk (clk), .r (Fresh[654]), .c ({new_AGEMA_signal_6305, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M57_U1 ( .a ({new_AGEMA_signal_6203, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_5154, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}), .clk (clk), .r (Fresh[655]), .c ({new_AGEMA_signal_6306, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M58_U1 ( .a ({new_AGEMA_signal_6299, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_4955, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .clk (clk), .r (Fresh[656]), .c ({new_AGEMA_signal_6543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M59_U1 ( .a ({new_AGEMA_signal_6202, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_5155, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}), .clk (clk), .r (Fresh[657]), .c ({new_AGEMA_signal_6307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M60_U1 ( .a ({new_AGEMA_signal_6201, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_5323, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}), .clk (clk), .r (Fresh[658]), .c ({new_AGEMA_signal_6308, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M61_U1 ( .a ({new_AGEMA_signal_6298, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_4953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .clk (clk), .r (Fresh[659]), .c ({new_AGEMA_signal_6544, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M62_U1 ( .a ({new_AGEMA_signal_6537, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_4956, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}), .clk (clk), .r (Fresh[660]), .c ({new_AGEMA_signal_6774, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M63_U1 ( .a ({new_AGEMA_signal_6297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_4954, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .clk (clk), .r (Fresh[661]), .c ({new_AGEMA_signal_6545, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L0_U1 ( .a ({new_AGEMA_signal_6544, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}), .b ({new_AGEMA_signal_6774, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62}), .c ({new_AGEMA_signal_6971, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L1_U1 ( .a ({new_AGEMA_signal_6303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_6305, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56}), .c ({new_AGEMA_signal_6546, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L2_U1 ( .a ({new_AGEMA_signal_6538, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_6302, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48}), .c ({new_AGEMA_signal_6775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L3_U1 ( .a ({new_AGEMA_signal_6301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47}), .b ({new_AGEMA_signal_6542, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55}), .c ({new_AGEMA_signal_6776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L4_U1 ( .a ({new_AGEMA_signal_6541, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54}), .b ({new_AGEMA_signal_6543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58}), .c ({new_AGEMA_signal_6777, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L5_U1 ( .a ({new_AGEMA_signal_6539, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49}), .b ({new_AGEMA_signal_6544, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_6778, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L6_U1 ( .a ({new_AGEMA_signal_6774, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62}), .b ({new_AGEMA_signal_6778, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5}), .c ({new_AGEMA_signal_6972, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L7_U1 ( .a ({new_AGEMA_signal_6538, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_6776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3}), .c ({new_AGEMA_signal_6973, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L8_U1 ( .a ({new_AGEMA_signal_6304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51}), .b ({new_AGEMA_signal_6307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59}), .c ({new_AGEMA_signal_6547, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L9_U1 ( .a ({new_AGEMA_signal_6540, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_6773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53}), .c ({new_AGEMA_signal_6974, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L10_U1 ( .a ({new_AGEMA_signal_6773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53}), .b ({new_AGEMA_signal_6777, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_6975, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L11_U1 ( .a ({new_AGEMA_signal_6308, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60}), .b ({new_AGEMA_signal_6775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_6976, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L12_U1 ( .a ({new_AGEMA_signal_6302, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48}), .b ({new_AGEMA_signal_6304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51}), .c ({new_AGEMA_signal_6548, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L13_U1 ( .a ({new_AGEMA_signal_6303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_6971, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_7155, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L14_U1 ( .a ({new_AGEMA_signal_6540, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_6544, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_6779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L15_U1 ( .a ({new_AGEMA_signal_6542, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55}), .b ({new_AGEMA_signal_6546, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_6780, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L16_U1 ( .a ({new_AGEMA_signal_6305, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56}), .b ({new_AGEMA_signal_6971, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_7156, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L17_U1 ( .a ({new_AGEMA_signal_6306, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57}), .b ({new_AGEMA_signal_6546, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_6781, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L18_U1 ( .a ({new_AGEMA_signal_6543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58}), .b ({new_AGEMA_signal_6547, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8}), .c ({new_AGEMA_signal_6782, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L19_U1 ( .a ({new_AGEMA_signal_6545, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63}), .b ({new_AGEMA_signal_6777, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_6977, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L20_U1 ( .a ({new_AGEMA_signal_6971, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}), .b ({new_AGEMA_signal_6546, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_7157, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L21_U1 ( .a ({new_AGEMA_signal_6546, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .b ({new_AGEMA_signal_6973, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7}), .c ({new_AGEMA_signal_7158, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L22_U1 ( .a ({new_AGEMA_signal_6776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3}), .b ({new_AGEMA_signal_6548, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12}), .c ({new_AGEMA_signal_6978, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L23_U1 ( .a ({new_AGEMA_signal_6782, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18}), .b ({new_AGEMA_signal_6775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_6979, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L24_U1 ( .a ({new_AGEMA_signal_6780, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15}), .b ({new_AGEMA_signal_6974, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_7159, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L25_U1 ( .a ({new_AGEMA_signal_6972, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_6975, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_7160, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L26_U1 ( .a ({new_AGEMA_signal_6973, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7}), .b ({new_AGEMA_signal_6974, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_7161, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L27_U1 ( .a ({new_AGEMA_signal_6547, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8}), .b ({new_AGEMA_signal_6975, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_7162, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L28_U1 ( .a ({new_AGEMA_signal_6976, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_6779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14}), .c ({new_AGEMA_signal_7163, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L29_U1 ( .a ({new_AGEMA_signal_6976, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_6781, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17}), .c ({new_AGEMA_signal_7164, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S0_U1 ( .a ({new_AGEMA_signal_6972, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_7159, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24}), .c ({new_AGEMA_signal_7371, KeyExpansionIns_tmp[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S1_U1 ( .a ({new_AGEMA_signal_7156, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16}), .b ({new_AGEMA_signal_7161, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26}), .c ({new_AGEMA_signal_7372, KeyExpansionIns_tmp[14]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S2_U1 ( .a ({new_AGEMA_signal_6977, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19}), .b ({new_AGEMA_signal_7163, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28}), .c ({new_AGEMA_signal_7373, KeyExpansionIns_tmp[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S3_U1 ( .a ({new_AGEMA_signal_6972, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_7158, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21}), .c ({new_AGEMA_signal_7374, KeyExpansionIns_tmp[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S4_U1 ( .a ({new_AGEMA_signal_7157, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20}), .b ({new_AGEMA_signal_6978, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22}), .c ({new_AGEMA_signal_7375, KeyExpansionIns_tmp[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S5_U1 ( .a ({new_AGEMA_signal_7160, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25}), .b ({new_AGEMA_signal_7164, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29}), .c ({new_AGEMA_signal_7376, KeyExpansionIns_tmp[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S6_U1 ( .a ({new_AGEMA_signal_7155, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13}), .b ({new_AGEMA_signal_7162, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27}), .c ({new_AGEMA_signal_7377, KeyExpansionIns_tmp[9]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S7_U1 ( .a ({new_AGEMA_signal_6972, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_6979, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23}), .c ({new_AGEMA_signal_7165, KeyExpansionIns_tmp[8]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M46_U1 ( .a ({new_AGEMA_signal_6312, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_5157, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .clk (clk), .r (Fresh[662]), .c ({new_AGEMA_signal_6550, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M47_U1 ( .a ({new_AGEMA_signal_6208, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_5332, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8}), .clk (clk), .r (Fresh[663]), .c ({new_AGEMA_signal_6313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M48_U1 ( .a ({new_AGEMA_signal_6207, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_4682, RoundKey[24]}), .clk (clk), .r (Fresh[664]), .c ({new_AGEMA_signal_6314, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M49_U1 ( .a ({new_AGEMA_signal_6311, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_5161, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .clk (clk), .r (Fresh[665]), .c ({new_AGEMA_signal_6551, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M50_U1 ( .a ({new_AGEMA_signal_6206, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_5158, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}), .clk (clk), .r (Fresh[666]), .c ({new_AGEMA_signal_6315, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M51_U1 ( .a ({new_AGEMA_signal_6205, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_5335, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}), .clk (clk), .r (Fresh[667]), .c ({new_AGEMA_signal_6316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M52_U1 ( .a ({new_AGEMA_signal_6310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_5160, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15}), .clk (clk), .r (Fresh[668]), .c ({new_AGEMA_signal_6552, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M53_U1 ( .a ({new_AGEMA_signal_6549, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_5164, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27}), .clk (clk), .r (Fresh[669]), .c ({new_AGEMA_signal_6783, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M54_U1 ( .a ({new_AGEMA_signal_6309, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_5333, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}), .clk (clk), .r (Fresh[670]), .c ({new_AGEMA_signal_6553, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M55_U1 ( .a ({new_AGEMA_signal_6312, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_5159, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13}), .clk (clk), .r (Fresh[671]), .c ({new_AGEMA_signal_6554, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M56_U1 ( .a ({new_AGEMA_signal_6208, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_5337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23}), .clk (clk), .r (Fresh[672]), .c ({new_AGEMA_signal_6317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M57_U1 ( .a ({new_AGEMA_signal_6207, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_5162, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}), .clk (clk), .r (Fresh[673]), .c ({new_AGEMA_signal_6318, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M58_U1 ( .a ({new_AGEMA_signal_6311, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_4965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .clk (clk), .r (Fresh[674]), .c ({new_AGEMA_signal_6555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M59_U1 ( .a ({new_AGEMA_signal_6206, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_5163, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}), .clk (clk), .r (Fresh[675]), .c ({new_AGEMA_signal_6319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M60_U1 ( .a ({new_AGEMA_signal_6205, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_5336, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}), .clk (clk), .r (Fresh[676]), .c ({new_AGEMA_signal_6320, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M61_U1 ( .a ({new_AGEMA_signal_6310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_4963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .clk (clk), .r (Fresh[677]), .c ({new_AGEMA_signal_6556, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M62_U1 ( .a ({new_AGEMA_signal_6549, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_4966, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}), .clk (clk), .r (Fresh[678]), .c ({new_AGEMA_signal_6784, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M63_U1 ( .a ({new_AGEMA_signal_6309, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_4964, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .clk (clk), .r (Fresh[679]), .c ({new_AGEMA_signal_6557, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L0_U1 ( .a ({new_AGEMA_signal_6556, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}), .b ({new_AGEMA_signal_6784, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62}), .c ({new_AGEMA_signal_6980, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L1_U1 ( .a ({new_AGEMA_signal_6315, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_6317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56}), .c ({new_AGEMA_signal_6558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L2_U1 ( .a ({new_AGEMA_signal_6550, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_6314, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48}), .c ({new_AGEMA_signal_6785, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L3_U1 ( .a ({new_AGEMA_signal_6313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47}), .b ({new_AGEMA_signal_6554, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55}), .c ({new_AGEMA_signal_6786, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L4_U1 ( .a ({new_AGEMA_signal_6553, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54}), .b ({new_AGEMA_signal_6555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58}), .c ({new_AGEMA_signal_6787, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L5_U1 ( .a ({new_AGEMA_signal_6551, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49}), .b ({new_AGEMA_signal_6556, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_6788, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L6_U1 ( .a ({new_AGEMA_signal_6784, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62}), .b ({new_AGEMA_signal_6788, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5}), .c ({new_AGEMA_signal_6981, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L7_U1 ( .a ({new_AGEMA_signal_6550, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_6786, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3}), .c ({new_AGEMA_signal_6982, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L8_U1 ( .a ({new_AGEMA_signal_6316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51}), .b ({new_AGEMA_signal_6319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59}), .c ({new_AGEMA_signal_6559, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L9_U1 ( .a ({new_AGEMA_signal_6552, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_6783, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53}), .c ({new_AGEMA_signal_6983, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L10_U1 ( .a ({new_AGEMA_signal_6783, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53}), .b ({new_AGEMA_signal_6787, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_6984, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L11_U1 ( .a ({new_AGEMA_signal_6320, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60}), .b ({new_AGEMA_signal_6785, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_6985, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L12_U1 ( .a ({new_AGEMA_signal_6314, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48}), .b ({new_AGEMA_signal_6316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51}), .c ({new_AGEMA_signal_6560, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L13_U1 ( .a ({new_AGEMA_signal_6315, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_6980, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_7166, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L14_U1 ( .a ({new_AGEMA_signal_6552, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_6556, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_6789, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L15_U1 ( .a ({new_AGEMA_signal_6554, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55}), .b ({new_AGEMA_signal_6558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_6790, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L16_U1 ( .a ({new_AGEMA_signal_6317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56}), .b ({new_AGEMA_signal_6980, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_7167, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L17_U1 ( .a ({new_AGEMA_signal_6318, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57}), .b ({new_AGEMA_signal_6558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_6791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L18_U1 ( .a ({new_AGEMA_signal_6555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58}), .b ({new_AGEMA_signal_6559, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8}), .c ({new_AGEMA_signal_6792, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L19_U1 ( .a ({new_AGEMA_signal_6557, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63}), .b ({new_AGEMA_signal_6787, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_6986, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L20_U1 ( .a ({new_AGEMA_signal_6980, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}), .b ({new_AGEMA_signal_6558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_7168, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L21_U1 ( .a ({new_AGEMA_signal_6558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .b ({new_AGEMA_signal_6982, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7}), .c ({new_AGEMA_signal_7169, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L22_U1 ( .a ({new_AGEMA_signal_6786, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3}), .b ({new_AGEMA_signal_6560, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12}), .c ({new_AGEMA_signal_6987, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L23_U1 ( .a ({new_AGEMA_signal_6792, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18}), .b ({new_AGEMA_signal_6785, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_6988, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L24_U1 ( .a ({new_AGEMA_signal_6790, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15}), .b ({new_AGEMA_signal_6983, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_7170, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L25_U1 ( .a ({new_AGEMA_signal_6981, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_6984, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_7171, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L26_U1 ( .a ({new_AGEMA_signal_6982, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7}), .b ({new_AGEMA_signal_6983, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_7172, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L27_U1 ( .a ({new_AGEMA_signal_6559, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8}), .b ({new_AGEMA_signal_6984, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_7173, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L28_U1 ( .a ({new_AGEMA_signal_6985, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_6789, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14}), .c ({new_AGEMA_signal_7174, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L29_U1 ( .a ({new_AGEMA_signal_6985, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_6791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17}), .c ({new_AGEMA_signal_7175, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S0_U1 ( .a ({new_AGEMA_signal_6981, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_7170, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24}), .c ({new_AGEMA_signal_7378, KeyExpansionIns_tmp[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S1_U1 ( .a ({new_AGEMA_signal_7167, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16}), .b ({new_AGEMA_signal_7172, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26}), .c ({new_AGEMA_signal_7379, KeyExpansionIns_tmp[6]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S2_U1 ( .a ({new_AGEMA_signal_6986, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19}), .b ({new_AGEMA_signal_7174, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28}), .c ({new_AGEMA_signal_7380, KeyExpansionIns_tmp[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S3_U1 ( .a ({new_AGEMA_signal_6981, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_7169, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21}), .c ({new_AGEMA_signal_7381, KeyExpansionIns_tmp[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S4_U1 ( .a ({new_AGEMA_signal_7168, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20}), .b ({new_AGEMA_signal_6987, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22}), .c ({new_AGEMA_signal_7382, KeyExpansionIns_tmp[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S5_U1 ( .a ({new_AGEMA_signal_7171, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25}), .b ({new_AGEMA_signal_7175, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29}), .c ({new_AGEMA_signal_7383, KeyExpansionIns_tmp[2]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S6_U1 ( .a ({new_AGEMA_signal_7166, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13}), .b ({new_AGEMA_signal_7173, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27}), .c ({new_AGEMA_signal_7384, KeyExpansionIns_tmp[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S7_U1 ( .a ({new_AGEMA_signal_6981, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_6988, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23}), .c ({new_AGEMA_signal_7176, KeyExpansionIns_tmp[0]}) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8432, RoundReg_Inst_ff_SDE_0_next_state}), .Q ({new_AGEMA_signal_4549, RoundInput[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8606, RoundReg_Inst_ff_SDE_1_next_state}), .Q ({new_AGEMA_signal_4666, RoundInput[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8434, RoundReg_Inst_ff_SDE_2_next_state}), .Q ({new_AGEMA_signal_4699, RoundInput[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8608, RoundReg_Inst_ff_SDE_3_next_state}), .Q ({new_AGEMA_signal_4732, RoundInput[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8610, RoundReg_Inst_ff_SDE_4_next_state}), .Q ({new_AGEMA_signal_4765, RoundInput[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8436, RoundReg_Inst_ff_SDE_5_next_state}), .Q ({new_AGEMA_signal_4798, RoundInput[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8438, RoundReg_Inst_ff_SDE_6_next_state}), .Q ({new_AGEMA_signal_4831, RoundInput[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8440, RoundReg_Inst_ff_SDE_7_next_state}), .Q ({new_AGEMA_signal_4864, RoundInput[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8442, RoundReg_Inst_ff_SDE_8_next_state}), .Q ({new_AGEMA_signal_4897, RoundInput[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8612, RoundReg_Inst_ff_SDE_9_next_state}), .Q ({new_AGEMA_signal_4930, RoundInput[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8444, RoundReg_Inst_ff_SDE_10_next_state}), .Q ({new_AGEMA_signal_4582, RoundInput[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8614, RoundReg_Inst_ff_SDE_11_next_state}), .Q ({new_AGEMA_signal_4615, RoundInput[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8616, RoundReg_Inst_ff_SDE_12_next_state}), .Q ({new_AGEMA_signal_4642, RoundInput[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8446, RoundReg_Inst_ff_SDE_13_next_state}), .Q ({new_AGEMA_signal_4645, RoundInput[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8448, RoundReg_Inst_ff_SDE_14_next_state}), .Q ({new_AGEMA_signal_4648, RoundInput[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8450, RoundReg_Inst_ff_SDE_15_next_state}), .Q ({new_AGEMA_signal_4651, RoundInput[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8452, RoundReg_Inst_ff_SDE_16_next_state}), .Q ({new_AGEMA_signal_4654, RoundInput[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8618, RoundReg_Inst_ff_SDE_17_next_state}), .Q ({new_AGEMA_signal_4657, RoundInput[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8454, RoundReg_Inst_ff_SDE_18_next_state}), .Q ({new_AGEMA_signal_4660, RoundInput[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8620, RoundReg_Inst_ff_SDE_19_next_state}), .Q ({new_AGEMA_signal_4663, RoundInput[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8622, RoundReg_Inst_ff_SDE_20_next_state}), .Q ({new_AGEMA_signal_4669, RoundInput[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8456, RoundReg_Inst_ff_SDE_21_next_state}), .Q ({new_AGEMA_signal_4672, RoundInput[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8458, RoundReg_Inst_ff_SDE_22_next_state}), .Q ({new_AGEMA_signal_4675, RoundInput[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8460, RoundReg_Inst_ff_SDE_23_next_state}), .Q ({new_AGEMA_signal_4678, RoundInput[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8462, RoundReg_Inst_ff_SDE_24_next_state}), .Q ({new_AGEMA_signal_4681, RoundInput[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8624, RoundReg_Inst_ff_SDE_25_next_state}), .Q ({new_AGEMA_signal_4684, RoundInput[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8464, RoundReg_Inst_ff_SDE_26_next_state}), .Q ({new_AGEMA_signal_4687, RoundInput[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8626, RoundReg_Inst_ff_SDE_27_next_state}), .Q ({new_AGEMA_signal_4690, RoundInput[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8628, RoundReg_Inst_ff_SDE_28_next_state}), .Q ({new_AGEMA_signal_4693, RoundInput[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8466, RoundReg_Inst_ff_SDE_29_next_state}), .Q ({new_AGEMA_signal_4696, RoundInput[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8468, RoundReg_Inst_ff_SDE_30_next_state}), .Q ({new_AGEMA_signal_4702, RoundInput[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8470, RoundReg_Inst_ff_SDE_31_next_state}), .Q ({new_AGEMA_signal_4705, RoundInput[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8472, RoundReg_Inst_ff_SDE_32_next_state}), .Q ({new_AGEMA_signal_4708, RoundInput[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8630, RoundReg_Inst_ff_SDE_33_next_state}), .Q ({new_AGEMA_signal_4711, RoundInput[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8474, RoundReg_Inst_ff_SDE_34_next_state}), .Q ({new_AGEMA_signal_4714, RoundInput[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8632, RoundReg_Inst_ff_SDE_35_next_state}), .Q ({new_AGEMA_signal_4717, RoundInput[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8634, RoundReg_Inst_ff_SDE_36_next_state}), .Q ({new_AGEMA_signal_4720, RoundInput[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8476, RoundReg_Inst_ff_SDE_37_next_state}), .Q ({new_AGEMA_signal_4723, RoundInput[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8478, RoundReg_Inst_ff_SDE_38_next_state}), .Q ({new_AGEMA_signal_4726, RoundInput[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8480, RoundReg_Inst_ff_SDE_39_next_state}), .Q ({new_AGEMA_signal_4729, RoundInput[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8482, RoundReg_Inst_ff_SDE_40_next_state}), .Q ({new_AGEMA_signal_4735, RoundInput[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8636, RoundReg_Inst_ff_SDE_41_next_state}), .Q ({new_AGEMA_signal_4738, RoundInput[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8484, RoundReg_Inst_ff_SDE_42_next_state}), .Q ({new_AGEMA_signal_4741, RoundInput[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8638, RoundReg_Inst_ff_SDE_43_next_state}), .Q ({new_AGEMA_signal_4744, RoundInput[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8640, RoundReg_Inst_ff_SDE_44_next_state}), .Q ({new_AGEMA_signal_4747, RoundInput[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8486, RoundReg_Inst_ff_SDE_45_next_state}), .Q ({new_AGEMA_signal_4750, RoundInput[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8488, RoundReg_Inst_ff_SDE_46_next_state}), .Q ({new_AGEMA_signal_4753, RoundInput[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8490, RoundReg_Inst_ff_SDE_47_next_state}), .Q ({new_AGEMA_signal_4756, RoundInput[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8492, RoundReg_Inst_ff_SDE_48_next_state}), .Q ({new_AGEMA_signal_4759, RoundInput[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8642, RoundReg_Inst_ff_SDE_49_next_state}), .Q ({new_AGEMA_signal_4762, RoundInput[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8494, RoundReg_Inst_ff_SDE_50_next_state}), .Q ({new_AGEMA_signal_4768, RoundInput[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8644, RoundReg_Inst_ff_SDE_51_next_state}), .Q ({new_AGEMA_signal_4771, RoundInput[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8646, RoundReg_Inst_ff_SDE_52_next_state}), .Q ({new_AGEMA_signal_4774, RoundInput[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8496, RoundReg_Inst_ff_SDE_53_next_state}), .Q ({new_AGEMA_signal_4777, RoundInput[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8498, RoundReg_Inst_ff_SDE_54_next_state}), .Q ({new_AGEMA_signal_4780, RoundInput[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8500, RoundReg_Inst_ff_SDE_55_next_state}), .Q ({new_AGEMA_signal_4783, RoundInput[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8502, RoundReg_Inst_ff_SDE_56_next_state}), .Q ({new_AGEMA_signal_4786, RoundInput[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8648, RoundReg_Inst_ff_SDE_57_next_state}), .Q ({new_AGEMA_signal_4789, RoundInput[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8504, RoundReg_Inst_ff_SDE_58_next_state}), .Q ({new_AGEMA_signal_4792, RoundInput[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8650, RoundReg_Inst_ff_SDE_59_next_state}), .Q ({new_AGEMA_signal_4795, RoundInput[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8652, RoundReg_Inst_ff_SDE_60_next_state}), .Q ({new_AGEMA_signal_4801, RoundInput[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8506, RoundReg_Inst_ff_SDE_61_next_state}), .Q ({new_AGEMA_signal_4804, RoundInput[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8508, RoundReg_Inst_ff_SDE_62_next_state}), .Q ({new_AGEMA_signal_4807, RoundInput[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8510, RoundReg_Inst_ff_SDE_63_next_state}), .Q ({new_AGEMA_signal_4810, RoundInput[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8512, RoundReg_Inst_ff_SDE_64_next_state}), .Q ({new_AGEMA_signal_4813, RoundInput[64]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8654, RoundReg_Inst_ff_SDE_65_next_state}), .Q ({new_AGEMA_signal_4816, RoundInput[65]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8514, RoundReg_Inst_ff_SDE_66_next_state}), .Q ({new_AGEMA_signal_4819, RoundInput[66]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8656, RoundReg_Inst_ff_SDE_67_next_state}), .Q ({new_AGEMA_signal_4822, RoundInput[67]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8658, RoundReg_Inst_ff_SDE_68_next_state}), .Q ({new_AGEMA_signal_4825, RoundInput[68]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8516, RoundReg_Inst_ff_SDE_69_next_state}), .Q ({new_AGEMA_signal_4828, RoundInput[69]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8518, RoundReg_Inst_ff_SDE_70_next_state}), .Q ({new_AGEMA_signal_4834, RoundInput[70]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8520, RoundReg_Inst_ff_SDE_71_next_state}), .Q ({new_AGEMA_signal_4837, RoundInput[71]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8522, RoundReg_Inst_ff_SDE_72_next_state}), .Q ({new_AGEMA_signal_4840, RoundInput[72]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8660, RoundReg_Inst_ff_SDE_73_next_state}), .Q ({new_AGEMA_signal_4843, RoundInput[73]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8524, RoundReg_Inst_ff_SDE_74_next_state}), .Q ({new_AGEMA_signal_4846, RoundInput[74]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8662, RoundReg_Inst_ff_SDE_75_next_state}), .Q ({new_AGEMA_signal_4849, RoundInput[75]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8664, RoundReg_Inst_ff_SDE_76_next_state}), .Q ({new_AGEMA_signal_4852, RoundInput[76]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8526, RoundReg_Inst_ff_SDE_77_next_state}), .Q ({new_AGEMA_signal_4855, RoundInput[77]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8528, RoundReg_Inst_ff_SDE_78_next_state}), .Q ({new_AGEMA_signal_4858, RoundInput[78]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8530, RoundReg_Inst_ff_SDE_79_next_state}), .Q ({new_AGEMA_signal_4861, RoundInput[79]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8532, RoundReg_Inst_ff_SDE_80_next_state}), .Q ({new_AGEMA_signal_4867, RoundInput[80]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8666, RoundReg_Inst_ff_SDE_81_next_state}), .Q ({new_AGEMA_signal_4870, RoundInput[81]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8534, RoundReg_Inst_ff_SDE_82_next_state}), .Q ({new_AGEMA_signal_4873, RoundInput[82]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8668, RoundReg_Inst_ff_SDE_83_next_state}), .Q ({new_AGEMA_signal_4876, RoundInput[83]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8670, RoundReg_Inst_ff_SDE_84_next_state}), .Q ({new_AGEMA_signal_4879, RoundInput[84]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8536, RoundReg_Inst_ff_SDE_85_next_state}), .Q ({new_AGEMA_signal_4882, RoundInput[85]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8538, RoundReg_Inst_ff_SDE_86_next_state}), .Q ({new_AGEMA_signal_4885, RoundInput[86]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8540, RoundReg_Inst_ff_SDE_87_next_state}), .Q ({new_AGEMA_signal_4888, RoundInput[87]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8542, RoundReg_Inst_ff_SDE_88_next_state}), .Q ({new_AGEMA_signal_4891, RoundInput[88]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8672, RoundReg_Inst_ff_SDE_89_next_state}), .Q ({new_AGEMA_signal_4894, RoundInput[89]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8544, RoundReg_Inst_ff_SDE_90_next_state}), .Q ({new_AGEMA_signal_4900, RoundInput[90]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8674, RoundReg_Inst_ff_SDE_91_next_state}), .Q ({new_AGEMA_signal_4903, RoundInput[91]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8676, RoundReg_Inst_ff_SDE_92_next_state}), .Q ({new_AGEMA_signal_4906, RoundInput[92]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8546, RoundReg_Inst_ff_SDE_93_next_state}), .Q ({new_AGEMA_signal_4909, RoundInput[93]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8548, RoundReg_Inst_ff_SDE_94_next_state}), .Q ({new_AGEMA_signal_4912, RoundInput[94]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8550, RoundReg_Inst_ff_SDE_95_next_state}), .Q ({new_AGEMA_signal_4915, RoundInput[95]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8552, RoundReg_Inst_ff_SDE_96_next_state}), .Q ({new_AGEMA_signal_4918, RoundInput[96]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8678, RoundReg_Inst_ff_SDE_97_next_state}), .Q ({new_AGEMA_signal_4921, RoundInput[97]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8554, RoundReg_Inst_ff_SDE_98_next_state}), .Q ({new_AGEMA_signal_4924, RoundInput[98]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8680, RoundReg_Inst_ff_SDE_99_next_state}), .Q ({new_AGEMA_signal_4927, RoundInput[99]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8682, RoundReg_Inst_ff_SDE_100_next_state}), .Q ({new_AGEMA_signal_4552, RoundInput[100]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8556, RoundReg_Inst_ff_SDE_101_next_state}), .Q ({new_AGEMA_signal_4555, RoundInput[101]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8558, RoundReg_Inst_ff_SDE_102_next_state}), .Q ({new_AGEMA_signal_4558, RoundInput[102]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8560, RoundReg_Inst_ff_SDE_103_next_state}), .Q ({new_AGEMA_signal_4561, RoundInput[103]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8562, RoundReg_Inst_ff_SDE_104_next_state}), .Q ({new_AGEMA_signal_4564, RoundInput[104]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8684, RoundReg_Inst_ff_SDE_105_next_state}), .Q ({new_AGEMA_signal_4567, RoundInput[105]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8564, RoundReg_Inst_ff_SDE_106_next_state}), .Q ({new_AGEMA_signal_4570, RoundInput[106]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8686, RoundReg_Inst_ff_SDE_107_next_state}), .Q ({new_AGEMA_signal_4573, RoundInput[107]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8688, RoundReg_Inst_ff_SDE_108_next_state}), .Q ({new_AGEMA_signal_4576, RoundInput[108]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8566, RoundReg_Inst_ff_SDE_109_next_state}), .Q ({new_AGEMA_signal_4579, RoundInput[109]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8568, RoundReg_Inst_ff_SDE_110_next_state}), .Q ({new_AGEMA_signal_4585, RoundInput[110]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8570, RoundReg_Inst_ff_SDE_111_next_state}), .Q ({new_AGEMA_signal_4588, RoundInput[111]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8572, RoundReg_Inst_ff_SDE_112_next_state}), .Q ({new_AGEMA_signal_4591, RoundInput[112]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8690, RoundReg_Inst_ff_SDE_113_next_state}), .Q ({new_AGEMA_signal_4594, RoundInput[113]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8574, RoundReg_Inst_ff_SDE_114_next_state}), .Q ({new_AGEMA_signal_4597, RoundInput[114]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8692, RoundReg_Inst_ff_SDE_115_next_state}), .Q ({new_AGEMA_signal_4600, RoundInput[115]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8694, RoundReg_Inst_ff_SDE_116_next_state}), .Q ({new_AGEMA_signal_4603, RoundInput[116]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8576, RoundReg_Inst_ff_SDE_117_next_state}), .Q ({new_AGEMA_signal_4606, RoundInput[117]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8578, RoundReg_Inst_ff_SDE_118_next_state}), .Q ({new_AGEMA_signal_4609, RoundInput[118]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8580, RoundReg_Inst_ff_SDE_119_next_state}), .Q ({new_AGEMA_signal_4612, RoundInput[119]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8582, RoundReg_Inst_ff_SDE_120_next_state}), .Q ({new_AGEMA_signal_4618, RoundInput[120]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8696, RoundReg_Inst_ff_SDE_121_next_state}), .Q ({new_AGEMA_signal_4621, RoundInput[121]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8584, RoundReg_Inst_ff_SDE_122_next_state}), .Q ({new_AGEMA_signal_4624, RoundInput[122]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8698, RoundReg_Inst_ff_SDE_123_next_state}), .Q ({new_AGEMA_signal_4627, RoundInput[123]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8700, RoundReg_Inst_ff_SDE_124_next_state}), .Q ({new_AGEMA_signal_4630, RoundInput[124]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8586, RoundReg_Inst_ff_SDE_125_next_state}), .Q ({new_AGEMA_signal_4633, RoundInput[125]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8588, RoundReg_Inst_ff_SDE_126_next_state}), .Q ({new_AGEMA_signal_4636, RoundInput[126]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) RoundReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8590, RoundReg_Inst_ff_SDE_127_next_state}), .Q ({new_AGEMA_signal_4639, RoundInput[127]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8098, KeyReg_Inst_ff_SDE_0_next_state}), .Q ({new_AGEMA_signal_4550, RoundKey[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8319, KeyReg_Inst_ff_SDE_1_next_state}), .Q ({new_AGEMA_signal_4667, RoundKey[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8321, KeyReg_Inst_ff_SDE_2_next_state}), .Q ({new_AGEMA_signal_4700, RoundKey[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8323, KeyReg_Inst_ff_SDE_3_next_state}), .Q ({new_AGEMA_signal_4733, RoundKey[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8325, KeyReg_Inst_ff_SDE_4_next_state}), .Q ({new_AGEMA_signal_4766, RoundKey[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8327, KeyReg_Inst_ff_SDE_5_next_state}), .Q ({new_AGEMA_signal_4799, RoundKey[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8329, KeyReg_Inst_ff_SDE_6_next_state}), .Q ({new_AGEMA_signal_4832, RoundKey[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8331, KeyReg_Inst_ff_SDE_7_next_state}), .Q ({new_AGEMA_signal_4865, RoundKey[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8100, KeyReg_Inst_ff_SDE_8_next_state}), .Q ({new_AGEMA_signal_4898, RoundKey[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8333, KeyReg_Inst_ff_SDE_9_next_state}), .Q ({new_AGEMA_signal_4931, RoundKey[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8335, KeyReg_Inst_ff_SDE_10_next_state}), .Q ({new_AGEMA_signal_4583, RoundKey[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8337, KeyReg_Inst_ff_SDE_11_next_state}), .Q ({new_AGEMA_signal_4616, RoundKey[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8339, KeyReg_Inst_ff_SDE_12_next_state}), .Q ({new_AGEMA_signal_4643, RoundKey[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8341, KeyReg_Inst_ff_SDE_13_next_state}), .Q ({new_AGEMA_signal_4646, RoundKey[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8343, KeyReg_Inst_ff_SDE_14_next_state}), .Q ({new_AGEMA_signal_4649, RoundKey[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8345, KeyReg_Inst_ff_SDE_15_next_state}), .Q ({new_AGEMA_signal_4652, RoundKey[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8102, KeyReg_Inst_ff_SDE_16_next_state}), .Q ({new_AGEMA_signal_4655, RoundKey[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8347, KeyReg_Inst_ff_SDE_17_next_state}), .Q ({new_AGEMA_signal_4658, RoundKey[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8349, KeyReg_Inst_ff_SDE_18_next_state}), .Q ({new_AGEMA_signal_4661, RoundKey[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8351, KeyReg_Inst_ff_SDE_19_next_state}), .Q ({new_AGEMA_signal_4664, RoundKey[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8353, KeyReg_Inst_ff_SDE_20_next_state}), .Q ({new_AGEMA_signal_4670, RoundKey[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8355, KeyReg_Inst_ff_SDE_21_next_state}), .Q ({new_AGEMA_signal_4673, RoundKey[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8357, KeyReg_Inst_ff_SDE_22_next_state}), .Q ({new_AGEMA_signal_4676, RoundKey[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8359, KeyReg_Inst_ff_SDE_23_next_state}), .Q ({new_AGEMA_signal_4679, RoundKey[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8361, KeyReg_Inst_ff_SDE_24_next_state}), .Q ({new_AGEMA_signal_4682, RoundKey[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8592, KeyReg_Inst_ff_SDE_25_next_state}), .Q ({new_AGEMA_signal_4685, RoundKey[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8594, KeyReg_Inst_ff_SDE_26_next_state}), .Q ({new_AGEMA_signal_4688, RoundKey[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8596, KeyReg_Inst_ff_SDE_27_next_state}), .Q ({new_AGEMA_signal_4691, RoundKey[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8598, KeyReg_Inst_ff_SDE_28_next_state}), .Q ({new_AGEMA_signal_4694, RoundKey[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8600, KeyReg_Inst_ff_SDE_29_next_state}), .Q ({new_AGEMA_signal_4697, RoundKey[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8602, KeyReg_Inst_ff_SDE_30_next_state}), .Q ({new_AGEMA_signal_4703, RoundKey[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8604, KeyReg_Inst_ff_SDE_31_next_state}), .Q ({new_AGEMA_signal_4706, RoundKey[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7874, KeyReg_Inst_ff_SDE_32_next_state}), .Q ({new_AGEMA_signal_4709, RoundKey[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8104, KeyReg_Inst_ff_SDE_33_next_state}), .Q ({new_AGEMA_signal_4712, RoundKey[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8106, KeyReg_Inst_ff_SDE_34_next_state}), .Q ({new_AGEMA_signal_4715, RoundKey[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8108, KeyReg_Inst_ff_SDE_35_next_state}), .Q ({new_AGEMA_signal_4718, RoundKey[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8110, KeyReg_Inst_ff_SDE_36_next_state}), .Q ({new_AGEMA_signal_4721, RoundKey[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8112, KeyReg_Inst_ff_SDE_37_next_state}), .Q ({new_AGEMA_signal_4724, RoundKey[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8114, KeyReg_Inst_ff_SDE_38_next_state}), .Q ({new_AGEMA_signal_4727, RoundKey[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8116, KeyReg_Inst_ff_SDE_39_next_state}), .Q ({new_AGEMA_signal_4730, RoundKey[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7876, KeyReg_Inst_ff_SDE_40_next_state}), .Q ({new_AGEMA_signal_4736, RoundKey[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8118, KeyReg_Inst_ff_SDE_41_next_state}), .Q ({new_AGEMA_signal_4739, RoundKey[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8120, KeyReg_Inst_ff_SDE_42_next_state}), .Q ({new_AGEMA_signal_4742, RoundKey[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8122, KeyReg_Inst_ff_SDE_43_next_state}), .Q ({new_AGEMA_signal_4745, RoundKey[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8124, KeyReg_Inst_ff_SDE_44_next_state}), .Q ({new_AGEMA_signal_4748, RoundKey[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8126, KeyReg_Inst_ff_SDE_45_next_state}), .Q ({new_AGEMA_signal_4751, RoundKey[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8128, KeyReg_Inst_ff_SDE_46_next_state}), .Q ({new_AGEMA_signal_4754, RoundKey[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8130, KeyReg_Inst_ff_SDE_47_next_state}), .Q ({new_AGEMA_signal_4757, RoundKey[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7878, KeyReg_Inst_ff_SDE_48_next_state}), .Q ({new_AGEMA_signal_4760, RoundKey[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8132, KeyReg_Inst_ff_SDE_49_next_state}), .Q ({new_AGEMA_signal_4763, RoundKey[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8134, KeyReg_Inst_ff_SDE_50_next_state}), .Q ({new_AGEMA_signal_4769, RoundKey[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8136, KeyReg_Inst_ff_SDE_51_next_state}), .Q ({new_AGEMA_signal_4772, RoundKey[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8138, KeyReg_Inst_ff_SDE_52_next_state}), .Q ({new_AGEMA_signal_4775, RoundKey[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8140, KeyReg_Inst_ff_SDE_53_next_state}), .Q ({new_AGEMA_signal_4778, RoundKey[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8142, KeyReg_Inst_ff_SDE_54_next_state}), .Q ({new_AGEMA_signal_4781, RoundKey[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8144, KeyReg_Inst_ff_SDE_55_next_state}), .Q ({new_AGEMA_signal_4784, RoundKey[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8146, KeyReg_Inst_ff_SDE_56_next_state}), .Q ({new_AGEMA_signal_4787, RoundKey[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8363, KeyReg_Inst_ff_SDE_57_next_state}), .Q ({new_AGEMA_signal_4790, RoundKey[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8365, KeyReg_Inst_ff_SDE_58_next_state}), .Q ({new_AGEMA_signal_4793, RoundKey[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8367, KeyReg_Inst_ff_SDE_59_next_state}), .Q ({new_AGEMA_signal_4796, RoundKey[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8369, KeyReg_Inst_ff_SDE_60_next_state}), .Q ({new_AGEMA_signal_4802, RoundKey[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8371, KeyReg_Inst_ff_SDE_61_next_state}), .Q ({new_AGEMA_signal_4805, RoundKey[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8373, KeyReg_Inst_ff_SDE_62_next_state}), .Q ({new_AGEMA_signal_4808, RoundKey[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8375, KeyReg_Inst_ff_SDE_63_next_state}), .Q ({new_AGEMA_signal_4811, RoundKey[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7664, KeyReg_Inst_ff_SDE_64_next_state}), .Q ({new_AGEMA_signal_4814, RoundKey[64]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7880, KeyReg_Inst_ff_SDE_65_next_state}), .Q ({new_AGEMA_signal_4817, RoundKey[65]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7882, KeyReg_Inst_ff_SDE_66_next_state}), .Q ({new_AGEMA_signal_4820, RoundKey[66]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7884, KeyReg_Inst_ff_SDE_67_next_state}), .Q ({new_AGEMA_signal_4823, RoundKey[67]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7886, KeyReg_Inst_ff_SDE_68_next_state}), .Q ({new_AGEMA_signal_4826, RoundKey[68]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7888, KeyReg_Inst_ff_SDE_69_next_state}), .Q ({new_AGEMA_signal_4829, RoundKey[69]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7890, KeyReg_Inst_ff_SDE_70_next_state}), .Q ({new_AGEMA_signal_4835, RoundKey[70]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7892, KeyReg_Inst_ff_SDE_71_next_state}), .Q ({new_AGEMA_signal_4838, RoundKey[71]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7666, KeyReg_Inst_ff_SDE_72_next_state}), .Q ({new_AGEMA_signal_4841, RoundKey[72]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7894, KeyReg_Inst_ff_SDE_73_next_state}), .Q ({new_AGEMA_signal_4844, RoundKey[73]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7896, KeyReg_Inst_ff_SDE_74_next_state}), .Q ({new_AGEMA_signal_4847, RoundKey[74]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7898, KeyReg_Inst_ff_SDE_75_next_state}), .Q ({new_AGEMA_signal_4850, RoundKey[75]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7900, KeyReg_Inst_ff_SDE_76_next_state}), .Q ({new_AGEMA_signal_4853, RoundKey[76]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7902, KeyReg_Inst_ff_SDE_77_next_state}), .Q ({new_AGEMA_signal_4856, RoundKey[77]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7904, KeyReg_Inst_ff_SDE_78_next_state}), .Q ({new_AGEMA_signal_4859, RoundKey[78]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7906, KeyReg_Inst_ff_SDE_79_next_state}), .Q ({new_AGEMA_signal_4862, RoundKey[79]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7668, KeyReg_Inst_ff_SDE_80_next_state}), .Q ({new_AGEMA_signal_4868, RoundKey[80]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7908, KeyReg_Inst_ff_SDE_81_next_state}), .Q ({new_AGEMA_signal_4871, RoundKey[81]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7910, KeyReg_Inst_ff_SDE_82_next_state}), .Q ({new_AGEMA_signal_4874, RoundKey[82]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7912, KeyReg_Inst_ff_SDE_83_next_state}), .Q ({new_AGEMA_signal_4877, RoundKey[83]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7914, KeyReg_Inst_ff_SDE_84_next_state}), .Q ({new_AGEMA_signal_4880, RoundKey[84]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7916, KeyReg_Inst_ff_SDE_85_next_state}), .Q ({new_AGEMA_signal_4883, RoundKey[85]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7918, KeyReg_Inst_ff_SDE_86_next_state}), .Q ({new_AGEMA_signal_4886, RoundKey[86]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7920, KeyReg_Inst_ff_SDE_87_next_state}), .Q ({new_AGEMA_signal_4889, RoundKey[87]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7922, KeyReg_Inst_ff_SDE_88_next_state}), .Q ({new_AGEMA_signal_4892, RoundKey[88]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8148, KeyReg_Inst_ff_SDE_89_next_state}), .Q ({new_AGEMA_signal_4895, RoundKey[89]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8150, KeyReg_Inst_ff_SDE_90_next_state}), .Q ({new_AGEMA_signal_4901, RoundKey[90]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8152, KeyReg_Inst_ff_SDE_91_next_state}), .Q ({new_AGEMA_signal_4904, RoundKey[91]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8154, KeyReg_Inst_ff_SDE_92_next_state}), .Q ({new_AGEMA_signal_4907, RoundKey[92]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8156, KeyReg_Inst_ff_SDE_93_next_state}), .Q ({new_AGEMA_signal_4910, RoundKey[93]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8158, KeyReg_Inst_ff_SDE_94_next_state}), .Q ({new_AGEMA_signal_4913, RoundKey[94]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_8160, KeyReg_Inst_ff_SDE_95_next_state}), .Q ({new_AGEMA_signal_4916, RoundKey[95]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7498, KeyReg_Inst_ff_SDE_96_next_state}), .Q ({new_AGEMA_signal_4919, RoundKey[96]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7670, KeyReg_Inst_ff_SDE_97_next_state}), .Q ({new_AGEMA_signal_4922, RoundKey[97]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7672, KeyReg_Inst_ff_SDE_98_next_state}), .Q ({new_AGEMA_signal_4925, RoundKey[98]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7674, KeyReg_Inst_ff_SDE_99_next_state}), .Q ({new_AGEMA_signal_4928, RoundKey[99]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7676, KeyReg_Inst_ff_SDE_100_next_state}), .Q ({new_AGEMA_signal_4553, RoundKey[100]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7678, KeyReg_Inst_ff_SDE_101_next_state}), .Q ({new_AGEMA_signal_4556, RoundKey[101]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7680, KeyReg_Inst_ff_SDE_102_next_state}), .Q ({new_AGEMA_signal_4559, RoundKey[102]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7682, KeyReg_Inst_ff_SDE_103_next_state}), .Q ({new_AGEMA_signal_4562, RoundKey[103]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7500, KeyReg_Inst_ff_SDE_104_next_state}), .Q ({new_AGEMA_signal_4565, RoundKey[104]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7684, KeyReg_Inst_ff_SDE_105_next_state}), .Q ({new_AGEMA_signal_4568, RoundKey[105]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7686, KeyReg_Inst_ff_SDE_106_next_state}), .Q ({new_AGEMA_signal_4571, RoundKey[106]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7688, KeyReg_Inst_ff_SDE_107_next_state}), .Q ({new_AGEMA_signal_4574, RoundKey[107]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7690, KeyReg_Inst_ff_SDE_108_next_state}), .Q ({new_AGEMA_signal_4577, RoundKey[108]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7692, KeyReg_Inst_ff_SDE_109_next_state}), .Q ({new_AGEMA_signal_4580, RoundKey[109]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7694, KeyReg_Inst_ff_SDE_110_next_state}), .Q ({new_AGEMA_signal_4586, RoundKey[110]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7696, KeyReg_Inst_ff_SDE_111_next_state}), .Q ({new_AGEMA_signal_4589, RoundKey[111]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7502, KeyReg_Inst_ff_SDE_112_next_state}), .Q ({new_AGEMA_signal_4592, RoundKey[112]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7698, KeyReg_Inst_ff_SDE_113_next_state}), .Q ({new_AGEMA_signal_4595, RoundKey[113]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7700, KeyReg_Inst_ff_SDE_114_next_state}), .Q ({new_AGEMA_signal_4598, RoundKey[114]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7702, KeyReg_Inst_ff_SDE_115_next_state}), .Q ({new_AGEMA_signal_4601, RoundKey[115]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7704, KeyReg_Inst_ff_SDE_116_next_state}), .Q ({new_AGEMA_signal_4604, RoundKey[116]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7706, KeyReg_Inst_ff_SDE_117_next_state}), .Q ({new_AGEMA_signal_4607, RoundKey[117]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7708, KeyReg_Inst_ff_SDE_118_next_state}), .Q ({new_AGEMA_signal_4610, RoundKey[118]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7710, KeyReg_Inst_ff_SDE_119_next_state}), .Q ({new_AGEMA_signal_4613, RoundKey[119]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7712, KeyReg_Inst_ff_SDE_120_next_state}), .Q ({new_AGEMA_signal_4619, RoundKey[120]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7924, KeyReg_Inst_ff_SDE_121_next_state}), .Q ({new_AGEMA_signal_4622, RoundKey[121]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7926, KeyReg_Inst_ff_SDE_122_next_state}), .Q ({new_AGEMA_signal_4625, RoundKey[122]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7928, KeyReg_Inst_ff_SDE_123_next_state}), .Q ({new_AGEMA_signal_4628, RoundKey[123]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7930, KeyReg_Inst_ff_SDE_124_next_state}), .Q ({new_AGEMA_signal_4631, RoundKey[124]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7932, KeyReg_Inst_ff_SDE_125_next_state}), .Q ({new_AGEMA_signal_4634, RoundKey[125]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7934, KeyReg_Inst_ff_SDE_126_next_state}), .Q ({new_AGEMA_signal_4637, RoundKey[126]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_7936, KeyReg_Inst_ff_SDE_127_next_state}), .Q ({new_AGEMA_signal_4640, RoundKey[127]}) ) ;
    DFF_X1 RoundCounterIns_count_reg_0__FF_FF ( .CK (clk_gated), .D (RoundCounterIns_N7), .Q (RoundCounter[0]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_1__FF_FF ( .CK (clk_gated), .D (RoundCounterIns_N8), .Q (RoundCounter[1]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_2__FF_FF ( .CK (clk_gated), .D (RoundCounterIns_n1), .Q (RoundCounter[2]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_3__FF_FF ( .CK (clk_gated), .D (RoundCounterIns_N10), .Q (RoundCounter[3]), .QN () ) ;
endmodule
