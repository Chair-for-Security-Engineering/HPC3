////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module AES in file /AGEMA/Designs/AES_round-based/AGEMA/AES.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module AES_HPC2_ClockGating_d2 (plaintext_s0, key_s0, clk, reset, key_s1, key_s2, plaintext_s1, plaintext_s2, Fresh, ciphertext_s0, done, ciphertext_s1, ciphertext_s2, Synch);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] key_s1 ;
    input [127:0] key_s2 ;
    input [127:0] plaintext_s1 ;
    input [127:0] plaintext_s2 ;
    input [2039:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    output [127:0] ciphertext_s2 ;
    output Synch ;
    wire n283 ;
    wire n285 ;
    wire n314 ;
    wire n315 ;
    wire n316 ;
    wire n317 ;
    wire n318 ;
    wire n319 ;
    wire n320 ;
    wire n321 ;
    wire n322 ;
    wire n323 ;
    wire n324 ;
    wire n325 ;
    wire n326 ;
    wire n327 ;
    wire n328 ;
    wire n329 ;
    wire n330 ;
    wire n331 ;
    wire n332 ;
    wire n333 ;
    wire n334 ;
    wire n335 ;
    wire n336 ;
    wire n337 ;
    wire n338 ;
    wire n339 ;
    wire RoundReg_Inst_ff_SDE_0_next_state ;
    wire RoundReg_Inst_ff_SDE_1_next_state ;
    wire RoundReg_Inst_ff_SDE_2_next_state ;
    wire RoundReg_Inst_ff_SDE_3_next_state ;
    wire RoundReg_Inst_ff_SDE_4_next_state ;
    wire RoundReg_Inst_ff_SDE_5_next_state ;
    wire RoundReg_Inst_ff_SDE_6_next_state ;
    wire RoundReg_Inst_ff_SDE_7_next_state ;
    wire RoundReg_Inst_ff_SDE_8_next_state ;
    wire RoundReg_Inst_ff_SDE_9_next_state ;
    wire RoundReg_Inst_ff_SDE_10_next_state ;
    wire RoundReg_Inst_ff_SDE_11_next_state ;
    wire RoundReg_Inst_ff_SDE_12_next_state ;
    wire RoundReg_Inst_ff_SDE_13_next_state ;
    wire RoundReg_Inst_ff_SDE_14_next_state ;
    wire RoundReg_Inst_ff_SDE_15_next_state ;
    wire RoundReg_Inst_ff_SDE_16_next_state ;
    wire RoundReg_Inst_ff_SDE_17_next_state ;
    wire RoundReg_Inst_ff_SDE_18_next_state ;
    wire RoundReg_Inst_ff_SDE_19_next_state ;
    wire RoundReg_Inst_ff_SDE_20_next_state ;
    wire RoundReg_Inst_ff_SDE_21_next_state ;
    wire RoundReg_Inst_ff_SDE_22_next_state ;
    wire RoundReg_Inst_ff_SDE_23_next_state ;
    wire RoundReg_Inst_ff_SDE_24_next_state ;
    wire RoundReg_Inst_ff_SDE_25_next_state ;
    wire RoundReg_Inst_ff_SDE_26_next_state ;
    wire RoundReg_Inst_ff_SDE_27_next_state ;
    wire RoundReg_Inst_ff_SDE_28_next_state ;
    wire RoundReg_Inst_ff_SDE_29_next_state ;
    wire RoundReg_Inst_ff_SDE_30_next_state ;
    wire RoundReg_Inst_ff_SDE_31_next_state ;
    wire RoundReg_Inst_ff_SDE_32_next_state ;
    wire RoundReg_Inst_ff_SDE_33_next_state ;
    wire RoundReg_Inst_ff_SDE_34_next_state ;
    wire RoundReg_Inst_ff_SDE_35_next_state ;
    wire RoundReg_Inst_ff_SDE_36_next_state ;
    wire RoundReg_Inst_ff_SDE_37_next_state ;
    wire RoundReg_Inst_ff_SDE_38_next_state ;
    wire RoundReg_Inst_ff_SDE_39_next_state ;
    wire RoundReg_Inst_ff_SDE_40_next_state ;
    wire RoundReg_Inst_ff_SDE_41_next_state ;
    wire RoundReg_Inst_ff_SDE_42_next_state ;
    wire RoundReg_Inst_ff_SDE_43_next_state ;
    wire RoundReg_Inst_ff_SDE_44_next_state ;
    wire RoundReg_Inst_ff_SDE_45_next_state ;
    wire RoundReg_Inst_ff_SDE_46_next_state ;
    wire RoundReg_Inst_ff_SDE_47_next_state ;
    wire RoundReg_Inst_ff_SDE_48_next_state ;
    wire RoundReg_Inst_ff_SDE_49_next_state ;
    wire RoundReg_Inst_ff_SDE_50_next_state ;
    wire RoundReg_Inst_ff_SDE_51_next_state ;
    wire RoundReg_Inst_ff_SDE_52_next_state ;
    wire RoundReg_Inst_ff_SDE_53_next_state ;
    wire RoundReg_Inst_ff_SDE_54_next_state ;
    wire RoundReg_Inst_ff_SDE_55_next_state ;
    wire RoundReg_Inst_ff_SDE_56_next_state ;
    wire RoundReg_Inst_ff_SDE_57_next_state ;
    wire RoundReg_Inst_ff_SDE_58_next_state ;
    wire RoundReg_Inst_ff_SDE_59_next_state ;
    wire RoundReg_Inst_ff_SDE_60_next_state ;
    wire RoundReg_Inst_ff_SDE_61_next_state ;
    wire RoundReg_Inst_ff_SDE_62_next_state ;
    wire RoundReg_Inst_ff_SDE_63_next_state ;
    wire RoundReg_Inst_ff_SDE_64_next_state ;
    wire RoundReg_Inst_ff_SDE_65_next_state ;
    wire RoundReg_Inst_ff_SDE_66_next_state ;
    wire RoundReg_Inst_ff_SDE_67_next_state ;
    wire RoundReg_Inst_ff_SDE_68_next_state ;
    wire RoundReg_Inst_ff_SDE_69_next_state ;
    wire RoundReg_Inst_ff_SDE_70_next_state ;
    wire RoundReg_Inst_ff_SDE_71_next_state ;
    wire RoundReg_Inst_ff_SDE_72_next_state ;
    wire RoundReg_Inst_ff_SDE_73_next_state ;
    wire RoundReg_Inst_ff_SDE_74_next_state ;
    wire RoundReg_Inst_ff_SDE_75_next_state ;
    wire RoundReg_Inst_ff_SDE_76_next_state ;
    wire RoundReg_Inst_ff_SDE_77_next_state ;
    wire RoundReg_Inst_ff_SDE_78_next_state ;
    wire RoundReg_Inst_ff_SDE_79_next_state ;
    wire RoundReg_Inst_ff_SDE_80_next_state ;
    wire RoundReg_Inst_ff_SDE_81_next_state ;
    wire RoundReg_Inst_ff_SDE_82_next_state ;
    wire RoundReg_Inst_ff_SDE_83_next_state ;
    wire RoundReg_Inst_ff_SDE_84_next_state ;
    wire RoundReg_Inst_ff_SDE_85_next_state ;
    wire RoundReg_Inst_ff_SDE_86_next_state ;
    wire RoundReg_Inst_ff_SDE_87_next_state ;
    wire RoundReg_Inst_ff_SDE_88_next_state ;
    wire RoundReg_Inst_ff_SDE_89_next_state ;
    wire RoundReg_Inst_ff_SDE_90_next_state ;
    wire RoundReg_Inst_ff_SDE_91_next_state ;
    wire RoundReg_Inst_ff_SDE_92_next_state ;
    wire RoundReg_Inst_ff_SDE_93_next_state ;
    wire RoundReg_Inst_ff_SDE_94_next_state ;
    wire RoundReg_Inst_ff_SDE_95_next_state ;
    wire RoundReg_Inst_ff_SDE_96_next_state ;
    wire RoundReg_Inst_ff_SDE_97_next_state ;
    wire RoundReg_Inst_ff_SDE_98_next_state ;
    wire RoundReg_Inst_ff_SDE_99_next_state ;
    wire RoundReg_Inst_ff_SDE_100_next_state ;
    wire RoundReg_Inst_ff_SDE_101_next_state ;
    wire RoundReg_Inst_ff_SDE_102_next_state ;
    wire RoundReg_Inst_ff_SDE_103_next_state ;
    wire RoundReg_Inst_ff_SDE_104_next_state ;
    wire RoundReg_Inst_ff_SDE_105_next_state ;
    wire RoundReg_Inst_ff_SDE_106_next_state ;
    wire RoundReg_Inst_ff_SDE_107_next_state ;
    wire RoundReg_Inst_ff_SDE_108_next_state ;
    wire RoundReg_Inst_ff_SDE_109_next_state ;
    wire RoundReg_Inst_ff_SDE_110_next_state ;
    wire RoundReg_Inst_ff_SDE_111_next_state ;
    wire RoundReg_Inst_ff_SDE_112_next_state ;
    wire RoundReg_Inst_ff_SDE_113_next_state ;
    wire RoundReg_Inst_ff_SDE_114_next_state ;
    wire RoundReg_Inst_ff_SDE_115_next_state ;
    wire RoundReg_Inst_ff_SDE_116_next_state ;
    wire RoundReg_Inst_ff_SDE_117_next_state ;
    wire RoundReg_Inst_ff_SDE_118_next_state ;
    wire RoundReg_Inst_ff_SDE_119_next_state ;
    wire RoundReg_Inst_ff_SDE_120_next_state ;
    wire RoundReg_Inst_ff_SDE_121_next_state ;
    wire RoundReg_Inst_ff_SDE_122_next_state ;
    wire RoundReg_Inst_ff_SDE_123_next_state ;
    wire RoundReg_Inst_ff_SDE_124_next_state ;
    wire RoundReg_Inst_ff_SDE_125_next_state ;
    wire RoundReg_Inst_ff_SDE_126_next_state ;
    wire RoundReg_Inst_ff_SDE_127_next_state ;
    wire SubBytesIns_Inst_Sbox_0_L29 ;
    wire SubBytesIns_Inst_Sbox_0_L28 ;
    wire SubBytesIns_Inst_Sbox_0_L27 ;
    wire SubBytesIns_Inst_Sbox_0_L26 ;
    wire SubBytesIns_Inst_Sbox_0_L25 ;
    wire SubBytesIns_Inst_Sbox_0_L24 ;
    wire SubBytesIns_Inst_Sbox_0_L23 ;
    wire SubBytesIns_Inst_Sbox_0_L22 ;
    wire SubBytesIns_Inst_Sbox_0_L21 ;
    wire SubBytesIns_Inst_Sbox_0_L20 ;
    wire SubBytesIns_Inst_Sbox_0_L19 ;
    wire SubBytesIns_Inst_Sbox_0_L18 ;
    wire SubBytesIns_Inst_Sbox_0_L17 ;
    wire SubBytesIns_Inst_Sbox_0_L16 ;
    wire SubBytesIns_Inst_Sbox_0_L15 ;
    wire SubBytesIns_Inst_Sbox_0_L14 ;
    wire SubBytesIns_Inst_Sbox_0_L13 ;
    wire SubBytesIns_Inst_Sbox_0_L12 ;
    wire SubBytesIns_Inst_Sbox_0_L11 ;
    wire SubBytesIns_Inst_Sbox_0_L10 ;
    wire SubBytesIns_Inst_Sbox_0_L9 ;
    wire SubBytesIns_Inst_Sbox_0_L8 ;
    wire SubBytesIns_Inst_Sbox_0_L7 ;
    wire SubBytesIns_Inst_Sbox_0_L6 ;
    wire SubBytesIns_Inst_Sbox_0_L5 ;
    wire SubBytesIns_Inst_Sbox_0_L4 ;
    wire SubBytesIns_Inst_Sbox_0_L3 ;
    wire SubBytesIns_Inst_Sbox_0_L2 ;
    wire SubBytesIns_Inst_Sbox_0_L1 ;
    wire SubBytesIns_Inst_Sbox_0_L0 ;
    wire SubBytesIns_Inst_Sbox_0_M63 ;
    wire SubBytesIns_Inst_Sbox_0_M62 ;
    wire SubBytesIns_Inst_Sbox_0_M61 ;
    wire SubBytesIns_Inst_Sbox_0_M60 ;
    wire SubBytesIns_Inst_Sbox_0_M59 ;
    wire SubBytesIns_Inst_Sbox_0_M58 ;
    wire SubBytesIns_Inst_Sbox_0_M57 ;
    wire SubBytesIns_Inst_Sbox_0_M56 ;
    wire SubBytesIns_Inst_Sbox_0_M55 ;
    wire SubBytesIns_Inst_Sbox_0_M54 ;
    wire SubBytesIns_Inst_Sbox_0_M53 ;
    wire SubBytesIns_Inst_Sbox_0_M52 ;
    wire SubBytesIns_Inst_Sbox_0_M51 ;
    wire SubBytesIns_Inst_Sbox_0_M50 ;
    wire SubBytesIns_Inst_Sbox_0_M49 ;
    wire SubBytesIns_Inst_Sbox_0_M48 ;
    wire SubBytesIns_Inst_Sbox_0_M47 ;
    wire SubBytesIns_Inst_Sbox_0_M46 ;
    wire SubBytesIns_Inst_Sbox_0_M45 ;
    wire SubBytesIns_Inst_Sbox_0_M44 ;
    wire SubBytesIns_Inst_Sbox_0_M43 ;
    wire SubBytesIns_Inst_Sbox_0_M42 ;
    wire SubBytesIns_Inst_Sbox_0_M41 ;
    wire SubBytesIns_Inst_Sbox_0_M40 ;
    wire SubBytesIns_Inst_Sbox_0_M39 ;
    wire SubBytesIns_Inst_Sbox_0_M38 ;
    wire SubBytesIns_Inst_Sbox_0_M37 ;
    wire SubBytesIns_Inst_Sbox_0_M36 ;
    wire SubBytesIns_Inst_Sbox_0_M35 ;
    wire SubBytesIns_Inst_Sbox_0_M34 ;
    wire SubBytesIns_Inst_Sbox_0_M33 ;
    wire SubBytesIns_Inst_Sbox_0_M32 ;
    wire SubBytesIns_Inst_Sbox_0_M31 ;
    wire SubBytesIns_Inst_Sbox_0_M30 ;
    wire SubBytesIns_Inst_Sbox_0_M29 ;
    wire SubBytesIns_Inst_Sbox_0_M28 ;
    wire SubBytesIns_Inst_Sbox_0_M27 ;
    wire SubBytesIns_Inst_Sbox_0_M26 ;
    wire SubBytesIns_Inst_Sbox_0_M25 ;
    wire SubBytesIns_Inst_Sbox_0_M24 ;
    wire SubBytesIns_Inst_Sbox_0_M23 ;
    wire SubBytesIns_Inst_Sbox_0_M22 ;
    wire SubBytesIns_Inst_Sbox_0_M21 ;
    wire SubBytesIns_Inst_Sbox_0_M20 ;
    wire SubBytesIns_Inst_Sbox_0_M19 ;
    wire SubBytesIns_Inst_Sbox_0_M18 ;
    wire SubBytesIns_Inst_Sbox_0_M17 ;
    wire SubBytesIns_Inst_Sbox_0_M16 ;
    wire SubBytesIns_Inst_Sbox_0_M15 ;
    wire SubBytesIns_Inst_Sbox_0_M14 ;
    wire SubBytesIns_Inst_Sbox_0_M13 ;
    wire SubBytesIns_Inst_Sbox_0_M12 ;
    wire SubBytesIns_Inst_Sbox_0_M11 ;
    wire SubBytesIns_Inst_Sbox_0_M10 ;
    wire SubBytesIns_Inst_Sbox_0_M9 ;
    wire SubBytesIns_Inst_Sbox_0_M8 ;
    wire SubBytesIns_Inst_Sbox_0_M7 ;
    wire SubBytesIns_Inst_Sbox_0_M6 ;
    wire SubBytesIns_Inst_Sbox_0_M5 ;
    wire SubBytesIns_Inst_Sbox_0_M4 ;
    wire SubBytesIns_Inst_Sbox_0_M3 ;
    wire SubBytesIns_Inst_Sbox_0_M2 ;
    wire SubBytesIns_Inst_Sbox_0_M1 ;
    wire SubBytesIns_Inst_Sbox_0_T27 ;
    wire SubBytesIns_Inst_Sbox_0_T26 ;
    wire SubBytesIns_Inst_Sbox_0_T25 ;
    wire SubBytesIns_Inst_Sbox_0_T24 ;
    wire SubBytesIns_Inst_Sbox_0_T23 ;
    wire SubBytesIns_Inst_Sbox_0_T22 ;
    wire SubBytesIns_Inst_Sbox_0_T21 ;
    wire SubBytesIns_Inst_Sbox_0_T20 ;
    wire SubBytesIns_Inst_Sbox_0_T19 ;
    wire SubBytesIns_Inst_Sbox_0_T18 ;
    wire SubBytesIns_Inst_Sbox_0_T17 ;
    wire SubBytesIns_Inst_Sbox_0_T16 ;
    wire SubBytesIns_Inst_Sbox_0_T15 ;
    wire SubBytesIns_Inst_Sbox_0_T14 ;
    wire SubBytesIns_Inst_Sbox_0_T13 ;
    wire SubBytesIns_Inst_Sbox_0_T12 ;
    wire SubBytesIns_Inst_Sbox_0_T11 ;
    wire SubBytesIns_Inst_Sbox_0_T10 ;
    wire SubBytesIns_Inst_Sbox_0_T9 ;
    wire SubBytesIns_Inst_Sbox_0_T8 ;
    wire SubBytesIns_Inst_Sbox_0_T7 ;
    wire SubBytesIns_Inst_Sbox_0_T6 ;
    wire SubBytesIns_Inst_Sbox_0_T5 ;
    wire SubBytesIns_Inst_Sbox_0_T4 ;
    wire SubBytesIns_Inst_Sbox_0_T3 ;
    wire SubBytesIns_Inst_Sbox_0_T2 ;
    wire SubBytesIns_Inst_Sbox_0_T1 ;
    wire SubBytesIns_Inst_Sbox_1_L29 ;
    wire SubBytesIns_Inst_Sbox_1_L28 ;
    wire SubBytesIns_Inst_Sbox_1_L27 ;
    wire SubBytesIns_Inst_Sbox_1_L26 ;
    wire SubBytesIns_Inst_Sbox_1_L25 ;
    wire SubBytesIns_Inst_Sbox_1_L24 ;
    wire SubBytesIns_Inst_Sbox_1_L23 ;
    wire SubBytesIns_Inst_Sbox_1_L22 ;
    wire SubBytesIns_Inst_Sbox_1_L21 ;
    wire SubBytesIns_Inst_Sbox_1_L20 ;
    wire SubBytesIns_Inst_Sbox_1_L19 ;
    wire SubBytesIns_Inst_Sbox_1_L18 ;
    wire SubBytesIns_Inst_Sbox_1_L17 ;
    wire SubBytesIns_Inst_Sbox_1_L16 ;
    wire SubBytesIns_Inst_Sbox_1_L15 ;
    wire SubBytesIns_Inst_Sbox_1_L14 ;
    wire SubBytesIns_Inst_Sbox_1_L13 ;
    wire SubBytesIns_Inst_Sbox_1_L12 ;
    wire SubBytesIns_Inst_Sbox_1_L11 ;
    wire SubBytesIns_Inst_Sbox_1_L10 ;
    wire SubBytesIns_Inst_Sbox_1_L9 ;
    wire SubBytesIns_Inst_Sbox_1_L8 ;
    wire SubBytesIns_Inst_Sbox_1_L7 ;
    wire SubBytesIns_Inst_Sbox_1_L6 ;
    wire SubBytesIns_Inst_Sbox_1_L5 ;
    wire SubBytesIns_Inst_Sbox_1_L4 ;
    wire SubBytesIns_Inst_Sbox_1_L3 ;
    wire SubBytesIns_Inst_Sbox_1_L2 ;
    wire SubBytesIns_Inst_Sbox_1_L1 ;
    wire SubBytesIns_Inst_Sbox_1_L0 ;
    wire SubBytesIns_Inst_Sbox_1_M63 ;
    wire SubBytesIns_Inst_Sbox_1_M62 ;
    wire SubBytesIns_Inst_Sbox_1_M61 ;
    wire SubBytesIns_Inst_Sbox_1_M60 ;
    wire SubBytesIns_Inst_Sbox_1_M59 ;
    wire SubBytesIns_Inst_Sbox_1_M58 ;
    wire SubBytesIns_Inst_Sbox_1_M57 ;
    wire SubBytesIns_Inst_Sbox_1_M56 ;
    wire SubBytesIns_Inst_Sbox_1_M55 ;
    wire SubBytesIns_Inst_Sbox_1_M54 ;
    wire SubBytesIns_Inst_Sbox_1_M53 ;
    wire SubBytesIns_Inst_Sbox_1_M52 ;
    wire SubBytesIns_Inst_Sbox_1_M51 ;
    wire SubBytesIns_Inst_Sbox_1_M50 ;
    wire SubBytesIns_Inst_Sbox_1_M49 ;
    wire SubBytesIns_Inst_Sbox_1_M48 ;
    wire SubBytesIns_Inst_Sbox_1_M47 ;
    wire SubBytesIns_Inst_Sbox_1_M46 ;
    wire SubBytesIns_Inst_Sbox_1_M45 ;
    wire SubBytesIns_Inst_Sbox_1_M44 ;
    wire SubBytesIns_Inst_Sbox_1_M43 ;
    wire SubBytesIns_Inst_Sbox_1_M42 ;
    wire SubBytesIns_Inst_Sbox_1_M41 ;
    wire SubBytesIns_Inst_Sbox_1_M40 ;
    wire SubBytesIns_Inst_Sbox_1_M39 ;
    wire SubBytesIns_Inst_Sbox_1_M38 ;
    wire SubBytesIns_Inst_Sbox_1_M37 ;
    wire SubBytesIns_Inst_Sbox_1_M36 ;
    wire SubBytesIns_Inst_Sbox_1_M35 ;
    wire SubBytesIns_Inst_Sbox_1_M34 ;
    wire SubBytesIns_Inst_Sbox_1_M33 ;
    wire SubBytesIns_Inst_Sbox_1_M32 ;
    wire SubBytesIns_Inst_Sbox_1_M31 ;
    wire SubBytesIns_Inst_Sbox_1_M30 ;
    wire SubBytesIns_Inst_Sbox_1_M29 ;
    wire SubBytesIns_Inst_Sbox_1_M28 ;
    wire SubBytesIns_Inst_Sbox_1_M27 ;
    wire SubBytesIns_Inst_Sbox_1_M26 ;
    wire SubBytesIns_Inst_Sbox_1_M25 ;
    wire SubBytesIns_Inst_Sbox_1_M24 ;
    wire SubBytesIns_Inst_Sbox_1_M23 ;
    wire SubBytesIns_Inst_Sbox_1_M22 ;
    wire SubBytesIns_Inst_Sbox_1_M21 ;
    wire SubBytesIns_Inst_Sbox_1_M20 ;
    wire SubBytesIns_Inst_Sbox_1_M19 ;
    wire SubBytesIns_Inst_Sbox_1_M18 ;
    wire SubBytesIns_Inst_Sbox_1_M17 ;
    wire SubBytesIns_Inst_Sbox_1_M16 ;
    wire SubBytesIns_Inst_Sbox_1_M15 ;
    wire SubBytesIns_Inst_Sbox_1_M14 ;
    wire SubBytesIns_Inst_Sbox_1_M13 ;
    wire SubBytesIns_Inst_Sbox_1_M12 ;
    wire SubBytesIns_Inst_Sbox_1_M11 ;
    wire SubBytesIns_Inst_Sbox_1_M10 ;
    wire SubBytesIns_Inst_Sbox_1_M9 ;
    wire SubBytesIns_Inst_Sbox_1_M8 ;
    wire SubBytesIns_Inst_Sbox_1_M7 ;
    wire SubBytesIns_Inst_Sbox_1_M6 ;
    wire SubBytesIns_Inst_Sbox_1_M5 ;
    wire SubBytesIns_Inst_Sbox_1_M4 ;
    wire SubBytesIns_Inst_Sbox_1_M3 ;
    wire SubBytesIns_Inst_Sbox_1_M2 ;
    wire SubBytesIns_Inst_Sbox_1_M1 ;
    wire SubBytesIns_Inst_Sbox_1_T27 ;
    wire SubBytesIns_Inst_Sbox_1_T26 ;
    wire SubBytesIns_Inst_Sbox_1_T25 ;
    wire SubBytesIns_Inst_Sbox_1_T24 ;
    wire SubBytesIns_Inst_Sbox_1_T23 ;
    wire SubBytesIns_Inst_Sbox_1_T22 ;
    wire SubBytesIns_Inst_Sbox_1_T21 ;
    wire SubBytesIns_Inst_Sbox_1_T20 ;
    wire SubBytesIns_Inst_Sbox_1_T19 ;
    wire SubBytesIns_Inst_Sbox_1_T18 ;
    wire SubBytesIns_Inst_Sbox_1_T17 ;
    wire SubBytesIns_Inst_Sbox_1_T16 ;
    wire SubBytesIns_Inst_Sbox_1_T15 ;
    wire SubBytesIns_Inst_Sbox_1_T14 ;
    wire SubBytesIns_Inst_Sbox_1_T13 ;
    wire SubBytesIns_Inst_Sbox_1_T12 ;
    wire SubBytesIns_Inst_Sbox_1_T11 ;
    wire SubBytesIns_Inst_Sbox_1_T10 ;
    wire SubBytesIns_Inst_Sbox_1_T9 ;
    wire SubBytesIns_Inst_Sbox_1_T8 ;
    wire SubBytesIns_Inst_Sbox_1_T7 ;
    wire SubBytesIns_Inst_Sbox_1_T6 ;
    wire SubBytesIns_Inst_Sbox_1_T5 ;
    wire SubBytesIns_Inst_Sbox_1_T4 ;
    wire SubBytesIns_Inst_Sbox_1_T3 ;
    wire SubBytesIns_Inst_Sbox_1_T2 ;
    wire SubBytesIns_Inst_Sbox_1_T1 ;
    wire SubBytesIns_Inst_Sbox_2_L29 ;
    wire SubBytesIns_Inst_Sbox_2_L28 ;
    wire SubBytesIns_Inst_Sbox_2_L27 ;
    wire SubBytesIns_Inst_Sbox_2_L26 ;
    wire SubBytesIns_Inst_Sbox_2_L25 ;
    wire SubBytesIns_Inst_Sbox_2_L24 ;
    wire SubBytesIns_Inst_Sbox_2_L23 ;
    wire SubBytesIns_Inst_Sbox_2_L22 ;
    wire SubBytesIns_Inst_Sbox_2_L21 ;
    wire SubBytesIns_Inst_Sbox_2_L20 ;
    wire SubBytesIns_Inst_Sbox_2_L19 ;
    wire SubBytesIns_Inst_Sbox_2_L18 ;
    wire SubBytesIns_Inst_Sbox_2_L17 ;
    wire SubBytesIns_Inst_Sbox_2_L16 ;
    wire SubBytesIns_Inst_Sbox_2_L15 ;
    wire SubBytesIns_Inst_Sbox_2_L14 ;
    wire SubBytesIns_Inst_Sbox_2_L13 ;
    wire SubBytesIns_Inst_Sbox_2_L12 ;
    wire SubBytesIns_Inst_Sbox_2_L11 ;
    wire SubBytesIns_Inst_Sbox_2_L10 ;
    wire SubBytesIns_Inst_Sbox_2_L9 ;
    wire SubBytesIns_Inst_Sbox_2_L8 ;
    wire SubBytesIns_Inst_Sbox_2_L7 ;
    wire SubBytesIns_Inst_Sbox_2_L6 ;
    wire SubBytesIns_Inst_Sbox_2_L5 ;
    wire SubBytesIns_Inst_Sbox_2_L4 ;
    wire SubBytesIns_Inst_Sbox_2_L3 ;
    wire SubBytesIns_Inst_Sbox_2_L2 ;
    wire SubBytesIns_Inst_Sbox_2_L1 ;
    wire SubBytesIns_Inst_Sbox_2_L0 ;
    wire SubBytesIns_Inst_Sbox_2_M63 ;
    wire SubBytesIns_Inst_Sbox_2_M62 ;
    wire SubBytesIns_Inst_Sbox_2_M61 ;
    wire SubBytesIns_Inst_Sbox_2_M60 ;
    wire SubBytesIns_Inst_Sbox_2_M59 ;
    wire SubBytesIns_Inst_Sbox_2_M58 ;
    wire SubBytesIns_Inst_Sbox_2_M57 ;
    wire SubBytesIns_Inst_Sbox_2_M56 ;
    wire SubBytesIns_Inst_Sbox_2_M55 ;
    wire SubBytesIns_Inst_Sbox_2_M54 ;
    wire SubBytesIns_Inst_Sbox_2_M53 ;
    wire SubBytesIns_Inst_Sbox_2_M52 ;
    wire SubBytesIns_Inst_Sbox_2_M51 ;
    wire SubBytesIns_Inst_Sbox_2_M50 ;
    wire SubBytesIns_Inst_Sbox_2_M49 ;
    wire SubBytesIns_Inst_Sbox_2_M48 ;
    wire SubBytesIns_Inst_Sbox_2_M47 ;
    wire SubBytesIns_Inst_Sbox_2_M46 ;
    wire SubBytesIns_Inst_Sbox_2_M45 ;
    wire SubBytesIns_Inst_Sbox_2_M44 ;
    wire SubBytesIns_Inst_Sbox_2_M43 ;
    wire SubBytesIns_Inst_Sbox_2_M42 ;
    wire SubBytesIns_Inst_Sbox_2_M41 ;
    wire SubBytesIns_Inst_Sbox_2_M40 ;
    wire SubBytesIns_Inst_Sbox_2_M39 ;
    wire SubBytesIns_Inst_Sbox_2_M38 ;
    wire SubBytesIns_Inst_Sbox_2_M37 ;
    wire SubBytesIns_Inst_Sbox_2_M36 ;
    wire SubBytesIns_Inst_Sbox_2_M35 ;
    wire SubBytesIns_Inst_Sbox_2_M34 ;
    wire SubBytesIns_Inst_Sbox_2_M33 ;
    wire SubBytesIns_Inst_Sbox_2_M32 ;
    wire SubBytesIns_Inst_Sbox_2_M31 ;
    wire SubBytesIns_Inst_Sbox_2_M30 ;
    wire SubBytesIns_Inst_Sbox_2_M29 ;
    wire SubBytesIns_Inst_Sbox_2_M28 ;
    wire SubBytesIns_Inst_Sbox_2_M27 ;
    wire SubBytesIns_Inst_Sbox_2_M26 ;
    wire SubBytesIns_Inst_Sbox_2_M25 ;
    wire SubBytesIns_Inst_Sbox_2_M24 ;
    wire SubBytesIns_Inst_Sbox_2_M23 ;
    wire SubBytesIns_Inst_Sbox_2_M22 ;
    wire SubBytesIns_Inst_Sbox_2_M21 ;
    wire SubBytesIns_Inst_Sbox_2_M20 ;
    wire SubBytesIns_Inst_Sbox_2_M19 ;
    wire SubBytesIns_Inst_Sbox_2_M18 ;
    wire SubBytesIns_Inst_Sbox_2_M17 ;
    wire SubBytesIns_Inst_Sbox_2_M16 ;
    wire SubBytesIns_Inst_Sbox_2_M15 ;
    wire SubBytesIns_Inst_Sbox_2_M14 ;
    wire SubBytesIns_Inst_Sbox_2_M13 ;
    wire SubBytesIns_Inst_Sbox_2_M12 ;
    wire SubBytesIns_Inst_Sbox_2_M11 ;
    wire SubBytesIns_Inst_Sbox_2_M10 ;
    wire SubBytesIns_Inst_Sbox_2_M9 ;
    wire SubBytesIns_Inst_Sbox_2_M8 ;
    wire SubBytesIns_Inst_Sbox_2_M7 ;
    wire SubBytesIns_Inst_Sbox_2_M6 ;
    wire SubBytesIns_Inst_Sbox_2_M5 ;
    wire SubBytesIns_Inst_Sbox_2_M4 ;
    wire SubBytesIns_Inst_Sbox_2_M3 ;
    wire SubBytesIns_Inst_Sbox_2_M2 ;
    wire SubBytesIns_Inst_Sbox_2_M1 ;
    wire SubBytesIns_Inst_Sbox_2_T27 ;
    wire SubBytesIns_Inst_Sbox_2_T26 ;
    wire SubBytesIns_Inst_Sbox_2_T25 ;
    wire SubBytesIns_Inst_Sbox_2_T24 ;
    wire SubBytesIns_Inst_Sbox_2_T23 ;
    wire SubBytesIns_Inst_Sbox_2_T22 ;
    wire SubBytesIns_Inst_Sbox_2_T21 ;
    wire SubBytesIns_Inst_Sbox_2_T20 ;
    wire SubBytesIns_Inst_Sbox_2_T19 ;
    wire SubBytesIns_Inst_Sbox_2_T18 ;
    wire SubBytesIns_Inst_Sbox_2_T17 ;
    wire SubBytesIns_Inst_Sbox_2_T16 ;
    wire SubBytesIns_Inst_Sbox_2_T15 ;
    wire SubBytesIns_Inst_Sbox_2_T14 ;
    wire SubBytesIns_Inst_Sbox_2_T13 ;
    wire SubBytesIns_Inst_Sbox_2_T12 ;
    wire SubBytesIns_Inst_Sbox_2_T11 ;
    wire SubBytesIns_Inst_Sbox_2_T10 ;
    wire SubBytesIns_Inst_Sbox_2_T9 ;
    wire SubBytesIns_Inst_Sbox_2_T8 ;
    wire SubBytesIns_Inst_Sbox_2_T7 ;
    wire SubBytesIns_Inst_Sbox_2_T6 ;
    wire SubBytesIns_Inst_Sbox_2_T5 ;
    wire SubBytesIns_Inst_Sbox_2_T4 ;
    wire SubBytesIns_Inst_Sbox_2_T3 ;
    wire SubBytesIns_Inst_Sbox_2_T2 ;
    wire SubBytesIns_Inst_Sbox_2_T1 ;
    wire SubBytesIns_Inst_Sbox_3_L29 ;
    wire SubBytesIns_Inst_Sbox_3_L28 ;
    wire SubBytesIns_Inst_Sbox_3_L27 ;
    wire SubBytesIns_Inst_Sbox_3_L26 ;
    wire SubBytesIns_Inst_Sbox_3_L25 ;
    wire SubBytesIns_Inst_Sbox_3_L24 ;
    wire SubBytesIns_Inst_Sbox_3_L23 ;
    wire SubBytesIns_Inst_Sbox_3_L22 ;
    wire SubBytesIns_Inst_Sbox_3_L21 ;
    wire SubBytesIns_Inst_Sbox_3_L20 ;
    wire SubBytesIns_Inst_Sbox_3_L19 ;
    wire SubBytesIns_Inst_Sbox_3_L18 ;
    wire SubBytesIns_Inst_Sbox_3_L17 ;
    wire SubBytesIns_Inst_Sbox_3_L16 ;
    wire SubBytesIns_Inst_Sbox_3_L15 ;
    wire SubBytesIns_Inst_Sbox_3_L14 ;
    wire SubBytesIns_Inst_Sbox_3_L13 ;
    wire SubBytesIns_Inst_Sbox_3_L12 ;
    wire SubBytesIns_Inst_Sbox_3_L11 ;
    wire SubBytesIns_Inst_Sbox_3_L10 ;
    wire SubBytesIns_Inst_Sbox_3_L9 ;
    wire SubBytesIns_Inst_Sbox_3_L8 ;
    wire SubBytesIns_Inst_Sbox_3_L7 ;
    wire SubBytesIns_Inst_Sbox_3_L6 ;
    wire SubBytesIns_Inst_Sbox_3_L5 ;
    wire SubBytesIns_Inst_Sbox_3_L4 ;
    wire SubBytesIns_Inst_Sbox_3_L3 ;
    wire SubBytesIns_Inst_Sbox_3_L2 ;
    wire SubBytesIns_Inst_Sbox_3_L1 ;
    wire SubBytesIns_Inst_Sbox_3_L0 ;
    wire SubBytesIns_Inst_Sbox_3_M63 ;
    wire SubBytesIns_Inst_Sbox_3_M62 ;
    wire SubBytesIns_Inst_Sbox_3_M61 ;
    wire SubBytesIns_Inst_Sbox_3_M60 ;
    wire SubBytesIns_Inst_Sbox_3_M59 ;
    wire SubBytesIns_Inst_Sbox_3_M58 ;
    wire SubBytesIns_Inst_Sbox_3_M57 ;
    wire SubBytesIns_Inst_Sbox_3_M56 ;
    wire SubBytesIns_Inst_Sbox_3_M55 ;
    wire SubBytesIns_Inst_Sbox_3_M54 ;
    wire SubBytesIns_Inst_Sbox_3_M53 ;
    wire SubBytesIns_Inst_Sbox_3_M52 ;
    wire SubBytesIns_Inst_Sbox_3_M51 ;
    wire SubBytesIns_Inst_Sbox_3_M50 ;
    wire SubBytesIns_Inst_Sbox_3_M49 ;
    wire SubBytesIns_Inst_Sbox_3_M48 ;
    wire SubBytesIns_Inst_Sbox_3_M47 ;
    wire SubBytesIns_Inst_Sbox_3_M46 ;
    wire SubBytesIns_Inst_Sbox_3_M45 ;
    wire SubBytesIns_Inst_Sbox_3_M44 ;
    wire SubBytesIns_Inst_Sbox_3_M43 ;
    wire SubBytesIns_Inst_Sbox_3_M42 ;
    wire SubBytesIns_Inst_Sbox_3_M41 ;
    wire SubBytesIns_Inst_Sbox_3_M40 ;
    wire SubBytesIns_Inst_Sbox_3_M39 ;
    wire SubBytesIns_Inst_Sbox_3_M38 ;
    wire SubBytesIns_Inst_Sbox_3_M37 ;
    wire SubBytesIns_Inst_Sbox_3_M36 ;
    wire SubBytesIns_Inst_Sbox_3_M35 ;
    wire SubBytesIns_Inst_Sbox_3_M34 ;
    wire SubBytesIns_Inst_Sbox_3_M33 ;
    wire SubBytesIns_Inst_Sbox_3_M32 ;
    wire SubBytesIns_Inst_Sbox_3_M31 ;
    wire SubBytesIns_Inst_Sbox_3_M30 ;
    wire SubBytesIns_Inst_Sbox_3_M29 ;
    wire SubBytesIns_Inst_Sbox_3_M28 ;
    wire SubBytesIns_Inst_Sbox_3_M27 ;
    wire SubBytesIns_Inst_Sbox_3_M26 ;
    wire SubBytesIns_Inst_Sbox_3_M25 ;
    wire SubBytesIns_Inst_Sbox_3_M24 ;
    wire SubBytesIns_Inst_Sbox_3_M23 ;
    wire SubBytesIns_Inst_Sbox_3_M22 ;
    wire SubBytesIns_Inst_Sbox_3_M21 ;
    wire SubBytesIns_Inst_Sbox_3_M20 ;
    wire SubBytesIns_Inst_Sbox_3_M19 ;
    wire SubBytesIns_Inst_Sbox_3_M18 ;
    wire SubBytesIns_Inst_Sbox_3_M17 ;
    wire SubBytesIns_Inst_Sbox_3_M16 ;
    wire SubBytesIns_Inst_Sbox_3_M15 ;
    wire SubBytesIns_Inst_Sbox_3_M14 ;
    wire SubBytesIns_Inst_Sbox_3_M13 ;
    wire SubBytesIns_Inst_Sbox_3_M12 ;
    wire SubBytesIns_Inst_Sbox_3_M11 ;
    wire SubBytesIns_Inst_Sbox_3_M10 ;
    wire SubBytesIns_Inst_Sbox_3_M9 ;
    wire SubBytesIns_Inst_Sbox_3_M8 ;
    wire SubBytesIns_Inst_Sbox_3_M7 ;
    wire SubBytesIns_Inst_Sbox_3_M6 ;
    wire SubBytesIns_Inst_Sbox_3_M5 ;
    wire SubBytesIns_Inst_Sbox_3_M4 ;
    wire SubBytesIns_Inst_Sbox_3_M3 ;
    wire SubBytesIns_Inst_Sbox_3_M2 ;
    wire SubBytesIns_Inst_Sbox_3_M1 ;
    wire SubBytesIns_Inst_Sbox_3_T27 ;
    wire SubBytesIns_Inst_Sbox_3_T26 ;
    wire SubBytesIns_Inst_Sbox_3_T25 ;
    wire SubBytesIns_Inst_Sbox_3_T24 ;
    wire SubBytesIns_Inst_Sbox_3_T23 ;
    wire SubBytesIns_Inst_Sbox_3_T22 ;
    wire SubBytesIns_Inst_Sbox_3_T21 ;
    wire SubBytesIns_Inst_Sbox_3_T20 ;
    wire SubBytesIns_Inst_Sbox_3_T19 ;
    wire SubBytesIns_Inst_Sbox_3_T18 ;
    wire SubBytesIns_Inst_Sbox_3_T17 ;
    wire SubBytesIns_Inst_Sbox_3_T16 ;
    wire SubBytesIns_Inst_Sbox_3_T15 ;
    wire SubBytesIns_Inst_Sbox_3_T14 ;
    wire SubBytesIns_Inst_Sbox_3_T13 ;
    wire SubBytesIns_Inst_Sbox_3_T12 ;
    wire SubBytesIns_Inst_Sbox_3_T11 ;
    wire SubBytesIns_Inst_Sbox_3_T10 ;
    wire SubBytesIns_Inst_Sbox_3_T9 ;
    wire SubBytesIns_Inst_Sbox_3_T8 ;
    wire SubBytesIns_Inst_Sbox_3_T7 ;
    wire SubBytesIns_Inst_Sbox_3_T6 ;
    wire SubBytesIns_Inst_Sbox_3_T5 ;
    wire SubBytesIns_Inst_Sbox_3_T4 ;
    wire SubBytesIns_Inst_Sbox_3_T3 ;
    wire SubBytesIns_Inst_Sbox_3_T2 ;
    wire SubBytesIns_Inst_Sbox_3_T1 ;
    wire SubBytesIns_Inst_Sbox_4_L29 ;
    wire SubBytesIns_Inst_Sbox_4_L28 ;
    wire SubBytesIns_Inst_Sbox_4_L27 ;
    wire SubBytesIns_Inst_Sbox_4_L26 ;
    wire SubBytesIns_Inst_Sbox_4_L25 ;
    wire SubBytesIns_Inst_Sbox_4_L24 ;
    wire SubBytesIns_Inst_Sbox_4_L23 ;
    wire SubBytesIns_Inst_Sbox_4_L22 ;
    wire SubBytesIns_Inst_Sbox_4_L21 ;
    wire SubBytesIns_Inst_Sbox_4_L20 ;
    wire SubBytesIns_Inst_Sbox_4_L19 ;
    wire SubBytesIns_Inst_Sbox_4_L18 ;
    wire SubBytesIns_Inst_Sbox_4_L17 ;
    wire SubBytesIns_Inst_Sbox_4_L16 ;
    wire SubBytesIns_Inst_Sbox_4_L15 ;
    wire SubBytesIns_Inst_Sbox_4_L14 ;
    wire SubBytesIns_Inst_Sbox_4_L13 ;
    wire SubBytesIns_Inst_Sbox_4_L12 ;
    wire SubBytesIns_Inst_Sbox_4_L11 ;
    wire SubBytesIns_Inst_Sbox_4_L10 ;
    wire SubBytesIns_Inst_Sbox_4_L9 ;
    wire SubBytesIns_Inst_Sbox_4_L8 ;
    wire SubBytesIns_Inst_Sbox_4_L7 ;
    wire SubBytesIns_Inst_Sbox_4_L6 ;
    wire SubBytesIns_Inst_Sbox_4_L5 ;
    wire SubBytesIns_Inst_Sbox_4_L4 ;
    wire SubBytesIns_Inst_Sbox_4_L3 ;
    wire SubBytesIns_Inst_Sbox_4_L2 ;
    wire SubBytesIns_Inst_Sbox_4_L1 ;
    wire SubBytesIns_Inst_Sbox_4_L0 ;
    wire SubBytesIns_Inst_Sbox_4_M63 ;
    wire SubBytesIns_Inst_Sbox_4_M62 ;
    wire SubBytesIns_Inst_Sbox_4_M61 ;
    wire SubBytesIns_Inst_Sbox_4_M60 ;
    wire SubBytesIns_Inst_Sbox_4_M59 ;
    wire SubBytesIns_Inst_Sbox_4_M58 ;
    wire SubBytesIns_Inst_Sbox_4_M57 ;
    wire SubBytesIns_Inst_Sbox_4_M56 ;
    wire SubBytesIns_Inst_Sbox_4_M55 ;
    wire SubBytesIns_Inst_Sbox_4_M54 ;
    wire SubBytesIns_Inst_Sbox_4_M53 ;
    wire SubBytesIns_Inst_Sbox_4_M52 ;
    wire SubBytesIns_Inst_Sbox_4_M51 ;
    wire SubBytesIns_Inst_Sbox_4_M50 ;
    wire SubBytesIns_Inst_Sbox_4_M49 ;
    wire SubBytesIns_Inst_Sbox_4_M48 ;
    wire SubBytesIns_Inst_Sbox_4_M47 ;
    wire SubBytesIns_Inst_Sbox_4_M46 ;
    wire SubBytesIns_Inst_Sbox_4_M45 ;
    wire SubBytesIns_Inst_Sbox_4_M44 ;
    wire SubBytesIns_Inst_Sbox_4_M43 ;
    wire SubBytesIns_Inst_Sbox_4_M42 ;
    wire SubBytesIns_Inst_Sbox_4_M41 ;
    wire SubBytesIns_Inst_Sbox_4_M40 ;
    wire SubBytesIns_Inst_Sbox_4_M39 ;
    wire SubBytesIns_Inst_Sbox_4_M38 ;
    wire SubBytesIns_Inst_Sbox_4_M37 ;
    wire SubBytesIns_Inst_Sbox_4_M36 ;
    wire SubBytesIns_Inst_Sbox_4_M35 ;
    wire SubBytesIns_Inst_Sbox_4_M34 ;
    wire SubBytesIns_Inst_Sbox_4_M33 ;
    wire SubBytesIns_Inst_Sbox_4_M32 ;
    wire SubBytesIns_Inst_Sbox_4_M31 ;
    wire SubBytesIns_Inst_Sbox_4_M30 ;
    wire SubBytesIns_Inst_Sbox_4_M29 ;
    wire SubBytesIns_Inst_Sbox_4_M28 ;
    wire SubBytesIns_Inst_Sbox_4_M27 ;
    wire SubBytesIns_Inst_Sbox_4_M26 ;
    wire SubBytesIns_Inst_Sbox_4_M25 ;
    wire SubBytesIns_Inst_Sbox_4_M24 ;
    wire SubBytesIns_Inst_Sbox_4_M23 ;
    wire SubBytesIns_Inst_Sbox_4_M22 ;
    wire SubBytesIns_Inst_Sbox_4_M21 ;
    wire SubBytesIns_Inst_Sbox_4_M20 ;
    wire SubBytesIns_Inst_Sbox_4_M19 ;
    wire SubBytesIns_Inst_Sbox_4_M18 ;
    wire SubBytesIns_Inst_Sbox_4_M17 ;
    wire SubBytesIns_Inst_Sbox_4_M16 ;
    wire SubBytesIns_Inst_Sbox_4_M15 ;
    wire SubBytesIns_Inst_Sbox_4_M14 ;
    wire SubBytesIns_Inst_Sbox_4_M13 ;
    wire SubBytesIns_Inst_Sbox_4_M12 ;
    wire SubBytesIns_Inst_Sbox_4_M11 ;
    wire SubBytesIns_Inst_Sbox_4_M10 ;
    wire SubBytesIns_Inst_Sbox_4_M9 ;
    wire SubBytesIns_Inst_Sbox_4_M8 ;
    wire SubBytesIns_Inst_Sbox_4_M7 ;
    wire SubBytesIns_Inst_Sbox_4_M6 ;
    wire SubBytesIns_Inst_Sbox_4_M5 ;
    wire SubBytesIns_Inst_Sbox_4_M4 ;
    wire SubBytesIns_Inst_Sbox_4_M3 ;
    wire SubBytesIns_Inst_Sbox_4_M2 ;
    wire SubBytesIns_Inst_Sbox_4_M1 ;
    wire SubBytesIns_Inst_Sbox_4_T27 ;
    wire SubBytesIns_Inst_Sbox_4_T26 ;
    wire SubBytesIns_Inst_Sbox_4_T25 ;
    wire SubBytesIns_Inst_Sbox_4_T24 ;
    wire SubBytesIns_Inst_Sbox_4_T23 ;
    wire SubBytesIns_Inst_Sbox_4_T22 ;
    wire SubBytesIns_Inst_Sbox_4_T21 ;
    wire SubBytesIns_Inst_Sbox_4_T20 ;
    wire SubBytesIns_Inst_Sbox_4_T19 ;
    wire SubBytesIns_Inst_Sbox_4_T18 ;
    wire SubBytesIns_Inst_Sbox_4_T17 ;
    wire SubBytesIns_Inst_Sbox_4_T16 ;
    wire SubBytesIns_Inst_Sbox_4_T15 ;
    wire SubBytesIns_Inst_Sbox_4_T14 ;
    wire SubBytesIns_Inst_Sbox_4_T13 ;
    wire SubBytesIns_Inst_Sbox_4_T12 ;
    wire SubBytesIns_Inst_Sbox_4_T11 ;
    wire SubBytesIns_Inst_Sbox_4_T10 ;
    wire SubBytesIns_Inst_Sbox_4_T9 ;
    wire SubBytesIns_Inst_Sbox_4_T8 ;
    wire SubBytesIns_Inst_Sbox_4_T7 ;
    wire SubBytesIns_Inst_Sbox_4_T6 ;
    wire SubBytesIns_Inst_Sbox_4_T5 ;
    wire SubBytesIns_Inst_Sbox_4_T4 ;
    wire SubBytesIns_Inst_Sbox_4_T3 ;
    wire SubBytesIns_Inst_Sbox_4_T2 ;
    wire SubBytesIns_Inst_Sbox_4_T1 ;
    wire SubBytesIns_Inst_Sbox_5_L29 ;
    wire SubBytesIns_Inst_Sbox_5_L28 ;
    wire SubBytesIns_Inst_Sbox_5_L27 ;
    wire SubBytesIns_Inst_Sbox_5_L26 ;
    wire SubBytesIns_Inst_Sbox_5_L25 ;
    wire SubBytesIns_Inst_Sbox_5_L24 ;
    wire SubBytesIns_Inst_Sbox_5_L23 ;
    wire SubBytesIns_Inst_Sbox_5_L22 ;
    wire SubBytesIns_Inst_Sbox_5_L21 ;
    wire SubBytesIns_Inst_Sbox_5_L20 ;
    wire SubBytesIns_Inst_Sbox_5_L19 ;
    wire SubBytesIns_Inst_Sbox_5_L18 ;
    wire SubBytesIns_Inst_Sbox_5_L17 ;
    wire SubBytesIns_Inst_Sbox_5_L16 ;
    wire SubBytesIns_Inst_Sbox_5_L15 ;
    wire SubBytesIns_Inst_Sbox_5_L14 ;
    wire SubBytesIns_Inst_Sbox_5_L13 ;
    wire SubBytesIns_Inst_Sbox_5_L12 ;
    wire SubBytesIns_Inst_Sbox_5_L11 ;
    wire SubBytesIns_Inst_Sbox_5_L10 ;
    wire SubBytesIns_Inst_Sbox_5_L9 ;
    wire SubBytesIns_Inst_Sbox_5_L8 ;
    wire SubBytesIns_Inst_Sbox_5_L7 ;
    wire SubBytesIns_Inst_Sbox_5_L6 ;
    wire SubBytesIns_Inst_Sbox_5_L5 ;
    wire SubBytesIns_Inst_Sbox_5_L4 ;
    wire SubBytesIns_Inst_Sbox_5_L3 ;
    wire SubBytesIns_Inst_Sbox_5_L2 ;
    wire SubBytesIns_Inst_Sbox_5_L1 ;
    wire SubBytesIns_Inst_Sbox_5_L0 ;
    wire SubBytesIns_Inst_Sbox_5_M63 ;
    wire SubBytesIns_Inst_Sbox_5_M62 ;
    wire SubBytesIns_Inst_Sbox_5_M61 ;
    wire SubBytesIns_Inst_Sbox_5_M60 ;
    wire SubBytesIns_Inst_Sbox_5_M59 ;
    wire SubBytesIns_Inst_Sbox_5_M58 ;
    wire SubBytesIns_Inst_Sbox_5_M57 ;
    wire SubBytesIns_Inst_Sbox_5_M56 ;
    wire SubBytesIns_Inst_Sbox_5_M55 ;
    wire SubBytesIns_Inst_Sbox_5_M54 ;
    wire SubBytesIns_Inst_Sbox_5_M53 ;
    wire SubBytesIns_Inst_Sbox_5_M52 ;
    wire SubBytesIns_Inst_Sbox_5_M51 ;
    wire SubBytesIns_Inst_Sbox_5_M50 ;
    wire SubBytesIns_Inst_Sbox_5_M49 ;
    wire SubBytesIns_Inst_Sbox_5_M48 ;
    wire SubBytesIns_Inst_Sbox_5_M47 ;
    wire SubBytesIns_Inst_Sbox_5_M46 ;
    wire SubBytesIns_Inst_Sbox_5_M45 ;
    wire SubBytesIns_Inst_Sbox_5_M44 ;
    wire SubBytesIns_Inst_Sbox_5_M43 ;
    wire SubBytesIns_Inst_Sbox_5_M42 ;
    wire SubBytesIns_Inst_Sbox_5_M41 ;
    wire SubBytesIns_Inst_Sbox_5_M40 ;
    wire SubBytesIns_Inst_Sbox_5_M39 ;
    wire SubBytesIns_Inst_Sbox_5_M38 ;
    wire SubBytesIns_Inst_Sbox_5_M37 ;
    wire SubBytesIns_Inst_Sbox_5_M36 ;
    wire SubBytesIns_Inst_Sbox_5_M35 ;
    wire SubBytesIns_Inst_Sbox_5_M34 ;
    wire SubBytesIns_Inst_Sbox_5_M33 ;
    wire SubBytesIns_Inst_Sbox_5_M32 ;
    wire SubBytesIns_Inst_Sbox_5_M31 ;
    wire SubBytesIns_Inst_Sbox_5_M30 ;
    wire SubBytesIns_Inst_Sbox_5_M29 ;
    wire SubBytesIns_Inst_Sbox_5_M28 ;
    wire SubBytesIns_Inst_Sbox_5_M27 ;
    wire SubBytesIns_Inst_Sbox_5_M26 ;
    wire SubBytesIns_Inst_Sbox_5_M25 ;
    wire SubBytesIns_Inst_Sbox_5_M24 ;
    wire SubBytesIns_Inst_Sbox_5_M23 ;
    wire SubBytesIns_Inst_Sbox_5_M22 ;
    wire SubBytesIns_Inst_Sbox_5_M21 ;
    wire SubBytesIns_Inst_Sbox_5_M20 ;
    wire SubBytesIns_Inst_Sbox_5_M19 ;
    wire SubBytesIns_Inst_Sbox_5_M18 ;
    wire SubBytesIns_Inst_Sbox_5_M17 ;
    wire SubBytesIns_Inst_Sbox_5_M16 ;
    wire SubBytesIns_Inst_Sbox_5_M15 ;
    wire SubBytesIns_Inst_Sbox_5_M14 ;
    wire SubBytesIns_Inst_Sbox_5_M13 ;
    wire SubBytesIns_Inst_Sbox_5_M12 ;
    wire SubBytesIns_Inst_Sbox_5_M11 ;
    wire SubBytesIns_Inst_Sbox_5_M10 ;
    wire SubBytesIns_Inst_Sbox_5_M9 ;
    wire SubBytesIns_Inst_Sbox_5_M8 ;
    wire SubBytesIns_Inst_Sbox_5_M7 ;
    wire SubBytesIns_Inst_Sbox_5_M6 ;
    wire SubBytesIns_Inst_Sbox_5_M5 ;
    wire SubBytesIns_Inst_Sbox_5_M4 ;
    wire SubBytesIns_Inst_Sbox_5_M3 ;
    wire SubBytesIns_Inst_Sbox_5_M2 ;
    wire SubBytesIns_Inst_Sbox_5_M1 ;
    wire SubBytesIns_Inst_Sbox_5_T27 ;
    wire SubBytesIns_Inst_Sbox_5_T26 ;
    wire SubBytesIns_Inst_Sbox_5_T25 ;
    wire SubBytesIns_Inst_Sbox_5_T24 ;
    wire SubBytesIns_Inst_Sbox_5_T23 ;
    wire SubBytesIns_Inst_Sbox_5_T22 ;
    wire SubBytesIns_Inst_Sbox_5_T21 ;
    wire SubBytesIns_Inst_Sbox_5_T20 ;
    wire SubBytesIns_Inst_Sbox_5_T19 ;
    wire SubBytesIns_Inst_Sbox_5_T18 ;
    wire SubBytesIns_Inst_Sbox_5_T17 ;
    wire SubBytesIns_Inst_Sbox_5_T16 ;
    wire SubBytesIns_Inst_Sbox_5_T15 ;
    wire SubBytesIns_Inst_Sbox_5_T14 ;
    wire SubBytesIns_Inst_Sbox_5_T13 ;
    wire SubBytesIns_Inst_Sbox_5_T12 ;
    wire SubBytesIns_Inst_Sbox_5_T11 ;
    wire SubBytesIns_Inst_Sbox_5_T10 ;
    wire SubBytesIns_Inst_Sbox_5_T9 ;
    wire SubBytesIns_Inst_Sbox_5_T8 ;
    wire SubBytesIns_Inst_Sbox_5_T7 ;
    wire SubBytesIns_Inst_Sbox_5_T6 ;
    wire SubBytesIns_Inst_Sbox_5_T5 ;
    wire SubBytesIns_Inst_Sbox_5_T4 ;
    wire SubBytesIns_Inst_Sbox_5_T3 ;
    wire SubBytesIns_Inst_Sbox_5_T2 ;
    wire SubBytesIns_Inst_Sbox_5_T1 ;
    wire SubBytesIns_Inst_Sbox_6_L29 ;
    wire SubBytesIns_Inst_Sbox_6_L28 ;
    wire SubBytesIns_Inst_Sbox_6_L27 ;
    wire SubBytesIns_Inst_Sbox_6_L26 ;
    wire SubBytesIns_Inst_Sbox_6_L25 ;
    wire SubBytesIns_Inst_Sbox_6_L24 ;
    wire SubBytesIns_Inst_Sbox_6_L23 ;
    wire SubBytesIns_Inst_Sbox_6_L22 ;
    wire SubBytesIns_Inst_Sbox_6_L21 ;
    wire SubBytesIns_Inst_Sbox_6_L20 ;
    wire SubBytesIns_Inst_Sbox_6_L19 ;
    wire SubBytesIns_Inst_Sbox_6_L18 ;
    wire SubBytesIns_Inst_Sbox_6_L17 ;
    wire SubBytesIns_Inst_Sbox_6_L16 ;
    wire SubBytesIns_Inst_Sbox_6_L15 ;
    wire SubBytesIns_Inst_Sbox_6_L14 ;
    wire SubBytesIns_Inst_Sbox_6_L13 ;
    wire SubBytesIns_Inst_Sbox_6_L12 ;
    wire SubBytesIns_Inst_Sbox_6_L11 ;
    wire SubBytesIns_Inst_Sbox_6_L10 ;
    wire SubBytesIns_Inst_Sbox_6_L9 ;
    wire SubBytesIns_Inst_Sbox_6_L8 ;
    wire SubBytesIns_Inst_Sbox_6_L7 ;
    wire SubBytesIns_Inst_Sbox_6_L6 ;
    wire SubBytesIns_Inst_Sbox_6_L5 ;
    wire SubBytesIns_Inst_Sbox_6_L4 ;
    wire SubBytesIns_Inst_Sbox_6_L3 ;
    wire SubBytesIns_Inst_Sbox_6_L2 ;
    wire SubBytesIns_Inst_Sbox_6_L1 ;
    wire SubBytesIns_Inst_Sbox_6_L0 ;
    wire SubBytesIns_Inst_Sbox_6_M63 ;
    wire SubBytesIns_Inst_Sbox_6_M62 ;
    wire SubBytesIns_Inst_Sbox_6_M61 ;
    wire SubBytesIns_Inst_Sbox_6_M60 ;
    wire SubBytesIns_Inst_Sbox_6_M59 ;
    wire SubBytesIns_Inst_Sbox_6_M58 ;
    wire SubBytesIns_Inst_Sbox_6_M57 ;
    wire SubBytesIns_Inst_Sbox_6_M56 ;
    wire SubBytesIns_Inst_Sbox_6_M55 ;
    wire SubBytesIns_Inst_Sbox_6_M54 ;
    wire SubBytesIns_Inst_Sbox_6_M53 ;
    wire SubBytesIns_Inst_Sbox_6_M52 ;
    wire SubBytesIns_Inst_Sbox_6_M51 ;
    wire SubBytesIns_Inst_Sbox_6_M50 ;
    wire SubBytesIns_Inst_Sbox_6_M49 ;
    wire SubBytesIns_Inst_Sbox_6_M48 ;
    wire SubBytesIns_Inst_Sbox_6_M47 ;
    wire SubBytesIns_Inst_Sbox_6_M46 ;
    wire SubBytesIns_Inst_Sbox_6_M45 ;
    wire SubBytesIns_Inst_Sbox_6_M44 ;
    wire SubBytesIns_Inst_Sbox_6_M43 ;
    wire SubBytesIns_Inst_Sbox_6_M42 ;
    wire SubBytesIns_Inst_Sbox_6_M41 ;
    wire SubBytesIns_Inst_Sbox_6_M40 ;
    wire SubBytesIns_Inst_Sbox_6_M39 ;
    wire SubBytesIns_Inst_Sbox_6_M38 ;
    wire SubBytesIns_Inst_Sbox_6_M37 ;
    wire SubBytesIns_Inst_Sbox_6_M36 ;
    wire SubBytesIns_Inst_Sbox_6_M35 ;
    wire SubBytesIns_Inst_Sbox_6_M34 ;
    wire SubBytesIns_Inst_Sbox_6_M33 ;
    wire SubBytesIns_Inst_Sbox_6_M32 ;
    wire SubBytesIns_Inst_Sbox_6_M31 ;
    wire SubBytesIns_Inst_Sbox_6_M30 ;
    wire SubBytesIns_Inst_Sbox_6_M29 ;
    wire SubBytesIns_Inst_Sbox_6_M28 ;
    wire SubBytesIns_Inst_Sbox_6_M27 ;
    wire SubBytesIns_Inst_Sbox_6_M26 ;
    wire SubBytesIns_Inst_Sbox_6_M25 ;
    wire SubBytesIns_Inst_Sbox_6_M24 ;
    wire SubBytesIns_Inst_Sbox_6_M23 ;
    wire SubBytesIns_Inst_Sbox_6_M22 ;
    wire SubBytesIns_Inst_Sbox_6_M21 ;
    wire SubBytesIns_Inst_Sbox_6_M20 ;
    wire SubBytesIns_Inst_Sbox_6_M19 ;
    wire SubBytesIns_Inst_Sbox_6_M18 ;
    wire SubBytesIns_Inst_Sbox_6_M17 ;
    wire SubBytesIns_Inst_Sbox_6_M16 ;
    wire SubBytesIns_Inst_Sbox_6_M15 ;
    wire SubBytesIns_Inst_Sbox_6_M14 ;
    wire SubBytesIns_Inst_Sbox_6_M13 ;
    wire SubBytesIns_Inst_Sbox_6_M12 ;
    wire SubBytesIns_Inst_Sbox_6_M11 ;
    wire SubBytesIns_Inst_Sbox_6_M10 ;
    wire SubBytesIns_Inst_Sbox_6_M9 ;
    wire SubBytesIns_Inst_Sbox_6_M8 ;
    wire SubBytesIns_Inst_Sbox_6_M7 ;
    wire SubBytesIns_Inst_Sbox_6_M6 ;
    wire SubBytesIns_Inst_Sbox_6_M5 ;
    wire SubBytesIns_Inst_Sbox_6_M4 ;
    wire SubBytesIns_Inst_Sbox_6_M3 ;
    wire SubBytesIns_Inst_Sbox_6_M2 ;
    wire SubBytesIns_Inst_Sbox_6_M1 ;
    wire SubBytesIns_Inst_Sbox_6_T27 ;
    wire SubBytesIns_Inst_Sbox_6_T26 ;
    wire SubBytesIns_Inst_Sbox_6_T25 ;
    wire SubBytesIns_Inst_Sbox_6_T24 ;
    wire SubBytesIns_Inst_Sbox_6_T23 ;
    wire SubBytesIns_Inst_Sbox_6_T22 ;
    wire SubBytesIns_Inst_Sbox_6_T21 ;
    wire SubBytesIns_Inst_Sbox_6_T20 ;
    wire SubBytesIns_Inst_Sbox_6_T19 ;
    wire SubBytesIns_Inst_Sbox_6_T18 ;
    wire SubBytesIns_Inst_Sbox_6_T17 ;
    wire SubBytesIns_Inst_Sbox_6_T16 ;
    wire SubBytesIns_Inst_Sbox_6_T15 ;
    wire SubBytesIns_Inst_Sbox_6_T14 ;
    wire SubBytesIns_Inst_Sbox_6_T13 ;
    wire SubBytesIns_Inst_Sbox_6_T12 ;
    wire SubBytesIns_Inst_Sbox_6_T11 ;
    wire SubBytesIns_Inst_Sbox_6_T10 ;
    wire SubBytesIns_Inst_Sbox_6_T9 ;
    wire SubBytesIns_Inst_Sbox_6_T8 ;
    wire SubBytesIns_Inst_Sbox_6_T7 ;
    wire SubBytesIns_Inst_Sbox_6_T6 ;
    wire SubBytesIns_Inst_Sbox_6_T5 ;
    wire SubBytesIns_Inst_Sbox_6_T4 ;
    wire SubBytesIns_Inst_Sbox_6_T3 ;
    wire SubBytesIns_Inst_Sbox_6_T2 ;
    wire SubBytesIns_Inst_Sbox_6_T1 ;
    wire SubBytesIns_Inst_Sbox_7_L29 ;
    wire SubBytesIns_Inst_Sbox_7_L28 ;
    wire SubBytesIns_Inst_Sbox_7_L27 ;
    wire SubBytesIns_Inst_Sbox_7_L26 ;
    wire SubBytesIns_Inst_Sbox_7_L25 ;
    wire SubBytesIns_Inst_Sbox_7_L24 ;
    wire SubBytesIns_Inst_Sbox_7_L23 ;
    wire SubBytesIns_Inst_Sbox_7_L22 ;
    wire SubBytesIns_Inst_Sbox_7_L21 ;
    wire SubBytesIns_Inst_Sbox_7_L20 ;
    wire SubBytesIns_Inst_Sbox_7_L19 ;
    wire SubBytesIns_Inst_Sbox_7_L18 ;
    wire SubBytesIns_Inst_Sbox_7_L17 ;
    wire SubBytesIns_Inst_Sbox_7_L16 ;
    wire SubBytesIns_Inst_Sbox_7_L15 ;
    wire SubBytesIns_Inst_Sbox_7_L14 ;
    wire SubBytesIns_Inst_Sbox_7_L13 ;
    wire SubBytesIns_Inst_Sbox_7_L12 ;
    wire SubBytesIns_Inst_Sbox_7_L11 ;
    wire SubBytesIns_Inst_Sbox_7_L10 ;
    wire SubBytesIns_Inst_Sbox_7_L9 ;
    wire SubBytesIns_Inst_Sbox_7_L8 ;
    wire SubBytesIns_Inst_Sbox_7_L7 ;
    wire SubBytesIns_Inst_Sbox_7_L6 ;
    wire SubBytesIns_Inst_Sbox_7_L5 ;
    wire SubBytesIns_Inst_Sbox_7_L4 ;
    wire SubBytesIns_Inst_Sbox_7_L3 ;
    wire SubBytesIns_Inst_Sbox_7_L2 ;
    wire SubBytesIns_Inst_Sbox_7_L1 ;
    wire SubBytesIns_Inst_Sbox_7_L0 ;
    wire SubBytesIns_Inst_Sbox_7_M63 ;
    wire SubBytesIns_Inst_Sbox_7_M62 ;
    wire SubBytesIns_Inst_Sbox_7_M61 ;
    wire SubBytesIns_Inst_Sbox_7_M60 ;
    wire SubBytesIns_Inst_Sbox_7_M59 ;
    wire SubBytesIns_Inst_Sbox_7_M58 ;
    wire SubBytesIns_Inst_Sbox_7_M57 ;
    wire SubBytesIns_Inst_Sbox_7_M56 ;
    wire SubBytesIns_Inst_Sbox_7_M55 ;
    wire SubBytesIns_Inst_Sbox_7_M54 ;
    wire SubBytesIns_Inst_Sbox_7_M53 ;
    wire SubBytesIns_Inst_Sbox_7_M52 ;
    wire SubBytesIns_Inst_Sbox_7_M51 ;
    wire SubBytesIns_Inst_Sbox_7_M50 ;
    wire SubBytesIns_Inst_Sbox_7_M49 ;
    wire SubBytesIns_Inst_Sbox_7_M48 ;
    wire SubBytesIns_Inst_Sbox_7_M47 ;
    wire SubBytesIns_Inst_Sbox_7_M46 ;
    wire SubBytesIns_Inst_Sbox_7_M45 ;
    wire SubBytesIns_Inst_Sbox_7_M44 ;
    wire SubBytesIns_Inst_Sbox_7_M43 ;
    wire SubBytesIns_Inst_Sbox_7_M42 ;
    wire SubBytesIns_Inst_Sbox_7_M41 ;
    wire SubBytesIns_Inst_Sbox_7_M40 ;
    wire SubBytesIns_Inst_Sbox_7_M39 ;
    wire SubBytesIns_Inst_Sbox_7_M38 ;
    wire SubBytesIns_Inst_Sbox_7_M37 ;
    wire SubBytesIns_Inst_Sbox_7_M36 ;
    wire SubBytesIns_Inst_Sbox_7_M35 ;
    wire SubBytesIns_Inst_Sbox_7_M34 ;
    wire SubBytesIns_Inst_Sbox_7_M33 ;
    wire SubBytesIns_Inst_Sbox_7_M32 ;
    wire SubBytesIns_Inst_Sbox_7_M31 ;
    wire SubBytesIns_Inst_Sbox_7_M30 ;
    wire SubBytesIns_Inst_Sbox_7_M29 ;
    wire SubBytesIns_Inst_Sbox_7_M28 ;
    wire SubBytesIns_Inst_Sbox_7_M27 ;
    wire SubBytesIns_Inst_Sbox_7_M26 ;
    wire SubBytesIns_Inst_Sbox_7_M25 ;
    wire SubBytesIns_Inst_Sbox_7_M24 ;
    wire SubBytesIns_Inst_Sbox_7_M23 ;
    wire SubBytesIns_Inst_Sbox_7_M22 ;
    wire SubBytesIns_Inst_Sbox_7_M21 ;
    wire SubBytesIns_Inst_Sbox_7_M20 ;
    wire SubBytesIns_Inst_Sbox_7_M19 ;
    wire SubBytesIns_Inst_Sbox_7_M18 ;
    wire SubBytesIns_Inst_Sbox_7_M17 ;
    wire SubBytesIns_Inst_Sbox_7_M16 ;
    wire SubBytesIns_Inst_Sbox_7_M15 ;
    wire SubBytesIns_Inst_Sbox_7_M14 ;
    wire SubBytesIns_Inst_Sbox_7_M13 ;
    wire SubBytesIns_Inst_Sbox_7_M12 ;
    wire SubBytesIns_Inst_Sbox_7_M11 ;
    wire SubBytesIns_Inst_Sbox_7_M10 ;
    wire SubBytesIns_Inst_Sbox_7_M9 ;
    wire SubBytesIns_Inst_Sbox_7_M8 ;
    wire SubBytesIns_Inst_Sbox_7_M7 ;
    wire SubBytesIns_Inst_Sbox_7_M6 ;
    wire SubBytesIns_Inst_Sbox_7_M5 ;
    wire SubBytesIns_Inst_Sbox_7_M4 ;
    wire SubBytesIns_Inst_Sbox_7_M3 ;
    wire SubBytesIns_Inst_Sbox_7_M2 ;
    wire SubBytesIns_Inst_Sbox_7_M1 ;
    wire SubBytesIns_Inst_Sbox_7_T27 ;
    wire SubBytesIns_Inst_Sbox_7_T26 ;
    wire SubBytesIns_Inst_Sbox_7_T25 ;
    wire SubBytesIns_Inst_Sbox_7_T24 ;
    wire SubBytesIns_Inst_Sbox_7_T23 ;
    wire SubBytesIns_Inst_Sbox_7_T22 ;
    wire SubBytesIns_Inst_Sbox_7_T21 ;
    wire SubBytesIns_Inst_Sbox_7_T20 ;
    wire SubBytesIns_Inst_Sbox_7_T19 ;
    wire SubBytesIns_Inst_Sbox_7_T18 ;
    wire SubBytesIns_Inst_Sbox_7_T17 ;
    wire SubBytesIns_Inst_Sbox_7_T16 ;
    wire SubBytesIns_Inst_Sbox_7_T15 ;
    wire SubBytesIns_Inst_Sbox_7_T14 ;
    wire SubBytesIns_Inst_Sbox_7_T13 ;
    wire SubBytesIns_Inst_Sbox_7_T12 ;
    wire SubBytesIns_Inst_Sbox_7_T11 ;
    wire SubBytesIns_Inst_Sbox_7_T10 ;
    wire SubBytesIns_Inst_Sbox_7_T9 ;
    wire SubBytesIns_Inst_Sbox_7_T8 ;
    wire SubBytesIns_Inst_Sbox_7_T7 ;
    wire SubBytesIns_Inst_Sbox_7_T6 ;
    wire SubBytesIns_Inst_Sbox_7_T5 ;
    wire SubBytesIns_Inst_Sbox_7_T4 ;
    wire SubBytesIns_Inst_Sbox_7_T3 ;
    wire SubBytesIns_Inst_Sbox_7_T2 ;
    wire SubBytesIns_Inst_Sbox_7_T1 ;
    wire SubBytesIns_Inst_Sbox_8_L29 ;
    wire SubBytesIns_Inst_Sbox_8_L28 ;
    wire SubBytesIns_Inst_Sbox_8_L27 ;
    wire SubBytesIns_Inst_Sbox_8_L26 ;
    wire SubBytesIns_Inst_Sbox_8_L25 ;
    wire SubBytesIns_Inst_Sbox_8_L24 ;
    wire SubBytesIns_Inst_Sbox_8_L23 ;
    wire SubBytesIns_Inst_Sbox_8_L22 ;
    wire SubBytesIns_Inst_Sbox_8_L21 ;
    wire SubBytesIns_Inst_Sbox_8_L20 ;
    wire SubBytesIns_Inst_Sbox_8_L19 ;
    wire SubBytesIns_Inst_Sbox_8_L18 ;
    wire SubBytesIns_Inst_Sbox_8_L17 ;
    wire SubBytesIns_Inst_Sbox_8_L16 ;
    wire SubBytesIns_Inst_Sbox_8_L15 ;
    wire SubBytesIns_Inst_Sbox_8_L14 ;
    wire SubBytesIns_Inst_Sbox_8_L13 ;
    wire SubBytesIns_Inst_Sbox_8_L12 ;
    wire SubBytesIns_Inst_Sbox_8_L11 ;
    wire SubBytesIns_Inst_Sbox_8_L10 ;
    wire SubBytesIns_Inst_Sbox_8_L9 ;
    wire SubBytesIns_Inst_Sbox_8_L8 ;
    wire SubBytesIns_Inst_Sbox_8_L7 ;
    wire SubBytesIns_Inst_Sbox_8_L6 ;
    wire SubBytesIns_Inst_Sbox_8_L5 ;
    wire SubBytesIns_Inst_Sbox_8_L4 ;
    wire SubBytesIns_Inst_Sbox_8_L3 ;
    wire SubBytesIns_Inst_Sbox_8_L2 ;
    wire SubBytesIns_Inst_Sbox_8_L1 ;
    wire SubBytesIns_Inst_Sbox_8_L0 ;
    wire SubBytesIns_Inst_Sbox_8_M63 ;
    wire SubBytesIns_Inst_Sbox_8_M62 ;
    wire SubBytesIns_Inst_Sbox_8_M61 ;
    wire SubBytesIns_Inst_Sbox_8_M60 ;
    wire SubBytesIns_Inst_Sbox_8_M59 ;
    wire SubBytesIns_Inst_Sbox_8_M58 ;
    wire SubBytesIns_Inst_Sbox_8_M57 ;
    wire SubBytesIns_Inst_Sbox_8_M56 ;
    wire SubBytesIns_Inst_Sbox_8_M55 ;
    wire SubBytesIns_Inst_Sbox_8_M54 ;
    wire SubBytesIns_Inst_Sbox_8_M53 ;
    wire SubBytesIns_Inst_Sbox_8_M52 ;
    wire SubBytesIns_Inst_Sbox_8_M51 ;
    wire SubBytesIns_Inst_Sbox_8_M50 ;
    wire SubBytesIns_Inst_Sbox_8_M49 ;
    wire SubBytesIns_Inst_Sbox_8_M48 ;
    wire SubBytesIns_Inst_Sbox_8_M47 ;
    wire SubBytesIns_Inst_Sbox_8_M46 ;
    wire SubBytesIns_Inst_Sbox_8_M45 ;
    wire SubBytesIns_Inst_Sbox_8_M44 ;
    wire SubBytesIns_Inst_Sbox_8_M43 ;
    wire SubBytesIns_Inst_Sbox_8_M42 ;
    wire SubBytesIns_Inst_Sbox_8_M41 ;
    wire SubBytesIns_Inst_Sbox_8_M40 ;
    wire SubBytesIns_Inst_Sbox_8_M39 ;
    wire SubBytesIns_Inst_Sbox_8_M38 ;
    wire SubBytesIns_Inst_Sbox_8_M37 ;
    wire SubBytesIns_Inst_Sbox_8_M36 ;
    wire SubBytesIns_Inst_Sbox_8_M35 ;
    wire SubBytesIns_Inst_Sbox_8_M34 ;
    wire SubBytesIns_Inst_Sbox_8_M33 ;
    wire SubBytesIns_Inst_Sbox_8_M32 ;
    wire SubBytesIns_Inst_Sbox_8_M31 ;
    wire SubBytesIns_Inst_Sbox_8_M30 ;
    wire SubBytesIns_Inst_Sbox_8_M29 ;
    wire SubBytesIns_Inst_Sbox_8_M28 ;
    wire SubBytesIns_Inst_Sbox_8_M27 ;
    wire SubBytesIns_Inst_Sbox_8_M26 ;
    wire SubBytesIns_Inst_Sbox_8_M25 ;
    wire SubBytesIns_Inst_Sbox_8_M24 ;
    wire SubBytesIns_Inst_Sbox_8_M23 ;
    wire SubBytesIns_Inst_Sbox_8_M22 ;
    wire SubBytesIns_Inst_Sbox_8_M21 ;
    wire SubBytesIns_Inst_Sbox_8_M20 ;
    wire SubBytesIns_Inst_Sbox_8_M19 ;
    wire SubBytesIns_Inst_Sbox_8_M18 ;
    wire SubBytesIns_Inst_Sbox_8_M17 ;
    wire SubBytesIns_Inst_Sbox_8_M16 ;
    wire SubBytesIns_Inst_Sbox_8_M15 ;
    wire SubBytesIns_Inst_Sbox_8_M14 ;
    wire SubBytesIns_Inst_Sbox_8_M13 ;
    wire SubBytesIns_Inst_Sbox_8_M12 ;
    wire SubBytesIns_Inst_Sbox_8_M11 ;
    wire SubBytesIns_Inst_Sbox_8_M10 ;
    wire SubBytesIns_Inst_Sbox_8_M9 ;
    wire SubBytesIns_Inst_Sbox_8_M8 ;
    wire SubBytesIns_Inst_Sbox_8_M7 ;
    wire SubBytesIns_Inst_Sbox_8_M6 ;
    wire SubBytesIns_Inst_Sbox_8_M5 ;
    wire SubBytesIns_Inst_Sbox_8_M4 ;
    wire SubBytesIns_Inst_Sbox_8_M3 ;
    wire SubBytesIns_Inst_Sbox_8_M2 ;
    wire SubBytesIns_Inst_Sbox_8_M1 ;
    wire SubBytesIns_Inst_Sbox_8_T27 ;
    wire SubBytesIns_Inst_Sbox_8_T26 ;
    wire SubBytesIns_Inst_Sbox_8_T25 ;
    wire SubBytesIns_Inst_Sbox_8_T24 ;
    wire SubBytesIns_Inst_Sbox_8_T23 ;
    wire SubBytesIns_Inst_Sbox_8_T22 ;
    wire SubBytesIns_Inst_Sbox_8_T21 ;
    wire SubBytesIns_Inst_Sbox_8_T20 ;
    wire SubBytesIns_Inst_Sbox_8_T19 ;
    wire SubBytesIns_Inst_Sbox_8_T18 ;
    wire SubBytesIns_Inst_Sbox_8_T17 ;
    wire SubBytesIns_Inst_Sbox_8_T16 ;
    wire SubBytesIns_Inst_Sbox_8_T15 ;
    wire SubBytesIns_Inst_Sbox_8_T14 ;
    wire SubBytesIns_Inst_Sbox_8_T13 ;
    wire SubBytesIns_Inst_Sbox_8_T12 ;
    wire SubBytesIns_Inst_Sbox_8_T11 ;
    wire SubBytesIns_Inst_Sbox_8_T10 ;
    wire SubBytesIns_Inst_Sbox_8_T9 ;
    wire SubBytesIns_Inst_Sbox_8_T8 ;
    wire SubBytesIns_Inst_Sbox_8_T7 ;
    wire SubBytesIns_Inst_Sbox_8_T6 ;
    wire SubBytesIns_Inst_Sbox_8_T5 ;
    wire SubBytesIns_Inst_Sbox_8_T4 ;
    wire SubBytesIns_Inst_Sbox_8_T3 ;
    wire SubBytesIns_Inst_Sbox_8_T2 ;
    wire SubBytesIns_Inst_Sbox_8_T1 ;
    wire SubBytesIns_Inst_Sbox_9_L29 ;
    wire SubBytesIns_Inst_Sbox_9_L28 ;
    wire SubBytesIns_Inst_Sbox_9_L27 ;
    wire SubBytesIns_Inst_Sbox_9_L26 ;
    wire SubBytesIns_Inst_Sbox_9_L25 ;
    wire SubBytesIns_Inst_Sbox_9_L24 ;
    wire SubBytesIns_Inst_Sbox_9_L23 ;
    wire SubBytesIns_Inst_Sbox_9_L22 ;
    wire SubBytesIns_Inst_Sbox_9_L21 ;
    wire SubBytesIns_Inst_Sbox_9_L20 ;
    wire SubBytesIns_Inst_Sbox_9_L19 ;
    wire SubBytesIns_Inst_Sbox_9_L18 ;
    wire SubBytesIns_Inst_Sbox_9_L17 ;
    wire SubBytesIns_Inst_Sbox_9_L16 ;
    wire SubBytesIns_Inst_Sbox_9_L15 ;
    wire SubBytesIns_Inst_Sbox_9_L14 ;
    wire SubBytesIns_Inst_Sbox_9_L13 ;
    wire SubBytesIns_Inst_Sbox_9_L12 ;
    wire SubBytesIns_Inst_Sbox_9_L11 ;
    wire SubBytesIns_Inst_Sbox_9_L10 ;
    wire SubBytesIns_Inst_Sbox_9_L9 ;
    wire SubBytesIns_Inst_Sbox_9_L8 ;
    wire SubBytesIns_Inst_Sbox_9_L7 ;
    wire SubBytesIns_Inst_Sbox_9_L6 ;
    wire SubBytesIns_Inst_Sbox_9_L5 ;
    wire SubBytesIns_Inst_Sbox_9_L4 ;
    wire SubBytesIns_Inst_Sbox_9_L3 ;
    wire SubBytesIns_Inst_Sbox_9_L2 ;
    wire SubBytesIns_Inst_Sbox_9_L1 ;
    wire SubBytesIns_Inst_Sbox_9_L0 ;
    wire SubBytesIns_Inst_Sbox_9_M63 ;
    wire SubBytesIns_Inst_Sbox_9_M62 ;
    wire SubBytesIns_Inst_Sbox_9_M61 ;
    wire SubBytesIns_Inst_Sbox_9_M60 ;
    wire SubBytesIns_Inst_Sbox_9_M59 ;
    wire SubBytesIns_Inst_Sbox_9_M58 ;
    wire SubBytesIns_Inst_Sbox_9_M57 ;
    wire SubBytesIns_Inst_Sbox_9_M56 ;
    wire SubBytesIns_Inst_Sbox_9_M55 ;
    wire SubBytesIns_Inst_Sbox_9_M54 ;
    wire SubBytesIns_Inst_Sbox_9_M53 ;
    wire SubBytesIns_Inst_Sbox_9_M52 ;
    wire SubBytesIns_Inst_Sbox_9_M51 ;
    wire SubBytesIns_Inst_Sbox_9_M50 ;
    wire SubBytesIns_Inst_Sbox_9_M49 ;
    wire SubBytesIns_Inst_Sbox_9_M48 ;
    wire SubBytesIns_Inst_Sbox_9_M47 ;
    wire SubBytesIns_Inst_Sbox_9_M46 ;
    wire SubBytesIns_Inst_Sbox_9_M45 ;
    wire SubBytesIns_Inst_Sbox_9_M44 ;
    wire SubBytesIns_Inst_Sbox_9_M43 ;
    wire SubBytesIns_Inst_Sbox_9_M42 ;
    wire SubBytesIns_Inst_Sbox_9_M41 ;
    wire SubBytesIns_Inst_Sbox_9_M40 ;
    wire SubBytesIns_Inst_Sbox_9_M39 ;
    wire SubBytesIns_Inst_Sbox_9_M38 ;
    wire SubBytesIns_Inst_Sbox_9_M37 ;
    wire SubBytesIns_Inst_Sbox_9_M36 ;
    wire SubBytesIns_Inst_Sbox_9_M35 ;
    wire SubBytesIns_Inst_Sbox_9_M34 ;
    wire SubBytesIns_Inst_Sbox_9_M33 ;
    wire SubBytesIns_Inst_Sbox_9_M32 ;
    wire SubBytesIns_Inst_Sbox_9_M31 ;
    wire SubBytesIns_Inst_Sbox_9_M30 ;
    wire SubBytesIns_Inst_Sbox_9_M29 ;
    wire SubBytesIns_Inst_Sbox_9_M28 ;
    wire SubBytesIns_Inst_Sbox_9_M27 ;
    wire SubBytesIns_Inst_Sbox_9_M26 ;
    wire SubBytesIns_Inst_Sbox_9_M25 ;
    wire SubBytesIns_Inst_Sbox_9_M24 ;
    wire SubBytesIns_Inst_Sbox_9_M23 ;
    wire SubBytesIns_Inst_Sbox_9_M22 ;
    wire SubBytesIns_Inst_Sbox_9_M21 ;
    wire SubBytesIns_Inst_Sbox_9_M20 ;
    wire SubBytesIns_Inst_Sbox_9_M19 ;
    wire SubBytesIns_Inst_Sbox_9_M18 ;
    wire SubBytesIns_Inst_Sbox_9_M17 ;
    wire SubBytesIns_Inst_Sbox_9_M16 ;
    wire SubBytesIns_Inst_Sbox_9_M15 ;
    wire SubBytesIns_Inst_Sbox_9_M14 ;
    wire SubBytesIns_Inst_Sbox_9_M13 ;
    wire SubBytesIns_Inst_Sbox_9_M12 ;
    wire SubBytesIns_Inst_Sbox_9_M11 ;
    wire SubBytesIns_Inst_Sbox_9_M10 ;
    wire SubBytesIns_Inst_Sbox_9_M9 ;
    wire SubBytesIns_Inst_Sbox_9_M8 ;
    wire SubBytesIns_Inst_Sbox_9_M7 ;
    wire SubBytesIns_Inst_Sbox_9_M6 ;
    wire SubBytesIns_Inst_Sbox_9_M5 ;
    wire SubBytesIns_Inst_Sbox_9_M4 ;
    wire SubBytesIns_Inst_Sbox_9_M3 ;
    wire SubBytesIns_Inst_Sbox_9_M2 ;
    wire SubBytesIns_Inst_Sbox_9_M1 ;
    wire SubBytesIns_Inst_Sbox_9_T27 ;
    wire SubBytesIns_Inst_Sbox_9_T26 ;
    wire SubBytesIns_Inst_Sbox_9_T25 ;
    wire SubBytesIns_Inst_Sbox_9_T24 ;
    wire SubBytesIns_Inst_Sbox_9_T23 ;
    wire SubBytesIns_Inst_Sbox_9_T22 ;
    wire SubBytesIns_Inst_Sbox_9_T21 ;
    wire SubBytesIns_Inst_Sbox_9_T20 ;
    wire SubBytesIns_Inst_Sbox_9_T19 ;
    wire SubBytesIns_Inst_Sbox_9_T18 ;
    wire SubBytesIns_Inst_Sbox_9_T17 ;
    wire SubBytesIns_Inst_Sbox_9_T16 ;
    wire SubBytesIns_Inst_Sbox_9_T15 ;
    wire SubBytesIns_Inst_Sbox_9_T14 ;
    wire SubBytesIns_Inst_Sbox_9_T13 ;
    wire SubBytesIns_Inst_Sbox_9_T12 ;
    wire SubBytesIns_Inst_Sbox_9_T11 ;
    wire SubBytesIns_Inst_Sbox_9_T10 ;
    wire SubBytesIns_Inst_Sbox_9_T9 ;
    wire SubBytesIns_Inst_Sbox_9_T8 ;
    wire SubBytesIns_Inst_Sbox_9_T7 ;
    wire SubBytesIns_Inst_Sbox_9_T6 ;
    wire SubBytesIns_Inst_Sbox_9_T5 ;
    wire SubBytesIns_Inst_Sbox_9_T4 ;
    wire SubBytesIns_Inst_Sbox_9_T3 ;
    wire SubBytesIns_Inst_Sbox_9_T2 ;
    wire SubBytesIns_Inst_Sbox_9_T1 ;
    wire SubBytesIns_Inst_Sbox_10_L29 ;
    wire SubBytesIns_Inst_Sbox_10_L28 ;
    wire SubBytesIns_Inst_Sbox_10_L27 ;
    wire SubBytesIns_Inst_Sbox_10_L26 ;
    wire SubBytesIns_Inst_Sbox_10_L25 ;
    wire SubBytesIns_Inst_Sbox_10_L24 ;
    wire SubBytesIns_Inst_Sbox_10_L23 ;
    wire SubBytesIns_Inst_Sbox_10_L22 ;
    wire SubBytesIns_Inst_Sbox_10_L21 ;
    wire SubBytesIns_Inst_Sbox_10_L20 ;
    wire SubBytesIns_Inst_Sbox_10_L19 ;
    wire SubBytesIns_Inst_Sbox_10_L18 ;
    wire SubBytesIns_Inst_Sbox_10_L17 ;
    wire SubBytesIns_Inst_Sbox_10_L16 ;
    wire SubBytesIns_Inst_Sbox_10_L15 ;
    wire SubBytesIns_Inst_Sbox_10_L14 ;
    wire SubBytesIns_Inst_Sbox_10_L13 ;
    wire SubBytesIns_Inst_Sbox_10_L12 ;
    wire SubBytesIns_Inst_Sbox_10_L11 ;
    wire SubBytesIns_Inst_Sbox_10_L10 ;
    wire SubBytesIns_Inst_Sbox_10_L9 ;
    wire SubBytesIns_Inst_Sbox_10_L8 ;
    wire SubBytesIns_Inst_Sbox_10_L7 ;
    wire SubBytesIns_Inst_Sbox_10_L6 ;
    wire SubBytesIns_Inst_Sbox_10_L5 ;
    wire SubBytesIns_Inst_Sbox_10_L4 ;
    wire SubBytesIns_Inst_Sbox_10_L3 ;
    wire SubBytesIns_Inst_Sbox_10_L2 ;
    wire SubBytesIns_Inst_Sbox_10_L1 ;
    wire SubBytesIns_Inst_Sbox_10_L0 ;
    wire SubBytesIns_Inst_Sbox_10_M63 ;
    wire SubBytesIns_Inst_Sbox_10_M62 ;
    wire SubBytesIns_Inst_Sbox_10_M61 ;
    wire SubBytesIns_Inst_Sbox_10_M60 ;
    wire SubBytesIns_Inst_Sbox_10_M59 ;
    wire SubBytesIns_Inst_Sbox_10_M58 ;
    wire SubBytesIns_Inst_Sbox_10_M57 ;
    wire SubBytesIns_Inst_Sbox_10_M56 ;
    wire SubBytesIns_Inst_Sbox_10_M55 ;
    wire SubBytesIns_Inst_Sbox_10_M54 ;
    wire SubBytesIns_Inst_Sbox_10_M53 ;
    wire SubBytesIns_Inst_Sbox_10_M52 ;
    wire SubBytesIns_Inst_Sbox_10_M51 ;
    wire SubBytesIns_Inst_Sbox_10_M50 ;
    wire SubBytesIns_Inst_Sbox_10_M49 ;
    wire SubBytesIns_Inst_Sbox_10_M48 ;
    wire SubBytesIns_Inst_Sbox_10_M47 ;
    wire SubBytesIns_Inst_Sbox_10_M46 ;
    wire SubBytesIns_Inst_Sbox_10_M45 ;
    wire SubBytesIns_Inst_Sbox_10_M44 ;
    wire SubBytesIns_Inst_Sbox_10_M43 ;
    wire SubBytesIns_Inst_Sbox_10_M42 ;
    wire SubBytesIns_Inst_Sbox_10_M41 ;
    wire SubBytesIns_Inst_Sbox_10_M40 ;
    wire SubBytesIns_Inst_Sbox_10_M39 ;
    wire SubBytesIns_Inst_Sbox_10_M38 ;
    wire SubBytesIns_Inst_Sbox_10_M37 ;
    wire SubBytesIns_Inst_Sbox_10_M36 ;
    wire SubBytesIns_Inst_Sbox_10_M35 ;
    wire SubBytesIns_Inst_Sbox_10_M34 ;
    wire SubBytesIns_Inst_Sbox_10_M33 ;
    wire SubBytesIns_Inst_Sbox_10_M32 ;
    wire SubBytesIns_Inst_Sbox_10_M31 ;
    wire SubBytesIns_Inst_Sbox_10_M30 ;
    wire SubBytesIns_Inst_Sbox_10_M29 ;
    wire SubBytesIns_Inst_Sbox_10_M28 ;
    wire SubBytesIns_Inst_Sbox_10_M27 ;
    wire SubBytesIns_Inst_Sbox_10_M26 ;
    wire SubBytesIns_Inst_Sbox_10_M25 ;
    wire SubBytesIns_Inst_Sbox_10_M24 ;
    wire SubBytesIns_Inst_Sbox_10_M23 ;
    wire SubBytesIns_Inst_Sbox_10_M22 ;
    wire SubBytesIns_Inst_Sbox_10_M21 ;
    wire SubBytesIns_Inst_Sbox_10_M20 ;
    wire SubBytesIns_Inst_Sbox_10_M19 ;
    wire SubBytesIns_Inst_Sbox_10_M18 ;
    wire SubBytesIns_Inst_Sbox_10_M17 ;
    wire SubBytesIns_Inst_Sbox_10_M16 ;
    wire SubBytesIns_Inst_Sbox_10_M15 ;
    wire SubBytesIns_Inst_Sbox_10_M14 ;
    wire SubBytesIns_Inst_Sbox_10_M13 ;
    wire SubBytesIns_Inst_Sbox_10_M12 ;
    wire SubBytesIns_Inst_Sbox_10_M11 ;
    wire SubBytesIns_Inst_Sbox_10_M10 ;
    wire SubBytesIns_Inst_Sbox_10_M9 ;
    wire SubBytesIns_Inst_Sbox_10_M8 ;
    wire SubBytesIns_Inst_Sbox_10_M7 ;
    wire SubBytesIns_Inst_Sbox_10_M6 ;
    wire SubBytesIns_Inst_Sbox_10_M5 ;
    wire SubBytesIns_Inst_Sbox_10_M4 ;
    wire SubBytesIns_Inst_Sbox_10_M3 ;
    wire SubBytesIns_Inst_Sbox_10_M2 ;
    wire SubBytesIns_Inst_Sbox_10_M1 ;
    wire SubBytesIns_Inst_Sbox_10_T27 ;
    wire SubBytesIns_Inst_Sbox_10_T26 ;
    wire SubBytesIns_Inst_Sbox_10_T25 ;
    wire SubBytesIns_Inst_Sbox_10_T24 ;
    wire SubBytesIns_Inst_Sbox_10_T23 ;
    wire SubBytesIns_Inst_Sbox_10_T22 ;
    wire SubBytesIns_Inst_Sbox_10_T21 ;
    wire SubBytesIns_Inst_Sbox_10_T20 ;
    wire SubBytesIns_Inst_Sbox_10_T19 ;
    wire SubBytesIns_Inst_Sbox_10_T18 ;
    wire SubBytesIns_Inst_Sbox_10_T17 ;
    wire SubBytesIns_Inst_Sbox_10_T16 ;
    wire SubBytesIns_Inst_Sbox_10_T15 ;
    wire SubBytesIns_Inst_Sbox_10_T14 ;
    wire SubBytesIns_Inst_Sbox_10_T13 ;
    wire SubBytesIns_Inst_Sbox_10_T12 ;
    wire SubBytesIns_Inst_Sbox_10_T11 ;
    wire SubBytesIns_Inst_Sbox_10_T10 ;
    wire SubBytesIns_Inst_Sbox_10_T9 ;
    wire SubBytesIns_Inst_Sbox_10_T8 ;
    wire SubBytesIns_Inst_Sbox_10_T7 ;
    wire SubBytesIns_Inst_Sbox_10_T6 ;
    wire SubBytesIns_Inst_Sbox_10_T5 ;
    wire SubBytesIns_Inst_Sbox_10_T4 ;
    wire SubBytesIns_Inst_Sbox_10_T3 ;
    wire SubBytesIns_Inst_Sbox_10_T2 ;
    wire SubBytesIns_Inst_Sbox_10_T1 ;
    wire SubBytesIns_Inst_Sbox_11_L29 ;
    wire SubBytesIns_Inst_Sbox_11_L28 ;
    wire SubBytesIns_Inst_Sbox_11_L27 ;
    wire SubBytesIns_Inst_Sbox_11_L26 ;
    wire SubBytesIns_Inst_Sbox_11_L25 ;
    wire SubBytesIns_Inst_Sbox_11_L24 ;
    wire SubBytesIns_Inst_Sbox_11_L23 ;
    wire SubBytesIns_Inst_Sbox_11_L22 ;
    wire SubBytesIns_Inst_Sbox_11_L21 ;
    wire SubBytesIns_Inst_Sbox_11_L20 ;
    wire SubBytesIns_Inst_Sbox_11_L19 ;
    wire SubBytesIns_Inst_Sbox_11_L18 ;
    wire SubBytesIns_Inst_Sbox_11_L17 ;
    wire SubBytesIns_Inst_Sbox_11_L16 ;
    wire SubBytesIns_Inst_Sbox_11_L15 ;
    wire SubBytesIns_Inst_Sbox_11_L14 ;
    wire SubBytesIns_Inst_Sbox_11_L13 ;
    wire SubBytesIns_Inst_Sbox_11_L12 ;
    wire SubBytesIns_Inst_Sbox_11_L11 ;
    wire SubBytesIns_Inst_Sbox_11_L10 ;
    wire SubBytesIns_Inst_Sbox_11_L9 ;
    wire SubBytesIns_Inst_Sbox_11_L8 ;
    wire SubBytesIns_Inst_Sbox_11_L7 ;
    wire SubBytesIns_Inst_Sbox_11_L6 ;
    wire SubBytesIns_Inst_Sbox_11_L5 ;
    wire SubBytesIns_Inst_Sbox_11_L4 ;
    wire SubBytesIns_Inst_Sbox_11_L3 ;
    wire SubBytesIns_Inst_Sbox_11_L2 ;
    wire SubBytesIns_Inst_Sbox_11_L1 ;
    wire SubBytesIns_Inst_Sbox_11_L0 ;
    wire SubBytesIns_Inst_Sbox_11_M63 ;
    wire SubBytesIns_Inst_Sbox_11_M62 ;
    wire SubBytesIns_Inst_Sbox_11_M61 ;
    wire SubBytesIns_Inst_Sbox_11_M60 ;
    wire SubBytesIns_Inst_Sbox_11_M59 ;
    wire SubBytesIns_Inst_Sbox_11_M58 ;
    wire SubBytesIns_Inst_Sbox_11_M57 ;
    wire SubBytesIns_Inst_Sbox_11_M56 ;
    wire SubBytesIns_Inst_Sbox_11_M55 ;
    wire SubBytesIns_Inst_Sbox_11_M54 ;
    wire SubBytesIns_Inst_Sbox_11_M53 ;
    wire SubBytesIns_Inst_Sbox_11_M52 ;
    wire SubBytesIns_Inst_Sbox_11_M51 ;
    wire SubBytesIns_Inst_Sbox_11_M50 ;
    wire SubBytesIns_Inst_Sbox_11_M49 ;
    wire SubBytesIns_Inst_Sbox_11_M48 ;
    wire SubBytesIns_Inst_Sbox_11_M47 ;
    wire SubBytesIns_Inst_Sbox_11_M46 ;
    wire SubBytesIns_Inst_Sbox_11_M45 ;
    wire SubBytesIns_Inst_Sbox_11_M44 ;
    wire SubBytesIns_Inst_Sbox_11_M43 ;
    wire SubBytesIns_Inst_Sbox_11_M42 ;
    wire SubBytesIns_Inst_Sbox_11_M41 ;
    wire SubBytesIns_Inst_Sbox_11_M40 ;
    wire SubBytesIns_Inst_Sbox_11_M39 ;
    wire SubBytesIns_Inst_Sbox_11_M38 ;
    wire SubBytesIns_Inst_Sbox_11_M37 ;
    wire SubBytesIns_Inst_Sbox_11_M36 ;
    wire SubBytesIns_Inst_Sbox_11_M35 ;
    wire SubBytesIns_Inst_Sbox_11_M34 ;
    wire SubBytesIns_Inst_Sbox_11_M33 ;
    wire SubBytesIns_Inst_Sbox_11_M32 ;
    wire SubBytesIns_Inst_Sbox_11_M31 ;
    wire SubBytesIns_Inst_Sbox_11_M30 ;
    wire SubBytesIns_Inst_Sbox_11_M29 ;
    wire SubBytesIns_Inst_Sbox_11_M28 ;
    wire SubBytesIns_Inst_Sbox_11_M27 ;
    wire SubBytesIns_Inst_Sbox_11_M26 ;
    wire SubBytesIns_Inst_Sbox_11_M25 ;
    wire SubBytesIns_Inst_Sbox_11_M24 ;
    wire SubBytesIns_Inst_Sbox_11_M23 ;
    wire SubBytesIns_Inst_Sbox_11_M22 ;
    wire SubBytesIns_Inst_Sbox_11_M21 ;
    wire SubBytesIns_Inst_Sbox_11_M20 ;
    wire SubBytesIns_Inst_Sbox_11_M19 ;
    wire SubBytesIns_Inst_Sbox_11_M18 ;
    wire SubBytesIns_Inst_Sbox_11_M17 ;
    wire SubBytesIns_Inst_Sbox_11_M16 ;
    wire SubBytesIns_Inst_Sbox_11_M15 ;
    wire SubBytesIns_Inst_Sbox_11_M14 ;
    wire SubBytesIns_Inst_Sbox_11_M13 ;
    wire SubBytesIns_Inst_Sbox_11_M12 ;
    wire SubBytesIns_Inst_Sbox_11_M11 ;
    wire SubBytesIns_Inst_Sbox_11_M10 ;
    wire SubBytesIns_Inst_Sbox_11_M9 ;
    wire SubBytesIns_Inst_Sbox_11_M8 ;
    wire SubBytesIns_Inst_Sbox_11_M7 ;
    wire SubBytesIns_Inst_Sbox_11_M6 ;
    wire SubBytesIns_Inst_Sbox_11_M5 ;
    wire SubBytesIns_Inst_Sbox_11_M4 ;
    wire SubBytesIns_Inst_Sbox_11_M3 ;
    wire SubBytesIns_Inst_Sbox_11_M2 ;
    wire SubBytesIns_Inst_Sbox_11_M1 ;
    wire SubBytesIns_Inst_Sbox_11_T27 ;
    wire SubBytesIns_Inst_Sbox_11_T26 ;
    wire SubBytesIns_Inst_Sbox_11_T25 ;
    wire SubBytesIns_Inst_Sbox_11_T24 ;
    wire SubBytesIns_Inst_Sbox_11_T23 ;
    wire SubBytesIns_Inst_Sbox_11_T22 ;
    wire SubBytesIns_Inst_Sbox_11_T21 ;
    wire SubBytesIns_Inst_Sbox_11_T20 ;
    wire SubBytesIns_Inst_Sbox_11_T19 ;
    wire SubBytesIns_Inst_Sbox_11_T18 ;
    wire SubBytesIns_Inst_Sbox_11_T17 ;
    wire SubBytesIns_Inst_Sbox_11_T16 ;
    wire SubBytesIns_Inst_Sbox_11_T15 ;
    wire SubBytesIns_Inst_Sbox_11_T14 ;
    wire SubBytesIns_Inst_Sbox_11_T13 ;
    wire SubBytesIns_Inst_Sbox_11_T12 ;
    wire SubBytesIns_Inst_Sbox_11_T11 ;
    wire SubBytesIns_Inst_Sbox_11_T10 ;
    wire SubBytesIns_Inst_Sbox_11_T9 ;
    wire SubBytesIns_Inst_Sbox_11_T8 ;
    wire SubBytesIns_Inst_Sbox_11_T7 ;
    wire SubBytesIns_Inst_Sbox_11_T6 ;
    wire SubBytesIns_Inst_Sbox_11_T5 ;
    wire SubBytesIns_Inst_Sbox_11_T4 ;
    wire SubBytesIns_Inst_Sbox_11_T3 ;
    wire SubBytesIns_Inst_Sbox_11_T2 ;
    wire SubBytesIns_Inst_Sbox_11_T1 ;
    wire SubBytesIns_Inst_Sbox_12_L29 ;
    wire SubBytesIns_Inst_Sbox_12_L28 ;
    wire SubBytesIns_Inst_Sbox_12_L27 ;
    wire SubBytesIns_Inst_Sbox_12_L26 ;
    wire SubBytesIns_Inst_Sbox_12_L25 ;
    wire SubBytesIns_Inst_Sbox_12_L24 ;
    wire SubBytesIns_Inst_Sbox_12_L23 ;
    wire SubBytesIns_Inst_Sbox_12_L22 ;
    wire SubBytesIns_Inst_Sbox_12_L21 ;
    wire SubBytesIns_Inst_Sbox_12_L20 ;
    wire SubBytesIns_Inst_Sbox_12_L19 ;
    wire SubBytesIns_Inst_Sbox_12_L18 ;
    wire SubBytesIns_Inst_Sbox_12_L17 ;
    wire SubBytesIns_Inst_Sbox_12_L16 ;
    wire SubBytesIns_Inst_Sbox_12_L15 ;
    wire SubBytesIns_Inst_Sbox_12_L14 ;
    wire SubBytesIns_Inst_Sbox_12_L13 ;
    wire SubBytesIns_Inst_Sbox_12_L12 ;
    wire SubBytesIns_Inst_Sbox_12_L11 ;
    wire SubBytesIns_Inst_Sbox_12_L10 ;
    wire SubBytesIns_Inst_Sbox_12_L9 ;
    wire SubBytesIns_Inst_Sbox_12_L8 ;
    wire SubBytesIns_Inst_Sbox_12_L7 ;
    wire SubBytesIns_Inst_Sbox_12_L6 ;
    wire SubBytesIns_Inst_Sbox_12_L5 ;
    wire SubBytesIns_Inst_Sbox_12_L4 ;
    wire SubBytesIns_Inst_Sbox_12_L3 ;
    wire SubBytesIns_Inst_Sbox_12_L2 ;
    wire SubBytesIns_Inst_Sbox_12_L1 ;
    wire SubBytesIns_Inst_Sbox_12_L0 ;
    wire SubBytesIns_Inst_Sbox_12_M63 ;
    wire SubBytesIns_Inst_Sbox_12_M62 ;
    wire SubBytesIns_Inst_Sbox_12_M61 ;
    wire SubBytesIns_Inst_Sbox_12_M60 ;
    wire SubBytesIns_Inst_Sbox_12_M59 ;
    wire SubBytesIns_Inst_Sbox_12_M58 ;
    wire SubBytesIns_Inst_Sbox_12_M57 ;
    wire SubBytesIns_Inst_Sbox_12_M56 ;
    wire SubBytesIns_Inst_Sbox_12_M55 ;
    wire SubBytesIns_Inst_Sbox_12_M54 ;
    wire SubBytesIns_Inst_Sbox_12_M53 ;
    wire SubBytesIns_Inst_Sbox_12_M52 ;
    wire SubBytesIns_Inst_Sbox_12_M51 ;
    wire SubBytesIns_Inst_Sbox_12_M50 ;
    wire SubBytesIns_Inst_Sbox_12_M49 ;
    wire SubBytesIns_Inst_Sbox_12_M48 ;
    wire SubBytesIns_Inst_Sbox_12_M47 ;
    wire SubBytesIns_Inst_Sbox_12_M46 ;
    wire SubBytesIns_Inst_Sbox_12_M45 ;
    wire SubBytesIns_Inst_Sbox_12_M44 ;
    wire SubBytesIns_Inst_Sbox_12_M43 ;
    wire SubBytesIns_Inst_Sbox_12_M42 ;
    wire SubBytesIns_Inst_Sbox_12_M41 ;
    wire SubBytesIns_Inst_Sbox_12_M40 ;
    wire SubBytesIns_Inst_Sbox_12_M39 ;
    wire SubBytesIns_Inst_Sbox_12_M38 ;
    wire SubBytesIns_Inst_Sbox_12_M37 ;
    wire SubBytesIns_Inst_Sbox_12_M36 ;
    wire SubBytesIns_Inst_Sbox_12_M35 ;
    wire SubBytesIns_Inst_Sbox_12_M34 ;
    wire SubBytesIns_Inst_Sbox_12_M33 ;
    wire SubBytesIns_Inst_Sbox_12_M32 ;
    wire SubBytesIns_Inst_Sbox_12_M31 ;
    wire SubBytesIns_Inst_Sbox_12_M30 ;
    wire SubBytesIns_Inst_Sbox_12_M29 ;
    wire SubBytesIns_Inst_Sbox_12_M28 ;
    wire SubBytesIns_Inst_Sbox_12_M27 ;
    wire SubBytesIns_Inst_Sbox_12_M26 ;
    wire SubBytesIns_Inst_Sbox_12_M25 ;
    wire SubBytesIns_Inst_Sbox_12_M24 ;
    wire SubBytesIns_Inst_Sbox_12_M23 ;
    wire SubBytesIns_Inst_Sbox_12_M22 ;
    wire SubBytesIns_Inst_Sbox_12_M21 ;
    wire SubBytesIns_Inst_Sbox_12_M20 ;
    wire SubBytesIns_Inst_Sbox_12_M19 ;
    wire SubBytesIns_Inst_Sbox_12_M18 ;
    wire SubBytesIns_Inst_Sbox_12_M17 ;
    wire SubBytesIns_Inst_Sbox_12_M16 ;
    wire SubBytesIns_Inst_Sbox_12_M15 ;
    wire SubBytesIns_Inst_Sbox_12_M14 ;
    wire SubBytesIns_Inst_Sbox_12_M13 ;
    wire SubBytesIns_Inst_Sbox_12_M12 ;
    wire SubBytesIns_Inst_Sbox_12_M11 ;
    wire SubBytesIns_Inst_Sbox_12_M10 ;
    wire SubBytesIns_Inst_Sbox_12_M9 ;
    wire SubBytesIns_Inst_Sbox_12_M8 ;
    wire SubBytesIns_Inst_Sbox_12_M7 ;
    wire SubBytesIns_Inst_Sbox_12_M6 ;
    wire SubBytesIns_Inst_Sbox_12_M5 ;
    wire SubBytesIns_Inst_Sbox_12_M4 ;
    wire SubBytesIns_Inst_Sbox_12_M3 ;
    wire SubBytesIns_Inst_Sbox_12_M2 ;
    wire SubBytesIns_Inst_Sbox_12_M1 ;
    wire SubBytesIns_Inst_Sbox_12_T27 ;
    wire SubBytesIns_Inst_Sbox_12_T26 ;
    wire SubBytesIns_Inst_Sbox_12_T25 ;
    wire SubBytesIns_Inst_Sbox_12_T24 ;
    wire SubBytesIns_Inst_Sbox_12_T23 ;
    wire SubBytesIns_Inst_Sbox_12_T22 ;
    wire SubBytesIns_Inst_Sbox_12_T21 ;
    wire SubBytesIns_Inst_Sbox_12_T20 ;
    wire SubBytesIns_Inst_Sbox_12_T19 ;
    wire SubBytesIns_Inst_Sbox_12_T18 ;
    wire SubBytesIns_Inst_Sbox_12_T17 ;
    wire SubBytesIns_Inst_Sbox_12_T16 ;
    wire SubBytesIns_Inst_Sbox_12_T15 ;
    wire SubBytesIns_Inst_Sbox_12_T14 ;
    wire SubBytesIns_Inst_Sbox_12_T13 ;
    wire SubBytesIns_Inst_Sbox_12_T12 ;
    wire SubBytesIns_Inst_Sbox_12_T11 ;
    wire SubBytesIns_Inst_Sbox_12_T10 ;
    wire SubBytesIns_Inst_Sbox_12_T9 ;
    wire SubBytesIns_Inst_Sbox_12_T8 ;
    wire SubBytesIns_Inst_Sbox_12_T7 ;
    wire SubBytesIns_Inst_Sbox_12_T6 ;
    wire SubBytesIns_Inst_Sbox_12_T5 ;
    wire SubBytesIns_Inst_Sbox_12_T4 ;
    wire SubBytesIns_Inst_Sbox_12_T3 ;
    wire SubBytesIns_Inst_Sbox_12_T2 ;
    wire SubBytesIns_Inst_Sbox_12_T1 ;
    wire SubBytesIns_Inst_Sbox_13_L29 ;
    wire SubBytesIns_Inst_Sbox_13_L28 ;
    wire SubBytesIns_Inst_Sbox_13_L27 ;
    wire SubBytesIns_Inst_Sbox_13_L26 ;
    wire SubBytesIns_Inst_Sbox_13_L25 ;
    wire SubBytesIns_Inst_Sbox_13_L24 ;
    wire SubBytesIns_Inst_Sbox_13_L23 ;
    wire SubBytesIns_Inst_Sbox_13_L22 ;
    wire SubBytesIns_Inst_Sbox_13_L21 ;
    wire SubBytesIns_Inst_Sbox_13_L20 ;
    wire SubBytesIns_Inst_Sbox_13_L19 ;
    wire SubBytesIns_Inst_Sbox_13_L18 ;
    wire SubBytesIns_Inst_Sbox_13_L17 ;
    wire SubBytesIns_Inst_Sbox_13_L16 ;
    wire SubBytesIns_Inst_Sbox_13_L15 ;
    wire SubBytesIns_Inst_Sbox_13_L14 ;
    wire SubBytesIns_Inst_Sbox_13_L13 ;
    wire SubBytesIns_Inst_Sbox_13_L12 ;
    wire SubBytesIns_Inst_Sbox_13_L11 ;
    wire SubBytesIns_Inst_Sbox_13_L10 ;
    wire SubBytesIns_Inst_Sbox_13_L9 ;
    wire SubBytesIns_Inst_Sbox_13_L8 ;
    wire SubBytesIns_Inst_Sbox_13_L7 ;
    wire SubBytesIns_Inst_Sbox_13_L6 ;
    wire SubBytesIns_Inst_Sbox_13_L5 ;
    wire SubBytesIns_Inst_Sbox_13_L4 ;
    wire SubBytesIns_Inst_Sbox_13_L3 ;
    wire SubBytesIns_Inst_Sbox_13_L2 ;
    wire SubBytesIns_Inst_Sbox_13_L1 ;
    wire SubBytesIns_Inst_Sbox_13_L0 ;
    wire SubBytesIns_Inst_Sbox_13_M63 ;
    wire SubBytesIns_Inst_Sbox_13_M62 ;
    wire SubBytesIns_Inst_Sbox_13_M61 ;
    wire SubBytesIns_Inst_Sbox_13_M60 ;
    wire SubBytesIns_Inst_Sbox_13_M59 ;
    wire SubBytesIns_Inst_Sbox_13_M58 ;
    wire SubBytesIns_Inst_Sbox_13_M57 ;
    wire SubBytesIns_Inst_Sbox_13_M56 ;
    wire SubBytesIns_Inst_Sbox_13_M55 ;
    wire SubBytesIns_Inst_Sbox_13_M54 ;
    wire SubBytesIns_Inst_Sbox_13_M53 ;
    wire SubBytesIns_Inst_Sbox_13_M52 ;
    wire SubBytesIns_Inst_Sbox_13_M51 ;
    wire SubBytesIns_Inst_Sbox_13_M50 ;
    wire SubBytesIns_Inst_Sbox_13_M49 ;
    wire SubBytesIns_Inst_Sbox_13_M48 ;
    wire SubBytesIns_Inst_Sbox_13_M47 ;
    wire SubBytesIns_Inst_Sbox_13_M46 ;
    wire SubBytesIns_Inst_Sbox_13_M45 ;
    wire SubBytesIns_Inst_Sbox_13_M44 ;
    wire SubBytesIns_Inst_Sbox_13_M43 ;
    wire SubBytesIns_Inst_Sbox_13_M42 ;
    wire SubBytesIns_Inst_Sbox_13_M41 ;
    wire SubBytesIns_Inst_Sbox_13_M40 ;
    wire SubBytesIns_Inst_Sbox_13_M39 ;
    wire SubBytesIns_Inst_Sbox_13_M38 ;
    wire SubBytesIns_Inst_Sbox_13_M37 ;
    wire SubBytesIns_Inst_Sbox_13_M36 ;
    wire SubBytesIns_Inst_Sbox_13_M35 ;
    wire SubBytesIns_Inst_Sbox_13_M34 ;
    wire SubBytesIns_Inst_Sbox_13_M33 ;
    wire SubBytesIns_Inst_Sbox_13_M32 ;
    wire SubBytesIns_Inst_Sbox_13_M31 ;
    wire SubBytesIns_Inst_Sbox_13_M30 ;
    wire SubBytesIns_Inst_Sbox_13_M29 ;
    wire SubBytesIns_Inst_Sbox_13_M28 ;
    wire SubBytesIns_Inst_Sbox_13_M27 ;
    wire SubBytesIns_Inst_Sbox_13_M26 ;
    wire SubBytesIns_Inst_Sbox_13_M25 ;
    wire SubBytesIns_Inst_Sbox_13_M24 ;
    wire SubBytesIns_Inst_Sbox_13_M23 ;
    wire SubBytesIns_Inst_Sbox_13_M22 ;
    wire SubBytesIns_Inst_Sbox_13_M21 ;
    wire SubBytesIns_Inst_Sbox_13_M20 ;
    wire SubBytesIns_Inst_Sbox_13_M19 ;
    wire SubBytesIns_Inst_Sbox_13_M18 ;
    wire SubBytesIns_Inst_Sbox_13_M17 ;
    wire SubBytesIns_Inst_Sbox_13_M16 ;
    wire SubBytesIns_Inst_Sbox_13_M15 ;
    wire SubBytesIns_Inst_Sbox_13_M14 ;
    wire SubBytesIns_Inst_Sbox_13_M13 ;
    wire SubBytesIns_Inst_Sbox_13_M12 ;
    wire SubBytesIns_Inst_Sbox_13_M11 ;
    wire SubBytesIns_Inst_Sbox_13_M10 ;
    wire SubBytesIns_Inst_Sbox_13_M9 ;
    wire SubBytesIns_Inst_Sbox_13_M8 ;
    wire SubBytesIns_Inst_Sbox_13_M7 ;
    wire SubBytesIns_Inst_Sbox_13_M6 ;
    wire SubBytesIns_Inst_Sbox_13_M5 ;
    wire SubBytesIns_Inst_Sbox_13_M4 ;
    wire SubBytesIns_Inst_Sbox_13_M3 ;
    wire SubBytesIns_Inst_Sbox_13_M2 ;
    wire SubBytesIns_Inst_Sbox_13_M1 ;
    wire SubBytesIns_Inst_Sbox_13_T27 ;
    wire SubBytesIns_Inst_Sbox_13_T26 ;
    wire SubBytesIns_Inst_Sbox_13_T25 ;
    wire SubBytesIns_Inst_Sbox_13_T24 ;
    wire SubBytesIns_Inst_Sbox_13_T23 ;
    wire SubBytesIns_Inst_Sbox_13_T22 ;
    wire SubBytesIns_Inst_Sbox_13_T21 ;
    wire SubBytesIns_Inst_Sbox_13_T20 ;
    wire SubBytesIns_Inst_Sbox_13_T19 ;
    wire SubBytesIns_Inst_Sbox_13_T18 ;
    wire SubBytesIns_Inst_Sbox_13_T17 ;
    wire SubBytesIns_Inst_Sbox_13_T16 ;
    wire SubBytesIns_Inst_Sbox_13_T15 ;
    wire SubBytesIns_Inst_Sbox_13_T14 ;
    wire SubBytesIns_Inst_Sbox_13_T13 ;
    wire SubBytesIns_Inst_Sbox_13_T12 ;
    wire SubBytesIns_Inst_Sbox_13_T11 ;
    wire SubBytesIns_Inst_Sbox_13_T10 ;
    wire SubBytesIns_Inst_Sbox_13_T9 ;
    wire SubBytesIns_Inst_Sbox_13_T8 ;
    wire SubBytesIns_Inst_Sbox_13_T7 ;
    wire SubBytesIns_Inst_Sbox_13_T6 ;
    wire SubBytesIns_Inst_Sbox_13_T5 ;
    wire SubBytesIns_Inst_Sbox_13_T4 ;
    wire SubBytesIns_Inst_Sbox_13_T3 ;
    wire SubBytesIns_Inst_Sbox_13_T2 ;
    wire SubBytesIns_Inst_Sbox_13_T1 ;
    wire SubBytesIns_Inst_Sbox_14_L29 ;
    wire SubBytesIns_Inst_Sbox_14_L28 ;
    wire SubBytesIns_Inst_Sbox_14_L27 ;
    wire SubBytesIns_Inst_Sbox_14_L26 ;
    wire SubBytesIns_Inst_Sbox_14_L25 ;
    wire SubBytesIns_Inst_Sbox_14_L24 ;
    wire SubBytesIns_Inst_Sbox_14_L23 ;
    wire SubBytesIns_Inst_Sbox_14_L22 ;
    wire SubBytesIns_Inst_Sbox_14_L21 ;
    wire SubBytesIns_Inst_Sbox_14_L20 ;
    wire SubBytesIns_Inst_Sbox_14_L19 ;
    wire SubBytesIns_Inst_Sbox_14_L18 ;
    wire SubBytesIns_Inst_Sbox_14_L17 ;
    wire SubBytesIns_Inst_Sbox_14_L16 ;
    wire SubBytesIns_Inst_Sbox_14_L15 ;
    wire SubBytesIns_Inst_Sbox_14_L14 ;
    wire SubBytesIns_Inst_Sbox_14_L13 ;
    wire SubBytesIns_Inst_Sbox_14_L12 ;
    wire SubBytesIns_Inst_Sbox_14_L11 ;
    wire SubBytesIns_Inst_Sbox_14_L10 ;
    wire SubBytesIns_Inst_Sbox_14_L9 ;
    wire SubBytesIns_Inst_Sbox_14_L8 ;
    wire SubBytesIns_Inst_Sbox_14_L7 ;
    wire SubBytesIns_Inst_Sbox_14_L6 ;
    wire SubBytesIns_Inst_Sbox_14_L5 ;
    wire SubBytesIns_Inst_Sbox_14_L4 ;
    wire SubBytesIns_Inst_Sbox_14_L3 ;
    wire SubBytesIns_Inst_Sbox_14_L2 ;
    wire SubBytesIns_Inst_Sbox_14_L1 ;
    wire SubBytesIns_Inst_Sbox_14_L0 ;
    wire SubBytesIns_Inst_Sbox_14_M63 ;
    wire SubBytesIns_Inst_Sbox_14_M62 ;
    wire SubBytesIns_Inst_Sbox_14_M61 ;
    wire SubBytesIns_Inst_Sbox_14_M60 ;
    wire SubBytesIns_Inst_Sbox_14_M59 ;
    wire SubBytesIns_Inst_Sbox_14_M58 ;
    wire SubBytesIns_Inst_Sbox_14_M57 ;
    wire SubBytesIns_Inst_Sbox_14_M56 ;
    wire SubBytesIns_Inst_Sbox_14_M55 ;
    wire SubBytesIns_Inst_Sbox_14_M54 ;
    wire SubBytesIns_Inst_Sbox_14_M53 ;
    wire SubBytesIns_Inst_Sbox_14_M52 ;
    wire SubBytesIns_Inst_Sbox_14_M51 ;
    wire SubBytesIns_Inst_Sbox_14_M50 ;
    wire SubBytesIns_Inst_Sbox_14_M49 ;
    wire SubBytesIns_Inst_Sbox_14_M48 ;
    wire SubBytesIns_Inst_Sbox_14_M47 ;
    wire SubBytesIns_Inst_Sbox_14_M46 ;
    wire SubBytesIns_Inst_Sbox_14_M45 ;
    wire SubBytesIns_Inst_Sbox_14_M44 ;
    wire SubBytesIns_Inst_Sbox_14_M43 ;
    wire SubBytesIns_Inst_Sbox_14_M42 ;
    wire SubBytesIns_Inst_Sbox_14_M41 ;
    wire SubBytesIns_Inst_Sbox_14_M40 ;
    wire SubBytesIns_Inst_Sbox_14_M39 ;
    wire SubBytesIns_Inst_Sbox_14_M38 ;
    wire SubBytesIns_Inst_Sbox_14_M37 ;
    wire SubBytesIns_Inst_Sbox_14_M36 ;
    wire SubBytesIns_Inst_Sbox_14_M35 ;
    wire SubBytesIns_Inst_Sbox_14_M34 ;
    wire SubBytesIns_Inst_Sbox_14_M33 ;
    wire SubBytesIns_Inst_Sbox_14_M32 ;
    wire SubBytesIns_Inst_Sbox_14_M31 ;
    wire SubBytesIns_Inst_Sbox_14_M30 ;
    wire SubBytesIns_Inst_Sbox_14_M29 ;
    wire SubBytesIns_Inst_Sbox_14_M28 ;
    wire SubBytesIns_Inst_Sbox_14_M27 ;
    wire SubBytesIns_Inst_Sbox_14_M26 ;
    wire SubBytesIns_Inst_Sbox_14_M25 ;
    wire SubBytesIns_Inst_Sbox_14_M24 ;
    wire SubBytesIns_Inst_Sbox_14_M23 ;
    wire SubBytesIns_Inst_Sbox_14_M22 ;
    wire SubBytesIns_Inst_Sbox_14_M21 ;
    wire SubBytesIns_Inst_Sbox_14_M20 ;
    wire SubBytesIns_Inst_Sbox_14_M19 ;
    wire SubBytesIns_Inst_Sbox_14_M18 ;
    wire SubBytesIns_Inst_Sbox_14_M17 ;
    wire SubBytesIns_Inst_Sbox_14_M16 ;
    wire SubBytesIns_Inst_Sbox_14_M15 ;
    wire SubBytesIns_Inst_Sbox_14_M14 ;
    wire SubBytesIns_Inst_Sbox_14_M13 ;
    wire SubBytesIns_Inst_Sbox_14_M12 ;
    wire SubBytesIns_Inst_Sbox_14_M11 ;
    wire SubBytesIns_Inst_Sbox_14_M10 ;
    wire SubBytesIns_Inst_Sbox_14_M9 ;
    wire SubBytesIns_Inst_Sbox_14_M8 ;
    wire SubBytesIns_Inst_Sbox_14_M7 ;
    wire SubBytesIns_Inst_Sbox_14_M6 ;
    wire SubBytesIns_Inst_Sbox_14_M5 ;
    wire SubBytesIns_Inst_Sbox_14_M4 ;
    wire SubBytesIns_Inst_Sbox_14_M3 ;
    wire SubBytesIns_Inst_Sbox_14_M2 ;
    wire SubBytesIns_Inst_Sbox_14_M1 ;
    wire SubBytesIns_Inst_Sbox_14_T27 ;
    wire SubBytesIns_Inst_Sbox_14_T26 ;
    wire SubBytesIns_Inst_Sbox_14_T25 ;
    wire SubBytesIns_Inst_Sbox_14_T24 ;
    wire SubBytesIns_Inst_Sbox_14_T23 ;
    wire SubBytesIns_Inst_Sbox_14_T22 ;
    wire SubBytesIns_Inst_Sbox_14_T21 ;
    wire SubBytesIns_Inst_Sbox_14_T20 ;
    wire SubBytesIns_Inst_Sbox_14_T19 ;
    wire SubBytesIns_Inst_Sbox_14_T18 ;
    wire SubBytesIns_Inst_Sbox_14_T17 ;
    wire SubBytesIns_Inst_Sbox_14_T16 ;
    wire SubBytesIns_Inst_Sbox_14_T15 ;
    wire SubBytesIns_Inst_Sbox_14_T14 ;
    wire SubBytesIns_Inst_Sbox_14_T13 ;
    wire SubBytesIns_Inst_Sbox_14_T12 ;
    wire SubBytesIns_Inst_Sbox_14_T11 ;
    wire SubBytesIns_Inst_Sbox_14_T10 ;
    wire SubBytesIns_Inst_Sbox_14_T9 ;
    wire SubBytesIns_Inst_Sbox_14_T8 ;
    wire SubBytesIns_Inst_Sbox_14_T7 ;
    wire SubBytesIns_Inst_Sbox_14_T6 ;
    wire SubBytesIns_Inst_Sbox_14_T5 ;
    wire SubBytesIns_Inst_Sbox_14_T4 ;
    wire SubBytesIns_Inst_Sbox_14_T3 ;
    wire SubBytesIns_Inst_Sbox_14_T2 ;
    wire SubBytesIns_Inst_Sbox_14_T1 ;
    wire SubBytesIns_Inst_Sbox_15_L29 ;
    wire SubBytesIns_Inst_Sbox_15_L28 ;
    wire SubBytesIns_Inst_Sbox_15_L27 ;
    wire SubBytesIns_Inst_Sbox_15_L26 ;
    wire SubBytesIns_Inst_Sbox_15_L25 ;
    wire SubBytesIns_Inst_Sbox_15_L24 ;
    wire SubBytesIns_Inst_Sbox_15_L23 ;
    wire SubBytesIns_Inst_Sbox_15_L22 ;
    wire SubBytesIns_Inst_Sbox_15_L21 ;
    wire SubBytesIns_Inst_Sbox_15_L20 ;
    wire SubBytesIns_Inst_Sbox_15_L19 ;
    wire SubBytesIns_Inst_Sbox_15_L18 ;
    wire SubBytesIns_Inst_Sbox_15_L17 ;
    wire SubBytesIns_Inst_Sbox_15_L16 ;
    wire SubBytesIns_Inst_Sbox_15_L15 ;
    wire SubBytesIns_Inst_Sbox_15_L14 ;
    wire SubBytesIns_Inst_Sbox_15_L13 ;
    wire SubBytesIns_Inst_Sbox_15_L12 ;
    wire SubBytesIns_Inst_Sbox_15_L11 ;
    wire SubBytesIns_Inst_Sbox_15_L10 ;
    wire SubBytesIns_Inst_Sbox_15_L9 ;
    wire SubBytesIns_Inst_Sbox_15_L8 ;
    wire SubBytesIns_Inst_Sbox_15_L7 ;
    wire SubBytesIns_Inst_Sbox_15_L6 ;
    wire SubBytesIns_Inst_Sbox_15_L5 ;
    wire SubBytesIns_Inst_Sbox_15_L4 ;
    wire SubBytesIns_Inst_Sbox_15_L3 ;
    wire SubBytesIns_Inst_Sbox_15_L2 ;
    wire SubBytesIns_Inst_Sbox_15_L1 ;
    wire SubBytesIns_Inst_Sbox_15_L0 ;
    wire SubBytesIns_Inst_Sbox_15_M63 ;
    wire SubBytesIns_Inst_Sbox_15_M62 ;
    wire SubBytesIns_Inst_Sbox_15_M61 ;
    wire SubBytesIns_Inst_Sbox_15_M60 ;
    wire SubBytesIns_Inst_Sbox_15_M59 ;
    wire SubBytesIns_Inst_Sbox_15_M58 ;
    wire SubBytesIns_Inst_Sbox_15_M57 ;
    wire SubBytesIns_Inst_Sbox_15_M56 ;
    wire SubBytesIns_Inst_Sbox_15_M55 ;
    wire SubBytesIns_Inst_Sbox_15_M54 ;
    wire SubBytesIns_Inst_Sbox_15_M53 ;
    wire SubBytesIns_Inst_Sbox_15_M52 ;
    wire SubBytesIns_Inst_Sbox_15_M51 ;
    wire SubBytesIns_Inst_Sbox_15_M50 ;
    wire SubBytesIns_Inst_Sbox_15_M49 ;
    wire SubBytesIns_Inst_Sbox_15_M48 ;
    wire SubBytesIns_Inst_Sbox_15_M47 ;
    wire SubBytesIns_Inst_Sbox_15_M46 ;
    wire SubBytesIns_Inst_Sbox_15_M45 ;
    wire SubBytesIns_Inst_Sbox_15_M44 ;
    wire SubBytesIns_Inst_Sbox_15_M43 ;
    wire SubBytesIns_Inst_Sbox_15_M42 ;
    wire SubBytesIns_Inst_Sbox_15_M41 ;
    wire SubBytesIns_Inst_Sbox_15_M40 ;
    wire SubBytesIns_Inst_Sbox_15_M39 ;
    wire SubBytesIns_Inst_Sbox_15_M38 ;
    wire SubBytesIns_Inst_Sbox_15_M37 ;
    wire SubBytesIns_Inst_Sbox_15_M36 ;
    wire SubBytesIns_Inst_Sbox_15_M35 ;
    wire SubBytesIns_Inst_Sbox_15_M34 ;
    wire SubBytesIns_Inst_Sbox_15_M33 ;
    wire SubBytesIns_Inst_Sbox_15_M32 ;
    wire SubBytesIns_Inst_Sbox_15_M31 ;
    wire SubBytesIns_Inst_Sbox_15_M30 ;
    wire SubBytesIns_Inst_Sbox_15_M29 ;
    wire SubBytesIns_Inst_Sbox_15_M28 ;
    wire SubBytesIns_Inst_Sbox_15_M27 ;
    wire SubBytesIns_Inst_Sbox_15_M26 ;
    wire SubBytesIns_Inst_Sbox_15_M25 ;
    wire SubBytesIns_Inst_Sbox_15_M24 ;
    wire SubBytesIns_Inst_Sbox_15_M23 ;
    wire SubBytesIns_Inst_Sbox_15_M22 ;
    wire SubBytesIns_Inst_Sbox_15_M21 ;
    wire SubBytesIns_Inst_Sbox_15_M20 ;
    wire SubBytesIns_Inst_Sbox_15_M19 ;
    wire SubBytesIns_Inst_Sbox_15_M18 ;
    wire SubBytesIns_Inst_Sbox_15_M17 ;
    wire SubBytesIns_Inst_Sbox_15_M16 ;
    wire SubBytesIns_Inst_Sbox_15_M15 ;
    wire SubBytesIns_Inst_Sbox_15_M14 ;
    wire SubBytesIns_Inst_Sbox_15_M13 ;
    wire SubBytesIns_Inst_Sbox_15_M12 ;
    wire SubBytesIns_Inst_Sbox_15_M11 ;
    wire SubBytesIns_Inst_Sbox_15_M10 ;
    wire SubBytesIns_Inst_Sbox_15_M9 ;
    wire SubBytesIns_Inst_Sbox_15_M8 ;
    wire SubBytesIns_Inst_Sbox_15_M7 ;
    wire SubBytesIns_Inst_Sbox_15_M6 ;
    wire SubBytesIns_Inst_Sbox_15_M5 ;
    wire SubBytesIns_Inst_Sbox_15_M4 ;
    wire SubBytesIns_Inst_Sbox_15_M3 ;
    wire SubBytesIns_Inst_Sbox_15_M2 ;
    wire SubBytesIns_Inst_Sbox_15_M1 ;
    wire SubBytesIns_Inst_Sbox_15_T27 ;
    wire SubBytesIns_Inst_Sbox_15_T26 ;
    wire SubBytesIns_Inst_Sbox_15_T25 ;
    wire SubBytesIns_Inst_Sbox_15_T24 ;
    wire SubBytesIns_Inst_Sbox_15_T23 ;
    wire SubBytesIns_Inst_Sbox_15_T22 ;
    wire SubBytesIns_Inst_Sbox_15_T21 ;
    wire SubBytesIns_Inst_Sbox_15_T20 ;
    wire SubBytesIns_Inst_Sbox_15_T19 ;
    wire SubBytesIns_Inst_Sbox_15_T18 ;
    wire SubBytesIns_Inst_Sbox_15_T17 ;
    wire SubBytesIns_Inst_Sbox_15_T16 ;
    wire SubBytesIns_Inst_Sbox_15_T15 ;
    wire SubBytesIns_Inst_Sbox_15_T14 ;
    wire SubBytesIns_Inst_Sbox_15_T13 ;
    wire SubBytesIns_Inst_Sbox_15_T12 ;
    wire SubBytesIns_Inst_Sbox_15_T11 ;
    wire SubBytesIns_Inst_Sbox_15_T10 ;
    wire SubBytesIns_Inst_Sbox_15_T9 ;
    wire SubBytesIns_Inst_Sbox_15_T8 ;
    wire SubBytesIns_Inst_Sbox_15_T7 ;
    wire SubBytesIns_Inst_Sbox_15_T6 ;
    wire SubBytesIns_Inst_Sbox_15_T5 ;
    wire SubBytesIns_Inst_Sbox_15_T4 ;
    wire SubBytesIns_Inst_Sbox_15_T3 ;
    wire SubBytesIns_Inst_Sbox_15_T2 ;
    wire SubBytesIns_Inst_Sbox_15_T1 ;
    wire MixColumnsIns_MixOneColumnInst_0_n64 ;
    wire MixColumnsIns_MixOneColumnInst_0_n63 ;
    wire MixColumnsIns_MixOneColumnInst_0_n62 ;
    wire MixColumnsIns_MixOneColumnInst_0_n61 ;
    wire MixColumnsIns_MixOneColumnInst_0_n60 ;
    wire MixColumnsIns_MixOneColumnInst_0_n59 ;
    wire MixColumnsIns_MixOneColumnInst_0_n58 ;
    wire MixColumnsIns_MixOneColumnInst_0_n57 ;
    wire MixColumnsIns_MixOneColumnInst_0_n56 ;
    wire MixColumnsIns_MixOneColumnInst_0_n55 ;
    wire MixColumnsIns_MixOneColumnInst_0_n54 ;
    wire MixColumnsIns_MixOneColumnInst_0_n53 ;
    wire MixColumnsIns_MixOneColumnInst_0_n52 ;
    wire MixColumnsIns_MixOneColumnInst_0_n51 ;
    wire MixColumnsIns_MixOneColumnInst_0_n50 ;
    wire MixColumnsIns_MixOneColumnInst_0_n49 ;
    wire MixColumnsIns_MixOneColumnInst_0_n48 ;
    wire MixColumnsIns_MixOneColumnInst_0_n47 ;
    wire MixColumnsIns_MixOneColumnInst_0_n46 ;
    wire MixColumnsIns_MixOneColumnInst_0_n45 ;
    wire MixColumnsIns_MixOneColumnInst_0_n44 ;
    wire MixColumnsIns_MixOneColumnInst_0_n43 ;
    wire MixColumnsIns_MixOneColumnInst_0_n42 ;
    wire MixColumnsIns_MixOneColumnInst_0_n41 ;
    wire MixColumnsIns_MixOneColumnInst_0_n40 ;
    wire MixColumnsIns_MixOneColumnInst_0_n39 ;
    wire MixColumnsIns_MixOneColumnInst_0_n38 ;
    wire MixColumnsIns_MixOneColumnInst_0_n37 ;
    wire MixColumnsIns_MixOneColumnInst_0_n36 ;
    wire MixColumnsIns_MixOneColumnInst_0_n35 ;
    wire MixColumnsIns_MixOneColumnInst_0_n34 ;
    wire MixColumnsIns_MixOneColumnInst_0_n33 ;
    wire MixColumnsIns_MixOneColumnInst_0_n32 ;
    wire MixColumnsIns_MixOneColumnInst_0_n31 ;
    wire MixColumnsIns_MixOneColumnInst_0_n30 ;
    wire MixColumnsIns_MixOneColumnInst_0_n29 ;
    wire MixColumnsIns_MixOneColumnInst_0_n28 ;
    wire MixColumnsIns_MixOneColumnInst_0_n27 ;
    wire MixColumnsIns_MixOneColumnInst_0_n26 ;
    wire MixColumnsIns_MixOneColumnInst_0_n25 ;
    wire MixColumnsIns_MixOneColumnInst_0_n24 ;
    wire MixColumnsIns_MixOneColumnInst_0_n23 ;
    wire MixColumnsIns_MixOneColumnInst_0_n22 ;
    wire MixColumnsIns_MixOneColumnInst_0_n21 ;
    wire MixColumnsIns_MixOneColumnInst_0_n20 ;
    wire MixColumnsIns_MixOneColumnInst_0_n19 ;
    wire MixColumnsIns_MixOneColumnInst_0_n18 ;
    wire MixColumnsIns_MixOneColumnInst_0_n17 ;
    wire MixColumnsIns_MixOneColumnInst_0_n16 ;
    wire MixColumnsIns_MixOneColumnInst_0_n15 ;
    wire MixColumnsIns_MixOneColumnInst_0_n14 ;
    wire MixColumnsIns_MixOneColumnInst_0_n13 ;
    wire MixColumnsIns_MixOneColumnInst_0_n12 ;
    wire MixColumnsIns_MixOneColumnInst_0_n11 ;
    wire MixColumnsIns_MixOneColumnInst_0_n10 ;
    wire MixColumnsIns_MixOneColumnInst_0_n9 ;
    wire MixColumnsIns_MixOneColumnInst_0_n8 ;
    wire MixColumnsIns_MixOneColumnInst_0_n7 ;
    wire MixColumnsIns_MixOneColumnInst_0_n6 ;
    wire MixColumnsIns_MixOneColumnInst_0_n5 ;
    wire MixColumnsIns_MixOneColumnInst_0_n4 ;
    wire MixColumnsIns_MixOneColumnInst_0_n3 ;
    wire MixColumnsIns_MixOneColumnInst_0_n2 ;
    wire MixColumnsIns_MixOneColumnInst_0_n1 ;
    wire MixColumnsIns_MixOneColumnInst_1_n64 ;
    wire MixColumnsIns_MixOneColumnInst_1_n63 ;
    wire MixColumnsIns_MixOneColumnInst_1_n62 ;
    wire MixColumnsIns_MixOneColumnInst_1_n61 ;
    wire MixColumnsIns_MixOneColumnInst_1_n60 ;
    wire MixColumnsIns_MixOneColumnInst_1_n59 ;
    wire MixColumnsIns_MixOneColumnInst_1_n58 ;
    wire MixColumnsIns_MixOneColumnInst_1_n57 ;
    wire MixColumnsIns_MixOneColumnInst_1_n56 ;
    wire MixColumnsIns_MixOneColumnInst_1_n55 ;
    wire MixColumnsIns_MixOneColumnInst_1_n54 ;
    wire MixColumnsIns_MixOneColumnInst_1_n53 ;
    wire MixColumnsIns_MixOneColumnInst_1_n52 ;
    wire MixColumnsIns_MixOneColumnInst_1_n51 ;
    wire MixColumnsIns_MixOneColumnInst_1_n50 ;
    wire MixColumnsIns_MixOneColumnInst_1_n49 ;
    wire MixColumnsIns_MixOneColumnInst_1_n48 ;
    wire MixColumnsIns_MixOneColumnInst_1_n47 ;
    wire MixColumnsIns_MixOneColumnInst_1_n46 ;
    wire MixColumnsIns_MixOneColumnInst_1_n45 ;
    wire MixColumnsIns_MixOneColumnInst_1_n44 ;
    wire MixColumnsIns_MixOneColumnInst_1_n43 ;
    wire MixColumnsIns_MixOneColumnInst_1_n42 ;
    wire MixColumnsIns_MixOneColumnInst_1_n41 ;
    wire MixColumnsIns_MixOneColumnInst_1_n40 ;
    wire MixColumnsIns_MixOneColumnInst_1_n39 ;
    wire MixColumnsIns_MixOneColumnInst_1_n38 ;
    wire MixColumnsIns_MixOneColumnInst_1_n37 ;
    wire MixColumnsIns_MixOneColumnInst_1_n36 ;
    wire MixColumnsIns_MixOneColumnInst_1_n35 ;
    wire MixColumnsIns_MixOneColumnInst_1_n34 ;
    wire MixColumnsIns_MixOneColumnInst_1_n33 ;
    wire MixColumnsIns_MixOneColumnInst_1_n32 ;
    wire MixColumnsIns_MixOneColumnInst_1_n31 ;
    wire MixColumnsIns_MixOneColumnInst_1_n30 ;
    wire MixColumnsIns_MixOneColumnInst_1_n29 ;
    wire MixColumnsIns_MixOneColumnInst_1_n28 ;
    wire MixColumnsIns_MixOneColumnInst_1_n27 ;
    wire MixColumnsIns_MixOneColumnInst_1_n26 ;
    wire MixColumnsIns_MixOneColumnInst_1_n25 ;
    wire MixColumnsIns_MixOneColumnInst_1_n24 ;
    wire MixColumnsIns_MixOneColumnInst_1_n23 ;
    wire MixColumnsIns_MixOneColumnInst_1_n22 ;
    wire MixColumnsIns_MixOneColumnInst_1_n21 ;
    wire MixColumnsIns_MixOneColumnInst_1_n20 ;
    wire MixColumnsIns_MixOneColumnInst_1_n19 ;
    wire MixColumnsIns_MixOneColumnInst_1_n18 ;
    wire MixColumnsIns_MixOneColumnInst_1_n17 ;
    wire MixColumnsIns_MixOneColumnInst_1_n16 ;
    wire MixColumnsIns_MixOneColumnInst_1_n15 ;
    wire MixColumnsIns_MixOneColumnInst_1_n14 ;
    wire MixColumnsIns_MixOneColumnInst_1_n13 ;
    wire MixColumnsIns_MixOneColumnInst_1_n12 ;
    wire MixColumnsIns_MixOneColumnInst_1_n11 ;
    wire MixColumnsIns_MixOneColumnInst_1_n10 ;
    wire MixColumnsIns_MixOneColumnInst_1_n9 ;
    wire MixColumnsIns_MixOneColumnInst_1_n8 ;
    wire MixColumnsIns_MixOneColumnInst_1_n7 ;
    wire MixColumnsIns_MixOneColumnInst_1_n6 ;
    wire MixColumnsIns_MixOneColumnInst_1_n5 ;
    wire MixColumnsIns_MixOneColumnInst_1_n4 ;
    wire MixColumnsIns_MixOneColumnInst_1_n3 ;
    wire MixColumnsIns_MixOneColumnInst_1_n2 ;
    wire MixColumnsIns_MixOneColumnInst_1_n1 ;
    wire MixColumnsIns_MixOneColumnInst_2_n64 ;
    wire MixColumnsIns_MixOneColumnInst_2_n63 ;
    wire MixColumnsIns_MixOneColumnInst_2_n62 ;
    wire MixColumnsIns_MixOneColumnInst_2_n61 ;
    wire MixColumnsIns_MixOneColumnInst_2_n60 ;
    wire MixColumnsIns_MixOneColumnInst_2_n59 ;
    wire MixColumnsIns_MixOneColumnInst_2_n58 ;
    wire MixColumnsIns_MixOneColumnInst_2_n57 ;
    wire MixColumnsIns_MixOneColumnInst_2_n56 ;
    wire MixColumnsIns_MixOneColumnInst_2_n55 ;
    wire MixColumnsIns_MixOneColumnInst_2_n54 ;
    wire MixColumnsIns_MixOneColumnInst_2_n53 ;
    wire MixColumnsIns_MixOneColumnInst_2_n52 ;
    wire MixColumnsIns_MixOneColumnInst_2_n51 ;
    wire MixColumnsIns_MixOneColumnInst_2_n50 ;
    wire MixColumnsIns_MixOneColumnInst_2_n49 ;
    wire MixColumnsIns_MixOneColumnInst_2_n48 ;
    wire MixColumnsIns_MixOneColumnInst_2_n47 ;
    wire MixColumnsIns_MixOneColumnInst_2_n46 ;
    wire MixColumnsIns_MixOneColumnInst_2_n45 ;
    wire MixColumnsIns_MixOneColumnInst_2_n44 ;
    wire MixColumnsIns_MixOneColumnInst_2_n43 ;
    wire MixColumnsIns_MixOneColumnInst_2_n42 ;
    wire MixColumnsIns_MixOneColumnInst_2_n41 ;
    wire MixColumnsIns_MixOneColumnInst_2_n40 ;
    wire MixColumnsIns_MixOneColumnInst_2_n39 ;
    wire MixColumnsIns_MixOneColumnInst_2_n38 ;
    wire MixColumnsIns_MixOneColumnInst_2_n37 ;
    wire MixColumnsIns_MixOneColumnInst_2_n36 ;
    wire MixColumnsIns_MixOneColumnInst_2_n35 ;
    wire MixColumnsIns_MixOneColumnInst_2_n34 ;
    wire MixColumnsIns_MixOneColumnInst_2_n33 ;
    wire MixColumnsIns_MixOneColumnInst_2_n32 ;
    wire MixColumnsIns_MixOneColumnInst_2_n31 ;
    wire MixColumnsIns_MixOneColumnInst_2_n30 ;
    wire MixColumnsIns_MixOneColumnInst_2_n29 ;
    wire MixColumnsIns_MixOneColumnInst_2_n28 ;
    wire MixColumnsIns_MixOneColumnInst_2_n27 ;
    wire MixColumnsIns_MixOneColumnInst_2_n26 ;
    wire MixColumnsIns_MixOneColumnInst_2_n25 ;
    wire MixColumnsIns_MixOneColumnInst_2_n24 ;
    wire MixColumnsIns_MixOneColumnInst_2_n23 ;
    wire MixColumnsIns_MixOneColumnInst_2_n22 ;
    wire MixColumnsIns_MixOneColumnInst_2_n21 ;
    wire MixColumnsIns_MixOneColumnInst_2_n20 ;
    wire MixColumnsIns_MixOneColumnInst_2_n19 ;
    wire MixColumnsIns_MixOneColumnInst_2_n18 ;
    wire MixColumnsIns_MixOneColumnInst_2_n17 ;
    wire MixColumnsIns_MixOneColumnInst_2_n16 ;
    wire MixColumnsIns_MixOneColumnInst_2_n15 ;
    wire MixColumnsIns_MixOneColumnInst_2_n14 ;
    wire MixColumnsIns_MixOneColumnInst_2_n13 ;
    wire MixColumnsIns_MixOneColumnInst_2_n12 ;
    wire MixColumnsIns_MixOneColumnInst_2_n11 ;
    wire MixColumnsIns_MixOneColumnInst_2_n10 ;
    wire MixColumnsIns_MixOneColumnInst_2_n9 ;
    wire MixColumnsIns_MixOneColumnInst_2_n8 ;
    wire MixColumnsIns_MixOneColumnInst_2_n7 ;
    wire MixColumnsIns_MixOneColumnInst_2_n6 ;
    wire MixColumnsIns_MixOneColumnInst_2_n5 ;
    wire MixColumnsIns_MixOneColumnInst_2_n4 ;
    wire MixColumnsIns_MixOneColumnInst_2_n3 ;
    wire MixColumnsIns_MixOneColumnInst_2_n2 ;
    wire MixColumnsIns_MixOneColumnInst_2_n1 ;
    wire MixColumnsIns_MixOneColumnInst_3_n64 ;
    wire MixColumnsIns_MixOneColumnInst_3_n63 ;
    wire MixColumnsIns_MixOneColumnInst_3_n62 ;
    wire MixColumnsIns_MixOneColumnInst_3_n61 ;
    wire MixColumnsIns_MixOneColumnInst_3_n60 ;
    wire MixColumnsIns_MixOneColumnInst_3_n59 ;
    wire MixColumnsIns_MixOneColumnInst_3_n58 ;
    wire MixColumnsIns_MixOneColumnInst_3_n57 ;
    wire MixColumnsIns_MixOneColumnInst_3_n56 ;
    wire MixColumnsIns_MixOneColumnInst_3_n55 ;
    wire MixColumnsIns_MixOneColumnInst_3_n54 ;
    wire MixColumnsIns_MixOneColumnInst_3_n53 ;
    wire MixColumnsIns_MixOneColumnInst_3_n52 ;
    wire MixColumnsIns_MixOneColumnInst_3_n51 ;
    wire MixColumnsIns_MixOneColumnInst_3_n50 ;
    wire MixColumnsIns_MixOneColumnInst_3_n49 ;
    wire MixColumnsIns_MixOneColumnInst_3_n48 ;
    wire MixColumnsIns_MixOneColumnInst_3_n47 ;
    wire MixColumnsIns_MixOneColumnInst_3_n46 ;
    wire MixColumnsIns_MixOneColumnInst_3_n45 ;
    wire MixColumnsIns_MixOneColumnInst_3_n44 ;
    wire MixColumnsIns_MixOneColumnInst_3_n43 ;
    wire MixColumnsIns_MixOneColumnInst_3_n42 ;
    wire MixColumnsIns_MixOneColumnInst_3_n41 ;
    wire MixColumnsIns_MixOneColumnInst_3_n40 ;
    wire MixColumnsIns_MixOneColumnInst_3_n39 ;
    wire MixColumnsIns_MixOneColumnInst_3_n38 ;
    wire MixColumnsIns_MixOneColumnInst_3_n37 ;
    wire MixColumnsIns_MixOneColumnInst_3_n36 ;
    wire MixColumnsIns_MixOneColumnInst_3_n35 ;
    wire MixColumnsIns_MixOneColumnInst_3_n34 ;
    wire MixColumnsIns_MixOneColumnInst_3_n33 ;
    wire MixColumnsIns_MixOneColumnInst_3_n32 ;
    wire MixColumnsIns_MixOneColumnInst_3_n31 ;
    wire MixColumnsIns_MixOneColumnInst_3_n30 ;
    wire MixColumnsIns_MixOneColumnInst_3_n29 ;
    wire MixColumnsIns_MixOneColumnInst_3_n28 ;
    wire MixColumnsIns_MixOneColumnInst_3_n27 ;
    wire MixColumnsIns_MixOneColumnInst_3_n26 ;
    wire MixColumnsIns_MixOneColumnInst_3_n25 ;
    wire MixColumnsIns_MixOneColumnInst_3_n24 ;
    wire MixColumnsIns_MixOneColumnInst_3_n23 ;
    wire MixColumnsIns_MixOneColumnInst_3_n22 ;
    wire MixColumnsIns_MixOneColumnInst_3_n21 ;
    wire MixColumnsIns_MixOneColumnInst_3_n20 ;
    wire MixColumnsIns_MixOneColumnInst_3_n19 ;
    wire MixColumnsIns_MixOneColumnInst_3_n18 ;
    wire MixColumnsIns_MixOneColumnInst_3_n17 ;
    wire MixColumnsIns_MixOneColumnInst_3_n16 ;
    wire MixColumnsIns_MixOneColumnInst_3_n15 ;
    wire MixColumnsIns_MixOneColumnInst_3_n14 ;
    wire MixColumnsIns_MixOneColumnInst_3_n13 ;
    wire MixColumnsIns_MixOneColumnInst_3_n12 ;
    wire MixColumnsIns_MixOneColumnInst_3_n11 ;
    wire MixColumnsIns_MixOneColumnInst_3_n10 ;
    wire MixColumnsIns_MixOneColumnInst_3_n9 ;
    wire MixColumnsIns_MixOneColumnInst_3_n8 ;
    wire MixColumnsIns_MixOneColumnInst_3_n7 ;
    wire MixColumnsIns_MixOneColumnInst_3_n6 ;
    wire MixColumnsIns_MixOneColumnInst_3_n5 ;
    wire MixColumnsIns_MixOneColumnInst_3_n4 ;
    wire MixColumnsIns_MixOneColumnInst_3_n3 ;
    wire MixColumnsIns_MixOneColumnInst_3_n2 ;
    wire MixColumnsIns_MixOneColumnInst_3_n1 ;
    wire KeyReg_Inst_ff_SDE_0_next_state ;
    wire KeyReg_Inst_ff_SDE_1_next_state ;
    wire KeyReg_Inst_ff_SDE_2_next_state ;
    wire KeyReg_Inst_ff_SDE_3_next_state ;
    wire KeyReg_Inst_ff_SDE_4_next_state ;
    wire KeyReg_Inst_ff_SDE_5_next_state ;
    wire KeyReg_Inst_ff_SDE_6_next_state ;
    wire KeyReg_Inst_ff_SDE_7_next_state ;
    wire KeyReg_Inst_ff_SDE_8_next_state ;
    wire KeyReg_Inst_ff_SDE_9_next_state ;
    wire KeyReg_Inst_ff_SDE_10_next_state ;
    wire KeyReg_Inst_ff_SDE_11_next_state ;
    wire KeyReg_Inst_ff_SDE_12_next_state ;
    wire KeyReg_Inst_ff_SDE_13_next_state ;
    wire KeyReg_Inst_ff_SDE_14_next_state ;
    wire KeyReg_Inst_ff_SDE_15_next_state ;
    wire KeyReg_Inst_ff_SDE_16_next_state ;
    wire KeyReg_Inst_ff_SDE_17_next_state ;
    wire KeyReg_Inst_ff_SDE_18_next_state ;
    wire KeyReg_Inst_ff_SDE_19_next_state ;
    wire KeyReg_Inst_ff_SDE_20_next_state ;
    wire KeyReg_Inst_ff_SDE_21_next_state ;
    wire KeyReg_Inst_ff_SDE_22_next_state ;
    wire KeyReg_Inst_ff_SDE_23_next_state ;
    wire KeyReg_Inst_ff_SDE_24_next_state ;
    wire KeyReg_Inst_ff_SDE_25_next_state ;
    wire KeyReg_Inst_ff_SDE_26_next_state ;
    wire KeyReg_Inst_ff_SDE_27_next_state ;
    wire KeyReg_Inst_ff_SDE_28_next_state ;
    wire KeyReg_Inst_ff_SDE_29_next_state ;
    wire KeyReg_Inst_ff_SDE_30_next_state ;
    wire KeyReg_Inst_ff_SDE_31_next_state ;
    wire KeyReg_Inst_ff_SDE_32_next_state ;
    wire KeyReg_Inst_ff_SDE_33_next_state ;
    wire KeyReg_Inst_ff_SDE_34_next_state ;
    wire KeyReg_Inst_ff_SDE_35_next_state ;
    wire KeyReg_Inst_ff_SDE_36_next_state ;
    wire KeyReg_Inst_ff_SDE_37_next_state ;
    wire KeyReg_Inst_ff_SDE_38_next_state ;
    wire KeyReg_Inst_ff_SDE_39_next_state ;
    wire KeyReg_Inst_ff_SDE_40_next_state ;
    wire KeyReg_Inst_ff_SDE_41_next_state ;
    wire KeyReg_Inst_ff_SDE_42_next_state ;
    wire KeyReg_Inst_ff_SDE_43_next_state ;
    wire KeyReg_Inst_ff_SDE_44_next_state ;
    wire KeyReg_Inst_ff_SDE_45_next_state ;
    wire KeyReg_Inst_ff_SDE_46_next_state ;
    wire KeyReg_Inst_ff_SDE_47_next_state ;
    wire KeyReg_Inst_ff_SDE_48_next_state ;
    wire KeyReg_Inst_ff_SDE_49_next_state ;
    wire KeyReg_Inst_ff_SDE_50_next_state ;
    wire KeyReg_Inst_ff_SDE_51_next_state ;
    wire KeyReg_Inst_ff_SDE_52_next_state ;
    wire KeyReg_Inst_ff_SDE_53_next_state ;
    wire KeyReg_Inst_ff_SDE_54_next_state ;
    wire KeyReg_Inst_ff_SDE_55_next_state ;
    wire KeyReg_Inst_ff_SDE_56_next_state ;
    wire KeyReg_Inst_ff_SDE_57_next_state ;
    wire KeyReg_Inst_ff_SDE_58_next_state ;
    wire KeyReg_Inst_ff_SDE_59_next_state ;
    wire KeyReg_Inst_ff_SDE_60_next_state ;
    wire KeyReg_Inst_ff_SDE_61_next_state ;
    wire KeyReg_Inst_ff_SDE_62_next_state ;
    wire KeyReg_Inst_ff_SDE_63_next_state ;
    wire KeyReg_Inst_ff_SDE_64_next_state ;
    wire KeyReg_Inst_ff_SDE_65_next_state ;
    wire KeyReg_Inst_ff_SDE_66_next_state ;
    wire KeyReg_Inst_ff_SDE_67_next_state ;
    wire KeyReg_Inst_ff_SDE_68_next_state ;
    wire KeyReg_Inst_ff_SDE_69_next_state ;
    wire KeyReg_Inst_ff_SDE_70_next_state ;
    wire KeyReg_Inst_ff_SDE_71_next_state ;
    wire KeyReg_Inst_ff_SDE_72_next_state ;
    wire KeyReg_Inst_ff_SDE_73_next_state ;
    wire KeyReg_Inst_ff_SDE_74_next_state ;
    wire KeyReg_Inst_ff_SDE_75_next_state ;
    wire KeyReg_Inst_ff_SDE_76_next_state ;
    wire KeyReg_Inst_ff_SDE_77_next_state ;
    wire KeyReg_Inst_ff_SDE_78_next_state ;
    wire KeyReg_Inst_ff_SDE_79_next_state ;
    wire KeyReg_Inst_ff_SDE_80_next_state ;
    wire KeyReg_Inst_ff_SDE_81_next_state ;
    wire KeyReg_Inst_ff_SDE_82_next_state ;
    wire KeyReg_Inst_ff_SDE_83_next_state ;
    wire KeyReg_Inst_ff_SDE_84_next_state ;
    wire KeyReg_Inst_ff_SDE_85_next_state ;
    wire KeyReg_Inst_ff_SDE_86_next_state ;
    wire KeyReg_Inst_ff_SDE_87_next_state ;
    wire KeyReg_Inst_ff_SDE_88_next_state ;
    wire KeyReg_Inst_ff_SDE_89_next_state ;
    wire KeyReg_Inst_ff_SDE_90_next_state ;
    wire KeyReg_Inst_ff_SDE_91_next_state ;
    wire KeyReg_Inst_ff_SDE_92_next_state ;
    wire KeyReg_Inst_ff_SDE_93_next_state ;
    wire KeyReg_Inst_ff_SDE_94_next_state ;
    wire KeyReg_Inst_ff_SDE_95_next_state ;
    wire KeyReg_Inst_ff_SDE_96_next_state ;
    wire KeyReg_Inst_ff_SDE_97_next_state ;
    wire KeyReg_Inst_ff_SDE_98_next_state ;
    wire KeyReg_Inst_ff_SDE_99_next_state ;
    wire KeyReg_Inst_ff_SDE_100_next_state ;
    wire KeyReg_Inst_ff_SDE_101_next_state ;
    wire KeyReg_Inst_ff_SDE_102_next_state ;
    wire KeyReg_Inst_ff_SDE_103_next_state ;
    wire KeyReg_Inst_ff_SDE_104_next_state ;
    wire KeyReg_Inst_ff_SDE_105_next_state ;
    wire KeyReg_Inst_ff_SDE_106_next_state ;
    wire KeyReg_Inst_ff_SDE_107_next_state ;
    wire KeyReg_Inst_ff_SDE_108_next_state ;
    wire KeyReg_Inst_ff_SDE_109_next_state ;
    wire KeyReg_Inst_ff_SDE_110_next_state ;
    wire KeyReg_Inst_ff_SDE_111_next_state ;
    wire KeyReg_Inst_ff_SDE_112_next_state ;
    wire KeyReg_Inst_ff_SDE_113_next_state ;
    wire KeyReg_Inst_ff_SDE_114_next_state ;
    wire KeyReg_Inst_ff_SDE_115_next_state ;
    wire KeyReg_Inst_ff_SDE_116_next_state ;
    wire KeyReg_Inst_ff_SDE_117_next_state ;
    wire KeyReg_Inst_ff_SDE_118_next_state ;
    wire KeyReg_Inst_ff_SDE_119_next_state ;
    wire KeyReg_Inst_ff_SDE_120_next_state ;
    wire KeyReg_Inst_ff_SDE_121_next_state ;
    wire KeyReg_Inst_ff_SDE_122_next_state ;
    wire KeyReg_Inst_ff_SDE_123_next_state ;
    wire KeyReg_Inst_ff_SDE_124_next_state ;
    wire KeyReg_Inst_ff_SDE_125_next_state ;
    wire KeyReg_Inst_ff_SDE_126_next_state ;
    wire KeyReg_Inst_ff_SDE_127_next_state ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_ ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1 ;
    wire RoundCounterIns_n13 ;
    wire RoundCounterIns_n12 ;
    wire RoundCounterIns_n11 ;
    wire RoundCounterIns_n10 ;
    wire RoundCounterIns_n9 ;
    wire RoundCounterIns_n8 ;
    wire RoundCounterIns_n7 ;
    wire RoundCounterIns_n4 ;
    wire RoundCounterIns_n3 ;
    wire RoundCounterIns_n2 ;
    wire RoundCounterIns_n1 ;
    wire RoundCounterIns_N10 ;
    wire RoundCounterIns_n5 ;
    wire RoundCounterIns_N8 ;
    wire RoundCounterIns_n6 ;
    wire RoundCounterIns_N7 ;
    wire [127:0] RoundOutput ;
    wire [127:0] RoundInput ;
    wire [123:0] MixColumnsInput ;
    wire [127:0] MixColumnsOutput ;
    wire [127:0] KeyExpansionOutput ;
    wire [127:0] RoundKey ;
    wire [5:0] Rcon ;
    wire [3:0] RoundCounter ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_0_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_1_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_2_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_3_DoubleBytes ;
    wire [31:0] KeyExpansionIns_tmp ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5203 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5239 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6654 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;
    wire new_AGEMA_signal_6672 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6677 ;
    wire new_AGEMA_signal_6678 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6682 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6688 ;
    wire new_AGEMA_signal_6689 ;
    wire new_AGEMA_signal_6690 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6695 ;
    wire new_AGEMA_signal_6696 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6700 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6706 ;
    wire new_AGEMA_signal_6707 ;
    wire new_AGEMA_signal_6708 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6713 ;
    wire new_AGEMA_signal_6714 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6718 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6724 ;
    wire new_AGEMA_signal_6725 ;
    wire new_AGEMA_signal_6726 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7036 ;
    wire new_AGEMA_signal_7037 ;
    wire new_AGEMA_signal_7038 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7042 ;
    wire new_AGEMA_signal_7043 ;
    wire new_AGEMA_signal_7044 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7048 ;
    wire new_AGEMA_signal_7049 ;
    wire new_AGEMA_signal_7050 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7054 ;
    wire new_AGEMA_signal_7055 ;
    wire new_AGEMA_signal_7056 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7060 ;
    wire new_AGEMA_signal_7061 ;
    wire new_AGEMA_signal_7062 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7066 ;
    wire new_AGEMA_signal_7067 ;
    wire new_AGEMA_signal_7068 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7072 ;
    wire new_AGEMA_signal_7073 ;
    wire new_AGEMA_signal_7074 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7078 ;
    wire new_AGEMA_signal_7079 ;
    wire new_AGEMA_signal_7080 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7084 ;
    wire new_AGEMA_signal_7085 ;
    wire new_AGEMA_signal_7086 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7090 ;
    wire new_AGEMA_signal_7091 ;
    wire new_AGEMA_signal_7092 ;
    wire new_AGEMA_signal_7093 ;
    wire new_AGEMA_signal_7094 ;
    wire new_AGEMA_signal_7095 ;
    wire new_AGEMA_signal_7096 ;
    wire new_AGEMA_signal_7097 ;
    wire new_AGEMA_signal_7098 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7102 ;
    wire new_AGEMA_signal_7103 ;
    wire new_AGEMA_signal_7104 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7108 ;
    wire new_AGEMA_signal_7109 ;
    wire new_AGEMA_signal_7110 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7114 ;
    wire new_AGEMA_signal_7115 ;
    wire new_AGEMA_signal_7116 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7120 ;
    wire new_AGEMA_signal_7121 ;
    wire new_AGEMA_signal_7122 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7126 ;
    wire new_AGEMA_signal_7127 ;
    wire new_AGEMA_signal_7128 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7132 ;
    wire new_AGEMA_signal_7133 ;
    wire new_AGEMA_signal_7134 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7138 ;
    wire new_AGEMA_signal_7139 ;
    wire new_AGEMA_signal_7140 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7144 ;
    wire new_AGEMA_signal_7145 ;
    wire new_AGEMA_signal_7146 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7150 ;
    wire new_AGEMA_signal_7151 ;
    wire new_AGEMA_signal_7152 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7156 ;
    wire new_AGEMA_signal_7157 ;
    wire new_AGEMA_signal_7158 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7162 ;
    wire new_AGEMA_signal_7163 ;
    wire new_AGEMA_signal_7164 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7168 ;
    wire new_AGEMA_signal_7169 ;
    wire new_AGEMA_signal_7170 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7174 ;
    wire new_AGEMA_signal_7175 ;
    wire new_AGEMA_signal_7176 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7180 ;
    wire new_AGEMA_signal_7181 ;
    wire new_AGEMA_signal_7182 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7186 ;
    wire new_AGEMA_signal_7187 ;
    wire new_AGEMA_signal_7188 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7192 ;
    wire new_AGEMA_signal_7193 ;
    wire new_AGEMA_signal_7194 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7198 ;
    wire new_AGEMA_signal_7199 ;
    wire new_AGEMA_signal_7200 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7204 ;
    wire new_AGEMA_signal_7205 ;
    wire new_AGEMA_signal_7206 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7489 ;
    wire new_AGEMA_signal_7490 ;
    wire new_AGEMA_signal_7491 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7495 ;
    wire new_AGEMA_signal_7496 ;
    wire new_AGEMA_signal_7497 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7499 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7501 ;
    wire new_AGEMA_signal_7502 ;
    wire new_AGEMA_signal_7503 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7507 ;
    wire new_AGEMA_signal_7508 ;
    wire new_AGEMA_signal_7509 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7513 ;
    wire new_AGEMA_signal_7514 ;
    wire new_AGEMA_signal_7515 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7519 ;
    wire new_AGEMA_signal_7520 ;
    wire new_AGEMA_signal_7521 ;
    wire new_AGEMA_signal_7522 ;
    wire new_AGEMA_signal_7523 ;
    wire new_AGEMA_signal_7524 ;
    wire new_AGEMA_signal_7525 ;
    wire new_AGEMA_signal_7526 ;
    wire new_AGEMA_signal_7527 ;
    wire new_AGEMA_signal_7528 ;
    wire new_AGEMA_signal_7529 ;
    wire new_AGEMA_signal_7530 ;
    wire new_AGEMA_signal_7531 ;
    wire new_AGEMA_signal_7532 ;
    wire new_AGEMA_signal_7533 ;
    wire new_AGEMA_signal_7534 ;
    wire new_AGEMA_signal_7535 ;
    wire new_AGEMA_signal_7536 ;
    wire new_AGEMA_signal_7537 ;
    wire new_AGEMA_signal_7538 ;
    wire new_AGEMA_signal_7539 ;
    wire new_AGEMA_signal_7540 ;
    wire new_AGEMA_signal_7541 ;
    wire new_AGEMA_signal_7542 ;
    wire new_AGEMA_signal_7543 ;
    wire new_AGEMA_signal_7544 ;
    wire new_AGEMA_signal_7545 ;
    wire new_AGEMA_signal_7546 ;
    wire new_AGEMA_signal_7547 ;
    wire new_AGEMA_signal_7548 ;
    wire new_AGEMA_signal_7549 ;
    wire new_AGEMA_signal_7550 ;
    wire new_AGEMA_signal_7551 ;
    wire new_AGEMA_signal_7552 ;
    wire new_AGEMA_signal_7553 ;
    wire new_AGEMA_signal_7554 ;
    wire new_AGEMA_signal_7555 ;
    wire new_AGEMA_signal_7556 ;
    wire new_AGEMA_signal_7557 ;
    wire new_AGEMA_signal_7558 ;
    wire new_AGEMA_signal_7559 ;
    wire new_AGEMA_signal_7560 ;
    wire new_AGEMA_signal_7561 ;
    wire new_AGEMA_signal_7562 ;
    wire new_AGEMA_signal_7563 ;
    wire new_AGEMA_signal_7564 ;
    wire new_AGEMA_signal_7565 ;
    wire new_AGEMA_signal_7566 ;
    wire new_AGEMA_signal_7567 ;
    wire new_AGEMA_signal_7568 ;
    wire new_AGEMA_signal_7569 ;
    wire new_AGEMA_signal_7570 ;
    wire new_AGEMA_signal_7571 ;
    wire new_AGEMA_signal_7572 ;
    wire new_AGEMA_signal_7573 ;
    wire new_AGEMA_signal_7574 ;
    wire new_AGEMA_signal_7575 ;
    wire new_AGEMA_signal_7576 ;
    wire new_AGEMA_signal_7577 ;
    wire new_AGEMA_signal_7578 ;
    wire new_AGEMA_signal_7579 ;
    wire new_AGEMA_signal_7580 ;
    wire new_AGEMA_signal_7581 ;
    wire new_AGEMA_signal_7582 ;
    wire new_AGEMA_signal_7583 ;
    wire new_AGEMA_signal_7584 ;
    wire new_AGEMA_signal_7585 ;
    wire new_AGEMA_signal_7586 ;
    wire new_AGEMA_signal_7587 ;
    wire new_AGEMA_signal_7588 ;
    wire new_AGEMA_signal_7589 ;
    wire new_AGEMA_signal_7590 ;
    wire new_AGEMA_signal_7591 ;
    wire new_AGEMA_signal_7592 ;
    wire new_AGEMA_signal_7593 ;
    wire new_AGEMA_signal_7594 ;
    wire new_AGEMA_signal_7595 ;
    wire new_AGEMA_signal_7596 ;
    wire new_AGEMA_signal_7597 ;
    wire new_AGEMA_signal_7598 ;
    wire new_AGEMA_signal_7599 ;
    wire new_AGEMA_signal_7600 ;
    wire new_AGEMA_signal_7601 ;
    wire new_AGEMA_signal_7602 ;
    wire new_AGEMA_signal_7603 ;
    wire new_AGEMA_signal_7604 ;
    wire new_AGEMA_signal_7605 ;
    wire new_AGEMA_signal_7606 ;
    wire new_AGEMA_signal_7607 ;
    wire new_AGEMA_signal_7608 ;
    wire new_AGEMA_signal_7609 ;
    wire new_AGEMA_signal_7610 ;
    wire new_AGEMA_signal_7611 ;
    wire new_AGEMA_signal_7612 ;
    wire new_AGEMA_signal_7613 ;
    wire new_AGEMA_signal_7614 ;
    wire new_AGEMA_signal_7615 ;
    wire new_AGEMA_signal_7616 ;
    wire new_AGEMA_signal_7617 ;
    wire new_AGEMA_signal_7618 ;
    wire new_AGEMA_signal_7619 ;
    wire new_AGEMA_signal_7620 ;
    wire new_AGEMA_signal_7621 ;
    wire new_AGEMA_signal_7622 ;
    wire new_AGEMA_signal_7623 ;
    wire new_AGEMA_signal_7624 ;
    wire new_AGEMA_signal_7625 ;
    wire new_AGEMA_signal_7626 ;
    wire new_AGEMA_signal_7627 ;
    wire new_AGEMA_signal_7628 ;
    wire new_AGEMA_signal_7629 ;
    wire new_AGEMA_signal_7630 ;
    wire new_AGEMA_signal_7631 ;
    wire new_AGEMA_signal_7632 ;
    wire new_AGEMA_signal_7633 ;
    wire new_AGEMA_signal_7634 ;
    wire new_AGEMA_signal_7635 ;
    wire new_AGEMA_signal_7636 ;
    wire new_AGEMA_signal_7637 ;
    wire new_AGEMA_signal_7638 ;
    wire new_AGEMA_signal_7639 ;
    wire new_AGEMA_signal_7640 ;
    wire new_AGEMA_signal_7641 ;
    wire new_AGEMA_signal_7642 ;
    wire new_AGEMA_signal_7643 ;
    wire new_AGEMA_signal_7644 ;
    wire new_AGEMA_signal_7645 ;
    wire new_AGEMA_signal_7646 ;
    wire new_AGEMA_signal_7647 ;
    wire new_AGEMA_signal_7648 ;
    wire new_AGEMA_signal_7649 ;
    wire new_AGEMA_signal_7650 ;
    wire new_AGEMA_signal_7651 ;
    wire new_AGEMA_signal_7652 ;
    wire new_AGEMA_signal_7653 ;
    wire new_AGEMA_signal_7654 ;
    wire new_AGEMA_signal_7655 ;
    wire new_AGEMA_signal_7656 ;
    wire new_AGEMA_signal_7657 ;
    wire new_AGEMA_signal_7658 ;
    wire new_AGEMA_signal_7659 ;
    wire new_AGEMA_signal_7660 ;
    wire new_AGEMA_signal_7661 ;
    wire new_AGEMA_signal_7662 ;
    wire new_AGEMA_signal_7663 ;
    wire new_AGEMA_signal_7664 ;
    wire new_AGEMA_signal_7665 ;
    wire new_AGEMA_signal_7666 ;
    wire new_AGEMA_signal_7667 ;
    wire new_AGEMA_signal_7668 ;
    wire new_AGEMA_signal_7669 ;
    wire new_AGEMA_signal_7670 ;
    wire new_AGEMA_signal_7671 ;
    wire new_AGEMA_signal_7672 ;
    wire new_AGEMA_signal_7673 ;
    wire new_AGEMA_signal_7674 ;
    wire new_AGEMA_signal_7675 ;
    wire new_AGEMA_signal_7676 ;
    wire new_AGEMA_signal_7677 ;
    wire new_AGEMA_signal_7678 ;
    wire new_AGEMA_signal_7679 ;
    wire new_AGEMA_signal_7680 ;
    wire new_AGEMA_signal_7681 ;
    wire new_AGEMA_signal_7682 ;
    wire new_AGEMA_signal_7683 ;
    wire new_AGEMA_signal_7684 ;
    wire new_AGEMA_signal_7685 ;
    wire new_AGEMA_signal_7686 ;
    wire new_AGEMA_signal_7687 ;
    wire new_AGEMA_signal_7688 ;
    wire new_AGEMA_signal_7689 ;
    wire new_AGEMA_signal_7690 ;
    wire new_AGEMA_signal_7691 ;
    wire new_AGEMA_signal_7692 ;
    wire new_AGEMA_signal_7693 ;
    wire new_AGEMA_signal_7694 ;
    wire new_AGEMA_signal_7695 ;
    wire new_AGEMA_signal_7696 ;
    wire new_AGEMA_signal_7697 ;
    wire new_AGEMA_signal_7698 ;
    wire new_AGEMA_signal_7699 ;
    wire new_AGEMA_signal_7700 ;
    wire new_AGEMA_signal_7701 ;
    wire new_AGEMA_signal_7702 ;
    wire new_AGEMA_signal_7703 ;
    wire new_AGEMA_signal_7704 ;
    wire new_AGEMA_signal_7705 ;
    wire new_AGEMA_signal_7706 ;
    wire new_AGEMA_signal_7707 ;
    wire new_AGEMA_signal_7708 ;
    wire new_AGEMA_signal_7709 ;
    wire new_AGEMA_signal_7710 ;
    wire new_AGEMA_signal_7711 ;
    wire new_AGEMA_signal_7712 ;
    wire new_AGEMA_signal_7713 ;
    wire new_AGEMA_signal_7714 ;
    wire new_AGEMA_signal_7715 ;
    wire new_AGEMA_signal_7716 ;
    wire new_AGEMA_signal_7717 ;
    wire new_AGEMA_signal_7718 ;
    wire new_AGEMA_signal_7719 ;
    wire new_AGEMA_signal_7720 ;
    wire new_AGEMA_signal_7721 ;
    wire new_AGEMA_signal_7722 ;
    wire new_AGEMA_signal_7723 ;
    wire new_AGEMA_signal_7724 ;
    wire new_AGEMA_signal_7725 ;
    wire new_AGEMA_signal_7726 ;
    wire new_AGEMA_signal_7727 ;
    wire new_AGEMA_signal_7728 ;
    wire new_AGEMA_signal_7729 ;
    wire new_AGEMA_signal_7730 ;
    wire new_AGEMA_signal_7731 ;
    wire new_AGEMA_signal_7732 ;
    wire new_AGEMA_signal_7733 ;
    wire new_AGEMA_signal_7734 ;
    wire new_AGEMA_signal_7735 ;
    wire new_AGEMA_signal_7736 ;
    wire new_AGEMA_signal_7737 ;
    wire new_AGEMA_signal_7738 ;
    wire new_AGEMA_signal_7739 ;
    wire new_AGEMA_signal_7740 ;
    wire new_AGEMA_signal_7741 ;
    wire new_AGEMA_signal_7742 ;
    wire new_AGEMA_signal_7743 ;
    wire new_AGEMA_signal_7744 ;
    wire new_AGEMA_signal_7745 ;
    wire new_AGEMA_signal_7746 ;
    wire new_AGEMA_signal_7747 ;
    wire new_AGEMA_signal_7748 ;
    wire new_AGEMA_signal_7749 ;
    wire new_AGEMA_signal_7750 ;
    wire new_AGEMA_signal_7751 ;
    wire new_AGEMA_signal_7752 ;
    wire new_AGEMA_signal_7753 ;
    wire new_AGEMA_signal_7754 ;
    wire new_AGEMA_signal_7755 ;
    wire new_AGEMA_signal_7756 ;
    wire new_AGEMA_signal_7757 ;
    wire new_AGEMA_signal_7758 ;
    wire new_AGEMA_signal_7759 ;
    wire new_AGEMA_signal_7760 ;
    wire new_AGEMA_signal_7761 ;
    wire new_AGEMA_signal_7762 ;
    wire new_AGEMA_signal_7763 ;
    wire new_AGEMA_signal_7764 ;
    wire new_AGEMA_signal_7765 ;
    wire new_AGEMA_signal_7766 ;
    wire new_AGEMA_signal_7767 ;
    wire new_AGEMA_signal_7768 ;
    wire new_AGEMA_signal_7769 ;
    wire new_AGEMA_signal_7770 ;
    wire new_AGEMA_signal_7771 ;
    wire new_AGEMA_signal_7772 ;
    wire new_AGEMA_signal_7773 ;
    wire new_AGEMA_signal_7774 ;
    wire new_AGEMA_signal_7775 ;
    wire new_AGEMA_signal_7776 ;
    wire new_AGEMA_signal_7777 ;
    wire new_AGEMA_signal_7778 ;
    wire new_AGEMA_signal_7779 ;
    wire new_AGEMA_signal_7780 ;
    wire new_AGEMA_signal_7781 ;
    wire new_AGEMA_signal_7782 ;
    wire new_AGEMA_signal_7783 ;
    wire new_AGEMA_signal_7784 ;
    wire new_AGEMA_signal_7785 ;
    wire new_AGEMA_signal_7786 ;
    wire new_AGEMA_signal_7787 ;
    wire new_AGEMA_signal_7788 ;
    wire new_AGEMA_signal_7789 ;
    wire new_AGEMA_signal_7790 ;
    wire new_AGEMA_signal_7791 ;
    wire new_AGEMA_signal_7792 ;
    wire new_AGEMA_signal_7793 ;
    wire new_AGEMA_signal_7794 ;
    wire new_AGEMA_signal_7795 ;
    wire new_AGEMA_signal_7796 ;
    wire new_AGEMA_signal_7797 ;
    wire new_AGEMA_signal_7798 ;
    wire new_AGEMA_signal_7799 ;
    wire new_AGEMA_signal_7800 ;
    wire new_AGEMA_signal_7801 ;
    wire new_AGEMA_signal_7802 ;
    wire new_AGEMA_signal_7803 ;
    wire new_AGEMA_signal_7804 ;
    wire new_AGEMA_signal_7805 ;
    wire new_AGEMA_signal_7806 ;
    wire new_AGEMA_signal_7807 ;
    wire new_AGEMA_signal_7808 ;
    wire new_AGEMA_signal_7809 ;
    wire new_AGEMA_signal_7810 ;
    wire new_AGEMA_signal_7811 ;
    wire new_AGEMA_signal_7812 ;
    wire new_AGEMA_signal_7813 ;
    wire new_AGEMA_signal_7814 ;
    wire new_AGEMA_signal_7815 ;
    wire new_AGEMA_signal_7816 ;
    wire new_AGEMA_signal_7817 ;
    wire new_AGEMA_signal_7818 ;
    wire new_AGEMA_signal_7819 ;
    wire new_AGEMA_signal_7820 ;
    wire new_AGEMA_signal_7821 ;
    wire new_AGEMA_signal_7822 ;
    wire new_AGEMA_signal_7823 ;
    wire new_AGEMA_signal_7824 ;
    wire new_AGEMA_signal_7825 ;
    wire new_AGEMA_signal_7826 ;
    wire new_AGEMA_signal_7827 ;
    wire new_AGEMA_signal_7828 ;
    wire new_AGEMA_signal_7829 ;
    wire new_AGEMA_signal_7830 ;
    wire new_AGEMA_signal_7831 ;
    wire new_AGEMA_signal_7832 ;
    wire new_AGEMA_signal_7833 ;
    wire new_AGEMA_signal_7834 ;
    wire new_AGEMA_signal_7835 ;
    wire new_AGEMA_signal_7836 ;
    wire new_AGEMA_signal_7837 ;
    wire new_AGEMA_signal_7838 ;
    wire new_AGEMA_signal_7839 ;
    wire new_AGEMA_signal_7840 ;
    wire new_AGEMA_signal_7841 ;
    wire new_AGEMA_signal_7842 ;
    wire new_AGEMA_signal_7843 ;
    wire new_AGEMA_signal_7844 ;
    wire new_AGEMA_signal_7845 ;
    wire new_AGEMA_signal_7846 ;
    wire new_AGEMA_signal_7847 ;
    wire new_AGEMA_signal_7848 ;
    wire new_AGEMA_signal_7849 ;
    wire new_AGEMA_signal_7850 ;
    wire new_AGEMA_signal_7851 ;
    wire new_AGEMA_signal_7852 ;
    wire new_AGEMA_signal_7853 ;
    wire new_AGEMA_signal_7854 ;
    wire new_AGEMA_signal_7855 ;
    wire new_AGEMA_signal_7856 ;
    wire new_AGEMA_signal_7857 ;
    wire new_AGEMA_signal_7858 ;
    wire new_AGEMA_signal_7859 ;
    wire new_AGEMA_signal_7860 ;
    wire new_AGEMA_signal_7861 ;
    wire new_AGEMA_signal_7862 ;
    wire new_AGEMA_signal_7863 ;
    wire new_AGEMA_signal_7864 ;
    wire new_AGEMA_signal_7865 ;
    wire new_AGEMA_signal_7866 ;
    wire new_AGEMA_signal_7867 ;
    wire new_AGEMA_signal_7868 ;
    wire new_AGEMA_signal_7869 ;
    wire new_AGEMA_signal_7870 ;
    wire new_AGEMA_signal_7871 ;
    wire new_AGEMA_signal_7872 ;
    wire new_AGEMA_signal_7873 ;
    wire new_AGEMA_signal_7874 ;
    wire new_AGEMA_signal_7875 ;
    wire new_AGEMA_signal_7876 ;
    wire new_AGEMA_signal_7877 ;
    wire new_AGEMA_signal_7878 ;
    wire new_AGEMA_signal_7879 ;
    wire new_AGEMA_signal_7880 ;
    wire new_AGEMA_signal_7881 ;
    wire new_AGEMA_signal_7882 ;
    wire new_AGEMA_signal_7883 ;
    wire new_AGEMA_signal_7884 ;
    wire new_AGEMA_signal_7885 ;
    wire new_AGEMA_signal_7886 ;
    wire new_AGEMA_signal_7887 ;
    wire new_AGEMA_signal_7888 ;
    wire new_AGEMA_signal_7889 ;
    wire new_AGEMA_signal_7890 ;
    wire new_AGEMA_signal_7891 ;
    wire new_AGEMA_signal_7892 ;
    wire new_AGEMA_signal_7893 ;
    wire new_AGEMA_signal_7894 ;
    wire new_AGEMA_signal_7895 ;
    wire new_AGEMA_signal_7896 ;
    wire new_AGEMA_signal_7897 ;
    wire new_AGEMA_signal_7898 ;
    wire new_AGEMA_signal_7899 ;
    wire new_AGEMA_signal_7900 ;
    wire new_AGEMA_signal_7901 ;
    wire new_AGEMA_signal_7902 ;
    wire new_AGEMA_signal_7903 ;
    wire new_AGEMA_signal_7904 ;
    wire new_AGEMA_signal_7905 ;
    wire new_AGEMA_signal_7906 ;
    wire new_AGEMA_signal_7907 ;
    wire new_AGEMA_signal_7908 ;
    wire new_AGEMA_signal_7909 ;
    wire new_AGEMA_signal_7910 ;
    wire new_AGEMA_signal_7911 ;
    wire new_AGEMA_signal_7912 ;
    wire new_AGEMA_signal_7913 ;
    wire new_AGEMA_signal_7914 ;
    wire new_AGEMA_signal_7915 ;
    wire new_AGEMA_signal_7916 ;
    wire new_AGEMA_signal_7917 ;
    wire new_AGEMA_signal_7918 ;
    wire new_AGEMA_signal_7919 ;
    wire new_AGEMA_signal_7920 ;
    wire new_AGEMA_signal_7921 ;
    wire new_AGEMA_signal_7922 ;
    wire new_AGEMA_signal_7923 ;
    wire new_AGEMA_signal_7924 ;
    wire new_AGEMA_signal_7925 ;
    wire new_AGEMA_signal_7926 ;
    wire new_AGEMA_signal_7927 ;
    wire new_AGEMA_signal_7928 ;
    wire new_AGEMA_signal_7929 ;
    wire new_AGEMA_signal_7930 ;
    wire new_AGEMA_signal_7931 ;
    wire new_AGEMA_signal_7932 ;
    wire new_AGEMA_signal_7933 ;
    wire new_AGEMA_signal_7934 ;
    wire new_AGEMA_signal_7935 ;
    wire new_AGEMA_signal_7936 ;
    wire new_AGEMA_signal_7937 ;
    wire new_AGEMA_signal_7938 ;
    wire new_AGEMA_signal_7939 ;
    wire new_AGEMA_signal_7940 ;
    wire new_AGEMA_signal_7941 ;
    wire new_AGEMA_signal_7942 ;
    wire new_AGEMA_signal_7943 ;
    wire new_AGEMA_signal_7944 ;
    wire new_AGEMA_signal_7945 ;
    wire new_AGEMA_signal_7946 ;
    wire new_AGEMA_signal_7947 ;
    wire new_AGEMA_signal_7948 ;
    wire new_AGEMA_signal_7949 ;
    wire new_AGEMA_signal_7950 ;
    wire new_AGEMA_signal_7951 ;
    wire new_AGEMA_signal_7952 ;
    wire new_AGEMA_signal_7953 ;
    wire new_AGEMA_signal_7954 ;
    wire new_AGEMA_signal_7955 ;
    wire new_AGEMA_signal_7956 ;
    wire new_AGEMA_signal_7957 ;
    wire new_AGEMA_signal_7958 ;
    wire new_AGEMA_signal_7959 ;
    wire new_AGEMA_signal_7960 ;
    wire new_AGEMA_signal_7961 ;
    wire new_AGEMA_signal_7962 ;
    wire new_AGEMA_signal_7963 ;
    wire new_AGEMA_signal_7964 ;
    wire new_AGEMA_signal_7965 ;
    wire new_AGEMA_signal_7966 ;
    wire new_AGEMA_signal_7967 ;
    wire new_AGEMA_signal_7968 ;
    wire new_AGEMA_signal_7969 ;
    wire new_AGEMA_signal_7970 ;
    wire new_AGEMA_signal_7971 ;
    wire new_AGEMA_signal_7972 ;
    wire new_AGEMA_signal_7973 ;
    wire new_AGEMA_signal_7974 ;
    wire new_AGEMA_signal_7975 ;
    wire new_AGEMA_signal_7976 ;
    wire new_AGEMA_signal_7977 ;
    wire new_AGEMA_signal_7978 ;
    wire new_AGEMA_signal_7979 ;
    wire new_AGEMA_signal_7980 ;
    wire new_AGEMA_signal_7981 ;
    wire new_AGEMA_signal_7982 ;
    wire new_AGEMA_signal_7983 ;
    wire new_AGEMA_signal_7984 ;
    wire new_AGEMA_signal_7985 ;
    wire new_AGEMA_signal_7986 ;
    wire new_AGEMA_signal_7987 ;
    wire new_AGEMA_signal_7988 ;
    wire new_AGEMA_signal_7989 ;
    wire new_AGEMA_signal_7990 ;
    wire new_AGEMA_signal_7991 ;
    wire new_AGEMA_signal_7992 ;
    wire new_AGEMA_signal_7993 ;
    wire new_AGEMA_signal_7994 ;
    wire new_AGEMA_signal_7995 ;
    wire new_AGEMA_signal_7996 ;
    wire new_AGEMA_signal_7997 ;
    wire new_AGEMA_signal_7998 ;
    wire new_AGEMA_signal_7999 ;
    wire new_AGEMA_signal_8000 ;
    wire new_AGEMA_signal_8001 ;
    wire new_AGEMA_signal_8002 ;
    wire new_AGEMA_signal_8003 ;
    wire new_AGEMA_signal_8004 ;
    wire new_AGEMA_signal_8005 ;
    wire new_AGEMA_signal_8006 ;
    wire new_AGEMA_signal_8007 ;
    wire new_AGEMA_signal_8008 ;
    wire new_AGEMA_signal_8009 ;
    wire new_AGEMA_signal_8010 ;
    wire new_AGEMA_signal_8011 ;
    wire new_AGEMA_signal_8012 ;
    wire new_AGEMA_signal_8013 ;
    wire new_AGEMA_signal_8014 ;
    wire new_AGEMA_signal_8015 ;
    wire new_AGEMA_signal_8016 ;
    wire new_AGEMA_signal_8017 ;
    wire new_AGEMA_signal_8018 ;
    wire new_AGEMA_signal_8019 ;
    wire new_AGEMA_signal_8020 ;
    wire new_AGEMA_signal_8021 ;
    wire new_AGEMA_signal_8022 ;
    wire new_AGEMA_signal_8023 ;
    wire new_AGEMA_signal_8024 ;
    wire new_AGEMA_signal_8025 ;
    wire new_AGEMA_signal_8026 ;
    wire new_AGEMA_signal_8027 ;
    wire new_AGEMA_signal_8028 ;
    wire new_AGEMA_signal_8029 ;
    wire new_AGEMA_signal_8030 ;
    wire new_AGEMA_signal_8031 ;
    wire new_AGEMA_signal_8032 ;
    wire new_AGEMA_signal_8033 ;
    wire new_AGEMA_signal_8034 ;
    wire new_AGEMA_signal_8035 ;
    wire new_AGEMA_signal_8036 ;
    wire new_AGEMA_signal_8037 ;
    wire new_AGEMA_signal_8038 ;
    wire new_AGEMA_signal_8039 ;
    wire new_AGEMA_signal_8040 ;
    wire new_AGEMA_signal_8041 ;
    wire new_AGEMA_signal_8042 ;
    wire new_AGEMA_signal_8043 ;
    wire new_AGEMA_signal_8044 ;
    wire new_AGEMA_signal_8045 ;
    wire new_AGEMA_signal_8046 ;
    wire new_AGEMA_signal_8047 ;
    wire new_AGEMA_signal_8048 ;
    wire new_AGEMA_signal_8049 ;
    wire new_AGEMA_signal_8050 ;
    wire new_AGEMA_signal_8051 ;
    wire new_AGEMA_signal_8052 ;
    wire new_AGEMA_signal_8053 ;
    wire new_AGEMA_signal_8054 ;
    wire new_AGEMA_signal_8055 ;
    wire new_AGEMA_signal_8056 ;
    wire new_AGEMA_signal_8057 ;
    wire new_AGEMA_signal_8058 ;
    wire new_AGEMA_signal_8059 ;
    wire new_AGEMA_signal_8060 ;
    wire new_AGEMA_signal_8061 ;
    wire new_AGEMA_signal_8062 ;
    wire new_AGEMA_signal_8063 ;
    wire new_AGEMA_signal_8064 ;
    wire new_AGEMA_signal_8065 ;
    wire new_AGEMA_signal_8066 ;
    wire new_AGEMA_signal_8067 ;
    wire new_AGEMA_signal_8068 ;
    wire new_AGEMA_signal_8069 ;
    wire new_AGEMA_signal_8070 ;
    wire new_AGEMA_signal_8071 ;
    wire new_AGEMA_signal_8072 ;
    wire new_AGEMA_signal_8073 ;
    wire new_AGEMA_signal_8074 ;
    wire new_AGEMA_signal_8075 ;
    wire new_AGEMA_signal_8076 ;
    wire new_AGEMA_signal_8077 ;
    wire new_AGEMA_signal_8078 ;
    wire new_AGEMA_signal_8079 ;
    wire new_AGEMA_signal_8080 ;
    wire new_AGEMA_signal_8081 ;
    wire new_AGEMA_signal_8082 ;
    wire new_AGEMA_signal_8083 ;
    wire new_AGEMA_signal_8084 ;
    wire new_AGEMA_signal_8085 ;
    wire new_AGEMA_signal_8086 ;
    wire new_AGEMA_signal_8087 ;
    wire new_AGEMA_signal_8088 ;
    wire new_AGEMA_signal_8089 ;
    wire new_AGEMA_signal_8090 ;
    wire new_AGEMA_signal_8091 ;
    wire new_AGEMA_signal_8092 ;
    wire new_AGEMA_signal_8093 ;
    wire new_AGEMA_signal_8094 ;
    wire new_AGEMA_signal_8095 ;
    wire new_AGEMA_signal_8096 ;
    wire new_AGEMA_signal_8097 ;
    wire new_AGEMA_signal_8098 ;
    wire new_AGEMA_signal_8099 ;
    wire new_AGEMA_signal_8100 ;
    wire new_AGEMA_signal_8101 ;
    wire new_AGEMA_signal_8102 ;
    wire new_AGEMA_signal_8103 ;
    wire new_AGEMA_signal_8104 ;
    wire new_AGEMA_signal_8105 ;
    wire new_AGEMA_signal_8106 ;
    wire new_AGEMA_signal_8107 ;
    wire new_AGEMA_signal_8108 ;
    wire new_AGEMA_signal_8109 ;
    wire new_AGEMA_signal_8110 ;
    wire new_AGEMA_signal_8111 ;
    wire new_AGEMA_signal_8112 ;
    wire new_AGEMA_signal_8113 ;
    wire new_AGEMA_signal_8114 ;
    wire new_AGEMA_signal_8115 ;
    wire new_AGEMA_signal_8116 ;
    wire new_AGEMA_signal_8117 ;
    wire new_AGEMA_signal_8118 ;
    wire new_AGEMA_signal_8119 ;
    wire new_AGEMA_signal_8120 ;
    wire new_AGEMA_signal_8121 ;
    wire new_AGEMA_signal_8122 ;
    wire new_AGEMA_signal_8123 ;
    wire new_AGEMA_signal_8124 ;
    wire new_AGEMA_signal_8125 ;
    wire new_AGEMA_signal_8126 ;
    wire new_AGEMA_signal_8127 ;
    wire new_AGEMA_signal_8128 ;
    wire new_AGEMA_signal_8129 ;
    wire new_AGEMA_signal_8130 ;
    wire new_AGEMA_signal_8131 ;
    wire new_AGEMA_signal_8132 ;
    wire new_AGEMA_signal_8133 ;
    wire new_AGEMA_signal_8134 ;
    wire new_AGEMA_signal_8135 ;
    wire new_AGEMA_signal_8136 ;
    wire new_AGEMA_signal_8137 ;
    wire new_AGEMA_signal_8138 ;
    wire new_AGEMA_signal_8139 ;
    wire new_AGEMA_signal_8140 ;
    wire new_AGEMA_signal_8141 ;
    wire new_AGEMA_signal_8142 ;
    wire new_AGEMA_signal_8143 ;
    wire new_AGEMA_signal_8144 ;
    wire new_AGEMA_signal_8145 ;
    wire new_AGEMA_signal_8146 ;
    wire new_AGEMA_signal_8147 ;
    wire new_AGEMA_signal_8148 ;
    wire new_AGEMA_signal_8149 ;
    wire new_AGEMA_signal_8150 ;
    wire new_AGEMA_signal_8151 ;
    wire new_AGEMA_signal_8152 ;
    wire new_AGEMA_signal_8153 ;
    wire new_AGEMA_signal_8154 ;
    wire new_AGEMA_signal_8155 ;
    wire new_AGEMA_signal_8156 ;
    wire new_AGEMA_signal_8157 ;
    wire new_AGEMA_signal_8158 ;
    wire new_AGEMA_signal_8159 ;
    wire new_AGEMA_signal_8160 ;
    wire new_AGEMA_signal_8161 ;
    wire new_AGEMA_signal_8162 ;
    wire new_AGEMA_signal_8163 ;
    wire new_AGEMA_signal_8164 ;
    wire new_AGEMA_signal_8165 ;
    wire new_AGEMA_signal_8166 ;
    wire new_AGEMA_signal_8167 ;
    wire new_AGEMA_signal_8168 ;
    wire new_AGEMA_signal_8169 ;
    wire new_AGEMA_signal_8170 ;
    wire new_AGEMA_signal_8171 ;
    wire new_AGEMA_signal_8172 ;
    wire new_AGEMA_signal_8173 ;
    wire new_AGEMA_signal_8174 ;
    wire new_AGEMA_signal_8175 ;
    wire new_AGEMA_signal_8176 ;
    wire new_AGEMA_signal_8177 ;
    wire new_AGEMA_signal_8178 ;
    wire new_AGEMA_signal_8179 ;
    wire new_AGEMA_signal_8180 ;
    wire new_AGEMA_signal_8181 ;
    wire new_AGEMA_signal_8182 ;
    wire new_AGEMA_signal_8183 ;
    wire new_AGEMA_signal_8184 ;
    wire new_AGEMA_signal_8185 ;
    wire new_AGEMA_signal_8186 ;
    wire new_AGEMA_signal_8187 ;
    wire new_AGEMA_signal_8188 ;
    wire new_AGEMA_signal_8189 ;
    wire new_AGEMA_signal_8190 ;
    wire new_AGEMA_signal_8191 ;
    wire new_AGEMA_signal_8192 ;
    wire new_AGEMA_signal_8193 ;
    wire new_AGEMA_signal_8194 ;
    wire new_AGEMA_signal_8195 ;
    wire new_AGEMA_signal_8196 ;
    wire new_AGEMA_signal_8197 ;
    wire new_AGEMA_signal_8198 ;
    wire new_AGEMA_signal_8199 ;
    wire new_AGEMA_signal_8200 ;
    wire new_AGEMA_signal_8201 ;
    wire new_AGEMA_signal_8202 ;
    wire new_AGEMA_signal_8203 ;
    wire new_AGEMA_signal_8204 ;
    wire new_AGEMA_signal_8205 ;
    wire new_AGEMA_signal_8206 ;
    wire new_AGEMA_signal_8207 ;
    wire new_AGEMA_signal_8208 ;
    wire new_AGEMA_signal_8209 ;
    wire new_AGEMA_signal_8210 ;
    wire new_AGEMA_signal_8211 ;
    wire new_AGEMA_signal_8212 ;
    wire new_AGEMA_signal_8213 ;
    wire new_AGEMA_signal_8214 ;
    wire new_AGEMA_signal_8215 ;
    wire new_AGEMA_signal_8216 ;
    wire new_AGEMA_signal_8217 ;
    wire new_AGEMA_signal_8218 ;
    wire new_AGEMA_signal_8219 ;
    wire new_AGEMA_signal_8220 ;
    wire new_AGEMA_signal_8221 ;
    wire new_AGEMA_signal_8222 ;
    wire new_AGEMA_signal_8223 ;
    wire new_AGEMA_signal_8224 ;
    wire new_AGEMA_signal_8225 ;
    wire new_AGEMA_signal_8226 ;
    wire new_AGEMA_signal_8227 ;
    wire new_AGEMA_signal_8228 ;
    wire new_AGEMA_signal_8229 ;
    wire new_AGEMA_signal_8230 ;
    wire new_AGEMA_signal_8231 ;
    wire new_AGEMA_signal_8232 ;
    wire new_AGEMA_signal_8233 ;
    wire new_AGEMA_signal_8234 ;
    wire new_AGEMA_signal_8235 ;
    wire new_AGEMA_signal_8236 ;
    wire new_AGEMA_signal_8237 ;
    wire new_AGEMA_signal_8238 ;
    wire new_AGEMA_signal_8239 ;
    wire new_AGEMA_signal_8240 ;
    wire new_AGEMA_signal_8241 ;
    wire new_AGEMA_signal_8242 ;
    wire new_AGEMA_signal_8243 ;
    wire new_AGEMA_signal_8244 ;
    wire new_AGEMA_signal_8245 ;
    wire new_AGEMA_signal_8246 ;
    wire new_AGEMA_signal_8247 ;
    wire new_AGEMA_signal_8248 ;
    wire new_AGEMA_signal_8249 ;
    wire new_AGEMA_signal_8250 ;
    wire new_AGEMA_signal_8251 ;
    wire new_AGEMA_signal_8252 ;
    wire new_AGEMA_signal_8253 ;
    wire new_AGEMA_signal_8254 ;
    wire new_AGEMA_signal_8255 ;
    wire new_AGEMA_signal_8256 ;
    wire new_AGEMA_signal_8257 ;
    wire new_AGEMA_signal_8258 ;
    wire new_AGEMA_signal_8259 ;
    wire new_AGEMA_signal_8260 ;
    wire new_AGEMA_signal_8261 ;
    wire new_AGEMA_signal_8262 ;
    wire new_AGEMA_signal_8263 ;
    wire new_AGEMA_signal_8264 ;
    wire new_AGEMA_signal_8265 ;
    wire new_AGEMA_signal_8266 ;
    wire new_AGEMA_signal_8267 ;
    wire new_AGEMA_signal_8268 ;
    wire new_AGEMA_signal_8269 ;
    wire new_AGEMA_signal_8270 ;
    wire new_AGEMA_signal_8271 ;
    wire new_AGEMA_signal_8272 ;
    wire new_AGEMA_signal_8273 ;
    wire new_AGEMA_signal_8274 ;
    wire new_AGEMA_signal_8275 ;
    wire new_AGEMA_signal_8276 ;
    wire new_AGEMA_signal_8277 ;
    wire new_AGEMA_signal_8278 ;
    wire new_AGEMA_signal_8279 ;
    wire new_AGEMA_signal_8280 ;
    wire new_AGEMA_signal_8281 ;
    wire new_AGEMA_signal_8282 ;
    wire new_AGEMA_signal_8283 ;
    wire new_AGEMA_signal_8284 ;
    wire new_AGEMA_signal_8285 ;
    wire new_AGEMA_signal_8286 ;
    wire new_AGEMA_signal_8287 ;
    wire new_AGEMA_signal_8288 ;
    wire new_AGEMA_signal_8289 ;
    wire new_AGEMA_signal_8290 ;
    wire new_AGEMA_signal_8291 ;
    wire new_AGEMA_signal_8292 ;
    wire new_AGEMA_signal_8293 ;
    wire new_AGEMA_signal_8294 ;
    wire new_AGEMA_signal_8295 ;
    wire new_AGEMA_signal_8296 ;
    wire new_AGEMA_signal_8297 ;
    wire new_AGEMA_signal_8298 ;
    wire new_AGEMA_signal_8299 ;
    wire new_AGEMA_signal_8300 ;
    wire new_AGEMA_signal_8301 ;
    wire new_AGEMA_signal_8302 ;
    wire new_AGEMA_signal_8303 ;
    wire new_AGEMA_signal_8304 ;
    wire new_AGEMA_signal_8305 ;
    wire new_AGEMA_signal_8306 ;
    wire new_AGEMA_signal_8307 ;
    wire new_AGEMA_signal_8308 ;
    wire new_AGEMA_signal_8309 ;
    wire new_AGEMA_signal_8310 ;
    wire new_AGEMA_signal_8311 ;
    wire new_AGEMA_signal_8312 ;
    wire new_AGEMA_signal_8313 ;
    wire new_AGEMA_signal_8314 ;
    wire new_AGEMA_signal_8315 ;
    wire new_AGEMA_signal_8316 ;
    wire new_AGEMA_signal_8317 ;
    wire new_AGEMA_signal_8318 ;
    wire new_AGEMA_signal_8319 ;
    wire new_AGEMA_signal_8320 ;
    wire new_AGEMA_signal_8321 ;
    wire new_AGEMA_signal_8322 ;
    wire new_AGEMA_signal_8323 ;
    wire new_AGEMA_signal_8324 ;
    wire new_AGEMA_signal_8325 ;
    wire new_AGEMA_signal_8326 ;
    wire new_AGEMA_signal_8327 ;
    wire new_AGEMA_signal_8328 ;
    wire new_AGEMA_signal_8329 ;
    wire new_AGEMA_signal_8330 ;
    wire new_AGEMA_signal_8331 ;
    wire new_AGEMA_signal_8332 ;
    wire new_AGEMA_signal_8333 ;
    wire new_AGEMA_signal_8334 ;
    wire new_AGEMA_signal_8335 ;
    wire new_AGEMA_signal_8336 ;
    wire new_AGEMA_signal_8337 ;
    wire new_AGEMA_signal_8338 ;
    wire new_AGEMA_signal_8339 ;
    wire new_AGEMA_signal_8340 ;
    wire new_AGEMA_signal_8341 ;
    wire new_AGEMA_signal_8342 ;
    wire new_AGEMA_signal_8343 ;
    wire new_AGEMA_signal_8344 ;
    wire new_AGEMA_signal_8345 ;
    wire new_AGEMA_signal_8346 ;
    wire new_AGEMA_signal_8347 ;
    wire new_AGEMA_signal_8348 ;
    wire new_AGEMA_signal_8349 ;
    wire new_AGEMA_signal_8350 ;
    wire new_AGEMA_signal_8351 ;
    wire new_AGEMA_signal_8352 ;
    wire new_AGEMA_signal_8353 ;
    wire new_AGEMA_signal_8354 ;
    wire new_AGEMA_signal_8355 ;
    wire new_AGEMA_signal_8356 ;
    wire new_AGEMA_signal_8357 ;
    wire new_AGEMA_signal_8358 ;
    wire new_AGEMA_signal_8359 ;
    wire new_AGEMA_signal_8360 ;
    wire new_AGEMA_signal_8361 ;
    wire new_AGEMA_signal_8362 ;
    wire new_AGEMA_signal_8363 ;
    wire new_AGEMA_signal_8364 ;
    wire new_AGEMA_signal_8365 ;
    wire new_AGEMA_signal_8366 ;
    wire new_AGEMA_signal_8367 ;
    wire new_AGEMA_signal_8368 ;
    wire new_AGEMA_signal_8369 ;
    wire new_AGEMA_signal_8370 ;
    wire new_AGEMA_signal_8371 ;
    wire new_AGEMA_signal_8372 ;
    wire new_AGEMA_signal_8373 ;
    wire new_AGEMA_signal_8374 ;
    wire new_AGEMA_signal_8375 ;
    wire new_AGEMA_signal_8376 ;
    wire new_AGEMA_signal_8377 ;
    wire new_AGEMA_signal_8378 ;
    wire new_AGEMA_signal_8379 ;
    wire new_AGEMA_signal_8380 ;
    wire new_AGEMA_signal_8381 ;
    wire new_AGEMA_signal_8382 ;
    wire new_AGEMA_signal_8383 ;
    wire new_AGEMA_signal_8384 ;
    wire new_AGEMA_signal_8385 ;
    wire new_AGEMA_signal_8386 ;
    wire new_AGEMA_signal_8387 ;
    wire new_AGEMA_signal_8388 ;
    wire new_AGEMA_signal_8389 ;
    wire new_AGEMA_signal_8390 ;
    wire new_AGEMA_signal_8391 ;
    wire new_AGEMA_signal_8392 ;
    wire new_AGEMA_signal_8393 ;
    wire new_AGEMA_signal_8394 ;
    wire new_AGEMA_signal_8395 ;
    wire new_AGEMA_signal_8396 ;
    wire new_AGEMA_signal_8397 ;
    wire new_AGEMA_signal_8398 ;
    wire new_AGEMA_signal_8399 ;
    wire new_AGEMA_signal_8400 ;
    wire new_AGEMA_signal_8401 ;
    wire new_AGEMA_signal_8402 ;
    wire new_AGEMA_signal_8403 ;
    wire new_AGEMA_signal_8404 ;
    wire new_AGEMA_signal_8405 ;
    wire new_AGEMA_signal_8406 ;
    wire new_AGEMA_signal_8407 ;
    wire new_AGEMA_signal_8408 ;
    wire new_AGEMA_signal_8409 ;
    wire new_AGEMA_signal_8410 ;
    wire new_AGEMA_signal_8411 ;
    wire new_AGEMA_signal_8412 ;
    wire new_AGEMA_signal_8413 ;
    wire new_AGEMA_signal_8414 ;
    wire new_AGEMA_signal_8415 ;
    wire new_AGEMA_signal_8416 ;
    wire new_AGEMA_signal_8417 ;
    wire new_AGEMA_signal_8418 ;
    wire new_AGEMA_signal_8419 ;
    wire new_AGEMA_signal_8420 ;
    wire new_AGEMA_signal_8421 ;
    wire new_AGEMA_signal_8422 ;
    wire new_AGEMA_signal_8423 ;
    wire new_AGEMA_signal_8424 ;
    wire new_AGEMA_signal_8425 ;
    wire new_AGEMA_signal_8426 ;
    wire new_AGEMA_signal_8427 ;
    wire new_AGEMA_signal_8428 ;
    wire new_AGEMA_signal_8429 ;
    wire new_AGEMA_signal_8430 ;
    wire new_AGEMA_signal_8431 ;
    wire new_AGEMA_signal_8432 ;
    wire new_AGEMA_signal_8433 ;
    wire new_AGEMA_signal_8434 ;
    wire new_AGEMA_signal_8435 ;
    wire new_AGEMA_signal_8436 ;
    wire new_AGEMA_signal_8437 ;
    wire new_AGEMA_signal_8438 ;
    wire new_AGEMA_signal_8439 ;
    wire new_AGEMA_signal_8440 ;
    wire new_AGEMA_signal_8441 ;
    wire new_AGEMA_signal_8442 ;
    wire new_AGEMA_signal_8443 ;
    wire new_AGEMA_signal_8444 ;
    wire new_AGEMA_signal_8445 ;
    wire new_AGEMA_signal_8446 ;
    wire new_AGEMA_signal_8447 ;
    wire new_AGEMA_signal_8448 ;
    wire new_AGEMA_signal_8449 ;
    wire new_AGEMA_signal_8450 ;
    wire new_AGEMA_signal_8451 ;
    wire new_AGEMA_signal_8452 ;
    wire new_AGEMA_signal_8453 ;
    wire new_AGEMA_signal_8454 ;
    wire new_AGEMA_signal_8455 ;
    wire new_AGEMA_signal_8456 ;
    wire new_AGEMA_signal_8457 ;
    wire new_AGEMA_signal_8458 ;
    wire new_AGEMA_signal_8459 ;
    wire new_AGEMA_signal_8460 ;
    wire new_AGEMA_signal_8461 ;
    wire new_AGEMA_signal_8462 ;
    wire new_AGEMA_signal_8463 ;
    wire new_AGEMA_signal_8464 ;
    wire new_AGEMA_signal_8465 ;
    wire new_AGEMA_signal_8466 ;
    wire new_AGEMA_signal_8467 ;
    wire new_AGEMA_signal_8468 ;
    wire new_AGEMA_signal_8469 ;
    wire new_AGEMA_signal_8470 ;
    wire new_AGEMA_signal_8471 ;
    wire new_AGEMA_signal_8472 ;
    wire new_AGEMA_signal_8473 ;
    wire new_AGEMA_signal_8474 ;
    wire new_AGEMA_signal_8475 ;
    wire new_AGEMA_signal_8476 ;
    wire new_AGEMA_signal_8477 ;
    wire new_AGEMA_signal_8478 ;
    wire new_AGEMA_signal_8479 ;
    wire new_AGEMA_signal_8480 ;
    wire new_AGEMA_signal_8481 ;
    wire new_AGEMA_signal_8482 ;
    wire new_AGEMA_signal_8483 ;
    wire new_AGEMA_signal_8484 ;
    wire new_AGEMA_signal_8485 ;
    wire new_AGEMA_signal_8486 ;
    wire new_AGEMA_signal_8487 ;
    wire new_AGEMA_signal_8488 ;
    wire new_AGEMA_signal_8489 ;
    wire new_AGEMA_signal_8490 ;
    wire new_AGEMA_signal_8491 ;
    wire new_AGEMA_signal_8492 ;
    wire new_AGEMA_signal_8493 ;
    wire new_AGEMA_signal_8494 ;
    wire new_AGEMA_signal_8495 ;
    wire new_AGEMA_signal_8496 ;
    wire new_AGEMA_signal_8497 ;
    wire new_AGEMA_signal_8498 ;
    wire new_AGEMA_signal_8499 ;
    wire new_AGEMA_signal_8500 ;
    wire new_AGEMA_signal_8501 ;
    wire new_AGEMA_signal_8502 ;
    wire new_AGEMA_signal_8503 ;
    wire new_AGEMA_signal_8504 ;
    wire new_AGEMA_signal_8505 ;
    wire new_AGEMA_signal_8506 ;
    wire new_AGEMA_signal_8507 ;
    wire new_AGEMA_signal_8508 ;
    wire new_AGEMA_signal_8509 ;
    wire new_AGEMA_signal_8510 ;
    wire new_AGEMA_signal_8511 ;
    wire new_AGEMA_signal_8512 ;
    wire new_AGEMA_signal_8513 ;
    wire new_AGEMA_signal_8514 ;
    wire new_AGEMA_signal_8515 ;
    wire new_AGEMA_signal_8516 ;
    wire new_AGEMA_signal_8517 ;
    wire new_AGEMA_signal_8518 ;
    wire new_AGEMA_signal_8519 ;
    wire new_AGEMA_signal_8520 ;
    wire new_AGEMA_signal_8521 ;
    wire new_AGEMA_signal_8522 ;
    wire new_AGEMA_signal_8523 ;
    wire new_AGEMA_signal_8524 ;
    wire new_AGEMA_signal_8525 ;
    wire new_AGEMA_signal_8526 ;
    wire new_AGEMA_signal_8527 ;
    wire new_AGEMA_signal_8528 ;
    wire new_AGEMA_signal_8529 ;
    wire new_AGEMA_signal_8530 ;
    wire new_AGEMA_signal_8531 ;
    wire new_AGEMA_signal_8532 ;
    wire new_AGEMA_signal_8533 ;
    wire new_AGEMA_signal_8534 ;
    wire new_AGEMA_signal_8535 ;
    wire new_AGEMA_signal_8536 ;
    wire new_AGEMA_signal_8537 ;
    wire new_AGEMA_signal_8538 ;
    wire new_AGEMA_signal_8539 ;
    wire new_AGEMA_signal_8540 ;
    wire new_AGEMA_signal_8541 ;
    wire new_AGEMA_signal_8542 ;
    wire new_AGEMA_signal_8543 ;
    wire new_AGEMA_signal_8544 ;
    wire new_AGEMA_signal_8545 ;
    wire new_AGEMA_signal_8546 ;
    wire new_AGEMA_signal_8547 ;
    wire new_AGEMA_signal_8548 ;
    wire new_AGEMA_signal_8549 ;
    wire new_AGEMA_signal_8550 ;
    wire new_AGEMA_signal_8551 ;
    wire new_AGEMA_signal_8552 ;
    wire new_AGEMA_signal_8553 ;
    wire new_AGEMA_signal_8554 ;
    wire new_AGEMA_signal_8555 ;
    wire new_AGEMA_signal_8556 ;
    wire new_AGEMA_signal_8557 ;
    wire new_AGEMA_signal_8558 ;
    wire new_AGEMA_signal_8559 ;
    wire new_AGEMA_signal_8560 ;
    wire new_AGEMA_signal_8561 ;
    wire new_AGEMA_signal_8562 ;
    wire new_AGEMA_signal_8563 ;
    wire new_AGEMA_signal_8564 ;
    wire new_AGEMA_signal_8565 ;
    wire new_AGEMA_signal_8566 ;
    wire new_AGEMA_signal_8567 ;
    wire new_AGEMA_signal_8568 ;
    wire new_AGEMA_signal_8569 ;
    wire new_AGEMA_signal_8570 ;
    wire new_AGEMA_signal_8571 ;
    wire new_AGEMA_signal_8572 ;
    wire new_AGEMA_signal_8573 ;
    wire new_AGEMA_signal_8574 ;
    wire new_AGEMA_signal_8575 ;
    wire new_AGEMA_signal_8576 ;
    wire new_AGEMA_signal_8577 ;
    wire new_AGEMA_signal_8578 ;
    wire new_AGEMA_signal_8579 ;
    wire new_AGEMA_signal_8580 ;
    wire new_AGEMA_signal_8581 ;
    wire new_AGEMA_signal_8582 ;
    wire new_AGEMA_signal_8583 ;
    wire new_AGEMA_signal_8584 ;
    wire new_AGEMA_signal_8585 ;
    wire new_AGEMA_signal_8586 ;
    wire new_AGEMA_signal_8587 ;
    wire new_AGEMA_signal_8588 ;
    wire new_AGEMA_signal_8589 ;
    wire new_AGEMA_signal_8590 ;
    wire new_AGEMA_signal_8591 ;
    wire new_AGEMA_signal_8592 ;
    wire new_AGEMA_signal_8593 ;
    wire new_AGEMA_signal_8594 ;
    wire new_AGEMA_signal_8595 ;
    wire new_AGEMA_signal_8596 ;
    wire new_AGEMA_signal_8597 ;
    wire new_AGEMA_signal_8598 ;
    wire new_AGEMA_signal_8599 ;
    wire new_AGEMA_signal_8600 ;
    wire new_AGEMA_signal_8601 ;
    wire new_AGEMA_signal_8602 ;
    wire new_AGEMA_signal_8603 ;
    wire new_AGEMA_signal_8604 ;
    wire new_AGEMA_signal_8605 ;
    wire new_AGEMA_signal_8606 ;
    wire new_AGEMA_signal_8607 ;
    wire new_AGEMA_signal_8608 ;
    wire new_AGEMA_signal_8609 ;
    wire new_AGEMA_signal_8610 ;
    wire new_AGEMA_signal_8611 ;
    wire new_AGEMA_signal_8612 ;
    wire new_AGEMA_signal_8613 ;
    wire new_AGEMA_signal_8614 ;
    wire new_AGEMA_signal_8615 ;
    wire new_AGEMA_signal_8616 ;
    wire new_AGEMA_signal_8617 ;
    wire new_AGEMA_signal_8618 ;
    wire new_AGEMA_signal_8619 ;
    wire new_AGEMA_signal_8620 ;
    wire new_AGEMA_signal_8621 ;
    wire new_AGEMA_signal_8622 ;
    wire new_AGEMA_signal_8623 ;
    wire new_AGEMA_signal_8624 ;
    wire new_AGEMA_signal_8625 ;
    wire new_AGEMA_signal_8626 ;
    wire new_AGEMA_signal_8627 ;
    wire new_AGEMA_signal_8628 ;
    wire new_AGEMA_signal_8629 ;
    wire new_AGEMA_signal_8630 ;
    wire new_AGEMA_signal_8631 ;
    wire new_AGEMA_signal_8632 ;
    wire new_AGEMA_signal_8633 ;
    wire new_AGEMA_signal_8634 ;
    wire new_AGEMA_signal_8635 ;
    wire new_AGEMA_signal_8636 ;
    wire new_AGEMA_signal_8637 ;
    wire new_AGEMA_signal_8638 ;
    wire new_AGEMA_signal_8639 ;
    wire new_AGEMA_signal_8640 ;
    wire new_AGEMA_signal_8641 ;
    wire new_AGEMA_signal_8642 ;
    wire new_AGEMA_signal_8643 ;
    wire new_AGEMA_signal_8644 ;
    wire new_AGEMA_signal_8645 ;
    wire new_AGEMA_signal_8646 ;
    wire new_AGEMA_signal_8647 ;
    wire new_AGEMA_signal_8648 ;
    wire new_AGEMA_signal_8649 ;
    wire new_AGEMA_signal_8650 ;
    wire new_AGEMA_signal_8651 ;
    wire new_AGEMA_signal_8652 ;
    wire new_AGEMA_signal_8653 ;
    wire new_AGEMA_signal_8654 ;
    wire new_AGEMA_signal_8655 ;
    wire new_AGEMA_signal_8656 ;
    wire new_AGEMA_signal_8657 ;
    wire new_AGEMA_signal_8658 ;
    wire new_AGEMA_signal_8659 ;
    wire new_AGEMA_signal_8660 ;
    wire new_AGEMA_signal_8661 ;
    wire new_AGEMA_signal_8662 ;
    wire new_AGEMA_signal_8663 ;
    wire new_AGEMA_signal_8664 ;
    wire new_AGEMA_signal_8665 ;
    wire new_AGEMA_signal_8666 ;
    wire new_AGEMA_signal_8667 ;
    wire new_AGEMA_signal_8668 ;
    wire new_AGEMA_signal_8669 ;
    wire new_AGEMA_signal_8670 ;
    wire new_AGEMA_signal_8671 ;
    wire new_AGEMA_signal_8672 ;
    wire new_AGEMA_signal_8673 ;
    wire new_AGEMA_signal_8674 ;
    wire new_AGEMA_signal_8675 ;
    wire new_AGEMA_signal_8676 ;
    wire new_AGEMA_signal_8677 ;
    wire new_AGEMA_signal_8678 ;
    wire new_AGEMA_signal_8679 ;
    wire new_AGEMA_signal_8680 ;
    wire new_AGEMA_signal_8681 ;
    wire new_AGEMA_signal_8682 ;
    wire new_AGEMA_signal_8683 ;
    wire new_AGEMA_signal_8684 ;
    wire new_AGEMA_signal_8685 ;
    wire new_AGEMA_signal_8686 ;
    wire new_AGEMA_signal_8687 ;
    wire new_AGEMA_signal_8688 ;
    wire new_AGEMA_signal_8689 ;
    wire new_AGEMA_signal_8690 ;
    wire new_AGEMA_signal_8691 ;
    wire new_AGEMA_signal_8692 ;
    wire new_AGEMA_signal_8693 ;
    wire new_AGEMA_signal_8694 ;
    wire new_AGEMA_signal_8695 ;
    wire new_AGEMA_signal_8696 ;
    wire new_AGEMA_signal_8697 ;
    wire new_AGEMA_signal_8698 ;
    wire new_AGEMA_signal_8699 ;
    wire new_AGEMA_signal_8700 ;
    wire new_AGEMA_signal_8701 ;
    wire new_AGEMA_signal_8702 ;
    wire new_AGEMA_signal_8703 ;
    wire new_AGEMA_signal_8704 ;
    wire new_AGEMA_signal_8705 ;
    wire new_AGEMA_signal_8706 ;
    wire new_AGEMA_signal_8707 ;
    wire new_AGEMA_signal_8708 ;
    wire new_AGEMA_signal_8709 ;
    wire new_AGEMA_signal_8710 ;
    wire new_AGEMA_signal_8711 ;
    wire new_AGEMA_signal_8712 ;
    wire new_AGEMA_signal_8713 ;
    wire new_AGEMA_signal_8714 ;
    wire new_AGEMA_signal_8715 ;
    wire new_AGEMA_signal_8716 ;
    wire new_AGEMA_signal_8717 ;
    wire new_AGEMA_signal_8718 ;
    wire new_AGEMA_signal_8719 ;
    wire new_AGEMA_signal_8720 ;
    wire new_AGEMA_signal_8721 ;
    wire new_AGEMA_signal_8722 ;
    wire new_AGEMA_signal_8723 ;
    wire new_AGEMA_signal_8724 ;
    wire new_AGEMA_signal_8725 ;
    wire new_AGEMA_signal_8726 ;
    wire new_AGEMA_signal_8727 ;
    wire new_AGEMA_signal_8728 ;
    wire new_AGEMA_signal_8729 ;
    wire new_AGEMA_signal_8730 ;
    wire new_AGEMA_signal_8731 ;
    wire new_AGEMA_signal_8732 ;
    wire new_AGEMA_signal_8733 ;
    wire new_AGEMA_signal_8734 ;
    wire new_AGEMA_signal_8735 ;
    wire new_AGEMA_signal_8736 ;
    wire new_AGEMA_signal_8737 ;
    wire new_AGEMA_signal_8738 ;
    wire new_AGEMA_signal_8739 ;
    wire new_AGEMA_signal_8740 ;
    wire new_AGEMA_signal_8741 ;
    wire new_AGEMA_signal_8742 ;
    wire new_AGEMA_signal_8743 ;
    wire new_AGEMA_signal_8744 ;
    wire new_AGEMA_signal_8745 ;
    wire new_AGEMA_signal_8746 ;
    wire new_AGEMA_signal_8747 ;
    wire new_AGEMA_signal_8748 ;
    wire new_AGEMA_signal_8749 ;
    wire new_AGEMA_signal_8750 ;
    wire new_AGEMA_signal_8751 ;
    wire new_AGEMA_signal_8752 ;
    wire new_AGEMA_signal_8753 ;
    wire new_AGEMA_signal_8754 ;
    wire new_AGEMA_signal_8755 ;
    wire new_AGEMA_signal_8756 ;
    wire new_AGEMA_signal_8757 ;
    wire new_AGEMA_signal_8758 ;
    wire new_AGEMA_signal_8759 ;
    wire new_AGEMA_signal_8760 ;
    wire new_AGEMA_signal_8761 ;
    wire new_AGEMA_signal_8762 ;
    wire new_AGEMA_signal_8763 ;
    wire new_AGEMA_signal_8764 ;
    wire new_AGEMA_signal_8765 ;
    wire new_AGEMA_signal_8766 ;
    wire new_AGEMA_signal_8767 ;
    wire new_AGEMA_signal_8768 ;
    wire new_AGEMA_signal_8769 ;
    wire new_AGEMA_signal_8770 ;
    wire new_AGEMA_signal_8771 ;
    wire new_AGEMA_signal_8772 ;
    wire new_AGEMA_signal_8773 ;
    wire new_AGEMA_signal_8774 ;
    wire new_AGEMA_signal_8775 ;
    wire new_AGEMA_signal_8776 ;
    wire new_AGEMA_signal_8777 ;
    wire new_AGEMA_signal_8778 ;
    wire new_AGEMA_signal_8779 ;
    wire new_AGEMA_signal_8780 ;
    wire new_AGEMA_signal_8781 ;
    wire new_AGEMA_signal_8782 ;
    wire new_AGEMA_signal_8783 ;
    wire new_AGEMA_signal_8784 ;
    wire new_AGEMA_signal_8785 ;
    wire new_AGEMA_signal_8786 ;
    wire new_AGEMA_signal_8787 ;
    wire new_AGEMA_signal_8788 ;
    wire new_AGEMA_signal_8789 ;
    wire new_AGEMA_signal_8790 ;
    wire new_AGEMA_signal_8791 ;
    wire new_AGEMA_signal_8792 ;
    wire new_AGEMA_signal_8793 ;
    wire new_AGEMA_signal_8794 ;
    wire new_AGEMA_signal_8795 ;
    wire new_AGEMA_signal_8796 ;
    wire new_AGEMA_signal_8797 ;
    wire new_AGEMA_signal_8798 ;
    wire new_AGEMA_signal_8799 ;
    wire new_AGEMA_signal_8800 ;
    wire new_AGEMA_signal_8801 ;
    wire new_AGEMA_signal_8802 ;
    wire new_AGEMA_signal_8803 ;
    wire new_AGEMA_signal_8804 ;
    wire new_AGEMA_signal_8805 ;
    wire new_AGEMA_signal_8806 ;
    wire new_AGEMA_signal_8807 ;
    wire new_AGEMA_signal_8808 ;
    wire new_AGEMA_signal_8809 ;
    wire new_AGEMA_signal_8810 ;
    wire new_AGEMA_signal_8811 ;
    wire new_AGEMA_signal_8812 ;
    wire new_AGEMA_signal_8813 ;
    wire new_AGEMA_signal_8814 ;
    wire new_AGEMA_signal_8815 ;
    wire new_AGEMA_signal_8816 ;
    wire new_AGEMA_signal_8817 ;
    wire new_AGEMA_signal_8818 ;
    wire new_AGEMA_signal_8819 ;
    wire new_AGEMA_signal_8820 ;
    wire new_AGEMA_signal_8821 ;
    wire new_AGEMA_signal_8822 ;
    wire new_AGEMA_signal_8823 ;
    wire new_AGEMA_signal_8824 ;
    wire new_AGEMA_signal_8825 ;
    wire new_AGEMA_signal_8826 ;
    wire new_AGEMA_signal_8827 ;
    wire new_AGEMA_signal_8828 ;
    wire new_AGEMA_signal_8829 ;
    wire new_AGEMA_signal_8830 ;
    wire new_AGEMA_signal_8831 ;
    wire new_AGEMA_signal_8832 ;
    wire new_AGEMA_signal_8833 ;
    wire new_AGEMA_signal_8834 ;
    wire new_AGEMA_signal_8835 ;
    wire new_AGEMA_signal_8836 ;
    wire new_AGEMA_signal_8837 ;
    wire new_AGEMA_signal_8838 ;
    wire new_AGEMA_signal_8839 ;
    wire new_AGEMA_signal_8840 ;
    wire new_AGEMA_signal_8841 ;
    wire new_AGEMA_signal_8842 ;
    wire new_AGEMA_signal_8843 ;
    wire new_AGEMA_signal_8844 ;
    wire new_AGEMA_signal_8845 ;
    wire new_AGEMA_signal_8846 ;
    wire new_AGEMA_signal_8847 ;
    wire new_AGEMA_signal_8848 ;
    wire new_AGEMA_signal_8849 ;
    wire new_AGEMA_signal_8850 ;
    wire new_AGEMA_signal_8851 ;
    wire new_AGEMA_signal_8852 ;
    wire new_AGEMA_signal_8853 ;
    wire new_AGEMA_signal_8854 ;
    wire new_AGEMA_signal_8855 ;
    wire new_AGEMA_signal_8856 ;
    wire new_AGEMA_signal_8857 ;
    wire new_AGEMA_signal_8858 ;
    wire new_AGEMA_signal_8859 ;
    wire new_AGEMA_signal_8860 ;
    wire new_AGEMA_signal_8861 ;
    wire new_AGEMA_signal_8862 ;
    wire new_AGEMA_signal_8863 ;
    wire new_AGEMA_signal_8864 ;
    wire new_AGEMA_signal_8865 ;
    wire new_AGEMA_signal_8866 ;
    wire new_AGEMA_signal_8867 ;
    wire new_AGEMA_signal_8868 ;
    wire new_AGEMA_signal_8869 ;
    wire new_AGEMA_signal_8870 ;
    wire new_AGEMA_signal_8871 ;
    wire new_AGEMA_signal_8872 ;
    wire new_AGEMA_signal_8873 ;
    wire new_AGEMA_signal_8874 ;
    wire new_AGEMA_signal_8875 ;
    wire new_AGEMA_signal_8876 ;
    wire new_AGEMA_signal_8877 ;
    wire new_AGEMA_signal_8878 ;
    wire new_AGEMA_signal_8879 ;
    wire new_AGEMA_signal_8880 ;
    wire new_AGEMA_signal_8881 ;
    wire new_AGEMA_signal_8882 ;
    wire new_AGEMA_signal_8883 ;
    wire new_AGEMA_signal_8884 ;
    wire new_AGEMA_signal_8885 ;
    wire new_AGEMA_signal_8886 ;
    wire new_AGEMA_signal_8887 ;
    wire new_AGEMA_signal_8888 ;
    wire new_AGEMA_signal_8889 ;
    wire new_AGEMA_signal_8890 ;
    wire new_AGEMA_signal_8891 ;
    wire new_AGEMA_signal_8892 ;
    wire new_AGEMA_signal_8893 ;
    wire new_AGEMA_signal_8894 ;
    wire new_AGEMA_signal_8895 ;
    wire new_AGEMA_signal_8896 ;
    wire new_AGEMA_signal_8897 ;
    wire new_AGEMA_signal_8898 ;
    wire new_AGEMA_signal_8899 ;
    wire new_AGEMA_signal_8900 ;
    wire new_AGEMA_signal_8901 ;
    wire new_AGEMA_signal_8902 ;
    wire new_AGEMA_signal_8903 ;
    wire new_AGEMA_signal_8904 ;
    wire new_AGEMA_signal_8905 ;
    wire new_AGEMA_signal_8906 ;
    wire new_AGEMA_signal_8907 ;
    wire new_AGEMA_signal_8908 ;
    wire new_AGEMA_signal_8909 ;
    wire new_AGEMA_signal_8910 ;
    wire new_AGEMA_signal_8911 ;
    wire new_AGEMA_signal_8912 ;
    wire new_AGEMA_signal_8913 ;
    wire new_AGEMA_signal_8914 ;
    wire new_AGEMA_signal_8915 ;
    wire new_AGEMA_signal_8916 ;
    wire new_AGEMA_signal_8917 ;
    wire new_AGEMA_signal_8918 ;
    wire new_AGEMA_signal_8919 ;
    wire new_AGEMA_signal_8920 ;
    wire new_AGEMA_signal_8921 ;
    wire new_AGEMA_signal_8922 ;
    wire new_AGEMA_signal_8923 ;
    wire new_AGEMA_signal_8924 ;
    wire new_AGEMA_signal_8925 ;
    wire new_AGEMA_signal_8926 ;
    wire new_AGEMA_signal_8927 ;
    wire new_AGEMA_signal_8928 ;
    wire new_AGEMA_signal_8929 ;
    wire new_AGEMA_signal_8930 ;
    wire new_AGEMA_signal_8931 ;
    wire new_AGEMA_signal_8932 ;
    wire new_AGEMA_signal_8933 ;
    wire new_AGEMA_signal_8934 ;
    wire new_AGEMA_signal_8935 ;
    wire new_AGEMA_signal_8936 ;
    wire new_AGEMA_signal_8937 ;
    wire new_AGEMA_signal_8938 ;
    wire new_AGEMA_signal_8939 ;
    wire new_AGEMA_signal_8940 ;
    wire new_AGEMA_signal_8941 ;
    wire new_AGEMA_signal_8942 ;
    wire new_AGEMA_signal_8943 ;
    wire new_AGEMA_signal_8944 ;
    wire new_AGEMA_signal_8945 ;
    wire new_AGEMA_signal_8946 ;
    wire new_AGEMA_signal_8947 ;
    wire new_AGEMA_signal_8948 ;
    wire new_AGEMA_signal_8949 ;
    wire new_AGEMA_signal_8950 ;
    wire new_AGEMA_signal_8951 ;
    wire new_AGEMA_signal_8952 ;
    wire new_AGEMA_signal_8953 ;
    wire new_AGEMA_signal_8954 ;
    wire new_AGEMA_signal_8955 ;
    wire new_AGEMA_signal_8956 ;
    wire new_AGEMA_signal_8957 ;
    wire new_AGEMA_signal_8958 ;
    wire new_AGEMA_signal_8959 ;
    wire new_AGEMA_signal_8960 ;
    wire new_AGEMA_signal_8961 ;
    wire new_AGEMA_signal_8962 ;
    wire new_AGEMA_signal_8963 ;
    wire new_AGEMA_signal_8964 ;
    wire new_AGEMA_signal_8965 ;
    wire new_AGEMA_signal_8966 ;
    wire new_AGEMA_signal_8967 ;
    wire new_AGEMA_signal_8968 ;
    wire new_AGEMA_signal_8969 ;
    wire new_AGEMA_signal_8970 ;
    wire new_AGEMA_signal_8971 ;
    wire new_AGEMA_signal_8972 ;
    wire new_AGEMA_signal_8973 ;
    wire new_AGEMA_signal_8974 ;
    wire new_AGEMA_signal_8975 ;
    wire new_AGEMA_signal_8976 ;
    wire new_AGEMA_signal_8977 ;
    wire new_AGEMA_signal_8978 ;
    wire new_AGEMA_signal_8979 ;
    wire new_AGEMA_signal_8980 ;
    wire new_AGEMA_signal_8981 ;
    wire new_AGEMA_signal_8982 ;
    wire new_AGEMA_signal_8983 ;
    wire new_AGEMA_signal_8984 ;
    wire new_AGEMA_signal_8985 ;
    wire new_AGEMA_signal_8986 ;
    wire new_AGEMA_signal_8987 ;
    wire new_AGEMA_signal_8988 ;
    wire new_AGEMA_signal_8989 ;
    wire new_AGEMA_signal_8990 ;
    wire new_AGEMA_signal_8991 ;
    wire new_AGEMA_signal_8992 ;
    wire new_AGEMA_signal_8993 ;
    wire new_AGEMA_signal_8994 ;
    wire new_AGEMA_signal_8995 ;
    wire new_AGEMA_signal_8996 ;
    wire new_AGEMA_signal_8997 ;
    wire new_AGEMA_signal_8998 ;
    wire new_AGEMA_signal_8999 ;
    wire new_AGEMA_signal_9000 ;
    wire new_AGEMA_signal_9001 ;
    wire new_AGEMA_signal_9002 ;
    wire new_AGEMA_signal_9003 ;
    wire new_AGEMA_signal_9004 ;
    wire new_AGEMA_signal_9005 ;
    wire new_AGEMA_signal_9006 ;
    wire new_AGEMA_signal_9007 ;
    wire new_AGEMA_signal_9008 ;
    wire new_AGEMA_signal_9009 ;
    wire new_AGEMA_signal_9010 ;
    wire new_AGEMA_signal_9011 ;
    wire new_AGEMA_signal_9012 ;
    wire new_AGEMA_signal_9013 ;
    wire new_AGEMA_signal_9014 ;
    wire new_AGEMA_signal_9015 ;
    wire new_AGEMA_signal_9016 ;
    wire new_AGEMA_signal_9017 ;
    wire new_AGEMA_signal_9018 ;
    wire new_AGEMA_signal_9019 ;
    wire new_AGEMA_signal_9020 ;
    wire new_AGEMA_signal_9021 ;
    wire new_AGEMA_signal_9022 ;
    wire new_AGEMA_signal_9023 ;
    wire new_AGEMA_signal_9024 ;
    wire new_AGEMA_signal_9025 ;
    wire new_AGEMA_signal_9026 ;
    wire new_AGEMA_signal_9027 ;
    wire new_AGEMA_signal_9028 ;
    wire new_AGEMA_signal_9029 ;
    wire new_AGEMA_signal_9030 ;
    wire new_AGEMA_signal_9031 ;
    wire new_AGEMA_signal_9032 ;
    wire new_AGEMA_signal_9033 ;
    wire new_AGEMA_signal_9034 ;
    wire new_AGEMA_signal_9035 ;
    wire new_AGEMA_signal_9036 ;
    wire new_AGEMA_signal_9037 ;
    wire new_AGEMA_signal_9038 ;
    wire new_AGEMA_signal_9039 ;
    wire new_AGEMA_signal_9040 ;
    wire new_AGEMA_signal_9041 ;
    wire new_AGEMA_signal_9042 ;
    wire new_AGEMA_signal_9043 ;
    wire new_AGEMA_signal_9044 ;
    wire new_AGEMA_signal_9045 ;
    wire new_AGEMA_signal_9046 ;
    wire new_AGEMA_signal_9047 ;
    wire new_AGEMA_signal_9048 ;
    wire new_AGEMA_signal_9049 ;
    wire new_AGEMA_signal_9050 ;
    wire new_AGEMA_signal_9051 ;
    wire new_AGEMA_signal_9052 ;
    wire new_AGEMA_signal_9053 ;
    wire new_AGEMA_signal_9054 ;
    wire new_AGEMA_signal_9055 ;
    wire new_AGEMA_signal_9056 ;
    wire new_AGEMA_signal_9057 ;
    wire new_AGEMA_signal_9058 ;
    wire new_AGEMA_signal_9059 ;
    wire new_AGEMA_signal_9060 ;
    wire new_AGEMA_signal_9061 ;
    wire new_AGEMA_signal_9062 ;
    wire new_AGEMA_signal_9063 ;
    wire new_AGEMA_signal_9064 ;
    wire new_AGEMA_signal_9065 ;
    wire new_AGEMA_signal_9066 ;
    wire new_AGEMA_signal_9067 ;
    wire new_AGEMA_signal_9068 ;
    wire new_AGEMA_signal_9069 ;
    wire new_AGEMA_signal_9070 ;
    wire new_AGEMA_signal_9071 ;
    wire new_AGEMA_signal_9072 ;
    wire new_AGEMA_signal_9073 ;
    wire new_AGEMA_signal_9074 ;
    wire new_AGEMA_signal_9075 ;
    wire new_AGEMA_signal_9076 ;
    wire new_AGEMA_signal_9077 ;
    wire new_AGEMA_signal_9078 ;
    wire new_AGEMA_signal_9079 ;
    wire new_AGEMA_signal_9080 ;
    wire new_AGEMA_signal_9081 ;
    wire new_AGEMA_signal_9082 ;
    wire new_AGEMA_signal_9083 ;
    wire new_AGEMA_signal_9084 ;
    wire new_AGEMA_signal_9085 ;
    wire new_AGEMA_signal_9086 ;
    wire new_AGEMA_signal_9087 ;
    wire new_AGEMA_signal_9088 ;
    wire new_AGEMA_signal_9089 ;
    wire new_AGEMA_signal_9090 ;
    wire new_AGEMA_signal_9091 ;
    wire new_AGEMA_signal_9092 ;
    wire new_AGEMA_signal_9093 ;
    wire new_AGEMA_signal_9094 ;
    wire new_AGEMA_signal_9095 ;
    wire new_AGEMA_signal_9096 ;
    wire new_AGEMA_signal_9097 ;
    wire new_AGEMA_signal_9098 ;
    wire new_AGEMA_signal_9099 ;
    wire new_AGEMA_signal_9100 ;
    wire new_AGEMA_signal_9101 ;
    wire new_AGEMA_signal_9102 ;
    wire new_AGEMA_signal_9103 ;
    wire new_AGEMA_signal_9104 ;
    wire new_AGEMA_signal_9105 ;
    wire new_AGEMA_signal_9106 ;
    wire new_AGEMA_signal_9107 ;
    wire new_AGEMA_signal_9108 ;
    wire new_AGEMA_signal_9109 ;
    wire new_AGEMA_signal_9110 ;
    wire new_AGEMA_signal_9111 ;
    wire new_AGEMA_signal_9112 ;
    wire new_AGEMA_signal_9113 ;
    wire new_AGEMA_signal_9114 ;
    wire new_AGEMA_signal_9115 ;
    wire new_AGEMA_signal_9116 ;
    wire new_AGEMA_signal_9117 ;
    wire new_AGEMA_signal_9118 ;
    wire new_AGEMA_signal_9119 ;
    wire new_AGEMA_signal_9120 ;
    wire new_AGEMA_signal_9121 ;
    wire new_AGEMA_signal_9122 ;
    wire new_AGEMA_signal_9123 ;
    wire new_AGEMA_signal_9124 ;
    wire new_AGEMA_signal_9125 ;
    wire new_AGEMA_signal_9126 ;
    wire new_AGEMA_signal_9127 ;
    wire new_AGEMA_signal_9128 ;
    wire new_AGEMA_signal_9129 ;
    wire new_AGEMA_signal_9130 ;
    wire new_AGEMA_signal_9131 ;
    wire new_AGEMA_signal_9132 ;
    wire new_AGEMA_signal_9133 ;
    wire new_AGEMA_signal_9134 ;
    wire new_AGEMA_signal_9135 ;
    wire new_AGEMA_signal_9136 ;
    wire new_AGEMA_signal_9137 ;
    wire new_AGEMA_signal_9138 ;
    wire new_AGEMA_signal_9139 ;
    wire new_AGEMA_signal_9140 ;
    wire new_AGEMA_signal_9141 ;
    wire new_AGEMA_signal_9142 ;
    wire new_AGEMA_signal_9143 ;
    wire new_AGEMA_signal_9144 ;
    wire new_AGEMA_signal_9145 ;
    wire new_AGEMA_signal_9146 ;
    wire new_AGEMA_signal_9147 ;
    wire new_AGEMA_signal_9148 ;
    wire new_AGEMA_signal_9149 ;
    wire new_AGEMA_signal_9150 ;
    wire new_AGEMA_signal_9151 ;
    wire new_AGEMA_signal_9152 ;
    wire new_AGEMA_signal_9153 ;
    wire new_AGEMA_signal_9154 ;
    wire new_AGEMA_signal_9155 ;
    wire new_AGEMA_signal_9156 ;
    wire new_AGEMA_signal_9157 ;
    wire new_AGEMA_signal_9158 ;
    wire new_AGEMA_signal_9159 ;
    wire new_AGEMA_signal_9160 ;
    wire new_AGEMA_signal_9161 ;
    wire new_AGEMA_signal_9162 ;
    wire new_AGEMA_signal_9163 ;
    wire new_AGEMA_signal_9164 ;
    wire new_AGEMA_signal_9165 ;
    wire new_AGEMA_signal_9166 ;
    wire new_AGEMA_signal_9167 ;
    wire new_AGEMA_signal_9168 ;
    wire new_AGEMA_signal_9169 ;
    wire new_AGEMA_signal_9170 ;
    wire new_AGEMA_signal_9171 ;
    wire new_AGEMA_signal_9172 ;
    wire new_AGEMA_signal_9173 ;
    wire new_AGEMA_signal_9174 ;
    wire new_AGEMA_signal_9175 ;
    wire new_AGEMA_signal_9176 ;
    wire new_AGEMA_signal_9177 ;
    wire new_AGEMA_signal_9178 ;
    wire new_AGEMA_signal_9179 ;
    wire new_AGEMA_signal_9180 ;
    wire new_AGEMA_signal_9181 ;
    wire new_AGEMA_signal_9182 ;
    wire new_AGEMA_signal_9183 ;
    wire new_AGEMA_signal_9184 ;
    wire new_AGEMA_signal_9185 ;
    wire new_AGEMA_signal_9186 ;
    wire new_AGEMA_signal_9187 ;
    wire new_AGEMA_signal_9188 ;
    wire new_AGEMA_signal_9189 ;
    wire new_AGEMA_signal_9190 ;
    wire new_AGEMA_signal_9191 ;
    wire new_AGEMA_signal_9192 ;
    wire new_AGEMA_signal_9193 ;
    wire new_AGEMA_signal_9194 ;
    wire new_AGEMA_signal_9195 ;
    wire new_AGEMA_signal_9196 ;
    wire new_AGEMA_signal_9197 ;
    wire new_AGEMA_signal_9198 ;
    wire new_AGEMA_signal_9199 ;
    wire new_AGEMA_signal_9200 ;
    wire new_AGEMA_signal_9201 ;
    wire new_AGEMA_signal_9202 ;
    wire new_AGEMA_signal_9203 ;
    wire new_AGEMA_signal_9204 ;
    wire new_AGEMA_signal_9205 ;
    wire new_AGEMA_signal_9206 ;
    wire new_AGEMA_signal_9207 ;
    wire new_AGEMA_signal_9208 ;
    wire new_AGEMA_signal_9209 ;
    wire new_AGEMA_signal_9210 ;
    wire new_AGEMA_signal_9211 ;
    wire new_AGEMA_signal_9212 ;
    wire new_AGEMA_signal_9213 ;
    wire new_AGEMA_signal_9214 ;
    wire new_AGEMA_signal_9215 ;
    wire new_AGEMA_signal_9216 ;
    wire new_AGEMA_signal_9217 ;
    wire new_AGEMA_signal_9218 ;
    wire new_AGEMA_signal_9219 ;
    wire new_AGEMA_signal_9220 ;
    wire new_AGEMA_signal_9221 ;
    wire new_AGEMA_signal_9222 ;
    wire new_AGEMA_signal_9223 ;
    wire new_AGEMA_signal_9224 ;
    wire new_AGEMA_signal_9225 ;
    wire new_AGEMA_signal_9226 ;
    wire new_AGEMA_signal_9227 ;
    wire new_AGEMA_signal_9228 ;
    wire new_AGEMA_signal_9229 ;
    wire new_AGEMA_signal_9230 ;
    wire new_AGEMA_signal_9231 ;
    wire new_AGEMA_signal_9232 ;
    wire new_AGEMA_signal_9233 ;
    wire new_AGEMA_signal_9234 ;
    wire new_AGEMA_signal_9235 ;
    wire new_AGEMA_signal_9236 ;
    wire new_AGEMA_signal_9237 ;
    wire new_AGEMA_signal_9238 ;
    wire new_AGEMA_signal_9239 ;
    wire new_AGEMA_signal_9240 ;
    wire new_AGEMA_signal_9241 ;
    wire new_AGEMA_signal_9242 ;
    wire new_AGEMA_signal_9243 ;
    wire new_AGEMA_signal_9244 ;
    wire new_AGEMA_signal_9245 ;
    wire new_AGEMA_signal_9246 ;
    wire new_AGEMA_signal_9247 ;
    wire new_AGEMA_signal_9248 ;
    wire new_AGEMA_signal_9249 ;
    wire new_AGEMA_signal_9250 ;
    wire new_AGEMA_signal_9251 ;
    wire new_AGEMA_signal_9252 ;
    wire new_AGEMA_signal_9253 ;
    wire new_AGEMA_signal_9254 ;
    wire new_AGEMA_signal_9255 ;
    wire new_AGEMA_signal_9256 ;
    wire new_AGEMA_signal_9257 ;
    wire new_AGEMA_signal_9258 ;
    wire new_AGEMA_signal_9259 ;
    wire new_AGEMA_signal_9260 ;
    wire new_AGEMA_signal_9261 ;
    wire new_AGEMA_signal_9262 ;
    wire new_AGEMA_signal_9263 ;
    wire new_AGEMA_signal_9264 ;
    wire new_AGEMA_signal_9265 ;
    wire new_AGEMA_signal_9266 ;
    wire new_AGEMA_signal_9267 ;
    wire new_AGEMA_signal_9268 ;
    wire new_AGEMA_signal_9269 ;
    wire new_AGEMA_signal_9270 ;
    wire new_AGEMA_signal_9271 ;
    wire new_AGEMA_signal_9272 ;
    wire new_AGEMA_signal_9273 ;
    wire new_AGEMA_signal_9274 ;
    wire new_AGEMA_signal_9275 ;
    wire new_AGEMA_signal_9276 ;
    wire new_AGEMA_signal_9277 ;
    wire new_AGEMA_signal_9278 ;
    wire new_AGEMA_signal_9279 ;
    wire new_AGEMA_signal_9280 ;
    wire new_AGEMA_signal_9281 ;
    wire new_AGEMA_signal_9282 ;
    wire new_AGEMA_signal_9283 ;
    wire new_AGEMA_signal_9284 ;
    wire new_AGEMA_signal_9285 ;
    wire new_AGEMA_signal_9286 ;
    wire new_AGEMA_signal_9287 ;
    wire new_AGEMA_signal_9288 ;
    wire new_AGEMA_signal_9289 ;
    wire new_AGEMA_signal_9290 ;
    wire new_AGEMA_signal_9291 ;
    wire new_AGEMA_signal_9292 ;
    wire new_AGEMA_signal_9293 ;
    wire new_AGEMA_signal_9294 ;
    wire new_AGEMA_signal_9295 ;
    wire new_AGEMA_signal_9296 ;
    wire new_AGEMA_signal_9297 ;
    wire new_AGEMA_signal_9298 ;
    wire new_AGEMA_signal_9299 ;
    wire new_AGEMA_signal_9300 ;
    wire new_AGEMA_signal_9301 ;
    wire new_AGEMA_signal_9302 ;
    wire new_AGEMA_signal_9303 ;
    wire new_AGEMA_signal_9304 ;
    wire new_AGEMA_signal_9305 ;
    wire new_AGEMA_signal_9306 ;
    wire new_AGEMA_signal_9307 ;
    wire new_AGEMA_signal_9308 ;
    wire new_AGEMA_signal_9309 ;
    wire new_AGEMA_signal_9310 ;
    wire new_AGEMA_signal_9311 ;
    wire new_AGEMA_signal_9312 ;
    wire new_AGEMA_signal_9313 ;
    wire new_AGEMA_signal_9314 ;
    wire new_AGEMA_signal_9315 ;
    wire new_AGEMA_signal_9316 ;
    wire new_AGEMA_signal_9317 ;
    wire new_AGEMA_signal_9318 ;
    wire new_AGEMA_signal_9319 ;
    wire new_AGEMA_signal_9320 ;
    wire new_AGEMA_signal_9321 ;
    wire new_AGEMA_signal_9322 ;
    wire new_AGEMA_signal_9323 ;
    wire new_AGEMA_signal_9324 ;
    wire new_AGEMA_signal_9325 ;
    wire new_AGEMA_signal_9326 ;
    wire new_AGEMA_signal_9327 ;
    wire new_AGEMA_signal_9328 ;
    wire new_AGEMA_signal_9329 ;
    wire new_AGEMA_signal_9330 ;
    wire new_AGEMA_signal_9331 ;
    wire new_AGEMA_signal_9332 ;
    wire new_AGEMA_signal_9333 ;
    wire new_AGEMA_signal_9334 ;
    wire new_AGEMA_signal_9335 ;
    wire new_AGEMA_signal_9336 ;
    wire new_AGEMA_signal_9337 ;
    wire new_AGEMA_signal_9338 ;
    wire new_AGEMA_signal_9339 ;
    wire new_AGEMA_signal_9340 ;
    wire new_AGEMA_signal_9341 ;
    wire new_AGEMA_signal_9342 ;
    wire new_AGEMA_signal_9343 ;
    wire new_AGEMA_signal_9344 ;
    wire new_AGEMA_signal_9345 ;
    wire new_AGEMA_signal_9346 ;
    wire new_AGEMA_signal_9347 ;
    wire new_AGEMA_signal_9348 ;
    wire new_AGEMA_signal_9349 ;
    wire new_AGEMA_signal_9350 ;
    wire new_AGEMA_signal_9351 ;
    wire new_AGEMA_signal_9352 ;
    wire new_AGEMA_signal_9353 ;
    wire new_AGEMA_signal_9354 ;
    wire new_AGEMA_signal_9355 ;
    wire new_AGEMA_signal_9356 ;
    wire new_AGEMA_signal_9357 ;
    wire new_AGEMA_signal_9358 ;
    wire new_AGEMA_signal_9359 ;
    wire new_AGEMA_signal_9360 ;
    wire new_AGEMA_signal_9361 ;
    wire new_AGEMA_signal_9362 ;
    wire new_AGEMA_signal_9363 ;
    wire new_AGEMA_signal_9364 ;
    wire new_AGEMA_signal_9365 ;
    wire new_AGEMA_signal_9366 ;
    wire new_AGEMA_signal_9367 ;
    wire new_AGEMA_signal_9368 ;
    wire new_AGEMA_signal_9369 ;
    wire new_AGEMA_signal_9370 ;
    wire new_AGEMA_signal_9371 ;
    wire new_AGEMA_signal_9372 ;
    wire new_AGEMA_signal_9373 ;
    wire new_AGEMA_signal_9374 ;
    wire new_AGEMA_signal_9375 ;
    wire new_AGEMA_signal_9376 ;
    wire new_AGEMA_signal_9377 ;
    wire new_AGEMA_signal_9378 ;
    wire new_AGEMA_signal_9379 ;
    wire new_AGEMA_signal_9380 ;
    wire new_AGEMA_signal_9381 ;
    wire new_AGEMA_signal_9382 ;
    wire new_AGEMA_signal_9383 ;
    wire new_AGEMA_signal_9384 ;
    wire new_AGEMA_signal_9385 ;
    wire new_AGEMA_signal_9386 ;
    wire new_AGEMA_signal_9387 ;
    wire new_AGEMA_signal_9388 ;
    wire new_AGEMA_signal_9389 ;
    wire new_AGEMA_signal_9390 ;
    wire new_AGEMA_signal_9391 ;
    wire new_AGEMA_signal_9392 ;
    wire new_AGEMA_signal_9393 ;
    wire new_AGEMA_signal_9394 ;
    wire new_AGEMA_signal_9395 ;
    wire new_AGEMA_signal_9396 ;
    wire new_AGEMA_signal_9397 ;
    wire new_AGEMA_signal_9398 ;
    wire new_AGEMA_signal_9399 ;
    wire new_AGEMA_signal_9400 ;
    wire new_AGEMA_signal_9401 ;
    wire new_AGEMA_signal_9402 ;
    wire new_AGEMA_signal_9403 ;
    wire new_AGEMA_signal_9404 ;
    wire new_AGEMA_signal_9405 ;
    wire new_AGEMA_signal_9406 ;
    wire new_AGEMA_signal_9407 ;
    wire new_AGEMA_signal_9408 ;
    wire new_AGEMA_signal_9409 ;
    wire new_AGEMA_signal_9410 ;
    wire new_AGEMA_signal_9411 ;
    wire new_AGEMA_signal_9412 ;
    wire new_AGEMA_signal_9413 ;
    wire new_AGEMA_signal_9414 ;
    wire new_AGEMA_signal_9415 ;
    wire new_AGEMA_signal_9416 ;
    wire new_AGEMA_signal_9417 ;
    wire new_AGEMA_signal_9418 ;
    wire new_AGEMA_signal_9419 ;
    wire new_AGEMA_signal_9420 ;
    wire new_AGEMA_signal_9421 ;
    wire new_AGEMA_signal_9422 ;
    wire new_AGEMA_signal_9423 ;
    wire new_AGEMA_signal_9424 ;
    wire new_AGEMA_signal_9425 ;
    wire new_AGEMA_signal_9426 ;
    wire new_AGEMA_signal_9427 ;
    wire new_AGEMA_signal_9428 ;
    wire new_AGEMA_signal_9429 ;
    wire new_AGEMA_signal_9430 ;
    wire new_AGEMA_signal_9431 ;
    wire new_AGEMA_signal_9432 ;
    wire new_AGEMA_signal_9433 ;
    wire new_AGEMA_signal_9434 ;
    wire new_AGEMA_signal_9435 ;
    wire new_AGEMA_signal_9436 ;
    wire new_AGEMA_signal_9437 ;
    wire new_AGEMA_signal_9438 ;
    wire new_AGEMA_signal_9439 ;
    wire new_AGEMA_signal_9440 ;
    wire new_AGEMA_signal_9441 ;
    wire new_AGEMA_signal_9442 ;
    wire new_AGEMA_signal_9443 ;
    wire new_AGEMA_signal_9444 ;
    wire new_AGEMA_signal_9445 ;
    wire new_AGEMA_signal_9446 ;
    wire new_AGEMA_signal_9447 ;
    wire new_AGEMA_signal_9448 ;
    wire new_AGEMA_signal_9449 ;
    wire new_AGEMA_signal_9450 ;
    wire new_AGEMA_signal_9451 ;
    wire new_AGEMA_signal_9452 ;
    wire new_AGEMA_signal_9453 ;
    wire new_AGEMA_signal_9454 ;
    wire new_AGEMA_signal_9455 ;
    wire new_AGEMA_signal_9456 ;
    wire new_AGEMA_signal_9457 ;
    wire new_AGEMA_signal_9458 ;
    wire new_AGEMA_signal_9459 ;
    wire new_AGEMA_signal_9460 ;
    wire new_AGEMA_signal_9461 ;
    wire new_AGEMA_signal_9462 ;
    wire new_AGEMA_signal_9463 ;
    wire new_AGEMA_signal_9464 ;
    wire new_AGEMA_signal_9465 ;
    wire new_AGEMA_signal_9466 ;
    wire new_AGEMA_signal_9467 ;
    wire new_AGEMA_signal_9468 ;
    wire new_AGEMA_signal_9469 ;
    wire new_AGEMA_signal_9470 ;
    wire new_AGEMA_signal_9471 ;
    wire new_AGEMA_signal_9472 ;
    wire new_AGEMA_signal_9473 ;
    wire new_AGEMA_signal_9474 ;
    wire new_AGEMA_signal_9475 ;
    wire new_AGEMA_signal_9476 ;
    wire new_AGEMA_signal_9477 ;
    wire new_AGEMA_signal_9478 ;
    wire new_AGEMA_signal_9479 ;
    wire new_AGEMA_signal_9480 ;
    wire new_AGEMA_signal_9481 ;
    wire new_AGEMA_signal_9482 ;
    wire new_AGEMA_signal_9483 ;
    wire new_AGEMA_signal_9484 ;
    wire new_AGEMA_signal_9485 ;
    wire new_AGEMA_signal_9486 ;
    wire new_AGEMA_signal_9487 ;
    wire new_AGEMA_signal_9488 ;
    wire new_AGEMA_signal_9489 ;
    wire new_AGEMA_signal_9490 ;
    wire new_AGEMA_signal_9491 ;
    wire new_AGEMA_signal_9492 ;
    wire new_AGEMA_signal_9493 ;
    wire new_AGEMA_signal_9494 ;
    wire new_AGEMA_signal_9495 ;
    wire new_AGEMA_signal_9496 ;
    wire new_AGEMA_signal_9497 ;
    wire new_AGEMA_signal_9498 ;
    wire new_AGEMA_signal_9499 ;
    wire new_AGEMA_signal_9500 ;
    wire new_AGEMA_signal_9501 ;
    wire new_AGEMA_signal_9502 ;
    wire new_AGEMA_signal_9503 ;
    wire new_AGEMA_signal_9504 ;
    wire new_AGEMA_signal_9505 ;
    wire new_AGEMA_signal_9506 ;
    wire new_AGEMA_signal_9507 ;
    wire new_AGEMA_signal_9508 ;
    wire new_AGEMA_signal_9509 ;
    wire new_AGEMA_signal_9510 ;
    wire new_AGEMA_signal_9511 ;
    wire new_AGEMA_signal_9512 ;
    wire new_AGEMA_signal_9513 ;
    wire new_AGEMA_signal_9514 ;
    wire new_AGEMA_signal_9515 ;
    wire new_AGEMA_signal_9516 ;
    wire new_AGEMA_signal_9517 ;
    wire new_AGEMA_signal_9518 ;
    wire new_AGEMA_signal_9519 ;
    wire new_AGEMA_signal_9520 ;
    wire new_AGEMA_signal_9521 ;
    wire new_AGEMA_signal_9522 ;
    wire new_AGEMA_signal_9523 ;
    wire new_AGEMA_signal_9524 ;
    wire new_AGEMA_signal_9525 ;
    wire new_AGEMA_signal_9526 ;
    wire new_AGEMA_signal_9527 ;
    wire new_AGEMA_signal_9528 ;
    wire new_AGEMA_signal_9529 ;
    wire new_AGEMA_signal_9530 ;
    wire new_AGEMA_signal_9531 ;
    wire new_AGEMA_signal_9532 ;
    wire new_AGEMA_signal_9533 ;
    wire new_AGEMA_signal_9534 ;
    wire new_AGEMA_signal_9535 ;
    wire new_AGEMA_signal_9536 ;
    wire new_AGEMA_signal_9537 ;
    wire new_AGEMA_signal_9538 ;
    wire new_AGEMA_signal_9539 ;
    wire new_AGEMA_signal_9540 ;
    wire new_AGEMA_signal_9541 ;
    wire new_AGEMA_signal_9542 ;
    wire new_AGEMA_signal_9543 ;
    wire new_AGEMA_signal_9544 ;
    wire new_AGEMA_signal_9545 ;
    wire new_AGEMA_signal_9546 ;
    wire new_AGEMA_signal_9547 ;
    wire new_AGEMA_signal_9548 ;
    wire new_AGEMA_signal_9549 ;
    wire new_AGEMA_signal_9550 ;
    wire new_AGEMA_signal_9551 ;
    wire new_AGEMA_signal_9552 ;
    wire new_AGEMA_signal_9553 ;
    wire new_AGEMA_signal_9554 ;
    wire new_AGEMA_signal_9555 ;
    wire new_AGEMA_signal_9556 ;
    wire new_AGEMA_signal_9557 ;
    wire new_AGEMA_signal_9558 ;
    wire new_AGEMA_signal_9559 ;
    wire new_AGEMA_signal_9560 ;
    wire new_AGEMA_signal_9561 ;
    wire new_AGEMA_signal_9562 ;
    wire new_AGEMA_signal_9563 ;
    wire new_AGEMA_signal_9564 ;
    wire new_AGEMA_signal_9565 ;
    wire new_AGEMA_signal_9566 ;
    wire new_AGEMA_signal_9567 ;
    wire new_AGEMA_signal_9568 ;
    wire new_AGEMA_signal_9569 ;
    wire new_AGEMA_signal_9570 ;
    wire new_AGEMA_signal_9571 ;
    wire new_AGEMA_signal_9572 ;
    wire new_AGEMA_signal_9573 ;
    wire new_AGEMA_signal_9574 ;
    wire new_AGEMA_signal_9575 ;
    wire new_AGEMA_signal_9576 ;
    wire new_AGEMA_signal_9577 ;
    wire new_AGEMA_signal_9578 ;
    wire new_AGEMA_signal_9579 ;
    wire new_AGEMA_signal_9580 ;
    wire new_AGEMA_signal_9581 ;
    wire new_AGEMA_signal_9582 ;
    wire new_AGEMA_signal_9583 ;
    wire new_AGEMA_signal_9584 ;
    wire new_AGEMA_signal_9585 ;
    wire new_AGEMA_signal_9586 ;
    wire new_AGEMA_signal_9587 ;
    wire new_AGEMA_signal_9588 ;
    wire new_AGEMA_signal_9589 ;
    wire new_AGEMA_signal_9590 ;
    wire new_AGEMA_signal_9591 ;
    wire new_AGEMA_signal_9592 ;
    wire new_AGEMA_signal_9593 ;
    wire new_AGEMA_signal_9594 ;
    wire new_AGEMA_signal_9595 ;
    wire new_AGEMA_signal_9596 ;
    wire new_AGEMA_signal_9597 ;
    wire new_AGEMA_signal_9598 ;
    wire new_AGEMA_signal_9599 ;
    wire new_AGEMA_signal_9600 ;
    wire new_AGEMA_signal_9601 ;
    wire new_AGEMA_signal_9602 ;
    wire new_AGEMA_signal_9603 ;
    wire new_AGEMA_signal_9604 ;
    wire new_AGEMA_signal_9605 ;
    wire new_AGEMA_signal_9606 ;
    wire new_AGEMA_signal_9607 ;
    wire new_AGEMA_signal_9608 ;
    wire new_AGEMA_signal_9609 ;
    wire new_AGEMA_signal_9610 ;
    wire new_AGEMA_signal_9611 ;
    wire new_AGEMA_signal_9612 ;
    wire new_AGEMA_signal_9613 ;
    wire new_AGEMA_signal_9614 ;
    wire new_AGEMA_signal_9615 ;
    wire new_AGEMA_signal_9616 ;
    wire new_AGEMA_signal_9617 ;
    wire new_AGEMA_signal_9618 ;
    wire new_AGEMA_signal_9619 ;
    wire new_AGEMA_signal_9620 ;
    wire new_AGEMA_signal_9621 ;
    wire new_AGEMA_signal_9622 ;
    wire new_AGEMA_signal_9623 ;
    wire new_AGEMA_signal_9624 ;
    wire new_AGEMA_signal_9625 ;
    wire new_AGEMA_signal_9626 ;
    wire new_AGEMA_signal_9627 ;
    wire new_AGEMA_signal_9628 ;
    wire new_AGEMA_signal_9629 ;
    wire new_AGEMA_signal_9630 ;
    wire new_AGEMA_signal_9631 ;
    wire new_AGEMA_signal_9632 ;
    wire new_AGEMA_signal_9633 ;
    wire new_AGEMA_signal_9634 ;
    wire new_AGEMA_signal_9635 ;
    wire new_AGEMA_signal_9636 ;
    wire new_AGEMA_signal_9637 ;
    wire new_AGEMA_signal_9638 ;
    wire new_AGEMA_signal_9639 ;
    wire new_AGEMA_signal_9640 ;
    wire new_AGEMA_signal_9641 ;
    wire new_AGEMA_signal_9642 ;
    wire new_AGEMA_signal_9643 ;
    wire new_AGEMA_signal_9644 ;
    wire new_AGEMA_signal_9645 ;
    wire new_AGEMA_signal_9646 ;
    wire new_AGEMA_signal_9647 ;
    wire new_AGEMA_signal_9648 ;
    wire new_AGEMA_signal_9649 ;
    wire new_AGEMA_signal_9650 ;
    wire new_AGEMA_signal_9651 ;
    wire new_AGEMA_signal_9652 ;
    wire new_AGEMA_signal_9653 ;
    wire new_AGEMA_signal_9654 ;
    wire new_AGEMA_signal_9655 ;
    wire new_AGEMA_signal_9656 ;
    wire new_AGEMA_signal_9657 ;
    wire new_AGEMA_signal_9658 ;
    wire new_AGEMA_signal_9659 ;
    wire new_AGEMA_signal_9660 ;
    wire new_AGEMA_signal_9661 ;
    wire new_AGEMA_signal_9662 ;
    wire new_AGEMA_signal_9663 ;
    wire new_AGEMA_signal_9664 ;
    wire new_AGEMA_signal_9665 ;
    wire new_AGEMA_signal_9666 ;
    wire new_AGEMA_signal_9667 ;
    wire new_AGEMA_signal_9668 ;
    wire new_AGEMA_signal_9669 ;
    wire new_AGEMA_signal_9670 ;
    wire new_AGEMA_signal_9671 ;
    wire new_AGEMA_signal_9672 ;
    wire new_AGEMA_signal_9673 ;
    wire new_AGEMA_signal_9674 ;
    wire new_AGEMA_signal_9675 ;
    wire new_AGEMA_signal_9676 ;
    wire new_AGEMA_signal_9677 ;
    wire new_AGEMA_signal_9678 ;
    wire new_AGEMA_signal_9679 ;
    wire new_AGEMA_signal_9680 ;
    wire new_AGEMA_signal_9681 ;
    wire new_AGEMA_signal_9682 ;
    wire new_AGEMA_signal_9683 ;
    wire new_AGEMA_signal_9684 ;
    wire new_AGEMA_signal_9685 ;
    wire new_AGEMA_signal_9686 ;
    wire new_AGEMA_signal_9687 ;
    wire new_AGEMA_signal_9688 ;
    wire new_AGEMA_signal_9689 ;
    wire new_AGEMA_signal_9690 ;
    wire new_AGEMA_signal_9691 ;
    wire new_AGEMA_signal_9692 ;
    wire new_AGEMA_signal_9693 ;
    wire new_AGEMA_signal_9694 ;
    wire new_AGEMA_signal_9695 ;
    wire new_AGEMA_signal_9696 ;
    wire new_AGEMA_signal_9697 ;
    wire new_AGEMA_signal_9698 ;
    wire new_AGEMA_signal_9699 ;
    wire new_AGEMA_signal_9700 ;
    wire new_AGEMA_signal_9701 ;
    wire new_AGEMA_signal_9702 ;
    wire new_AGEMA_signal_9703 ;
    wire new_AGEMA_signal_9704 ;
    wire new_AGEMA_signal_9705 ;
    wire new_AGEMA_signal_9706 ;
    wire new_AGEMA_signal_9707 ;
    wire new_AGEMA_signal_9708 ;
    wire new_AGEMA_signal_9709 ;
    wire new_AGEMA_signal_9710 ;
    wire new_AGEMA_signal_9711 ;
    wire new_AGEMA_signal_9712 ;
    wire new_AGEMA_signal_9713 ;
    wire new_AGEMA_signal_9714 ;
    wire new_AGEMA_signal_9715 ;
    wire new_AGEMA_signal_9716 ;
    wire new_AGEMA_signal_9717 ;
    wire new_AGEMA_signal_9718 ;
    wire new_AGEMA_signal_9719 ;
    wire new_AGEMA_signal_9720 ;
    wire new_AGEMA_signal_9721 ;
    wire new_AGEMA_signal_9722 ;
    wire new_AGEMA_signal_9723 ;
    wire new_AGEMA_signal_9724 ;
    wire new_AGEMA_signal_9725 ;
    wire new_AGEMA_signal_9726 ;
    wire new_AGEMA_signal_9727 ;
    wire new_AGEMA_signal_9728 ;
    wire new_AGEMA_signal_9729 ;
    wire new_AGEMA_signal_9730 ;
    wire new_AGEMA_signal_9731 ;
    wire new_AGEMA_signal_9732 ;
    wire new_AGEMA_signal_9733 ;
    wire new_AGEMA_signal_9734 ;
    wire new_AGEMA_signal_9735 ;
    wire new_AGEMA_signal_9736 ;
    wire new_AGEMA_signal_9737 ;
    wire new_AGEMA_signal_9738 ;
    wire new_AGEMA_signal_9739 ;
    wire new_AGEMA_signal_9740 ;
    wire new_AGEMA_signal_9741 ;
    wire new_AGEMA_signal_9742 ;
    wire new_AGEMA_signal_9743 ;
    wire new_AGEMA_signal_9744 ;
    wire new_AGEMA_signal_9745 ;
    wire new_AGEMA_signal_9746 ;
    wire new_AGEMA_signal_9747 ;
    wire new_AGEMA_signal_9748 ;
    wire new_AGEMA_signal_9749 ;
    wire new_AGEMA_signal_9750 ;
    wire new_AGEMA_signal_9751 ;
    wire new_AGEMA_signal_9752 ;
    wire new_AGEMA_signal_9753 ;
    wire new_AGEMA_signal_9754 ;
    wire new_AGEMA_signal_9755 ;
    wire new_AGEMA_signal_9756 ;
    wire new_AGEMA_signal_9757 ;
    wire new_AGEMA_signal_9758 ;
    wire new_AGEMA_signal_9759 ;
    wire new_AGEMA_signal_9760 ;
    wire new_AGEMA_signal_9761 ;
    wire new_AGEMA_signal_9762 ;
    wire new_AGEMA_signal_9763 ;
    wire new_AGEMA_signal_9764 ;
    wire new_AGEMA_signal_9765 ;
    wire new_AGEMA_signal_9766 ;
    wire new_AGEMA_signal_9767 ;
    wire new_AGEMA_signal_9768 ;
    wire new_AGEMA_signal_9769 ;
    wire new_AGEMA_signal_9770 ;
    wire new_AGEMA_signal_9771 ;
    wire new_AGEMA_signal_9772 ;
    wire new_AGEMA_signal_9773 ;
    wire new_AGEMA_signal_9774 ;
    wire new_AGEMA_signal_9775 ;
    wire new_AGEMA_signal_9776 ;
    wire new_AGEMA_signal_9777 ;
    wire new_AGEMA_signal_9778 ;
    wire new_AGEMA_signal_9779 ;
    wire new_AGEMA_signal_9780 ;
    wire new_AGEMA_signal_9781 ;
    wire new_AGEMA_signal_9782 ;
    wire new_AGEMA_signal_9783 ;
    wire new_AGEMA_signal_9784 ;
    wire new_AGEMA_signal_9785 ;
    wire new_AGEMA_signal_9786 ;
    wire new_AGEMA_signal_9787 ;
    wire new_AGEMA_signal_9788 ;
    wire new_AGEMA_signal_9789 ;
    wire new_AGEMA_signal_9790 ;
    wire new_AGEMA_signal_9791 ;
    wire new_AGEMA_signal_9792 ;
    wire new_AGEMA_signal_9793 ;
    wire new_AGEMA_signal_9794 ;
    wire new_AGEMA_signal_9795 ;
    wire new_AGEMA_signal_9796 ;
    wire new_AGEMA_signal_9797 ;
    wire new_AGEMA_signal_9798 ;
    wire new_AGEMA_signal_9799 ;
    wire new_AGEMA_signal_9800 ;
    wire new_AGEMA_signal_9801 ;
    wire new_AGEMA_signal_9802 ;
    wire new_AGEMA_signal_9803 ;
    wire new_AGEMA_signal_9804 ;
    wire new_AGEMA_signal_9805 ;
    wire new_AGEMA_signal_9806 ;
    wire new_AGEMA_signal_9807 ;
    wire new_AGEMA_signal_9808 ;
    wire new_AGEMA_signal_9809 ;
    wire new_AGEMA_signal_9810 ;
    wire new_AGEMA_signal_9811 ;
    wire new_AGEMA_signal_9812 ;
    wire new_AGEMA_signal_9813 ;
    wire new_AGEMA_signal_9814 ;
    wire new_AGEMA_signal_9815 ;
    wire new_AGEMA_signal_9816 ;
    wire new_AGEMA_signal_9817 ;
    wire new_AGEMA_signal_9818 ;
    wire new_AGEMA_signal_9819 ;
    wire new_AGEMA_signal_9820 ;
    wire new_AGEMA_signal_9821 ;
    wire new_AGEMA_signal_9822 ;
    wire new_AGEMA_signal_9823 ;
    wire new_AGEMA_signal_9824 ;
    wire new_AGEMA_signal_9825 ;
    wire new_AGEMA_signal_9826 ;
    wire new_AGEMA_signal_9827 ;
    wire new_AGEMA_signal_9828 ;
    wire new_AGEMA_signal_9829 ;
    wire new_AGEMA_signal_9830 ;
    wire new_AGEMA_signal_9831 ;
    wire new_AGEMA_signal_9832 ;
    wire new_AGEMA_signal_9833 ;
    wire new_AGEMA_signal_9834 ;
    wire new_AGEMA_signal_9835 ;
    wire new_AGEMA_signal_9836 ;
    wire new_AGEMA_signal_9837 ;
    wire new_AGEMA_signal_9838 ;
    wire new_AGEMA_signal_9839 ;
    wire new_AGEMA_signal_9840 ;
    wire new_AGEMA_signal_9841 ;
    wire new_AGEMA_signal_9842 ;
    wire new_AGEMA_signal_9843 ;
    wire new_AGEMA_signal_9844 ;
    wire new_AGEMA_signal_9845 ;
    wire new_AGEMA_signal_9846 ;
    wire new_AGEMA_signal_9847 ;
    wire new_AGEMA_signal_9848 ;
    wire new_AGEMA_signal_9849 ;
    wire new_AGEMA_signal_9850 ;
    wire new_AGEMA_signal_9851 ;
    wire new_AGEMA_signal_9852 ;
    wire new_AGEMA_signal_9853 ;
    wire new_AGEMA_signal_9854 ;
    wire new_AGEMA_signal_9855 ;
    wire new_AGEMA_signal_9856 ;
    wire new_AGEMA_signal_9857 ;
    wire new_AGEMA_signal_9858 ;
    wire new_AGEMA_signal_9859 ;
    wire new_AGEMA_signal_9860 ;
    wire new_AGEMA_signal_9861 ;
    wire new_AGEMA_signal_9862 ;
    wire new_AGEMA_signal_9863 ;
    wire new_AGEMA_signal_9864 ;
    wire new_AGEMA_signal_9865 ;
    wire new_AGEMA_signal_9866 ;
    wire new_AGEMA_signal_9867 ;
    wire new_AGEMA_signal_9868 ;
    wire new_AGEMA_signal_9869 ;
    wire new_AGEMA_signal_9870 ;
    wire new_AGEMA_signal_9871 ;
    wire new_AGEMA_signal_9872 ;
    wire new_AGEMA_signal_9873 ;
    wire new_AGEMA_signal_9874 ;
    wire new_AGEMA_signal_9875 ;
    wire new_AGEMA_signal_9876 ;
    wire new_AGEMA_signal_9877 ;
    wire new_AGEMA_signal_9878 ;
    wire new_AGEMA_signal_9879 ;
    wire new_AGEMA_signal_9880 ;
    wire new_AGEMA_signal_9881 ;
    wire new_AGEMA_signal_9882 ;
    wire new_AGEMA_signal_9883 ;
    wire new_AGEMA_signal_9884 ;
    wire new_AGEMA_signal_9885 ;
    wire new_AGEMA_signal_9886 ;
    wire new_AGEMA_signal_9887 ;
    wire new_AGEMA_signal_9888 ;
    wire new_AGEMA_signal_9889 ;
    wire new_AGEMA_signal_9890 ;
    wire new_AGEMA_signal_9891 ;
    wire new_AGEMA_signal_9892 ;
    wire new_AGEMA_signal_9893 ;
    wire new_AGEMA_signal_9894 ;
    wire new_AGEMA_signal_9895 ;
    wire new_AGEMA_signal_9896 ;
    wire new_AGEMA_signal_9897 ;
    wire new_AGEMA_signal_9898 ;
    wire new_AGEMA_signal_9899 ;
    wire new_AGEMA_signal_9900 ;
    wire new_AGEMA_signal_9901 ;
    wire new_AGEMA_signal_9902 ;
    wire new_AGEMA_signal_9903 ;
    wire new_AGEMA_signal_9904 ;
    wire new_AGEMA_signal_9905 ;
    wire new_AGEMA_signal_9906 ;
    wire new_AGEMA_signal_9907 ;
    wire new_AGEMA_signal_9908 ;
    wire new_AGEMA_signal_9909 ;
    wire new_AGEMA_signal_9910 ;
    wire new_AGEMA_signal_9911 ;
    wire new_AGEMA_signal_9912 ;
    wire new_AGEMA_signal_9913 ;
    wire new_AGEMA_signal_9914 ;
    wire new_AGEMA_signal_9915 ;
    wire new_AGEMA_signal_9916 ;
    wire new_AGEMA_signal_9917 ;
    wire new_AGEMA_signal_9918 ;
    wire new_AGEMA_signal_9919 ;
    wire new_AGEMA_signal_9920 ;
    wire new_AGEMA_signal_9921 ;
    wire new_AGEMA_signal_9922 ;
    wire new_AGEMA_signal_9923 ;
    wire new_AGEMA_signal_9924 ;
    wire new_AGEMA_signal_9925 ;
    wire new_AGEMA_signal_9926 ;
    wire new_AGEMA_signal_9927 ;
    wire new_AGEMA_signal_9928 ;
    wire new_AGEMA_signal_9929 ;
    wire new_AGEMA_signal_9930 ;
    wire new_AGEMA_signal_9931 ;
    wire new_AGEMA_signal_9932 ;
    wire new_AGEMA_signal_9933 ;
    wire new_AGEMA_signal_9934 ;
    wire new_AGEMA_signal_9935 ;
    wire new_AGEMA_signal_9936 ;
    wire new_AGEMA_signal_9937 ;
    wire new_AGEMA_signal_9938 ;
    wire new_AGEMA_signal_9939 ;
    wire new_AGEMA_signal_9940 ;
    wire new_AGEMA_signal_9941 ;
    wire new_AGEMA_signal_9942 ;
    wire new_AGEMA_signal_9943 ;
    wire new_AGEMA_signal_9944 ;
    wire new_AGEMA_signal_9945 ;
    wire new_AGEMA_signal_9946 ;
    wire new_AGEMA_signal_9947 ;
    wire new_AGEMA_signal_9948 ;
    wire new_AGEMA_signal_9949 ;
    wire new_AGEMA_signal_9950 ;
    wire new_AGEMA_signal_9951 ;
    wire new_AGEMA_signal_9952 ;
    wire new_AGEMA_signal_9953 ;
    wire new_AGEMA_signal_9954 ;
    wire new_AGEMA_signal_9955 ;
    wire new_AGEMA_signal_9956 ;
    wire new_AGEMA_signal_9957 ;
    wire new_AGEMA_signal_9958 ;
    wire new_AGEMA_signal_9959 ;
    wire new_AGEMA_signal_9960 ;
    wire new_AGEMA_signal_9961 ;
    wire new_AGEMA_signal_9962 ;
    wire new_AGEMA_signal_9963 ;
    wire new_AGEMA_signal_9964 ;
    wire new_AGEMA_signal_9965 ;
    wire new_AGEMA_signal_9966 ;
    wire new_AGEMA_signal_9967 ;
    wire new_AGEMA_signal_9968 ;
    wire new_AGEMA_signal_9969 ;
    wire new_AGEMA_signal_9970 ;
    wire new_AGEMA_signal_9971 ;
    wire new_AGEMA_signal_9972 ;
    wire new_AGEMA_signal_9973 ;
    wire new_AGEMA_signal_9974 ;
    wire new_AGEMA_signal_9975 ;
    wire new_AGEMA_signal_9976 ;
    wire new_AGEMA_signal_9977 ;
    wire new_AGEMA_signal_9978 ;
    wire new_AGEMA_signal_9979 ;
    wire new_AGEMA_signal_9980 ;
    wire new_AGEMA_signal_9981 ;
    wire new_AGEMA_signal_9982 ;
    wire new_AGEMA_signal_9983 ;
    wire new_AGEMA_signal_9984 ;
    wire new_AGEMA_signal_9985 ;
    wire new_AGEMA_signal_9986 ;
    wire new_AGEMA_signal_9987 ;
    wire new_AGEMA_signal_9988 ;
    wire new_AGEMA_signal_9989 ;
    wire new_AGEMA_signal_9990 ;
    wire new_AGEMA_signal_9991 ;
    wire new_AGEMA_signal_9992 ;
    wire new_AGEMA_signal_9993 ;
    wire new_AGEMA_signal_9994 ;
    wire new_AGEMA_signal_9995 ;
    wire new_AGEMA_signal_9996 ;
    wire new_AGEMA_signal_9997 ;
    wire new_AGEMA_signal_9998 ;
    wire new_AGEMA_signal_9999 ;
    wire new_AGEMA_signal_10000 ;
    wire new_AGEMA_signal_10001 ;
    wire new_AGEMA_signal_10002 ;
    wire new_AGEMA_signal_10003 ;
    wire new_AGEMA_signal_10004 ;
    wire new_AGEMA_signal_10005 ;
    wire new_AGEMA_signal_10006 ;
    wire new_AGEMA_signal_10007 ;
    wire new_AGEMA_signal_10008 ;
    wire new_AGEMA_signal_10009 ;
    wire new_AGEMA_signal_10010 ;
    wire new_AGEMA_signal_10011 ;
    wire new_AGEMA_signal_10012 ;
    wire new_AGEMA_signal_10013 ;
    wire new_AGEMA_signal_10014 ;
    wire new_AGEMA_signal_10015 ;
    wire new_AGEMA_signal_10016 ;
    wire new_AGEMA_signal_10017 ;
    wire new_AGEMA_signal_10018 ;
    wire new_AGEMA_signal_10019 ;
    wire new_AGEMA_signal_10020 ;
    wire new_AGEMA_signal_10021 ;
    wire new_AGEMA_signal_10022 ;
    wire new_AGEMA_signal_10023 ;
    wire new_AGEMA_signal_10024 ;
    wire new_AGEMA_signal_10025 ;
    wire new_AGEMA_signal_10026 ;
    wire new_AGEMA_signal_10027 ;
    wire new_AGEMA_signal_10028 ;
    wire new_AGEMA_signal_10029 ;
    wire new_AGEMA_signal_10030 ;
    wire new_AGEMA_signal_10031 ;
    wire new_AGEMA_signal_10032 ;
    wire new_AGEMA_signal_10033 ;
    wire new_AGEMA_signal_10034 ;
    wire new_AGEMA_signal_10035 ;
    wire new_AGEMA_signal_10036 ;
    wire new_AGEMA_signal_10037 ;
    wire new_AGEMA_signal_10038 ;
    wire new_AGEMA_signal_10039 ;
    wire new_AGEMA_signal_10040 ;
    wire new_AGEMA_signal_10041 ;
    wire new_AGEMA_signal_10042 ;
    wire new_AGEMA_signal_10043 ;
    wire new_AGEMA_signal_10044 ;
    wire new_AGEMA_signal_10045 ;
    wire new_AGEMA_signal_10046 ;
    wire new_AGEMA_signal_10047 ;
    wire new_AGEMA_signal_10048 ;
    wire new_AGEMA_signal_10049 ;
    wire new_AGEMA_signal_10050 ;
    wire new_AGEMA_signal_10051 ;
    wire new_AGEMA_signal_10052 ;
    wire new_AGEMA_signal_10053 ;
    wire new_AGEMA_signal_10054 ;
    wire new_AGEMA_signal_10055 ;
    wire new_AGEMA_signal_10056 ;
    wire new_AGEMA_signal_10057 ;
    wire new_AGEMA_signal_10058 ;
    wire new_AGEMA_signal_10059 ;
    wire new_AGEMA_signal_10060 ;
    wire new_AGEMA_signal_10061 ;
    wire new_AGEMA_signal_10062 ;
    wire new_AGEMA_signal_10063 ;
    wire new_AGEMA_signal_10064 ;
    wire new_AGEMA_signal_10065 ;
    wire new_AGEMA_signal_10066 ;
    wire new_AGEMA_signal_10067 ;
    wire new_AGEMA_signal_10068 ;
    wire new_AGEMA_signal_10069 ;
    wire new_AGEMA_signal_10070 ;
    wire new_AGEMA_signal_10071 ;
    wire new_AGEMA_signal_10072 ;
    wire new_AGEMA_signal_10073 ;
    wire new_AGEMA_signal_10074 ;
    wire new_AGEMA_signal_10075 ;
    wire new_AGEMA_signal_10076 ;
    wire new_AGEMA_signal_10077 ;
    wire new_AGEMA_signal_10078 ;
    wire new_AGEMA_signal_10079 ;
    wire new_AGEMA_signal_10080 ;
    wire new_AGEMA_signal_10081 ;
    wire new_AGEMA_signal_10082 ;
    wire new_AGEMA_signal_10083 ;
    wire new_AGEMA_signal_10084 ;
    wire new_AGEMA_signal_10085 ;
    wire new_AGEMA_signal_10086 ;
    wire new_AGEMA_signal_10087 ;
    wire new_AGEMA_signal_10088 ;
    wire new_AGEMA_signal_10089 ;
    wire new_AGEMA_signal_10090 ;
    wire new_AGEMA_signal_10091 ;
    wire new_AGEMA_signal_10092 ;
    wire new_AGEMA_signal_10093 ;
    wire new_AGEMA_signal_10094 ;
    wire new_AGEMA_signal_10095 ;
    wire new_AGEMA_signal_10096 ;
    wire new_AGEMA_signal_10097 ;
    wire new_AGEMA_signal_10098 ;
    wire new_AGEMA_signal_10099 ;
    wire new_AGEMA_signal_10100 ;
    wire new_AGEMA_signal_10101 ;
    wire new_AGEMA_signal_10102 ;
    wire new_AGEMA_signal_10103 ;
    wire new_AGEMA_signal_10104 ;
    wire new_AGEMA_signal_10105 ;
    wire new_AGEMA_signal_10106 ;
    wire new_AGEMA_signal_10107 ;
    wire new_AGEMA_signal_10108 ;
    wire new_AGEMA_signal_10109 ;
    wire new_AGEMA_signal_10110 ;
    wire new_AGEMA_signal_10111 ;
    wire new_AGEMA_signal_10112 ;
    wire new_AGEMA_signal_10113 ;
    wire new_AGEMA_signal_10114 ;
    wire new_AGEMA_signal_10115 ;
    wire new_AGEMA_signal_10116 ;
    wire new_AGEMA_signal_10117 ;
    wire new_AGEMA_signal_10118 ;
    wire new_AGEMA_signal_10119 ;
    wire new_AGEMA_signal_10120 ;
    wire new_AGEMA_signal_10121 ;
    wire new_AGEMA_signal_10122 ;
    wire new_AGEMA_signal_10123 ;
    wire new_AGEMA_signal_10124 ;
    wire new_AGEMA_signal_10125 ;
    wire new_AGEMA_signal_10126 ;
    wire new_AGEMA_signal_10127 ;
    wire new_AGEMA_signal_10128 ;
    wire new_AGEMA_signal_10129 ;
    wire new_AGEMA_signal_10130 ;
    wire new_AGEMA_signal_10131 ;
    wire new_AGEMA_signal_10132 ;
    wire new_AGEMA_signal_10133 ;
    wire new_AGEMA_signal_10134 ;
    wire new_AGEMA_signal_10135 ;
    wire new_AGEMA_signal_10136 ;
    wire new_AGEMA_signal_10137 ;
    wire new_AGEMA_signal_10138 ;
    wire new_AGEMA_signal_10139 ;
    wire new_AGEMA_signal_10140 ;
    wire new_AGEMA_signal_10141 ;
    wire new_AGEMA_signal_10142 ;
    wire new_AGEMA_signal_10143 ;
    wire new_AGEMA_signal_10144 ;
    wire new_AGEMA_signal_10145 ;
    wire new_AGEMA_signal_10146 ;
    wire new_AGEMA_signal_10147 ;
    wire new_AGEMA_signal_10148 ;
    wire new_AGEMA_signal_10149 ;
    wire new_AGEMA_signal_10150 ;
    wire new_AGEMA_signal_10151 ;
    wire new_AGEMA_signal_10152 ;
    wire new_AGEMA_signal_10153 ;
    wire new_AGEMA_signal_10154 ;
    wire new_AGEMA_signal_10155 ;
    wire new_AGEMA_signal_10156 ;
    wire new_AGEMA_signal_10157 ;
    wire new_AGEMA_signal_10158 ;
    wire new_AGEMA_signal_10159 ;
    wire new_AGEMA_signal_10160 ;
    wire new_AGEMA_signal_10161 ;
    wire new_AGEMA_signal_10162 ;
    wire new_AGEMA_signal_10163 ;
    wire new_AGEMA_signal_10164 ;
    wire new_AGEMA_signal_10165 ;
    wire new_AGEMA_signal_10166 ;
    wire new_AGEMA_signal_10167 ;
    wire new_AGEMA_signal_10168 ;
    wire new_AGEMA_signal_10169 ;
    wire new_AGEMA_signal_10170 ;
    wire new_AGEMA_signal_10171 ;
    wire new_AGEMA_signal_10172 ;
    wire new_AGEMA_signal_10173 ;
    wire new_AGEMA_signal_10174 ;
    wire new_AGEMA_signal_10175 ;
    wire new_AGEMA_signal_10176 ;
    wire new_AGEMA_signal_10177 ;
    wire new_AGEMA_signal_10178 ;
    wire new_AGEMA_signal_10179 ;
    wire new_AGEMA_signal_10180 ;
    wire new_AGEMA_signal_10181 ;
    wire new_AGEMA_signal_10182 ;
    wire new_AGEMA_signal_10183 ;
    wire new_AGEMA_signal_10184 ;
    wire new_AGEMA_signal_10185 ;
    wire new_AGEMA_signal_10186 ;
    wire new_AGEMA_signal_10187 ;
    wire new_AGEMA_signal_10188 ;
    wire new_AGEMA_signal_10189 ;
    wire new_AGEMA_signal_10190 ;
    wire new_AGEMA_signal_10191 ;
    wire new_AGEMA_signal_10192 ;
    wire new_AGEMA_signal_10193 ;
    wire new_AGEMA_signal_10194 ;
    wire new_AGEMA_signal_10195 ;
    wire new_AGEMA_signal_10196 ;
    wire new_AGEMA_signal_10197 ;
    wire new_AGEMA_signal_10198 ;
    wire new_AGEMA_signal_10199 ;
    wire new_AGEMA_signal_10200 ;
    wire new_AGEMA_signal_10201 ;
    wire new_AGEMA_signal_10202 ;
    wire new_AGEMA_signal_10203 ;
    wire new_AGEMA_signal_10204 ;
    wire new_AGEMA_signal_10205 ;
    wire new_AGEMA_signal_10206 ;
    wire new_AGEMA_signal_10207 ;
    wire new_AGEMA_signal_10208 ;
    wire new_AGEMA_signal_10209 ;
    wire new_AGEMA_signal_10210 ;
    wire new_AGEMA_signal_10211 ;
    wire new_AGEMA_signal_10212 ;
    wire new_AGEMA_signal_10213 ;
    wire new_AGEMA_signal_10214 ;
    wire new_AGEMA_signal_10215 ;
    wire new_AGEMA_signal_10216 ;
    wire new_AGEMA_signal_10217 ;
    wire new_AGEMA_signal_10218 ;
    wire new_AGEMA_signal_10219 ;
    wire new_AGEMA_signal_10220 ;
    wire new_AGEMA_signal_10221 ;
    wire new_AGEMA_signal_10222 ;
    wire new_AGEMA_signal_10223 ;
    wire new_AGEMA_signal_10224 ;
    wire new_AGEMA_signal_10225 ;
    wire new_AGEMA_signal_10226 ;
    wire new_AGEMA_signal_10227 ;
    wire new_AGEMA_signal_10228 ;
    wire new_AGEMA_signal_10229 ;
    wire new_AGEMA_signal_10230 ;
    wire new_AGEMA_signal_10231 ;
    wire new_AGEMA_signal_10232 ;
    wire new_AGEMA_signal_10233 ;
    wire new_AGEMA_signal_10234 ;
    wire new_AGEMA_signal_10235 ;
    wire new_AGEMA_signal_10236 ;
    wire new_AGEMA_signal_10237 ;
    wire new_AGEMA_signal_10238 ;
    wire new_AGEMA_signal_10239 ;
    wire new_AGEMA_signal_10240 ;
    wire new_AGEMA_signal_10241 ;
    wire new_AGEMA_signal_10242 ;
    wire new_AGEMA_signal_10243 ;
    wire new_AGEMA_signal_10244 ;
    wire new_AGEMA_signal_10245 ;
    wire new_AGEMA_signal_10246 ;
    wire new_AGEMA_signal_10247 ;
    wire new_AGEMA_signal_10248 ;
    wire new_AGEMA_signal_10249 ;
    wire new_AGEMA_signal_10250 ;
    wire new_AGEMA_signal_10251 ;
    wire new_AGEMA_signal_10252 ;
    wire new_AGEMA_signal_10253 ;
    wire new_AGEMA_signal_10254 ;
    wire new_AGEMA_signal_10255 ;
    wire new_AGEMA_signal_10256 ;
    wire new_AGEMA_signal_10257 ;
    wire new_AGEMA_signal_10258 ;
    wire new_AGEMA_signal_10259 ;
    wire new_AGEMA_signal_10260 ;
    wire new_AGEMA_signal_10261 ;
    wire new_AGEMA_signal_10262 ;
    wire new_AGEMA_signal_10263 ;
    wire new_AGEMA_signal_10264 ;
    wire new_AGEMA_signal_10265 ;
    wire new_AGEMA_signal_10266 ;
    wire new_AGEMA_signal_10267 ;
    wire new_AGEMA_signal_10268 ;
    wire new_AGEMA_signal_10269 ;
    wire new_AGEMA_signal_10270 ;
    wire new_AGEMA_signal_10271 ;
    wire new_AGEMA_signal_10272 ;
    wire new_AGEMA_signal_10273 ;
    wire new_AGEMA_signal_10274 ;
    wire new_AGEMA_signal_10275 ;
    wire new_AGEMA_signal_10276 ;
    wire new_AGEMA_signal_10277 ;
    wire new_AGEMA_signal_10278 ;
    wire new_AGEMA_signal_10279 ;
    wire new_AGEMA_signal_10280 ;
    wire new_AGEMA_signal_10281 ;
    wire new_AGEMA_signal_10282 ;
    wire new_AGEMA_signal_10283 ;
    wire new_AGEMA_signal_10284 ;
    wire new_AGEMA_signal_10285 ;
    wire new_AGEMA_signal_10286 ;
    wire new_AGEMA_signal_10287 ;
    wire new_AGEMA_signal_10288 ;
    wire new_AGEMA_signal_10289 ;
    wire new_AGEMA_signal_10290 ;
    wire new_AGEMA_signal_10291 ;
    wire new_AGEMA_signal_10292 ;
    wire new_AGEMA_signal_10293 ;
    wire new_AGEMA_signal_10294 ;
    wire new_AGEMA_signal_10295 ;
    wire new_AGEMA_signal_10296 ;
    wire new_AGEMA_signal_10297 ;
    wire new_AGEMA_signal_10298 ;
    wire new_AGEMA_signal_10299 ;
    wire new_AGEMA_signal_10300 ;
    wire new_AGEMA_signal_10301 ;
    wire new_AGEMA_signal_10302 ;
    wire new_AGEMA_signal_10303 ;
    wire new_AGEMA_signal_10304 ;
    wire new_AGEMA_signal_10305 ;
    wire new_AGEMA_signal_10306 ;
    wire new_AGEMA_signal_10307 ;
    wire new_AGEMA_signal_10308 ;
    wire new_AGEMA_signal_10309 ;
    wire new_AGEMA_signal_10310 ;
    wire new_AGEMA_signal_10311 ;
    wire new_AGEMA_signal_10312 ;
    wire new_AGEMA_signal_10313 ;
    wire new_AGEMA_signal_10314 ;
    wire new_AGEMA_signal_10315 ;
    wire new_AGEMA_signal_10316 ;
    wire new_AGEMA_signal_10317 ;
    wire new_AGEMA_signal_10318 ;
    wire new_AGEMA_signal_10319 ;
    wire new_AGEMA_signal_10320 ;
    wire new_AGEMA_signal_10321 ;
    wire new_AGEMA_signal_10322 ;
    wire new_AGEMA_signal_10323 ;
    wire new_AGEMA_signal_10324 ;
    wire new_AGEMA_signal_10325 ;
    wire new_AGEMA_signal_10326 ;
    wire new_AGEMA_signal_10327 ;
    wire new_AGEMA_signal_10328 ;
    wire new_AGEMA_signal_10329 ;
    wire new_AGEMA_signal_10330 ;
    wire new_AGEMA_signal_10331 ;
    wire new_AGEMA_signal_10332 ;
    wire new_AGEMA_signal_10333 ;
    wire new_AGEMA_signal_10334 ;
    wire new_AGEMA_signal_10335 ;
    wire new_AGEMA_signal_10336 ;
    wire new_AGEMA_signal_10337 ;
    wire new_AGEMA_signal_10338 ;
    wire new_AGEMA_signal_10339 ;
    wire new_AGEMA_signal_10340 ;
    wire new_AGEMA_signal_10341 ;
    wire new_AGEMA_signal_10342 ;
    wire new_AGEMA_signal_10343 ;
    wire new_AGEMA_signal_10344 ;
    wire new_AGEMA_signal_10345 ;
    wire new_AGEMA_signal_10346 ;
    wire new_AGEMA_signal_10347 ;
    wire new_AGEMA_signal_10348 ;
    wire new_AGEMA_signal_10349 ;
    wire new_AGEMA_signal_10350 ;
    wire new_AGEMA_signal_10351 ;
    wire new_AGEMA_signal_10352 ;
    wire new_AGEMA_signal_10353 ;
    wire new_AGEMA_signal_10354 ;
    wire new_AGEMA_signal_10355 ;
    wire new_AGEMA_signal_10356 ;
    wire new_AGEMA_signal_10357 ;
    wire new_AGEMA_signal_10358 ;
    wire new_AGEMA_signal_10359 ;
    wire new_AGEMA_signal_10360 ;
    wire new_AGEMA_signal_10361 ;
    wire new_AGEMA_signal_10362 ;
    wire new_AGEMA_signal_10363 ;
    wire new_AGEMA_signal_10364 ;
    wire new_AGEMA_signal_10365 ;
    wire new_AGEMA_signal_10366 ;
    wire new_AGEMA_signal_10367 ;
    wire new_AGEMA_signal_10368 ;
    wire new_AGEMA_signal_10369 ;
    wire new_AGEMA_signal_10370 ;
    wire new_AGEMA_signal_10371 ;
    wire new_AGEMA_signal_10372 ;
    wire new_AGEMA_signal_10373 ;
    wire new_AGEMA_signal_10374 ;
    wire new_AGEMA_signal_10375 ;
    wire new_AGEMA_signal_10376 ;
    wire new_AGEMA_signal_10377 ;
    wire new_AGEMA_signal_10378 ;
    wire new_AGEMA_signal_10379 ;
    wire new_AGEMA_signal_10380 ;
    wire new_AGEMA_signal_10381 ;
    wire new_AGEMA_signal_10382 ;
    wire new_AGEMA_signal_10383 ;
    wire new_AGEMA_signal_10384 ;
    wire new_AGEMA_signal_10385 ;
    wire new_AGEMA_signal_10386 ;
    wire new_AGEMA_signal_10387 ;
    wire new_AGEMA_signal_10388 ;
    wire new_AGEMA_signal_10389 ;
    wire new_AGEMA_signal_10390 ;
    wire new_AGEMA_signal_10391 ;
    wire new_AGEMA_signal_10392 ;
    wire new_AGEMA_signal_10393 ;
    wire new_AGEMA_signal_10394 ;
    wire new_AGEMA_signal_10395 ;
    wire new_AGEMA_signal_10396 ;
    wire new_AGEMA_signal_10397 ;
    wire new_AGEMA_signal_10398 ;
    wire new_AGEMA_signal_10399 ;
    wire new_AGEMA_signal_10400 ;
    wire new_AGEMA_signal_10401 ;
    wire new_AGEMA_signal_10402 ;
    wire new_AGEMA_signal_10403 ;
    wire new_AGEMA_signal_10404 ;
    wire new_AGEMA_signal_10405 ;
    wire new_AGEMA_signal_10406 ;
    wire new_AGEMA_signal_10407 ;
    wire new_AGEMA_signal_10408 ;
    wire new_AGEMA_signal_10409 ;
    wire new_AGEMA_signal_10410 ;
    wire new_AGEMA_signal_10411 ;
    wire new_AGEMA_signal_10412 ;
    wire new_AGEMA_signal_10413 ;
    wire new_AGEMA_signal_10414 ;
    wire new_AGEMA_signal_10415 ;
    wire new_AGEMA_signal_10416 ;
    wire new_AGEMA_signal_10417 ;
    wire new_AGEMA_signal_10418 ;
    wire new_AGEMA_signal_10419 ;
    wire new_AGEMA_signal_10420 ;
    wire new_AGEMA_signal_10421 ;
    wire new_AGEMA_signal_10422 ;
    wire new_AGEMA_signal_10423 ;
    wire new_AGEMA_signal_10424 ;
    wire new_AGEMA_signal_10425 ;
    wire new_AGEMA_signal_10426 ;
    wire new_AGEMA_signal_10427 ;
    wire new_AGEMA_signal_10428 ;
    wire new_AGEMA_signal_10429 ;
    wire new_AGEMA_signal_10430 ;
    wire new_AGEMA_signal_10431 ;
    wire new_AGEMA_signal_10432 ;
    wire new_AGEMA_signal_10433 ;
    wire new_AGEMA_signal_10434 ;
    wire new_AGEMA_signal_10435 ;
    wire new_AGEMA_signal_10436 ;
    wire new_AGEMA_signal_10437 ;
    wire new_AGEMA_signal_10438 ;
    wire new_AGEMA_signal_10439 ;
    wire new_AGEMA_signal_10440 ;
    wire new_AGEMA_signal_10441 ;
    wire new_AGEMA_signal_10442 ;
    wire new_AGEMA_signal_10443 ;
    wire new_AGEMA_signal_10444 ;
    wire new_AGEMA_signal_10447 ;
    wire new_AGEMA_signal_10448 ;
    wire new_AGEMA_signal_10451 ;
    wire new_AGEMA_signal_10452 ;
    wire new_AGEMA_signal_10455 ;
    wire new_AGEMA_signal_10456 ;
    wire new_AGEMA_signal_10457 ;
    wire new_AGEMA_signal_10458 ;
    wire new_AGEMA_signal_10459 ;
    wire new_AGEMA_signal_10460 ;
    wire new_AGEMA_signal_10461 ;
    wire new_AGEMA_signal_10462 ;
    wire new_AGEMA_signal_10463 ;
    wire new_AGEMA_signal_10464 ;
    wire new_AGEMA_signal_10465 ;
    wire new_AGEMA_signal_10466 ;
    wire new_AGEMA_signal_10467 ;
    wire new_AGEMA_signal_10468 ;
    wire new_AGEMA_signal_10469 ;
    wire new_AGEMA_signal_10470 ;
    wire new_AGEMA_signal_10471 ;
    wire new_AGEMA_signal_10472 ;
    wire new_AGEMA_signal_10473 ;
    wire new_AGEMA_signal_10474 ;
    wire new_AGEMA_signal_10475 ;
    wire new_AGEMA_signal_10476 ;
    wire new_AGEMA_signal_10477 ;
    wire new_AGEMA_signal_10478 ;
    wire new_AGEMA_signal_10479 ;
    wire new_AGEMA_signal_10480 ;
    wire new_AGEMA_signal_10481 ;
    wire new_AGEMA_signal_10482 ;
    wire new_AGEMA_signal_10483 ;
    wire new_AGEMA_signal_10484 ;
    wire new_AGEMA_signal_10485 ;
    wire new_AGEMA_signal_10486 ;
    wire new_AGEMA_signal_10487 ;
    wire new_AGEMA_signal_10488 ;
    wire new_AGEMA_signal_10489 ;
    wire new_AGEMA_signal_10490 ;
    wire new_AGEMA_signal_10491 ;
    wire new_AGEMA_signal_10492 ;
    wire new_AGEMA_signal_10493 ;
    wire new_AGEMA_signal_10494 ;
    wire new_AGEMA_signal_10495 ;
    wire new_AGEMA_signal_10496 ;
    wire new_AGEMA_signal_10497 ;
    wire new_AGEMA_signal_10498 ;
    wire new_AGEMA_signal_10499 ;
    wire new_AGEMA_signal_10500 ;
    wire new_AGEMA_signal_10501 ;
    wire new_AGEMA_signal_10502 ;
    wire new_AGEMA_signal_10503 ;
    wire new_AGEMA_signal_10504 ;
    wire new_AGEMA_signal_10505 ;
    wire new_AGEMA_signal_10506 ;
    wire new_AGEMA_signal_10507 ;
    wire new_AGEMA_signal_10508 ;
    wire new_AGEMA_signal_10509 ;
    wire new_AGEMA_signal_10510 ;
    wire new_AGEMA_signal_10511 ;
    wire new_AGEMA_signal_10512 ;
    wire new_AGEMA_signal_10513 ;
    wire new_AGEMA_signal_10514 ;
    wire new_AGEMA_signal_10515 ;
    wire new_AGEMA_signal_10516 ;
    wire new_AGEMA_signal_10517 ;
    wire new_AGEMA_signal_10518 ;
    wire new_AGEMA_signal_10519 ;
    wire new_AGEMA_signal_10520 ;
    wire new_AGEMA_signal_10521 ;
    wire new_AGEMA_signal_10522 ;
    wire new_AGEMA_signal_10523 ;
    wire new_AGEMA_signal_10524 ;
    wire new_AGEMA_signal_10525 ;
    wire new_AGEMA_signal_10526 ;
    wire new_AGEMA_signal_10527 ;
    wire new_AGEMA_signal_10528 ;
    wire new_AGEMA_signal_10529 ;
    wire new_AGEMA_signal_10530 ;
    wire new_AGEMA_signal_10531 ;
    wire new_AGEMA_signal_10532 ;
    wire new_AGEMA_signal_10533 ;
    wire new_AGEMA_signal_10534 ;
    wire new_AGEMA_signal_10535 ;
    wire new_AGEMA_signal_10536 ;
    wire new_AGEMA_signal_10537 ;
    wire new_AGEMA_signal_10538 ;
    wire new_AGEMA_signal_10539 ;
    wire new_AGEMA_signal_10540 ;
    wire new_AGEMA_signal_10541 ;
    wire new_AGEMA_signal_10542 ;
    wire new_AGEMA_signal_10543 ;
    wire new_AGEMA_signal_10544 ;
    wire new_AGEMA_signal_10545 ;
    wire new_AGEMA_signal_10546 ;
    wire new_AGEMA_signal_10547 ;
    wire new_AGEMA_signal_10548 ;
    wire new_AGEMA_signal_10549 ;
    wire new_AGEMA_signal_10550 ;
    wire new_AGEMA_signal_10551 ;
    wire new_AGEMA_signal_10552 ;
    wire new_AGEMA_signal_10553 ;
    wire new_AGEMA_signal_10554 ;
    wire new_AGEMA_signal_10555 ;
    wire new_AGEMA_signal_10556 ;
    wire new_AGEMA_signal_10557 ;
    wire new_AGEMA_signal_10558 ;
    wire new_AGEMA_signal_10559 ;
    wire new_AGEMA_signal_10560 ;
    wire new_AGEMA_signal_10561 ;
    wire new_AGEMA_signal_10562 ;
    wire new_AGEMA_signal_10563 ;
    wire new_AGEMA_signal_10564 ;
    wire new_AGEMA_signal_10565 ;
    wire new_AGEMA_signal_10566 ;
    wire new_AGEMA_signal_10567 ;
    wire new_AGEMA_signal_10568 ;
    wire new_AGEMA_signal_10569 ;
    wire new_AGEMA_signal_10570 ;
    wire new_AGEMA_signal_10571 ;
    wire new_AGEMA_signal_10572 ;
    wire new_AGEMA_signal_10573 ;
    wire new_AGEMA_signal_10574 ;
    wire new_AGEMA_signal_10575 ;
    wire new_AGEMA_signal_10576 ;
    wire new_AGEMA_signal_10577 ;
    wire new_AGEMA_signal_10578 ;
    wire new_AGEMA_signal_10579 ;
    wire new_AGEMA_signal_10580 ;
    wire new_AGEMA_signal_10581 ;
    wire new_AGEMA_signal_10582 ;
    wire new_AGEMA_signal_10583 ;
    wire new_AGEMA_signal_10584 ;
    wire new_AGEMA_signal_10585 ;
    wire new_AGEMA_signal_10586 ;
    wire new_AGEMA_signal_10587 ;
    wire new_AGEMA_signal_10588 ;
    wire new_AGEMA_signal_10589 ;
    wire new_AGEMA_signal_10590 ;
    wire new_AGEMA_signal_10591 ;
    wire new_AGEMA_signal_10592 ;
    wire new_AGEMA_signal_10593 ;
    wire new_AGEMA_signal_10594 ;
    wire new_AGEMA_signal_10595 ;
    wire new_AGEMA_signal_10596 ;
    wire new_AGEMA_signal_10597 ;
    wire new_AGEMA_signal_10598 ;
    wire new_AGEMA_signal_10599 ;
    wire new_AGEMA_signal_10600 ;
    wire new_AGEMA_signal_10601 ;
    wire new_AGEMA_signal_10602 ;
    wire new_AGEMA_signal_10603 ;
    wire new_AGEMA_signal_10604 ;
    wire new_AGEMA_signal_10605 ;
    wire new_AGEMA_signal_10606 ;
    wire new_AGEMA_signal_10607 ;
    wire new_AGEMA_signal_10608 ;
    wire new_AGEMA_signal_10609 ;
    wire new_AGEMA_signal_10610 ;
    wire new_AGEMA_signal_10611 ;
    wire new_AGEMA_signal_10612 ;
    wire new_AGEMA_signal_10613 ;
    wire new_AGEMA_signal_10614 ;
    wire new_AGEMA_signal_10615 ;
    wire new_AGEMA_signal_10616 ;
    wire new_AGEMA_signal_10617 ;
    wire new_AGEMA_signal_10618 ;
    wire new_AGEMA_signal_10619 ;
    wire new_AGEMA_signal_10620 ;
    wire new_AGEMA_signal_10621 ;
    wire new_AGEMA_signal_10622 ;
    wire new_AGEMA_signal_10623 ;
    wire new_AGEMA_signal_10624 ;
    wire new_AGEMA_signal_10625 ;
    wire new_AGEMA_signal_10626 ;
    wire new_AGEMA_signal_10627 ;
    wire new_AGEMA_signal_10628 ;
    wire new_AGEMA_signal_10629 ;
    wire new_AGEMA_signal_10630 ;
    wire new_AGEMA_signal_10631 ;
    wire new_AGEMA_signal_10632 ;
    wire new_AGEMA_signal_10633 ;
    wire new_AGEMA_signal_10634 ;
    wire new_AGEMA_signal_10635 ;
    wire new_AGEMA_signal_10636 ;
    wire new_AGEMA_signal_10637 ;
    wire new_AGEMA_signal_10638 ;
    wire new_AGEMA_signal_10639 ;
    wire new_AGEMA_signal_10640 ;
    wire new_AGEMA_signal_10641 ;
    wire new_AGEMA_signal_10642 ;
    wire new_AGEMA_signal_10643 ;
    wire new_AGEMA_signal_10644 ;
    wire new_AGEMA_signal_10645 ;
    wire new_AGEMA_signal_10646 ;
    wire new_AGEMA_signal_10647 ;
    wire new_AGEMA_signal_10648 ;
    wire new_AGEMA_signal_10649 ;
    wire new_AGEMA_signal_10650 ;
    wire new_AGEMA_signal_10651 ;
    wire new_AGEMA_signal_10652 ;
    wire new_AGEMA_signal_10653 ;
    wire new_AGEMA_signal_10654 ;
    wire new_AGEMA_signal_10655 ;
    wire new_AGEMA_signal_10656 ;
    wire new_AGEMA_signal_10657 ;
    wire new_AGEMA_signal_10658 ;
    wire new_AGEMA_signal_10659 ;
    wire new_AGEMA_signal_10660 ;
    wire new_AGEMA_signal_10661 ;
    wire new_AGEMA_signal_10662 ;
    wire new_AGEMA_signal_10663 ;
    wire new_AGEMA_signal_10664 ;
    wire new_AGEMA_signal_10665 ;
    wire new_AGEMA_signal_10666 ;
    wire new_AGEMA_signal_10667 ;
    wire new_AGEMA_signal_10668 ;
    wire new_AGEMA_signal_10669 ;
    wire new_AGEMA_signal_10670 ;
    wire new_AGEMA_signal_10671 ;
    wire new_AGEMA_signal_10672 ;
    wire new_AGEMA_signal_10673 ;
    wire new_AGEMA_signal_10674 ;
    wire new_AGEMA_signal_10675 ;
    wire new_AGEMA_signal_10676 ;
    wire new_AGEMA_signal_10677 ;
    wire new_AGEMA_signal_10678 ;
    wire new_AGEMA_signal_10679 ;
    wire new_AGEMA_signal_10680 ;
    wire new_AGEMA_signal_10681 ;
    wire new_AGEMA_signal_10682 ;
    wire new_AGEMA_signal_10683 ;
    wire new_AGEMA_signal_10684 ;
    wire new_AGEMA_signal_10685 ;
    wire new_AGEMA_signal_10686 ;
    wire new_AGEMA_signal_10687 ;
    wire new_AGEMA_signal_10688 ;
    wire new_AGEMA_signal_10689 ;
    wire new_AGEMA_signal_10690 ;
    wire new_AGEMA_signal_10691 ;
    wire new_AGEMA_signal_10692 ;
    wire new_AGEMA_signal_10693 ;
    wire new_AGEMA_signal_10694 ;
    wire new_AGEMA_signal_10695 ;
    wire new_AGEMA_signal_10696 ;
    wire new_AGEMA_signal_10697 ;
    wire new_AGEMA_signal_10698 ;
    wire new_AGEMA_signal_10699 ;
    wire new_AGEMA_signal_10700 ;
    wire new_AGEMA_signal_10701 ;
    wire new_AGEMA_signal_10702 ;
    wire new_AGEMA_signal_10703 ;
    wire new_AGEMA_signal_10704 ;
    wire new_AGEMA_signal_10705 ;
    wire new_AGEMA_signal_10706 ;
    wire new_AGEMA_signal_10707 ;
    wire new_AGEMA_signal_10708 ;
    wire new_AGEMA_signal_10709 ;
    wire new_AGEMA_signal_10710 ;
    wire new_AGEMA_signal_10711 ;
    wire new_AGEMA_signal_10712 ;
    wire new_AGEMA_signal_10713 ;
    wire new_AGEMA_signal_10714 ;
    wire new_AGEMA_signal_10715 ;
    wire new_AGEMA_signal_10716 ;
    wire new_AGEMA_signal_10717 ;
    wire new_AGEMA_signal_10718 ;
    wire new_AGEMA_signal_10719 ;
    wire new_AGEMA_signal_10720 ;
    wire new_AGEMA_signal_10721 ;
    wire new_AGEMA_signal_10722 ;
    wire new_AGEMA_signal_10723 ;
    wire new_AGEMA_signal_10724 ;
    wire new_AGEMA_signal_10725 ;
    wire new_AGEMA_signal_10726 ;
    wire new_AGEMA_signal_10727 ;
    wire new_AGEMA_signal_10728 ;
    wire new_AGEMA_signal_10729 ;
    wire new_AGEMA_signal_10730 ;
    wire new_AGEMA_signal_10731 ;
    wire new_AGEMA_signal_10732 ;
    wire new_AGEMA_signal_10733 ;
    wire new_AGEMA_signal_10734 ;
    wire new_AGEMA_signal_10735 ;
    wire new_AGEMA_signal_10736 ;
    wire new_AGEMA_signal_10737 ;
    wire new_AGEMA_signal_10738 ;
    wire new_AGEMA_signal_10739 ;
    wire new_AGEMA_signal_10740 ;
    wire new_AGEMA_signal_10741 ;
    wire new_AGEMA_signal_10742 ;
    wire new_AGEMA_signal_10743 ;
    wire new_AGEMA_signal_10744 ;
    wire new_AGEMA_signal_10745 ;
    wire new_AGEMA_signal_10746 ;
    wire new_AGEMA_signal_10747 ;
    wire new_AGEMA_signal_10748 ;
    wire new_AGEMA_signal_10749 ;
    wire new_AGEMA_signal_10750 ;
    wire new_AGEMA_signal_10751 ;
    wire new_AGEMA_signal_10752 ;
    wire new_AGEMA_signal_10753 ;
    wire new_AGEMA_signal_10754 ;
    wire new_AGEMA_signal_10755 ;
    wire new_AGEMA_signal_10756 ;
    wire new_AGEMA_signal_10757 ;
    wire new_AGEMA_signal_10758 ;
    wire new_AGEMA_signal_10759 ;
    wire new_AGEMA_signal_10760 ;
    wire new_AGEMA_signal_10761 ;
    wire new_AGEMA_signal_10762 ;
    wire new_AGEMA_signal_10763 ;
    wire new_AGEMA_signal_10764 ;
    wire new_AGEMA_signal_10765 ;
    wire new_AGEMA_signal_10766 ;
    wire new_AGEMA_signal_10767 ;
    wire new_AGEMA_signal_10768 ;
    wire new_AGEMA_signal_10769 ;
    wire new_AGEMA_signal_10770 ;
    wire new_AGEMA_signal_10771 ;
    wire new_AGEMA_signal_10772 ;
    wire new_AGEMA_signal_10773 ;
    wire new_AGEMA_signal_10774 ;
    wire new_AGEMA_signal_10775 ;
    wire new_AGEMA_signal_10776 ;
    wire new_AGEMA_signal_10779 ;
    wire new_AGEMA_signal_10780 ;
    wire new_AGEMA_signal_10783 ;
    wire new_AGEMA_signal_10784 ;
    wire new_AGEMA_signal_10787 ;
    wire new_AGEMA_signal_10788 ;
    wire new_AGEMA_signal_10791 ;
    wire new_AGEMA_signal_10792 ;
    wire new_AGEMA_signal_10795 ;
    wire new_AGEMA_signal_10796 ;
    wire new_AGEMA_signal_10799 ;
    wire new_AGEMA_signal_10800 ;
    wire new_AGEMA_signal_10803 ;
    wire new_AGEMA_signal_10804 ;
    wire new_AGEMA_signal_10807 ;
    wire new_AGEMA_signal_10808 ;
    wire new_AGEMA_signal_10811 ;
    wire new_AGEMA_signal_10812 ;
    wire new_AGEMA_signal_10815 ;
    wire new_AGEMA_signal_10816 ;
    wire new_AGEMA_signal_10819 ;
    wire new_AGEMA_signal_10820 ;
    wire new_AGEMA_signal_10823 ;
    wire new_AGEMA_signal_10824 ;
    wire new_AGEMA_signal_10827 ;
    wire new_AGEMA_signal_10828 ;
    wire new_AGEMA_signal_10831 ;
    wire new_AGEMA_signal_10832 ;
    wire new_AGEMA_signal_10835 ;
    wire new_AGEMA_signal_10836 ;
    wire new_AGEMA_signal_10839 ;
    wire new_AGEMA_signal_10840 ;
    wire new_AGEMA_signal_10843 ;
    wire new_AGEMA_signal_10844 ;
    wire new_AGEMA_signal_10847 ;
    wire new_AGEMA_signal_10848 ;
    wire new_AGEMA_signal_10851 ;
    wire new_AGEMA_signal_10852 ;
    wire new_AGEMA_signal_10855 ;
    wire new_AGEMA_signal_10856 ;
    wire new_AGEMA_signal_10859 ;
    wire new_AGEMA_signal_10860 ;
    wire new_AGEMA_signal_10863 ;
    wire new_AGEMA_signal_10864 ;
    wire new_AGEMA_signal_10867 ;
    wire new_AGEMA_signal_10868 ;
    wire new_AGEMA_signal_10871 ;
    wire new_AGEMA_signal_10872 ;
    wire new_AGEMA_signal_10875 ;
    wire new_AGEMA_signal_10876 ;
    wire new_AGEMA_signal_10877 ;
    wire new_AGEMA_signal_10878 ;
    wire new_AGEMA_signal_10879 ;
    wire new_AGEMA_signal_10880 ;
    wire new_AGEMA_signal_10881 ;
    wire new_AGEMA_signal_10882 ;
    wire new_AGEMA_signal_10883 ;
    wire new_AGEMA_signal_10884 ;
    wire new_AGEMA_signal_10885 ;
    wire new_AGEMA_signal_10886 ;
    wire new_AGEMA_signal_10887 ;
    wire new_AGEMA_signal_10888 ;
    wire new_AGEMA_signal_10889 ;
    wire new_AGEMA_signal_10890 ;
    wire new_AGEMA_signal_10891 ;
    wire new_AGEMA_signal_10892 ;
    wire new_AGEMA_signal_10893 ;
    wire new_AGEMA_signal_10894 ;
    wire new_AGEMA_signal_10895 ;
    wire new_AGEMA_signal_10896 ;
    wire new_AGEMA_signal_10897 ;
    wire new_AGEMA_signal_10898 ;
    wire new_AGEMA_signal_10899 ;
    wire new_AGEMA_signal_10900 ;
    wire new_AGEMA_signal_10901 ;
    wire new_AGEMA_signal_10902 ;
    wire new_AGEMA_signal_10903 ;
    wire new_AGEMA_signal_10904 ;
    wire new_AGEMA_signal_10905 ;
    wire new_AGEMA_signal_10906 ;
    wire new_AGEMA_signal_10907 ;
    wire new_AGEMA_signal_10908 ;
    wire new_AGEMA_signal_10909 ;
    wire new_AGEMA_signal_10910 ;
    wire new_AGEMA_signal_10911 ;
    wire new_AGEMA_signal_10912 ;
    wire new_AGEMA_signal_10913 ;
    wire new_AGEMA_signal_10914 ;
    wire new_AGEMA_signal_10915 ;
    wire new_AGEMA_signal_10916 ;
    wire new_AGEMA_signal_10917 ;
    wire new_AGEMA_signal_10918 ;
    wire new_AGEMA_signal_10919 ;
    wire new_AGEMA_signal_10920 ;
    wire new_AGEMA_signal_10921 ;
    wire new_AGEMA_signal_10922 ;
    wire new_AGEMA_signal_10923 ;
    wire new_AGEMA_signal_10924 ;
    wire new_AGEMA_signal_10925 ;
    wire new_AGEMA_signal_10926 ;
    wire new_AGEMA_signal_10927 ;
    wire new_AGEMA_signal_10928 ;
    wire new_AGEMA_signal_10929 ;
    wire new_AGEMA_signal_10930 ;
    wire new_AGEMA_signal_10931 ;
    wire new_AGEMA_signal_10932 ;
    wire new_AGEMA_signal_10933 ;
    wire new_AGEMA_signal_10934 ;
    wire new_AGEMA_signal_10935 ;
    wire new_AGEMA_signal_10936 ;
    wire new_AGEMA_signal_10937 ;
    wire new_AGEMA_signal_10938 ;
    wire new_AGEMA_signal_10939 ;
    wire new_AGEMA_signal_10940 ;
    wire new_AGEMA_signal_10941 ;
    wire new_AGEMA_signal_10942 ;
    wire new_AGEMA_signal_10943 ;
    wire new_AGEMA_signal_10944 ;
    wire new_AGEMA_signal_10945 ;
    wire new_AGEMA_signal_10946 ;
    wire new_AGEMA_signal_10947 ;
    wire new_AGEMA_signal_10948 ;
    wire new_AGEMA_signal_10949 ;
    wire new_AGEMA_signal_10950 ;
    wire new_AGEMA_signal_10951 ;
    wire new_AGEMA_signal_10952 ;
    wire new_AGEMA_signal_10953 ;
    wire new_AGEMA_signal_10954 ;
    wire new_AGEMA_signal_10955 ;
    wire new_AGEMA_signal_10956 ;
    wire new_AGEMA_signal_10957 ;
    wire new_AGEMA_signal_10958 ;
    wire new_AGEMA_signal_10959 ;
    wire new_AGEMA_signal_10960 ;
    wire new_AGEMA_signal_10961 ;
    wire new_AGEMA_signal_10962 ;
    wire new_AGEMA_signal_10963 ;
    wire new_AGEMA_signal_10964 ;
    wire new_AGEMA_signal_10965 ;
    wire new_AGEMA_signal_10966 ;
    wire new_AGEMA_signal_10967 ;
    wire new_AGEMA_signal_10968 ;
    wire new_AGEMA_signal_10969 ;
    wire new_AGEMA_signal_10970 ;
    wire new_AGEMA_signal_10971 ;
    wire new_AGEMA_signal_10972 ;
    wire new_AGEMA_signal_10973 ;
    wire new_AGEMA_signal_10974 ;
    wire new_AGEMA_signal_10975 ;
    wire new_AGEMA_signal_10976 ;
    wire new_AGEMA_signal_10977 ;
    wire new_AGEMA_signal_10978 ;
    wire new_AGEMA_signal_10979 ;
    wire new_AGEMA_signal_10980 ;
    wire new_AGEMA_signal_10981 ;
    wire new_AGEMA_signal_10982 ;
    wire new_AGEMA_signal_10983 ;
    wire new_AGEMA_signal_10984 ;
    wire new_AGEMA_signal_10985 ;
    wire new_AGEMA_signal_10986 ;
    wire new_AGEMA_signal_10987 ;
    wire new_AGEMA_signal_10988 ;
    wire new_AGEMA_signal_10989 ;
    wire new_AGEMA_signal_10990 ;
    wire new_AGEMA_signal_10991 ;
    wire new_AGEMA_signal_10992 ;
    wire new_AGEMA_signal_10993 ;
    wire new_AGEMA_signal_10994 ;
    wire new_AGEMA_signal_10995 ;
    wire new_AGEMA_signal_10996 ;
    wire new_AGEMA_signal_10997 ;
    wire new_AGEMA_signal_10998 ;
    wire new_AGEMA_signal_10999 ;
    wire new_AGEMA_signal_11000 ;
    wire new_AGEMA_signal_11001 ;
    wire new_AGEMA_signal_11002 ;
    wire new_AGEMA_signal_11003 ;
    wire new_AGEMA_signal_11004 ;
    wire new_AGEMA_signal_11005 ;
    wire new_AGEMA_signal_11006 ;
    wire new_AGEMA_signal_11007 ;
    wire new_AGEMA_signal_11008 ;
    wire new_AGEMA_signal_11009 ;
    wire new_AGEMA_signal_11010 ;
    wire new_AGEMA_signal_11011 ;
    wire new_AGEMA_signal_11012 ;
    wire new_AGEMA_signal_11013 ;
    wire new_AGEMA_signal_11014 ;
    wire new_AGEMA_signal_11015 ;
    wire new_AGEMA_signal_11016 ;
    wire new_AGEMA_signal_11017 ;
    wire new_AGEMA_signal_11018 ;
    wire new_AGEMA_signal_11019 ;
    wire new_AGEMA_signal_11020 ;
    wire new_AGEMA_signal_11021 ;
    wire new_AGEMA_signal_11022 ;
    wire new_AGEMA_signal_11023 ;
    wire new_AGEMA_signal_11024 ;
    wire new_AGEMA_signal_11025 ;
    wire new_AGEMA_signal_11026 ;
    wire new_AGEMA_signal_11027 ;
    wire new_AGEMA_signal_11028 ;
    wire new_AGEMA_signal_11029 ;
    wire new_AGEMA_signal_11030 ;
    wire new_AGEMA_signal_11031 ;
    wire new_AGEMA_signal_11032 ;
    wire new_AGEMA_signal_11033 ;
    wire new_AGEMA_signal_11034 ;
    wire new_AGEMA_signal_11035 ;
    wire new_AGEMA_signal_11036 ;
    wire new_AGEMA_signal_11037 ;
    wire new_AGEMA_signal_11038 ;
    wire new_AGEMA_signal_11039 ;
    wire new_AGEMA_signal_11040 ;
    wire new_AGEMA_signal_11041 ;
    wire new_AGEMA_signal_11042 ;
    wire new_AGEMA_signal_11043 ;
    wire new_AGEMA_signal_11044 ;
    wire new_AGEMA_signal_11045 ;
    wire new_AGEMA_signal_11046 ;
    wire new_AGEMA_signal_11047 ;
    wire new_AGEMA_signal_11048 ;
    wire new_AGEMA_signal_11049 ;
    wire new_AGEMA_signal_11050 ;
    wire new_AGEMA_signal_11051 ;
    wire new_AGEMA_signal_11052 ;
    wire new_AGEMA_signal_11053 ;
    wire new_AGEMA_signal_11054 ;
    wire new_AGEMA_signal_11055 ;
    wire new_AGEMA_signal_11056 ;
    wire new_AGEMA_signal_11057 ;
    wire new_AGEMA_signal_11058 ;
    wire new_AGEMA_signal_11059 ;
    wire new_AGEMA_signal_11060 ;
    wire new_AGEMA_signal_11061 ;
    wire new_AGEMA_signal_11062 ;
    wire new_AGEMA_signal_11063 ;
    wire new_AGEMA_signal_11064 ;
    wire new_AGEMA_signal_11065 ;
    wire new_AGEMA_signal_11066 ;
    wire new_AGEMA_signal_11067 ;
    wire new_AGEMA_signal_11068 ;
    wire new_AGEMA_signal_11069 ;
    wire new_AGEMA_signal_11070 ;
    wire new_AGEMA_signal_11071 ;
    wire new_AGEMA_signal_11072 ;
    wire new_AGEMA_signal_11073 ;
    wire new_AGEMA_signal_11074 ;
    wire new_AGEMA_signal_11075 ;
    wire new_AGEMA_signal_11076 ;
    wire new_AGEMA_signal_11077 ;
    wire new_AGEMA_signal_11078 ;
    wire new_AGEMA_signal_11079 ;
    wire new_AGEMA_signal_11080 ;
    wire new_AGEMA_signal_11081 ;
    wire new_AGEMA_signal_11082 ;
    wire new_AGEMA_signal_11083 ;
    wire new_AGEMA_signal_11084 ;
    wire new_AGEMA_signal_11085 ;
    wire new_AGEMA_signal_11086 ;
    wire new_AGEMA_signal_11087 ;
    wire new_AGEMA_signal_11088 ;
    wire new_AGEMA_signal_11089 ;
    wire new_AGEMA_signal_11090 ;
    wire new_AGEMA_signal_11091 ;
    wire new_AGEMA_signal_11092 ;
    wire new_AGEMA_signal_11093 ;
    wire new_AGEMA_signal_11094 ;
    wire new_AGEMA_signal_11095 ;
    wire new_AGEMA_signal_11096 ;
    wire new_AGEMA_signal_11097 ;
    wire new_AGEMA_signal_11098 ;
    wire new_AGEMA_signal_11099 ;
    wire new_AGEMA_signal_11100 ;
    wire new_AGEMA_signal_11101 ;
    wire new_AGEMA_signal_11102 ;
    wire new_AGEMA_signal_11103 ;
    wire new_AGEMA_signal_11104 ;
    wire new_AGEMA_signal_11105 ;
    wire new_AGEMA_signal_11106 ;
    wire new_AGEMA_signal_11107 ;
    wire new_AGEMA_signal_11108 ;
    wire new_AGEMA_signal_11109 ;
    wire new_AGEMA_signal_11110 ;
    wire new_AGEMA_signal_11111 ;
    wire new_AGEMA_signal_11112 ;
    wire new_AGEMA_signal_11113 ;
    wire new_AGEMA_signal_11114 ;
    wire new_AGEMA_signal_11115 ;
    wire new_AGEMA_signal_11116 ;
    wire new_AGEMA_signal_11117 ;
    wire new_AGEMA_signal_11118 ;
    wire new_AGEMA_signal_11119 ;
    wire new_AGEMA_signal_11120 ;
    wire new_AGEMA_signal_11121 ;
    wire new_AGEMA_signal_11122 ;
    wire new_AGEMA_signal_11123 ;
    wire new_AGEMA_signal_11124 ;
    wire new_AGEMA_signal_11125 ;
    wire new_AGEMA_signal_11126 ;
    wire new_AGEMA_signal_11127 ;
    wire new_AGEMA_signal_11128 ;
    wire new_AGEMA_signal_11129 ;
    wire new_AGEMA_signal_11130 ;
    wire new_AGEMA_signal_11131 ;
    wire new_AGEMA_signal_11132 ;
    wire new_AGEMA_signal_11133 ;
    wire new_AGEMA_signal_11134 ;
    wire new_AGEMA_signal_11135 ;
    wire new_AGEMA_signal_11136 ;
    wire new_AGEMA_signal_11137 ;
    wire new_AGEMA_signal_11138 ;
    wire new_AGEMA_signal_11139 ;
    wire new_AGEMA_signal_11140 ;
    wire new_AGEMA_signal_11141 ;
    wire new_AGEMA_signal_11142 ;
    wire new_AGEMA_signal_11143 ;
    wire new_AGEMA_signal_11144 ;
    wire new_AGEMA_signal_11145 ;
    wire new_AGEMA_signal_11146 ;
    wire new_AGEMA_signal_11147 ;
    wire new_AGEMA_signal_11148 ;
    wire new_AGEMA_signal_11149 ;
    wire new_AGEMA_signal_11150 ;
    wire new_AGEMA_signal_11151 ;
    wire new_AGEMA_signal_11152 ;
    wire new_AGEMA_signal_11153 ;
    wire new_AGEMA_signal_11154 ;
    wire new_AGEMA_signal_11155 ;
    wire new_AGEMA_signal_11156 ;
    wire new_AGEMA_signal_11157 ;
    wire new_AGEMA_signal_11158 ;
    wire new_AGEMA_signal_11159 ;
    wire new_AGEMA_signal_11160 ;
    wire new_AGEMA_signal_11161 ;
    wire new_AGEMA_signal_11162 ;
    wire new_AGEMA_signal_11163 ;
    wire new_AGEMA_signal_11164 ;
    wire new_AGEMA_signal_11165 ;
    wire new_AGEMA_signal_11166 ;
    wire new_AGEMA_signal_11167 ;
    wire new_AGEMA_signal_11168 ;
    wire new_AGEMA_signal_11169 ;
    wire new_AGEMA_signal_11170 ;
    wire new_AGEMA_signal_11171 ;
    wire new_AGEMA_signal_11172 ;
    wire new_AGEMA_signal_11173 ;
    wire new_AGEMA_signal_11174 ;
    wire new_AGEMA_signal_11175 ;
    wire new_AGEMA_signal_11176 ;
    wire new_AGEMA_signal_11177 ;
    wire new_AGEMA_signal_11178 ;
    wire new_AGEMA_signal_11179 ;
    wire new_AGEMA_signal_11180 ;
    wire new_AGEMA_signal_11181 ;
    wire new_AGEMA_signal_11182 ;
    wire new_AGEMA_signal_11183 ;
    wire new_AGEMA_signal_11184 ;
    wire new_AGEMA_signal_11185 ;
    wire new_AGEMA_signal_11186 ;
    wire new_AGEMA_signal_11187 ;
    wire new_AGEMA_signal_11188 ;
    wire new_AGEMA_signal_11189 ;
    wire new_AGEMA_signal_11190 ;
    wire new_AGEMA_signal_11191 ;
    wire new_AGEMA_signal_11192 ;
    wire new_AGEMA_signal_11193 ;
    wire new_AGEMA_signal_11194 ;
    wire new_AGEMA_signal_11195 ;
    wire new_AGEMA_signal_11196 ;
    wire new_AGEMA_signal_11199 ;
    wire new_AGEMA_signal_11200 ;
    wire new_AGEMA_signal_11203 ;
    wire new_AGEMA_signal_11204 ;
    wire new_AGEMA_signal_11207 ;
    wire new_AGEMA_signal_11208 ;
    wire new_AGEMA_signal_11211 ;
    wire new_AGEMA_signal_11212 ;
    wire new_AGEMA_signal_11215 ;
    wire new_AGEMA_signal_11216 ;
    wire new_AGEMA_signal_11219 ;
    wire new_AGEMA_signal_11220 ;
    wire new_AGEMA_signal_11223 ;
    wire new_AGEMA_signal_11224 ;
    wire new_AGEMA_signal_11227 ;
    wire new_AGEMA_signal_11228 ;
    wire new_AGEMA_signal_11231 ;
    wire new_AGEMA_signal_11232 ;
    wire new_AGEMA_signal_11235 ;
    wire new_AGEMA_signal_11236 ;
    wire new_AGEMA_signal_11239 ;
    wire new_AGEMA_signal_11240 ;
    wire new_AGEMA_signal_11243 ;
    wire new_AGEMA_signal_11244 ;
    wire new_AGEMA_signal_11247 ;
    wire new_AGEMA_signal_11248 ;
    wire new_AGEMA_signal_11251 ;
    wire new_AGEMA_signal_11252 ;
    wire new_AGEMA_signal_11255 ;
    wire new_AGEMA_signal_11256 ;
    wire new_AGEMA_signal_11259 ;
    wire new_AGEMA_signal_11260 ;
    wire new_AGEMA_signal_11263 ;
    wire new_AGEMA_signal_11264 ;
    wire new_AGEMA_signal_11267 ;
    wire new_AGEMA_signal_11268 ;
    wire new_AGEMA_signal_11271 ;
    wire new_AGEMA_signal_11272 ;
    wire new_AGEMA_signal_11275 ;
    wire new_AGEMA_signal_11276 ;
    wire new_AGEMA_signal_11279 ;
    wire new_AGEMA_signal_11280 ;
    wire new_AGEMA_signal_11283 ;
    wire new_AGEMA_signal_11284 ;
    wire new_AGEMA_signal_11287 ;
    wire new_AGEMA_signal_11288 ;
    wire new_AGEMA_signal_11291 ;
    wire new_AGEMA_signal_11292 ;
    wire new_AGEMA_signal_11295 ;
    wire new_AGEMA_signal_11296 ;
    wire new_AGEMA_signal_11299 ;
    wire new_AGEMA_signal_11300 ;
    wire new_AGEMA_signal_11303 ;
    wire new_AGEMA_signal_11304 ;
    wire new_AGEMA_signal_11307 ;
    wire new_AGEMA_signal_11308 ;
    wire new_AGEMA_signal_11311 ;
    wire new_AGEMA_signal_11312 ;
    wire new_AGEMA_signal_11315 ;
    wire new_AGEMA_signal_11316 ;
    wire new_AGEMA_signal_11319 ;
    wire new_AGEMA_signal_11320 ;
    wire new_AGEMA_signal_11323 ;
    wire new_AGEMA_signal_11324 ;
    wire new_AGEMA_signal_11325 ;
    wire new_AGEMA_signal_11326 ;
    wire new_AGEMA_signal_11327 ;
    wire new_AGEMA_signal_11328 ;
    wire new_AGEMA_signal_11329 ;
    wire new_AGEMA_signal_11330 ;
    wire new_AGEMA_signal_11331 ;
    wire new_AGEMA_signal_11332 ;
    wire new_AGEMA_signal_11333 ;
    wire new_AGEMA_signal_11334 ;
    wire new_AGEMA_signal_11335 ;
    wire new_AGEMA_signal_11336 ;
    wire new_AGEMA_signal_11337 ;
    wire new_AGEMA_signal_11338 ;
    wire new_AGEMA_signal_11339 ;
    wire new_AGEMA_signal_11340 ;
    wire new_AGEMA_signal_11341 ;
    wire new_AGEMA_signal_11342 ;
    wire new_AGEMA_signal_11343 ;
    wire new_AGEMA_signal_11344 ;
    wire new_AGEMA_signal_11345 ;
    wire new_AGEMA_signal_11346 ;
    wire new_AGEMA_signal_11347 ;
    wire new_AGEMA_signal_11348 ;
    wire new_AGEMA_signal_11349 ;
    wire new_AGEMA_signal_11350 ;
    wire new_AGEMA_signal_11351 ;
    wire new_AGEMA_signal_11352 ;
    wire new_AGEMA_signal_11353 ;
    wire new_AGEMA_signal_11354 ;
    wire new_AGEMA_signal_11355 ;
    wire new_AGEMA_signal_11356 ;
    wire new_AGEMA_signal_11357 ;
    wire new_AGEMA_signal_11358 ;
    wire new_AGEMA_signal_11359 ;
    wire new_AGEMA_signal_11360 ;
    wire new_AGEMA_signal_11361 ;
    wire new_AGEMA_signal_11362 ;
    wire new_AGEMA_signal_11363 ;
    wire new_AGEMA_signal_11364 ;
    wire new_AGEMA_signal_11365 ;
    wire new_AGEMA_signal_11366 ;
    wire new_AGEMA_signal_11367 ;
    wire new_AGEMA_signal_11368 ;
    wire new_AGEMA_signal_11369 ;
    wire new_AGEMA_signal_11370 ;
    wire new_AGEMA_signal_11371 ;
    wire new_AGEMA_signal_11372 ;
    wire new_AGEMA_signal_11373 ;
    wire new_AGEMA_signal_11374 ;
    wire new_AGEMA_signal_11375 ;
    wire new_AGEMA_signal_11376 ;
    wire new_AGEMA_signal_11377 ;
    wire new_AGEMA_signal_11378 ;
    wire new_AGEMA_signal_11379 ;
    wire new_AGEMA_signal_11380 ;
    wire new_AGEMA_signal_11381 ;
    wire new_AGEMA_signal_11382 ;
    wire new_AGEMA_signal_11383 ;
    wire new_AGEMA_signal_11384 ;
    wire new_AGEMA_signal_11385 ;
    wire new_AGEMA_signal_11386 ;
    wire new_AGEMA_signal_11387 ;
    wire new_AGEMA_signal_11388 ;
    wire new_AGEMA_signal_11389 ;
    wire new_AGEMA_signal_11390 ;
    wire new_AGEMA_signal_11391 ;
    wire new_AGEMA_signal_11392 ;
    wire new_AGEMA_signal_11393 ;
    wire new_AGEMA_signal_11394 ;
    wire new_AGEMA_signal_11395 ;
    wire new_AGEMA_signal_11396 ;
    wire new_AGEMA_signal_11397 ;
    wire new_AGEMA_signal_11398 ;
    wire new_AGEMA_signal_11399 ;
    wire new_AGEMA_signal_11400 ;
    wire new_AGEMA_signal_11401 ;
    wire new_AGEMA_signal_11402 ;
    wire new_AGEMA_signal_11403 ;
    wire new_AGEMA_signal_11404 ;
    wire new_AGEMA_signal_11405 ;
    wire new_AGEMA_signal_11406 ;
    wire new_AGEMA_signal_11407 ;
    wire new_AGEMA_signal_11408 ;
    wire new_AGEMA_signal_11409 ;
    wire new_AGEMA_signal_11410 ;
    wire new_AGEMA_signal_11411 ;
    wire new_AGEMA_signal_11412 ;
    wire new_AGEMA_signal_11413 ;
    wire new_AGEMA_signal_11414 ;
    wire new_AGEMA_signal_11415 ;
    wire new_AGEMA_signal_11416 ;
    wire new_AGEMA_signal_11417 ;
    wire new_AGEMA_signal_11418 ;
    wire new_AGEMA_signal_11419 ;
    wire new_AGEMA_signal_11420 ;
    wire new_AGEMA_signal_11421 ;
    wire new_AGEMA_signal_11422 ;
    wire new_AGEMA_signal_11423 ;
    wire new_AGEMA_signal_11424 ;
    wire new_AGEMA_signal_11425 ;
    wire new_AGEMA_signal_11426 ;
    wire new_AGEMA_signal_11427 ;
    wire new_AGEMA_signal_11428 ;
    wire new_AGEMA_signal_11429 ;
    wire new_AGEMA_signal_11430 ;
    wire new_AGEMA_signal_11431 ;
    wire new_AGEMA_signal_11432 ;
    wire new_AGEMA_signal_11433 ;
    wire new_AGEMA_signal_11434 ;
    wire new_AGEMA_signal_11435 ;
    wire new_AGEMA_signal_11436 ;
    wire new_AGEMA_signal_11437 ;
    wire new_AGEMA_signal_11438 ;
    wire new_AGEMA_signal_11439 ;
    wire new_AGEMA_signal_11440 ;
    wire new_AGEMA_signal_11441 ;
    wire new_AGEMA_signal_11442 ;
    wire new_AGEMA_signal_11443 ;
    wire new_AGEMA_signal_11444 ;
    wire new_AGEMA_signal_11445 ;
    wire new_AGEMA_signal_11446 ;
    wire new_AGEMA_signal_11447 ;
    wire new_AGEMA_signal_11448 ;
    wire new_AGEMA_signal_11449 ;
    wire new_AGEMA_signal_11450 ;
    wire new_AGEMA_signal_11451 ;
    wire new_AGEMA_signal_11452 ;
    wire new_AGEMA_signal_11453 ;
    wire new_AGEMA_signal_11454 ;
    wire new_AGEMA_signal_11455 ;
    wire new_AGEMA_signal_11456 ;
    wire new_AGEMA_signal_11457 ;
    wire new_AGEMA_signal_11458 ;
    wire new_AGEMA_signal_11459 ;
    wire new_AGEMA_signal_11460 ;
    wire new_AGEMA_signal_11461 ;
    wire new_AGEMA_signal_11462 ;
    wire new_AGEMA_signal_11463 ;
    wire new_AGEMA_signal_11464 ;
    wire new_AGEMA_signal_11465 ;
    wire new_AGEMA_signal_11466 ;
    wire new_AGEMA_signal_11467 ;
    wire new_AGEMA_signal_11468 ;
    wire new_AGEMA_signal_11469 ;
    wire new_AGEMA_signal_11470 ;
    wire new_AGEMA_signal_11471 ;
    wire new_AGEMA_signal_11472 ;
    wire new_AGEMA_signal_11473 ;
    wire new_AGEMA_signal_11474 ;
    wire new_AGEMA_signal_11475 ;
    wire new_AGEMA_signal_11476 ;
    wire new_AGEMA_signal_11477 ;
    wire new_AGEMA_signal_11478 ;
    wire new_AGEMA_signal_11479 ;
    wire new_AGEMA_signal_11480 ;
    wire new_AGEMA_signal_11481 ;
    wire new_AGEMA_signal_11482 ;
    wire new_AGEMA_signal_11483 ;
    wire new_AGEMA_signal_11484 ;
    wire new_AGEMA_signal_11485 ;
    wire new_AGEMA_signal_11486 ;
    wire new_AGEMA_signal_11487 ;
    wire new_AGEMA_signal_11488 ;
    wire new_AGEMA_signal_11489 ;
    wire new_AGEMA_signal_11490 ;
    wire new_AGEMA_signal_11491 ;
    wire new_AGEMA_signal_11492 ;
    wire new_AGEMA_signal_11493 ;
    wire new_AGEMA_signal_11494 ;
    wire new_AGEMA_signal_11495 ;
    wire new_AGEMA_signal_11496 ;
    wire new_AGEMA_signal_11497 ;
    wire new_AGEMA_signal_11498 ;
    wire new_AGEMA_signal_11499 ;
    wire new_AGEMA_signal_11500 ;
    wire new_AGEMA_signal_11501 ;
    wire new_AGEMA_signal_11502 ;
    wire new_AGEMA_signal_11503 ;
    wire new_AGEMA_signal_11504 ;
    wire new_AGEMA_signal_11505 ;
    wire new_AGEMA_signal_11506 ;
    wire new_AGEMA_signal_11507 ;
    wire new_AGEMA_signal_11508 ;
    wire new_AGEMA_signal_11509 ;
    wire new_AGEMA_signal_11510 ;
    wire new_AGEMA_signal_11511 ;
    wire new_AGEMA_signal_11512 ;
    wire new_AGEMA_signal_11513 ;
    wire new_AGEMA_signal_11514 ;
    wire new_AGEMA_signal_11515 ;
    wire new_AGEMA_signal_11516 ;
    wire new_AGEMA_signal_11517 ;
    wire new_AGEMA_signal_11518 ;
    wire new_AGEMA_signal_11519 ;
    wire new_AGEMA_signal_11520 ;
    wire new_AGEMA_signal_11521 ;
    wire new_AGEMA_signal_11522 ;
    wire new_AGEMA_signal_11523 ;
    wire new_AGEMA_signal_11524 ;
    wire new_AGEMA_signal_11525 ;
    wire new_AGEMA_signal_11526 ;
    wire new_AGEMA_signal_11527 ;
    wire new_AGEMA_signal_11528 ;
    wire new_AGEMA_signal_11529 ;
    wire new_AGEMA_signal_11530 ;
    wire new_AGEMA_signal_11531 ;
    wire new_AGEMA_signal_11532 ;
    wire new_AGEMA_signal_11533 ;
    wire new_AGEMA_signal_11534 ;
    wire new_AGEMA_signal_11535 ;
    wire new_AGEMA_signal_11536 ;
    wire new_AGEMA_signal_11537 ;
    wire new_AGEMA_signal_11538 ;
    wire new_AGEMA_signal_11539 ;
    wire new_AGEMA_signal_11540 ;
    wire new_AGEMA_signal_11541 ;
    wire new_AGEMA_signal_11542 ;
    wire new_AGEMA_signal_11543 ;
    wire new_AGEMA_signal_11544 ;
    wire new_AGEMA_signal_11545 ;
    wire new_AGEMA_signal_11546 ;
    wire new_AGEMA_signal_11547 ;
    wire new_AGEMA_signal_11548 ;
    wire new_AGEMA_signal_11549 ;
    wire new_AGEMA_signal_11550 ;
    wire new_AGEMA_signal_11551 ;
    wire new_AGEMA_signal_11552 ;
    wire new_AGEMA_signal_11553 ;
    wire new_AGEMA_signal_11554 ;
    wire new_AGEMA_signal_11555 ;
    wire new_AGEMA_signal_11556 ;
    wire new_AGEMA_signal_11557 ;
    wire new_AGEMA_signal_11558 ;
    wire new_AGEMA_signal_11559 ;
    wire new_AGEMA_signal_11560 ;
    wire new_AGEMA_signal_11561 ;
    wire new_AGEMA_signal_11562 ;
    wire new_AGEMA_signal_11563 ;
    wire new_AGEMA_signal_11564 ;
    wire new_AGEMA_signal_11565 ;
    wire new_AGEMA_signal_11566 ;
    wire new_AGEMA_signal_11567 ;
    wire new_AGEMA_signal_11568 ;
    wire new_AGEMA_signal_11569 ;
    wire new_AGEMA_signal_11570 ;
    wire new_AGEMA_signal_11571 ;
    wire new_AGEMA_signal_11572 ;
    wire new_AGEMA_signal_11573 ;
    wire new_AGEMA_signal_11574 ;
    wire new_AGEMA_signal_11575 ;
    wire new_AGEMA_signal_11576 ;
    wire new_AGEMA_signal_11577 ;
    wire new_AGEMA_signal_11578 ;
    wire new_AGEMA_signal_11579 ;
    wire new_AGEMA_signal_11580 ;
    wire new_AGEMA_signal_11581 ;
    wire new_AGEMA_signal_11582 ;
    wire new_AGEMA_signal_11583 ;
    wire new_AGEMA_signal_11584 ;
    wire new_AGEMA_signal_11585 ;
    wire new_AGEMA_signal_11586 ;
    wire new_AGEMA_signal_11587 ;
    wire new_AGEMA_signal_11588 ;
    wire new_AGEMA_signal_11589 ;
    wire new_AGEMA_signal_11590 ;
    wire new_AGEMA_signal_11591 ;
    wire new_AGEMA_signal_11592 ;
    wire new_AGEMA_signal_11593 ;
    wire new_AGEMA_signal_11594 ;
    wire new_AGEMA_signal_11595 ;
    wire new_AGEMA_signal_11596 ;
    wire new_AGEMA_signal_11597 ;
    wire new_AGEMA_signal_11598 ;
    wire new_AGEMA_signal_11599 ;
    wire new_AGEMA_signal_11600 ;
    wire new_AGEMA_signal_11601 ;
    wire new_AGEMA_signal_11602 ;
    wire new_AGEMA_signal_11603 ;
    wire new_AGEMA_signal_11604 ;
    wire new_AGEMA_signal_11605 ;
    wire new_AGEMA_signal_11606 ;
    wire new_AGEMA_signal_11607 ;
    wire new_AGEMA_signal_11608 ;
    wire new_AGEMA_signal_11609 ;
    wire new_AGEMA_signal_11610 ;
    wire new_AGEMA_signal_11611 ;
    wire new_AGEMA_signal_11612 ;
    wire new_AGEMA_signal_11613 ;
    wire new_AGEMA_signal_11614 ;
    wire new_AGEMA_signal_11615 ;
    wire new_AGEMA_signal_11616 ;
    wire new_AGEMA_signal_11617 ;
    wire new_AGEMA_signal_11618 ;
    wire new_AGEMA_signal_11619 ;
    wire new_AGEMA_signal_11620 ;
    wire new_AGEMA_signal_11621 ;
    wire new_AGEMA_signal_11622 ;
    wire new_AGEMA_signal_11623 ;
    wire new_AGEMA_signal_11624 ;
    wire new_AGEMA_signal_11625 ;
    wire new_AGEMA_signal_11626 ;
    wire new_AGEMA_signal_11627 ;
    wire new_AGEMA_signal_11628 ;
    wire new_AGEMA_signal_11629 ;
    wire new_AGEMA_signal_11630 ;
    wire new_AGEMA_signal_11631 ;
    wire new_AGEMA_signal_11632 ;
    wire new_AGEMA_signal_11633 ;
    wire new_AGEMA_signal_11634 ;
    wire new_AGEMA_signal_11635 ;
    wire new_AGEMA_signal_11636 ;
    wire new_AGEMA_signal_11637 ;
    wire new_AGEMA_signal_11638 ;
    wire new_AGEMA_signal_11639 ;
    wire new_AGEMA_signal_11640 ;
    wire new_AGEMA_signal_11641 ;
    wire new_AGEMA_signal_11642 ;
    wire new_AGEMA_signal_11643 ;
    wire new_AGEMA_signal_11644 ;
    wire new_AGEMA_signal_11647 ;
    wire new_AGEMA_signal_11648 ;
    wire new_AGEMA_signal_11651 ;
    wire new_AGEMA_signal_11652 ;
    wire new_AGEMA_signal_11655 ;
    wire new_AGEMA_signal_11656 ;
    wire new_AGEMA_signal_11659 ;
    wire new_AGEMA_signal_11660 ;
    wire new_AGEMA_signal_11663 ;
    wire new_AGEMA_signal_11664 ;
    wire new_AGEMA_signal_11667 ;
    wire new_AGEMA_signal_11668 ;
    wire new_AGEMA_signal_11671 ;
    wire new_AGEMA_signal_11672 ;
    wire new_AGEMA_signal_11675 ;
    wire new_AGEMA_signal_11676 ;
    wire new_AGEMA_signal_11679 ;
    wire new_AGEMA_signal_11680 ;
    wire new_AGEMA_signal_11683 ;
    wire new_AGEMA_signal_11684 ;
    wire new_AGEMA_signal_11687 ;
    wire new_AGEMA_signal_11688 ;
    wire new_AGEMA_signal_11691 ;
    wire new_AGEMA_signal_11692 ;
    wire new_AGEMA_signal_11695 ;
    wire new_AGEMA_signal_11696 ;
    wire new_AGEMA_signal_11699 ;
    wire new_AGEMA_signal_11700 ;
    wire new_AGEMA_signal_11703 ;
    wire new_AGEMA_signal_11704 ;
    wire new_AGEMA_signal_11707 ;
    wire new_AGEMA_signal_11708 ;
    wire new_AGEMA_signal_11711 ;
    wire new_AGEMA_signal_11712 ;
    wire new_AGEMA_signal_11715 ;
    wire new_AGEMA_signal_11716 ;
    wire new_AGEMA_signal_11719 ;
    wire new_AGEMA_signal_11720 ;
    wire new_AGEMA_signal_11723 ;
    wire new_AGEMA_signal_11724 ;
    wire new_AGEMA_signal_11727 ;
    wire new_AGEMA_signal_11728 ;
    wire new_AGEMA_signal_11731 ;
    wire new_AGEMA_signal_11732 ;
    wire new_AGEMA_signal_11735 ;
    wire new_AGEMA_signal_11736 ;
    wire new_AGEMA_signal_11739 ;
    wire new_AGEMA_signal_11740 ;
    wire new_AGEMA_signal_11743 ;
    wire new_AGEMA_signal_11744 ;
    wire new_AGEMA_signal_11747 ;
    wire new_AGEMA_signal_11748 ;
    wire new_AGEMA_signal_11751 ;
    wire new_AGEMA_signal_11752 ;
    wire new_AGEMA_signal_11755 ;
    wire new_AGEMA_signal_11756 ;
    wire new_AGEMA_signal_11759 ;
    wire new_AGEMA_signal_11760 ;
    wire new_AGEMA_signal_11763 ;
    wire new_AGEMA_signal_11764 ;
    wire new_AGEMA_signal_11767 ;
    wire new_AGEMA_signal_11768 ;
    wire new_AGEMA_signal_11771 ;
    wire new_AGEMA_signal_11772 ;
    wire new_AGEMA_signal_11773 ;
    wire new_AGEMA_signal_11774 ;
    wire new_AGEMA_signal_11775 ;
    wire new_AGEMA_signal_11776 ;
    wire new_AGEMA_signal_11777 ;
    wire new_AGEMA_signal_11778 ;
    wire new_AGEMA_signal_11779 ;
    wire new_AGEMA_signal_11780 ;
    wire new_AGEMA_signal_11781 ;
    wire new_AGEMA_signal_11782 ;
    wire new_AGEMA_signal_11783 ;
    wire new_AGEMA_signal_11784 ;
    wire new_AGEMA_signal_11785 ;
    wire new_AGEMA_signal_11786 ;
    wire new_AGEMA_signal_11787 ;
    wire new_AGEMA_signal_11788 ;
    wire new_AGEMA_signal_11789 ;
    wire new_AGEMA_signal_11790 ;
    wire new_AGEMA_signal_11791 ;
    wire new_AGEMA_signal_11792 ;
    wire new_AGEMA_signal_11793 ;
    wire new_AGEMA_signal_11794 ;
    wire new_AGEMA_signal_11795 ;
    wire new_AGEMA_signal_11796 ;
    wire new_AGEMA_signal_11797 ;
    wire new_AGEMA_signal_11798 ;
    wire new_AGEMA_signal_11799 ;
    wire new_AGEMA_signal_11800 ;
    wire new_AGEMA_signal_11801 ;
    wire new_AGEMA_signal_11802 ;
    wire new_AGEMA_signal_11803 ;
    wire new_AGEMA_signal_11804 ;
    wire new_AGEMA_signal_11805 ;
    wire new_AGEMA_signal_11806 ;
    wire new_AGEMA_signal_11807 ;
    wire new_AGEMA_signal_11808 ;
    wire new_AGEMA_signal_11809 ;
    wire new_AGEMA_signal_11810 ;
    wire new_AGEMA_signal_11811 ;
    wire new_AGEMA_signal_11812 ;
    wire new_AGEMA_signal_11813 ;
    wire new_AGEMA_signal_11814 ;
    wire new_AGEMA_signal_11815 ;
    wire new_AGEMA_signal_11816 ;
    wire new_AGEMA_signal_11817 ;
    wire new_AGEMA_signal_11818 ;
    wire new_AGEMA_signal_11819 ;
    wire new_AGEMA_signal_11820 ;
    wire new_AGEMA_signal_11821 ;
    wire new_AGEMA_signal_11822 ;
    wire new_AGEMA_signal_11823 ;
    wire new_AGEMA_signal_11824 ;
    wire new_AGEMA_signal_11825 ;
    wire new_AGEMA_signal_11826 ;
    wire new_AGEMA_signal_11827 ;
    wire new_AGEMA_signal_11828 ;
    wire new_AGEMA_signal_11829 ;
    wire new_AGEMA_signal_11830 ;
    wire new_AGEMA_signal_11831 ;
    wire new_AGEMA_signal_11832 ;
    wire new_AGEMA_signal_11833 ;
    wire new_AGEMA_signal_11834 ;
    wire new_AGEMA_signal_11835 ;
    wire new_AGEMA_signal_11836 ;
    wire new_AGEMA_signal_11837 ;
    wire new_AGEMA_signal_11838 ;
    wire new_AGEMA_signal_11839 ;
    wire new_AGEMA_signal_11840 ;
    wire new_AGEMA_signal_11841 ;
    wire new_AGEMA_signal_11842 ;
    wire new_AGEMA_signal_11843 ;
    wire new_AGEMA_signal_11844 ;
    wire new_AGEMA_signal_11845 ;
    wire new_AGEMA_signal_11846 ;
    wire new_AGEMA_signal_11847 ;
    wire new_AGEMA_signal_11848 ;
    wire new_AGEMA_signal_11849 ;
    wire new_AGEMA_signal_11850 ;
    wire new_AGEMA_signal_11851 ;
    wire new_AGEMA_signal_11852 ;
    wire new_AGEMA_signal_11853 ;
    wire new_AGEMA_signal_11854 ;
    wire new_AGEMA_signal_11855 ;
    wire new_AGEMA_signal_11856 ;
    wire new_AGEMA_signal_11857 ;
    wire new_AGEMA_signal_11858 ;
    wire new_AGEMA_signal_11859 ;
    wire new_AGEMA_signal_11860 ;
    wire new_AGEMA_signal_11861 ;
    wire new_AGEMA_signal_11862 ;
    wire new_AGEMA_signal_11863 ;
    wire new_AGEMA_signal_11864 ;
    wire new_AGEMA_signal_11865 ;
    wire new_AGEMA_signal_11866 ;
    wire new_AGEMA_signal_11867 ;
    wire new_AGEMA_signal_11868 ;
    wire new_AGEMA_signal_11869 ;
    wire new_AGEMA_signal_11870 ;
    wire new_AGEMA_signal_11871 ;
    wire new_AGEMA_signal_11872 ;
    wire new_AGEMA_signal_11873 ;
    wire new_AGEMA_signal_11874 ;
    wire new_AGEMA_signal_11875 ;
    wire new_AGEMA_signal_11876 ;
    wire new_AGEMA_signal_11877 ;
    wire new_AGEMA_signal_11878 ;
    wire new_AGEMA_signal_11879 ;
    wire new_AGEMA_signal_11880 ;
    wire new_AGEMA_signal_11881 ;
    wire new_AGEMA_signal_11882 ;
    wire new_AGEMA_signal_11883 ;
    wire new_AGEMA_signal_11884 ;
    wire new_AGEMA_signal_11885 ;
    wire new_AGEMA_signal_11886 ;
    wire new_AGEMA_signal_11887 ;
    wire new_AGEMA_signal_11888 ;
    wire new_AGEMA_signal_11889 ;
    wire new_AGEMA_signal_11890 ;
    wire new_AGEMA_signal_11891 ;
    wire new_AGEMA_signal_11892 ;
    wire new_AGEMA_signal_11893 ;
    wire new_AGEMA_signal_11894 ;
    wire new_AGEMA_signal_11895 ;
    wire new_AGEMA_signal_11896 ;
    wire new_AGEMA_signal_11897 ;
    wire new_AGEMA_signal_11898 ;
    wire new_AGEMA_signal_11899 ;
    wire new_AGEMA_signal_11900 ;
    wire new_AGEMA_signal_11901 ;
    wire new_AGEMA_signal_11902 ;
    wire new_AGEMA_signal_11903 ;
    wire new_AGEMA_signal_11904 ;
    wire new_AGEMA_signal_11905 ;
    wire new_AGEMA_signal_11906 ;
    wire new_AGEMA_signal_11907 ;
    wire new_AGEMA_signal_11908 ;
    wire new_AGEMA_signal_11909 ;
    wire new_AGEMA_signal_11910 ;
    wire new_AGEMA_signal_11911 ;
    wire new_AGEMA_signal_11912 ;
    wire new_AGEMA_signal_11913 ;
    wire new_AGEMA_signal_11914 ;
    wire new_AGEMA_signal_11915 ;
    wire new_AGEMA_signal_11916 ;
    wire new_AGEMA_signal_11917 ;
    wire new_AGEMA_signal_11918 ;
    wire new_AGEMA_signal_11919 ;
    wire new_AGEMA_signal_11920 ;
    wire new_AGEMA_signal_11921 ;
    wire new_AGEMA_signal_11922 ;
    wire new_AGEMA_signal_11923 ;
    wire new_AGEMA_signal_11924 ;
    wire new_AGEMA_signal_11925 ;
    wire new_AGEMA_signal_11926 ;
    wire new_AGEMA_signal_11927 ;
    wire new_AGEMA_signal_11928 ;
    wire new_AGEMA_signal_11929 ;
    wire new_AGEMA_signal_11930 ;
    wire new_AGEMA_signal_11931 ;
    wire new_AGEMA_signal_11932 ;
    wire new_AGEMA_signal_11933 ;
    wire new_AGEMA_signal_11934 ;
    wire new_AGEMA_signal_11935 ;
    wire new_AGEMA_signal_11936 ;
    wire new_AGEMA_signal_11937 ;
    wire new_AGEMA_signal_11938 ;
    wire new_AGEMA_signal_11939 ;
    wire new_AGEMA_signal_11940 ;
    wire new_AGEMA_signal_11941 ;
    wire new_AGEMA_signal_11942 ;
    wire new_AGEMA_signal_11943 ;
    wire new_AGEMA_signal_11944 ;
    wire new_AGEMA_signal_11945 ;
    wire new_AGEMA_signal_11946 ;
    wire new_AGEMA_signal_11947 ;
    wire new_AGEMA_signal_11948 ;
    wire new_AGEMA_signal_11949 ;
    wire new_AGEMA_signal_11950 ;
    wire new_AGEMA_signal_11951 ;
    wire new_AGEMA_signal_11952 ;
    wire new_AGEMA_signal_11953 ;
    wire new_AGEMA_signal_11954 ;
    wire new_AGEMA_signal_11955 ;
    wire new_AGEMA_signal_11956 ;
    wire new_AGEMA_signal_11957 ;
    wire new_AGEMA_signal_11958 ;
    wire new_AGEMA_signal_11959 ;
    wire new_AGEMA_signal_11960 ;
    wire new_AGEMA_signal_11961 ;
    wire new_AGEMA_signal_11962 ;
    wire new_AGEMA_signal_11963 ;
    wire new_AGEMA_signal_11964 ;
    wire new_AGEMA_signal_11965 ;
    wire new_AGEMA_signal_11966 ;
    wire new_AGEMA_signal_11967 ;
    wire new_AGEMA_signal_11968 ;
    wire new_AGEMA_signal_11969 ;
    wire new_AGEMA_signal_11970 ;
    wire new_AGEMA_signal_11971 ;
    wire new_AGEMA_signal_11972 ;
    wire new_AGEMA_signal_11973 ;
    wire new_AGEMA_signal_11974 ;
    wire new_AGEMA_signal_11975 ;
    wire new_AGEMA_signal_11976 ;
    wire new_AGEMA_signal_11977 ;
    wire new_AGEMA_signal_11978 ;
    wire new_AGEMA_signal_11979 ;
    wire new_AGEMA_signal_11980 ;
    wire new_AGEMA_signal_11981 ;
    wire new_AGEMA_signal_11982 ;
    wire new_AGEMA_signal_11983 ;
    wire new_AGEMA_signal_11984 ;
    wire new_AGEMA_signal_11985 ;
    wire new_AGEMA_signal_11986 ;
    wire new_AGEMA_signal_11987 ;
    wire new_AGEMA_signal_11988 ;
    wire new_AGEMA_signal_11989 ;
    wire new_AGEMA_signal_11990 ;
    wire new_AGEMA_signal_11991 ;
    wire new_AGEMA_signal_11992 ;
    wire new_AGEMA_signal_11993 ;
    wire new_AGEMA_signal_11994 ;
    wire new_AGEMA_signal_11995 ;
    wire new_AGEMA_signal_11996 ;
    wire new_AGEMA_signal_11997 ;
    wire new_AGEMA_signal_11998 ;
    wire new_AGEMA_signal_11999 ;
    wire new_AGEMA_signal_12000 ;
    wire new_AGEMA_signal_12001 ;
    wire new_AGEMA_signal_12002 ;
    wire new_AGEMA_signal_12003 ;
    wire new_AGEMA_signal_12004 ;
    wire new_AGEMA_signal_12005 ;
    wire new_AGEMA_signal_12006 ;
    wire new_AGEMA_signal_12007 ;
    wire new_AGEMA_signal_12008 ;
    wire new_AGEMA_signal_12009 ;
    wire new_AGEMA_signal_12010 ;
    wire new_AGEMA_signal_12011 ;
    wire new_AGEMA_signal_12012 ;
    wire new_AGEMA_signal_12013 ;
    wire new_AGEMA_signal_12014 ;
    wire new_AGEMA_signal_12015 ;
    wire new_AGEMA_signal_12016 ;
    wire new_AGEMA_signal_12017 ;
    wire new_AGEMA_signal_12018 ;
    wire new_AGEMA_signal_12019 ;
    wire new_AGEMA_signal_12020 ;
    wire new_AGEMA_signal_12021 ;
    wire new_AGEMA_signal_12022 ;
    wire new_AGEMA_signal_12023 ;
    wire new_AGEMA_signal_12024 ;
    wire new_AGEMA_signal_12025 ;
    wire new_AGEMA_signal_12026 ;
    wire new_AGEMA_signal_12027 ;
    wire new_AGEMA_signal_12028 ;
    wire new_AGEMA_signal_12029 ;
    wire new_AGEMA_signal_12030 ;
    wire new_AGEMA_signal_12031 ;
    wire new_AGEMA_signal_12032 ;
    wire new_AGEMA_signal_12033 ;
    wire new_AGEMA_signal_12034 ;
    wire new_AGEMA_signal_12035 ;
    wire new_AGEMA_signal_12036 ;
    wire new_AGEMA_signal_12037 ;
    wire new_AGEMA_signal_12038 ;
    wire new_AGEMA_signal_12039 ;
    wire new_AGEMA_signal_12040 ;
    wire new_AGEMA_signal_12041 ;
    wire new_AGEMA_signal_12042 ;
    wire new_AGEMA_signal_12043 ;
    wire new_AGEMA_signal_12044 ;
    wire new_AGEMA_signal_12045 ;
    wire new_AGEMA_signal_12046 ;
    wire new_AGEMA_signal_12047 ;
    wire new_AGEMA_signal_12048 ;
    wire new_AGEMA_signal_12049 ;
    wire new_AGEMA_signal_12050 ;
    wire new_AGEMA_signal_12051 ;
    wire new_AGEMA_signal_12052 ;
    wire new_AGEMA_signal_12053 ;
    wire new_AGEMA_signal_12054 ;
    wire new_AGEMA_signal_12055 ;
    wire new_AGEMA_signal_12056 ;
    wire new_AGEMA_signal_12057 ;
    wire new_AGEMA_signal_12058 ;
    wire new_AGEMA_signal_12059 ;
    wire new_AGEMA_signal_12060 ;
    wire new_AGEMA_signal_12061 ;
    wire new_AGEMA_signal_12062 ;
    wire new_AGEMA_signal_12063 ;
    wire new_AGEMA_signal_12064 ;
    wire new_AGEMA_signal_12065 ;
    wire new_AGEMA_signal_12066 ;
    wire new_AGEMA_signal_12067 ;
    wire new_AGEMA_signal_12068 ;
    wire new_AGEMA_signal_12069 ;
    wire new_AGEMA_signal_12070 ;
    wire new_AGEMA_signal_12071 ;
    wire new_AGEMA_signal_12072 ;
    wire new_AGEMA_signal_12073 ;
    wire new_AGEMA_signal_12074 ;
    wire new_AGEMA_signal_12075 ;
    wire new_AGEMA_signal_12076 ;
    wire new_AGEMA_signal_12077 ;
    wire new_AGEMA_signal_12078 ;
    wire new_AGEMA_signal_12079 ;
    wire new_AGEMA_signal_12080 ;
    wire new_AGEMA_signal_12081 ;
    wire new_AGEMA_signal_12082 ;
    wire new_AGEMA_signal_12083 ;
    wire new_AGEMA_signal_12084 ;
    wire new_AGEMA_signal_12085 ;
    wire new_AGEMA_signal_12086 ;
    wire new_AGEMA_signal_12089 ;
    wire new_AGEMA_signal_12090 ;
    wire new_AGEMA_signal_12093 ;
    wire new_AGEMA_signal_12094 ;
    wire new_AGEMA_signal_12097 ;
    wire new_AGEMA_signal_12098 ;
    wire new_AGEMA_signal_12101 ;
    wire new_AGEMA_signal_12102 ;
    wire new_AGEMA_signal_12105 ;
    wire new_AGEMA_signal_12106 ;
    wire new_AGEMA_signal_12109 ;
    wire new_AGEMA_signal_12110 ;
    wire new_AGEMA_signal_12113 ;
    wire new_AGEMA_signal_12114 ;
    wire new_AGEMA_signal_12117 ;
    wire new_AGEMA_signal_12118 ;
    wire new_AGEMA_signal_12121 ;
    wire new_AGEMA_signal_12122 ;
    wire new_AGEMA_signal_12125 ;
    wire new_AGEMA_signal_12126 ;
    wire new_AGEMA_signal_12129 ;
    wire new_AGEMA_signal_12130 ;
    wire new_AGEMA_signal_12133 ;
    wire new_AGEMA_signal_12134 ;
    wire new_AGEMA_signal_12137 ;
    wire new_AGEMA_signal_12138 ;
    wire new_AGEMA_signal_12141 ;
    wire new_AGEMA_signal_12142 ;
    wire new_AGEMA_signal_12145 ;
    wire new_AGEMA_signal_12146 ;
    wire new_AGEMA_signal_12149 ;
    wire new_AGEMA_signal_12150 ;
    wire new_AGEMA_signal_12153 ;
    wire new_AGEMA_signal_12154 ;
    wire new_AGEMA_signal_12157 ;
    wire new_AGEMA_signal_12158 ;
    wire new_AGEMA_signal_12161 ;
    wire new_AGEMA_signal_12162 ;
    wire new_AGEMA_signal_12165 ;
    wire new_AGEMA_signal_12166 ;
    wire new_AGEMA_signal_12169 ;
    wire new_AGEMA_signal_12170 ;
    wire new_AGEMA_signal_12173 ;
    wire new_AGEMA_signal_12174 ;
    wire new_AGEMA_signal_12177 ;
    wire new_AGEMA_signal_12178 ;
    wire new_AGEMA_signal_12181 ;
    wire new_AGEMA_signal_12182 ;
    wire new_AGEMA_signal_12185 ;
    wire new_AGEMA_signal_12186 ;
    wire new_AGEMA_signal_12189 ;
    wire new_AGEMA_signal_12190 ;
    wire new_AGEMA_signal_12193 ;
    wire new_AGEMA_signal_12194 ;
    wire new_AGEMA_signal_12197 ;
    wire new_AGEMA_signal_12198 ;
    wire new_AGEMA_signal_12201 ;
    wire new_AGEMA_signal_12202 ;
    wire new_AGEMA_signal_12203 ;
    wire new_AGEMA_signal_12204 ;
    wire new_AGEMA_signal_12205 ;
    wire new_AGEMA_signal_12206 ;
    wire new_AGEMA_signal_12207 ;
    wire new_AGEMA_signal_12208 ;
    wire new_AGEMA_signal_12209 ;
    wire new_AGEMA_signal_12210 ;
    wire new_AGEMA_signal_12211 ;
    wire new_AGEMA_signal_12212 ;
    wire new_AGEMA_signal_12213 ;
    wire new_AGEMA_signal_12214 ;
    wire new_AGEMA_signal_12215 ;
    wire new_AGEMA_signal_12216 ;
    wire new_AGEMA_signal_12217 ;
    wire new_AGEMA_signal_12218 ;
    wire new_AGEMA_signal_12219 ;
    wire new_AGEMA_signal_12220 ;
    wire new_AGEMA_signal_12221 ;
    wire new_AGEMA_signal_12222 ;
    wire new_AGEMA_signal_12223 ;
    wire new_AGEMA_signal_12224 ;
    wire new_AGEMA_signal_12225 ;
    wire new_AGEMA_signal_12226 ;
    wire new_AGEMA_signal_12227 ;
    wire new_AGEMA_signal_12228 ;
    wire new_AGEMA_signal_12229 ;
    wire new_AGEMA_signal_12230 ;
    wire new_AGEMA_signal_12231 ;
    wire new_AGEMA_signal_12232 ;
    wire new_AGEMA_signal_12233 ;
    wire new_AGEMA_signal_12234 ;
    wire new_AGEMA_signal_12235 ;
    wire new_AGEMA_signal_12236 ;
    wire new_AGEMA_signal_12237 ;
    wire new_AGEMA_signal_12238 ;
    wire new_AGEMA_signal_12239 ;
    wire new_AGEMA_signal_12240 ;
    wire new_AGEMA_signal_12241 ;
    wire new_AGEMA_signal_12242 ;
    wire new_AGEMA_signal_12243 ;
    wire new_AGEMA_signal_12244 ;
    wire new_AGEMA_signal_12245 ;
    wire new_AGEMA_signal_12246 ;
    wire new_AGEMA_signal_12247 ;
    wire new_AGEMA_signal_12248 ;
    wire new_AGEMA_signal_12249 ;
    wire new_AGEMA_signal_12250 ;
    wire new_AGEMA_signal_12251 ;
    wire new_AGEMA_signal_12252 ;
    wire new_AGEMA_signal_12253 ;
    wire new_AGEMA_signal_12254 ;
    wire new_AGEMA_signal_12255 ;
    wire new_AGEMA_signal_12256 ;
    wire new_AGEMA_signal_12257 ;
    wire new_AGEMA_signal_12258 ;
    wire new_AGEMA_signal_12259 ;
    wire new_AGEMA_signal_12260 ;
    wire new_AGEMA_signal_12261 ;
    wire new_AGEMA_signal_12262 ;
    wire new_AGEMA_signal_12263 ;
    wire new_AGEMA_signal_12264 ;
    wire new_AGEMA_signal_12265 ;
    wire new_AGEMA_signal_12266 ;
    wire new_AGEMA_signal_12267 ;
    wire new_AGEMA_signal_12268 ;
    wire new_AGEMA_signal_12269 ;
    wire new_AGEMA_signal_12270 ;
    wire new_AGEMA_signal_12271 ;
    wire new_AGEMA_signal_12272 ;
    wire new_AGEMA_signal_12273 ;
    wire new_AGEMA_signal_12274 ;
    wire new_AGEMA_signal_12275 ;
    wire new_AGEMA_signal_12276 ;
    wire new_AGEMA_signal_12277 ;
    wire new_AGEMA_signal_12278 ;
    wire new_AGEMA_signal_12279 ;
    wire new_AGEMA_signal_12280 ;
    wire new_AGEMA_signal_12281 ;
    wire new_AGEMA_signal_12282 ;
    wire new_AGEMA_signal_12283 ;
    wire new_AGEMA_signal_12284 ;
    wire new_AGEMA_signal_12285 ;
    wire new_AGEMA_signal_12286 ;
    wire new_AGEMA_signal_12287 ;
    wire new_AGEMA_signal_12288 ;
    wire new_AGEMA_signal_12289 ;
    wire new_AGEMA_signal_12290 ;
    wire new_AGEMA_signal_12291 ;
    wire new_AGEMA_signal_12292 ;
    wire new_AGEMA_signal_12293 ;
    wire new_AGEMA_signal_12294 ;
    wire new_AGEMA_signal_12295 ;
    wire new_AGEMA_signal_12296 ;
    wire new_AGEMA_signal_12297 ;
    wire new_AGEMA_signal_12298 ;
    wire new_AGEMA_signal_12299 ;
    wire new_AGEMA_signal_12300 ;
    wire new_AGEMA_signal_12301 ;
    wire new_AGEMA_signal_12302 ;
    wire new_AGEMA_signal_12303 ;
    wire new_AGEMA_signal_12304 ;
    wire new_AGEMA_signal_12305 ;
    wire new_AGEMA_signal_12306 ;
    wire new_AGEMA_signal_12307 ;
    wire new_AGEMA_signal_12308 ;
    wire new_AGEMA_signal_12309 ;
    wire new_AGEMA_signal_12310 ;
    wire new_AGEMA_signal_12311 ;
    wire new_AGEMA_signal_12312 ;
    wire new_AGEMA_signal_12315 ;
    wire new_AGEMA_signal_12316 ;
    wire new_AGEMA_signal_12319 ;
    wire new_AGEMA_signal_12320 ;
    wire new_AGEMA_signal_12323 ;
    wire new_AGEMA_signal_12324 ;
    wire new_AGEMA_signal_12327 ;
    wire new_AGEMA_signal_12328 ;
    wire new_AGEMA_signal_12331 ;
    wire new_AGEMA_signal_12332 ;
    wire new_AGEMA_signal_12335 ;
    wire new_AGEMA_signal_12336 ;
    wire new_AGEMA_signal_12339 ;
    wire new_AGEMA_signal_12340 ;
    wire new_AGEMA_signal_12343 ;
    wire new_AGEMA_signal_12344 ;
    wire new_AGEMA_signal_12347 ;
    wire new_AGEMA_signal_12348 ;
    wire new_AGEMA_signal_12351 ;
    wire new_AGEMA_signal_12352 ;
    wire new_AGEMA_signal_12355 ;
    wire new_AGEMA_signal_12356 ;
    wire new_AGEMA_signal_12359 ;
    wire new_AGEMA_signal_12360 ;
    wire new_AGEMA_signal_12363 ;
    wire new_AGEMA_signal_12364 ;
    wire new_AGEMA_signal_12367 ;
    wire new_AGEMA_signal_12368 ;
    wire new_AGEMA_signal_12371 ;
    wire new_AGEMA_signal_12372 ;
    wire new_AGEMA_signal_12375 ;
    wire new_AGEMA_signal_12376 ;
    wire new_AGEMA_signal_12379 ;
    wire new_AGEMA_signal_12380 ;
    wire new_AGEMA_signal_12383 ;
    wire new_AGEMA_signal_12384 ;
    wire new_AGEMA_signal_12387 ;
    wire new_AGEMA_signal_12388 ;
    wire new_AGEMA_signal_12391 ;
    wire new_AGEMA_signal_12392 ;
    wire new_AGEMA_signal_12395 ;
    wire new_AGEMA_signal_12396 ;
    wire new_AGEMA_signal_12399 ;
    wire new_AGEMA_signal_12400 ;
    wire new_AGEMA_signal_12403 ;
    wire new_AGEMA_signal_12404 ;
    wire new_AGEMA_signal_12407 ;
    wire new_AGEMA_signal_12408 ;
    wire new_AGEMA_signal_12411 ;
    wire new_AGEMA_signal_12412 ;
    wire new_AGEMA_signal_12415 ;
    wire new_AGEMA_signal_12416 ;
    wire new_AGEMA_signal_12419 ;
    wire new_AGEMA_signal_12420 ;
    wire new_AGEMA_signal_12423 ;
    wire new_AGEMA_signal_12424 ;
    wire new_AGEMA_signal_12427 ;
    wire new_AGEMA_signal_12428 ;
    wire new_AGEMA_signal_12431 ;
    wire new_AGEMA_signal_12432 ;
    wire new_AGEMA_signal_12435 ;
    wire new_AGEMA_signal_12436 ;
    wire new_AGEMA_signal_12439 ;
    wire new_AGEMA_signal_12440 ;
    wire new_AGEMA_signal_12443 ;
    wire new_AGEMA_signal_12444 ;
    wire new_AGEMA_signal_12447 ;
    wire new_AGEMA_signal_12448 ;
    wire new_AGEMA_signal_12451 ;
    wire new_AGEMA_signal_12452 ;
    wire new_AGEMA_signal_12455 ;
    wire new_AGEMA_signal_12456 ;
    wire new_AGEMA_signal_12459 ;
    wire new_AGEMA_signal_12460 ;
    wire new_AGEMA_signal_12463 ;
    wire new_AGEMA_signal_12464 ;
    wire new_AGEMA_signal_12467 ;
    wire new_AGEMA_signal_12468 ;
    wire new_AGEMA_signal_12471 ;
    wire new_AGEMA_signal_12472 ;
    wire new_AGEMA_signal_12475 ;
    wire new_AGEMA_signal_12476 ;
    wire new_AGEMA_signal_12479 ;
    wire new_AGEMA_signal_12480 ;
    wire new_AGEMA_signal_12483 ;
    wire new_AGEMA_signal_12484 ;
    wire new_AGEMA_signal_12487 ;
    wire new_AGEMA_signal_12488 ;
    wire new_AGEMA_signal_12491 ;
    wire new_AGEMA_signal_12492 ;
    wire new_AGEMA_signal_12495 ;
    wire new_AGEMA_signal_12496 ;
    wire new_AGEMA_signal_12499 ;
    wire new_AGEMA_signal_12500 ;
    wire new_AGEMA_signal_12503 ;
    wire new_AGEMA_signal_12504 ;
    wire new_AGEMA_signal_12507 ;
    wire new_AGEMA_signal_12508 ;
    wire new_AGEMA_signal_12511 ;
    wire new_AGEMA_signal_12512 ;
    wire new_AGEMA_signal_12515 ;
    wire new_AGEMA_signal_12516 ;
    wire new_AGEMA_signal_12519 ;
    wire new_AGEMA_signal_12520 ;
    wire new_AGEMA_signal_12523 ;
    wire new_AGEMA_signal_12524 ;
    wire new_AGEMA_signal_12527 ;
    wire new_AGEMA_signal_12528 ;
    wire new_AGEMA_signal_12531 ;
    wire new_AGEMA_signal_12532 ;
    wire new_AGEMA_signal_12535 ;
    wire new_AGEMA_signal_12536 ;
    wire new_AGEMA_signal_12539 ;
    wire new_AGEMA_signal_12540 ;
    wire new_AGEMA_signal_12543 ;
    wire new_AGEMA_signal_12544 ;
    wire new_AGEMA_signal_12547 ;
    wire new_AGEMA_signal_12548 ;
    wire new_AGEMA_signal_12551 ;
    wire new_AGEMA_signal_12552 ;
    wire new_AGEMA_signal_12555 ;
    wire new_AGEMA_signal_12556 ;
    wire new_AGEMA_signal_12559 ;
    wire new_AGEMA_signal_12560 ;
    wire new_AGEMA_signal_12563 ;
    wire new_AGEMA_signal_12564 ;
    wire new_AGEMA_signal_12567 ;
    wire new_AGEMA_signal_12568 ;
    wire new_AGEMA_signal_12571 ;
    wire new_AGEMA_signal_12572 ;
    wire new_AGEMA_signal_12575 ;
    wire new_AGEMA_signal_12576 ;
    wire new_AGEMA_signal_12579 ;
    wire new_AGEMA_signal_12580 ;
    wire new_AGEMA_signal_12583 ;
    wire new_AGEMA_signal_12584 ;
    wire new_AGEMA_signal_12587 ;
    wire new_AGEMA_signal_12588 ;
    wire new_AGEMA_signal_12591 ;
    wire new_AGEMA_signal_12592 ;
    wire new_AGEMA_signal_12595 ;
    wire new_AGEMA_signal_12596 ;
    wire new_AGEMA_signal_12599 ;
    wire new_AGEMA_signal_12600 ;
    wire new_AGEMA_signal_12603 ;
    wire new_AGEMA_signal_12604 ;
    wire new_AGEMA_signal_12607 ;
    wire new_AGEMA_signal_12608 ;
    wire new_AGEMA_signal_12611 ;
    wire new_AGEMA_signal_12612 ;
    wire new_AGEMA_signal_12615 ;
    wire new_AGEMA_signal_12616 ;
    wire new_AGEMA_signal_12619 ;
    wire new_AGEMA_signal_12620 ;
    wire new_AGEMA_signal_12623 ;
    wire new_AGEMA_signal_12624 ;
    wire new_AGEMA_signal_12627 ;
    wire new_AGEMA_signal_12628 ;
    wire new_AGEMA_signal_12631 ;
    wire new_AGEMA_signal_12632 ;
    wire new_AGEMA_signal_12635 ;
    wire new_AGEMA_signal_12636 ;
    wire new_AGEMA_signal_12639 ;
    wire new_AGEMA_signal_12640 ;
    wire new_AGEMA_signal_12643 ;
    wire new_AGEMA_signal_12644 ;
    wire new_AGEMA_signal_12647 ;
    wire new_AGEMA_signal_12648 ;
    wire new_AGEMA_signal_12651 ;
    wire new_AGEMA_signal_12652 ;
    wire new_AGEMA_signal_12655 ;
    wire new_AGEMA_signal_12656 ;
    wire new_AGEMA_signal_12659 ;
    wire new_AGEMA_signal_12660 ;
    wire new_AGEMA_signal_12663 ;
    wire new_AGEMA_signal_12664 ;
    wire new_AGEMA_signal_12667 ;
    wire new_AGEMA_signal_12668 ;
    wire new_AGEMA_signal_12671 ;
    wire new_AGEMA_signal_12672 ;
    wire new_AGEMA_signal_12675 ;
    wire new_AGEMA_signal_12676 ;
    wire new_AGEMA_signal_12679 ;
    wire new_AGEMA_signal_12680 ;
    wire new_AGEMA_signal_12683 ;
    wire new_AGEMA_signal_12684 ;
    wire new_AGEMA_signal_12687 ;
    wire new_AGEMA_signal_12688 ;
    wire new_AGEMA_signal_12691 ;
    wire new_AGEMA_signal_12692 ;
    wire new_AGEMA_signal_12695 ;
    wire new_AGEMA_signal_12696 ;
    wire new_AGEMA_signal_12699 ;
    wire new_AGEMA_signal_12700 ;
    wire new_AGEMA_signal_12703 ;
    wire new_AGEMA_signal_12704 ;
    wire new_AGEMA_signal_12707 ;
    wire new_AGEMA_signal_12708 ;
    wire new_AGEMA_signal_12711 ;
    wire new_AGEMA_signal_12712 ;
    wire new_AGEMA_signal_12715 ;
    wire new_AGEMA_signal_12716 ;
    wire new_AGEMA_signal_12719 ;
    wire new_AGEMA_signal_12720 ;
    wire new_AGEMA_signal_12723 ;
    wire new_AGEMA_signal_12724 ;
    wire new_AGEMA_signal_12727 ;
    wire new_AGEMA_signal_12728 ;
    wire new_AGEMA_signal_12731 ;
    wire new_AGEMA_signal_12732 ;
    wire new_AGEMA_signal_12735 ;
    wire new_AGEMA_signal_12736 ;
    wire new_AGEMA_signal_12739 ;
    wire new_AGEMA_signal_12740 ;
    wire new_AGEMA_signal_12743 ;
    wire new_AGEMA_signal_12744 ;
    wire new_AGEMA_signal_12747 ;
    wire new_AGEMA_signal_12748 ;
    wire new_AGEMA_signal_12751 ;
    wire new_AGEMA_signal_12752 ;
    wire new_AGEMA_signal_12755 ;
    wire new_AGEMA_signal_12756 ;
    wire new_AGEMA_signal_12759 ;
    wire new_AGEMA_signal_12760 ;
    wire new_AGEMA_signal_12763 ;
    wire new_AGEMA_signal_12764 ;
    wire new_AGEMA_signal_12767 ;
    wire new_AGEMA_signal_12768 ;
    wire new_AGEMA_signal_12771 ;
    wire new_AGEMA_signal_12772 ;
    wire new_AGEMA_signal_12775 ;
    wire new_AGEMA_signal_12776 ;
    wire new_AGEMA_signal_12779 ;
    wire new_AGEMA_signal_12780 ;
    wire new_AGEMA_signal_12783 ;
    wire new_AGEMA_signal_12784 ;
    wire new_AGEMA_signal_12787 ;
    wire new_AGEMA_signal_12788 ;
    wire new_AGEMA_signal_12791 ;
    wire new_AGEMA_signal_12792 ;
    wire new_AGEMA_signal_12795 ;
    wire new_AGEMA_signal_12796 ;
    wire new_AGEMA_signal_12799 ;
    wire new_AGEMA_signal_12800 ;
    wire new_AGEMA_signal_12803 ;
    wire new_AGEMA_signal_12804 ;
    wire new_AGEMA_signal_12807 ;
    wire new_AGEMA_signal_12808 ;
    wire new_AGEMA_signal_12811 ;
    wire new_AGEMA_signal_12812 ;
    wire new_AGEMA_signal_12815 ;
    wire new_AGEMA_signal_12816 ;
    wire new_AGEMA_signal_12819 ;
    wire new_AGEMA_signal_12820 ;
    wire new_AGEMA_signal_12823 ;
    wire new_AGEMA_signal_12824 ;
    wire new_AGEMA_signal_12827 ;
    wire new_AGEMA_signal_12828 ;
    wire new_AGEMA_signal_12831 ;
    wire new_AGEMA_signal_12832 ;
    wire new_AGEMA_signal_12835 ;
    wire new_AGEMA_signal_12836 ;
    wire new_AGEMA_signal_12839 ;
    wire new_AGEMA_signal_12840 ;
    wire new_AGEMA_signal_12843 ;
    wire new_AGEMA_signal_12844 ;
    wire new_AGEMA_signal_12847 ;
    wire new_AGEMA_signal_12848 ;
    wire new_AGEMA_signal_12851 ;
    wire new_AGEMA_signal_12852 ;
    wire clk_gated ;

    /* cells in depth 0 */
    INV_X1 U830 ( .A (n314), .ZN (n319) ) ;
    INV_X1 U831 ( .A (n314), .ZN (n320) ) ;
    INV_X1 U832 ( .A (n314), .ZN (n317) ) ;
    INV_X1 U833 ( .A (n314), .ZN (n315) ) ;
    INV_X1 U834 ( .A (n314), .ZN (n316) ) ;
    INV_X1 U835 ( .A (n314), .ZN (n318) ) ;
    NOR2_X1 U836 ( .A1 (n325), .A2 (n330), .ZN (n314) ) ;
    INV_X1 U837 ( .A (RoundCounter[0]), .ZN (n325) ) ;
    INV_X1 U838 ( .A (n314), .ZN (n321) ) ;
    NOR2_X1 U839 ( .A1 (RoundCounter[2]), .A2 (RoundCounter[1]), .ZN (n323) ) ;
    INV_X1 U840 ( .A (n323), .ZN (n322) ) ;
    NOR2_X1 U841 ( .A1 (RoundCounter[0]), .A2 (n322), .ZN (Rcon[0]) ) ;
    NOR2_X1 U842 ( .A1 (RoundCounter[0]), .A2 (RoundCounter[3]), .ZN (n337) ) ;
    NOR2_X1 U843 ( .A1 (n337), .A2 (n322), .ZN (Rcon[1]) ) ;
    NAND2_X1 U844 ( .A1 (RoundCounter[3]), .A2 (n323), .ZN (n330) ) ;
    INV_X1 U845 ( .A (RoundCounter[2]), .ZN (n328) ) ;
    AND2_X1 U846 ( .A1 (n328), .A2 (RoundCounter[1]), .ZN (n333) ) ;
    NAND2_X1 U847 ( .A1 (n337), .A2 (n333), .ZN (n324) ) ;
    NAND2_X1 U848 ( .A1 (n321), .A2 (n324), .ZN (Rcon[2]) ) ;
    NOR2_X1 U849 ( .A1 (RoundCounter[3]), .A2 (n325), .ZN (n335) ) ;
    NAND2_X1 U850 ( .A1 (n333), .A2 (n335), .ZN (n327) ) ;
    NAND2_X1 U851 ( .A1 (RoundCounter[3]), .A2 (Rcon[0]), .ZN (n326) ) ;
    NAND2_X1 U852 ( .A1 (n327), .A2 (n326), .ZN (Rcon[3]) ) ;
    NOR2_X1 U853 ( .A1 (RoundCounter[1]), .A2 (n328), .ZN (n331) ) ;
    NAND2_X1 U854 ( .A1 (n337), .A2 (n331), .ZN (n329) ) ;
    NAND2_X1 U855 ( .A1 (n330), .A2 (n329), .ZN (Rcon[4]) ) ;
    NAND2_X1 U856 ( .A1 (n335), .A2 (n331), .ZN (n332) ) ;
    NAND2_X1 U857 ( .A1 (n321), .A2 (n332), .ZN (Rcon[5]) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U986 ( .a ({new_AGEMA_signal_4550, new_AGEMA_signal_4549, RoundInput[0]}), .b ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, RoundKey[0]}), .c ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U987 ( .a ({new_AGEMA_signal_4556, new_AGEMA_signal_4555, RoundInput[100]}), .b ({new_AGEMA_signal_4558, new_AGEMA_signal_4557, RoundKey[100]}), .c ({ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U988 ( .a ({new_AGEMA_signal_4562, new_AGEMA_signal_4561, RoundInput[101]}), .b ({new_AGEMA_signal_4564, new_AGEMA_signal_4563, RoundKey[101]}), .c ({ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U989 ( .a ({new_AGEMA_signal_4568, new_AGEMA_signal_4567, RoundInput[102]}), .b ({new_AGEMA_signal_4570, new_AGEMA_signal_4569, RoundKey[102]}), .c ({ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U990 ( .a ({new_AGEMA_signal_4574, new_AGEMA_signal_4573, RoundInput[103]}), .b ({new_AGEMA_signal_4576, new_AGEMA_signal_4575, RoundKey[103]}), .c ({ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U991 ( .a ({new_AGEMA_signal_4580, new_AGEMA_signal_4579, RoundInput[104]}), .b ({new_AGEMA_signal_4582, new_AGEMA_signal_4581, RoundKey[104]}), .c ({ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U992 ( .a ({new_AGEMA_signal_4586, new_AGEMA_signal_4585, RoundInput[105]}), .b ({new_AGEMA_signal_4588, new_AGEMA_signal_4587, RoundKey[105]}), .c ({ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U993 ( .a ({new_AGEMA_signal_4592, new_AGEMA_signal_4591, RoundInput[106]}), .b ({new_AGEMA_signal_4594, new_AGEMA_signal_4593, RoundKey[106]}), .c ({ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U994 ( .a ({new_AGEMA_signal_4598, new_AGEMA_signal_4597, RoundInput[107]}), .b ({new_AGEMA_signal_4600, new_AGEMA_signal_4599, RoundKey[107]}), .c ({ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U995 ( .a ({new_AGEMA_signal_4604, new_AGEMA_signal_4603, RoundInput[108]}), .b ({new_AGEMA_signal_4606, new_AGEMA_signal_4605, RoundKey[108]}), .c ({ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U996 ( .a ({new_AGEMA_signal_4610, new_AGEMA_signal_4609, RoundInput[109]}), .b ({new_AGEMA_signal_4612, new_AGEMA_signal_4611, RoundKey[109]}), .c ({ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U997 ( .a ({new_AGEMA_signal_4616, new_AGEMA_signal_4615, RoundInput[10]}), .b ({new_AGEMA_signal_4618, new_AGEMA_signal_4617, RoundKey[10]}), .c ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U998 ( .a ({new_AGEMA_signal_4622, new_AGEMA_signal_4621, RoundInput[110]}), .b ({new_AGEMA_signal_4624, new_AGEMA_signal_4623, RoundKey[110]}), .c ({ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U999 ( .a ({new_AGEMA_signal_4628, new_AGEMA_signal_4627, RoundInput[111]}), .b ({new_AGEMA_signal_4630, new_AGEMA_signal_4629, RoundKey[111]}), .c ({ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1000 ( .a ({new_AGEMA_signal_4634, new_AGEMA_signal_4633, RoundInput[112]}), .b ({new_AGEMA_signal_4636, new_AGEMA_signal_4635, RoundKey[112]}), .c ({ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1001 ( .a ({new_AGEMA_signal_4640, new_AGEMA_signal_4639, RoundInput[113]}), .b ({new_AGEMA_signal_4642, new_AGEMA_signal_4641, RoundKey[113]}), .c ({ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1002 ( .a ({new_AGEMA_signal_4646, new_AGEMA_signal_4645, RoundInput[114]}), .b ({new_AGEMA_signal_4648, new_AGEMA_signal_4647, RoundKey[114]}), .c ({ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1003 ( .a ({new_AGEMA_signal_4652, new_AGEMA_signal_4651, RoundInput[115]}), .b ({new_AGEMA_signal_4654, new_AGEMA_signal_4653, RoundKey[115]}), .c ({ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1004 ( .a ({new_AGEMA_signal_4658, new_AGEMA_signal_4657, RoundInput[116]}), .b ({new_AGEMA_signal_4660, new_AGEMA_signal_4659, RoundKey[116]}), .c ({ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1005 ( .a ({new_AGEMA_signal_4664, new_AGEMA_signal_4663, RoundInput[117]}), .b ({new_AGEMA_signal_4666, new_AGEMA_signal_4665, RoundKey[117]}), .c ({ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1006 ( .a ({new_AGEMA_signal_4670, new_AGEMA_signal_4669, RoundInput[118]}), .b ({new_AGEMA_signal_4672, new_AGEMA_signal_4671, RoundKey[118]}), .c ({ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1007 ( .a ({new_AGEMA_signal_4676, new_AGEMA_signal_4675, RoundInput[119]}), .b ({new_AGEMA_signal_4678, new_AGEMA_signal_4677, RoundKey[119]}), .c ({ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1008 ( .a ({new_AGEMA_signal_4682, new_AGEMA_signal_4681, RoundInput[11]}), .b ({new_AGEMA_signal_4684, new_AGEMA_signal_4683, RoundKey[11]}), .c ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1009 ( .a ({new_AGEMA_signal_4688, new_AGEMA_signal_4687, RoundInput[120]}), .b ({new_AGEMA_signal_4690, new_AGEMA_signal_4689, RoundKey[120]}), .c ({ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1010 ( .a ({new_AGEMA_signal_4694, new_AGEMA_signal_4693, RoundInput[121]}), .b ({new_AGEMA_signal_4696, new_AGEMA_signal_4695, RoundKey[121]}), .c ({ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1011 ( .a ({new_AGEMA_signal_4700, new_AGEMA_signal_4699, RoundInput[122]}), .b ({new_AGEMA_signal_4702, new_AGEMA_signal_4701, RoundKey[122]}), .c ({ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1012 ( .a ({new_AGEMA_signal_4706, new_AGEMA_signal_4705, RoundInput[123]}), .b ({new_AGEMA_signal_4708, new_AGEMA_signal_4707, RoundKey[123]}), .c ({ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1013 ( .a ({new_AGEMA_signal_4712, new_AGEMA_signal_4711, RoundInput[124]}), .b ({new_AGEMA_signal_4714, new_AGEMA_signal_4713, RoundKey[124]}), .c ({ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1014 ( .a ({new_AGEMA_signal_4718, new_AGEMA_signal_4717, RoundInput[125]}), .b ({new_AGEMA_signal_4720, new_AGEMA_signal_4719, RoundKey[125]}), .c ({ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1015 ( .a ({new_AGEMA_signal_4724, new_AGEMA_signal_4723, RoundInput[126]}), .b ({new_AGEMA_signal_4726, new_AGEMA_signal_4725, RoundKey[126]}), .c ({ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1016 ( .a ({new_AGEMA_signal_4730, new_AGEMA_signal_4729, RoundInput[127]}), .b ({new_AGEMA_signal_4732, new_AGEMA_signal_4731, RoundKey[127]}), .c ({ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1017 ( .a ({new_AGEMA_signal_4736, new_AGEMA_signal_4735, RoundInput[12]}), .b ({new_AGEMA_signal_4738, new_AGEMA_signal_4737, RoundKey[12]}), .c ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1018 ( .a ({new_AGEMA_signal_4742, new_AGEMA_signal_4741, RoundInput[13]}), .b ({new_AGEMA_signal_4744, new_AGEMA_signal_4743, RoundKey[13]}), .c ({ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1019 ( .a ({new_AGEMA_signal_4748, new_AGEMA_signal_4747, RoundInput[14]}), .b ({new_AGEMA_signal_4750, new_AGEMA_signal_4749, RoundKey[14]}), .c ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1020 ( .a ({new_AGEMA_signal_4754, new_AGEMA_signal_4753, RoundInput[15]}), .b ({new_AGEMA_signal_4756, new_AGEMA_signal_4755, RoundKey[15]}), .c ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1021 ( .a ({new_AGEMA_signal_4760, new_AGEMA_signal_4759, RoundInput[16]}), .b ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, RoundKey[16]}), .c ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1022 ( .a ({new_AGEMA_signal_4766, new_AGEMA_signal_4765, RoundInput[17]}), .b ({new_AGEMA_signal_4768, new_AGEMA_signal_4767, RoundKey[17]}), .c ({ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1023 ( .a ({new_AGEMA_signal_4772, new_AGEMA_signal_4771, RoundInput[18]}), .b ({new_AGEMA_signal_4774, new_AGEMA_signal_4773, RoundKey[18]}), .c ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1024 ( .a ({new_AGEMA_signal_4778, new_AGEMA_signal_4777, RoundInput[19]}), .b ({new_AGEMA_signal_4780, new_AGEMA_signal_4779, RoundKey[19]}), .c ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1025 ( .a ({new_AGEMA_signal_4784, new_AGEMA_signal_4783, RoundInput[1]}), .b ({new_AGEMA_signal_4786, new_AGEMA_signal_4785, RoundKey[1]}), .c ({ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1026 ( .a ({new_AGEMA_signal_4790, new_AGEMA_signal_4789, RoundInput[20]}), .b ({new_AGEMA_signal_4792, new_AGEMA_signal_4791, RoundKey[20]}), .c ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1027 ( .a ({new_AGEMA_signal_4796, new_AGEMA_signal_4795, RoundInput[21]}), .b ({new_AGEMA_signal_4798, new_AGEMA_signal_4797, RoundKey[21]}), .c ({ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1028 ( .a ({new_AGEMA_signal_4802, new_AGEMA_signal_4801, RoundInput[22]}), .b ({new_AGEMA_signal_4804, new_AGEMA_signal_4803, RoundKey[22]}), .c ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1029 ( .a ({new_AGEMA_signal_4808, new_AGEMA_signal_4807, RoundInput[23]}), .b ({new_AGEMA_signal_4810, new_AGEMA_signal_4809, RoundKey[23]}), .c ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1030 ( .a ({new_AGEMA_signal_4814, new_AGEMA_signal_4813, RoundInput[24]}), .b ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, RoundKey[24]}), .c ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1031 ( .a ({new_AGEMA_signal_4820, new_AGEMA_signal_4819, RoundInput[25]}), .b ({new_AGEMA_signal_4822, new_AGEMA_signal_4821, RoundKey[25]}), .c ({ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1032 ( .a ({new_AGEMA_signal_4826, new_AGEMA_signal_4825, RoundInput[26]}), .b ({new_AGEMA_signal_4828, new_AGEMA_signal_4827, RoundKey[26]}), .c ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1033 ( .a ({new_AGEMA_signal_4832, new_AGEMA_signal_4831, RoundInput[27]}), .b ({new_AGEMA_signal_4834, new_AGEMA_signal_4833, RoundKey[27]}), .c ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1034 ( .a ({new_AGEMA_signal_4838, new_AGEMA_signal_4837, RoundInput[28]}), .b ({new_AGEMA_signal_4840, new_AGEMA_signal_4839, RoundKey[28]}), .c ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1035 ( .a ({new_AGEMA_signal_4844, new_AGEMA_signal_4843, RoundInput[29]}), .b ({new_AGEMA_signal_4846, new_AGEMA_signal_4845, RoundKey[29]}), .c ({ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1036 ( .a ({new_AGEMA_signal_4850, new_AGEMA_signal_4849, RoundInput[2]}), .b ({new_AGEMA_signal_4852, new_AGEMA_signal_4851, RoundKey[2]}), .c ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1037 ( .a ({new_AGEMA_signal_4856, new_AGEMA_signal_4855, RoundInput[30]}), .b ({new_AGEMA_signal_4858, new_AGEMA_signal_4857, RoundKey[30]}), .c ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1038 ( .a ({new_AGEMA_signal_4862, new_AGEMA_signal_4861, RoundInput[31]}), .b ({new_AGEMA_signal_4864, new_AGEMA_signal_4863, RoundKey[31]}), .c ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1039 ( .a ({new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundInput[32]}), .b ({new_AGEMA_signal_4870, new_AGEMA_signal_4869, RoundKey[32]}), .c ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1040 ( .a ({new_AGEMA_signal_4874, new_AGEMA_signal_4873, RoundInput[33]}), .b ({new_AGEMA_signal_4876, new_AGEMA_signal_4875, RoundKey[33]}), .c ({ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1041 ( .a ({new_AGEMA_signal_4880, new_AGEMA_signal_4879, RoundInput[34]}), .b ({new_AGEMA_signal_4882, new_AGEMA_signal_4881, RoundKey[34]}), .c ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1042 ( .a ({new_AGEMA_signal_4886, new_AGEMA_signal_4885, RoundInput[35]}), .b ({new_AGEMA_signal_4888, new_AGEMA_signal_4887, RoundKey[35]}), .c ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1043 ( .a ({new_AGEMA_signal_4892, new_AGEMA_signal_4891, RoundInput[36]}), .b ({new_AGEMA_signal_4894, new_AGEMA_signal_4893, RoundKey[36]}), .c ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1044 ( .a ({new_AGEMA_signal_4898, new_AGEMA_signal_4897, RoundInput[37]}), .b ({new_AGEMA_signal_4900, new_AGEMA_signal_4899, RoundKey[37]}), .c ({ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1045 ( .a ({new_AGEMA_signal_4904, new_AGEMA_signal_4903, RoundInput[38]}), .b ({new_AGEMA_signal_4906, new_AGEMA_signal_4905, RoundKey[38]}), .c ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1046 ( .a ({new_AGEMA_signal_4910, new_AGEMA_signal_4909, RoundInput[39]}), .b ({new_AGEMA_signal_4912, new_AGEMA_signal_4911, RoundKey[39]}), .c ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1047 ( .a ({new_AGEMA_signal_4916, new_AGEMA_signal_4915, RoundInput[3]}), .b ({new_AGEMA_signal_4918, new_AGEMA_signal_4917, RoundKey[3]}), .c ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1048 ( .a ({new_AGEMA_signal_4922, new_AGEMA_signal_4921, RoundInput[40]}), .b ({new_AGEMA_signal_4924, new_AGEMA_signal_4923, RoundKey[40]}), .c ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1049 ( .a ({new_AGEMA_signal_4928, new_AGEMA_signal_4927, RoundInput[41]}), .b ({new_AGEMA_signal_4930, new_AGEMA_signal_4929, RoundKey[41]}), .c ({ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1050 ( .a ({new_AGEMA_signal_4934, new_AGEMA_signal_4933, RoundInput[42]}), .b ({new_AGEMA_signal_4936, new_AGEMA_signal_4935, RoundKey[42]}), .c ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1051 ( .a ({new_AGEMA_signal_4940, new_AGEMA_signal_4939, RoundInput[43]}), .b ({new_AGEMA_signal_4942, new_AGEMA_signal_4941, RoundKey[43]}), .c ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1052 ( .a ({new_AGEMA_signal_4946, new_AGEMA_signal_4945, RoundInput[44]}), .b ({new_AGEMA_signal_4948, new_AGEMA_signal_4947, RoundKey[44]}), .c ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1053 ( .a ({new_AGEMA_signal_4952, new_AGEMA_signal_4951, RoundInput[45]}), .b ({new_AGEMA_signal_4954, new_AGEMA_signal_4953, RoundKey[45]}), .c ({ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1054 ( .a ({new_AGEMA_signal_4958, new_AGEMA_signal_4957, RoundInput[46]}), .b ({new_AGEMA_signal_4960, new_AGEMA_signal_4959, RoundKey[46]}), .c ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1055 ( .a ({new_AGEMA_signal_4964, new_AGEMA_signal_4963, RoundInput[47]}), .b ({new_AGEMA_signal_4966, new_AGEMA_signal_4965, RoundKey[47]}), .c ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1056 ( .a ({new_AGEMA_signal_4970, new_AGEMA_signal_4969, RoundInput[48]}), .b ({new_AGEMA_signal_4972, new_AGEMA_signal_4971, RoundKey[48]}), .c ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1057 ( .a ({new_AGEMA_signal_4976, new_AGEMA_signal_4975, RoundInput[49]}), .b ({new_AGEMA_signal_4978, new_AGEMA_signal_4977, RoundKey[49]}), .c ({ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1058 ( .a ({new_AGEMA_signal_4982, new_AGEMA_signal_4981, RoundInput[4]}), .b ({new_AGEMA_signal_4984, new_AGEMA_signal_4983, RoundKey[4]}), .c ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1059 ( .a ({new_AGEMA_signal_4988, new_AGEMA_signal_4987, RoundInput[50]}), .b ({new_AGEMA_signal_4990, new_AGEMA_signal_4989, RoundKey[50]}), .c ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1060 ( .a ({new_AGEMA_signal_4994, new_AGEMA_signal_4993, RoundInput[51]}), .b ({new_AGEMA_signal_4996, new_AGEMA_signal_4995, RoundKey[51]}), .c ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1061 ( .a ({new_AGEMA_signal_5000, new_AGEMA_signal_4999, RoundInput[52]}), .b ({new_AGEMA_signal_5002, new_AGEMA_signal_5001, RoundKey[52]}), .c ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1062 ( .a ({new_AGEMA_signal_5006, new_AGEMA_signal_5005, RoundInput[53]}), .b ({new_AGEMA_signal_5008, new_AGEMA_signal_5007, RoundKey[53]}), .c ({ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1063 ( .a ({new_AGEMA_signal_5012, new_AGEMA_signal_5011, RoundInput[54]}), .b ({new_AGEMA_signal_5014, new_AGEMA_signal_5013, RoundKey[54]}), .c ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1064 ( .a ({new_AGEMA_signal_5018, new_AGEMA_signal_5017, RoundInput[55]}), .b ({new_AGEMA_signal_5020, new_AGEMA_signal_5019, RoundKey[55]}), .c ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1065 ( .a ({new_AGEMA_signal_5024, new_AGEMA_signal_5023, RoundInput[56]}), .b ({new_AGEMA_signal_5026, new_AGEMA_signal_5025, RoundKey[56]}), .c ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1066 ( .a ({new_AGEMA_signal_5030, new_AGEMA_signal_5029, RoundInput[57]}), .b ({new_AGEMA_signal_5032, new_AGEMA_signal_5031, RoundKey[57]}), .c ({ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1067 ( .a ({new_AGEMA_signal_5036, new_AGEMA_signal_5035, RoundInput[58]}), .b ({new_AGEMA_signal_5038, new_AGEMA_signal_5037, RoundKey[58]}), .c ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1068 ( .a ({new_AGEMA_signal_5042, new_AGEMA_signal_5041, RoundInput[59]}), .b ({new_AGEMA_signal_5044, new_AGEMA_signal_5043, RoundKey[59]}), .c ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1069 ( .a ({new_AGEMA_signal_5048, new_AGEMA_signal_5047, RoundInput[5]}), .b ({new_AGEMA_signal_5050, new_AGEMA_signal_5049, RoundKey[5]}), .c ({ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1070 ( .a ({new_AGEMA_signal_5054, new_AGEMA_signal_5053, RoundInput[60]}), .b ({new_AGEMA_signal_5056, new_AGEMA_signal_5055, RoundKey[60]}), .c ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1071 ( .a ({new_AGEMA_signal_5060, new_AGEMA_signal_5059, RoundInput[61]}), .b ({new_AGEMA_signal_5062, new_AGEMA_signal_5061, RoundKey[61]}), .c ({ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1072 ( .a ({new_AGEMA_signal_5066, new_AGEMA_signal_5065, RoundInput[62]}), .b ({new_AGEMA_signal_5068, new_AGEMA_signal_5067, RoundKey[62]}), .c ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1073 ( .a ({new_AGEMA_signal_5072, new_AGEMA_signal_5071, RoundInput[63]}), .b ({new_AGEMA_signal_5074, new_AGEMA_signal_5073, RoundKey[63]}), .c ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1074 ( .a ({new_AGEMA_signal_5078, new_AGEMA_signal_5077, RoundInput[64]}), .b ({new_AGEMA_signal_5080, new_AGEMA_signal_5079, RoundKey[64]}), .c ({ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1075 ( .a ({new_AGEMA_signal_5084, new_AGEMA_signal_5083, RoundInput[65]}), .b ({new_AGEMA_signal_5086, new_AGEMA_signal_5085, RoundKey[65]}), .c ({ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1076 ( .a ({new_AGEMA_signal_5090, new_AGEMA_signal_5089, RoundInput[66]}), .b ({new_AGEMA_signal_5092, new_AGEMA_signal_5091, RoundKey[66]}), .c ({ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1077 ( .a ({new_AGEMA_signal_5096, new_AGEMA_signal_5095, RoundInput[67]}), .b ({new_AGEMA_signal_5098, new_AGEMA_signal_5097, RoundKey[67]}), .c ({ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1078 ( .a ({new_AGEMA_signal_5102, new_AGEMA_signal_5101, RoundInput[68]}), .b ({new_AGEMA_signal_5104, new_AGEMA_signal_5103, RoundKey[68]}), .c ({ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1079 ( .a ({new_AGEMA_signal_5108, new_AGEMA_signal_5107, RoundInput[69]}), .b ({new_AGEMA_signal_5110, new_AGEMA_signal_5109, RoundKey[69]}), .c ({ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1080 ( .a ({new_AGEMA_signal_5114, new_AGEMA_signal_5113, RoundInput[6]}), .b ({new_AGEMA_signal_5116, new_AGEMA_signal_5115, RoundKey[6]}), .c ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1081 ( .a ({new_AGEMA_signal_5120, new_AGEMA_signal_5119, RoundInput[70]}), .b ({new_AGEMA_signal_5122, new_AGEMA_signal_5121, RoundKey[70]}), .c ({ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1082 ( .a ({new_AGEMA_signal_5126, new_AGEMA_signal_5125, RoundInput[71]}), .b ({new_AGEMA_signal_5128, new_AGEMA_signal_5127, RoundKey[71]}), .c ({ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1083 ( .a ({new_AGEMA_signal_5132, new_AGEMA_signal_5131, RoundInput[72]}), .b ({new_AGEMA_signal_5134, new_AGEMA_signal_5133, RoundKey[72]}), .c ({ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1084 ( .a ({new_AGEMA_signal_5138, new_AGEMA_signal_5137, RoundInput[73]}), .b ({new_AGEMA_signal_5140, new_AGEMA_signal_5139, RoundKey[73]}), .c ({ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1085 ( .a ({new_AGEMA_signal_5144, new_AGEMA_signal_5143, RoundInput[74]}), .b ({new_AGEMA_signal_5146, new_AGEMA_signal_5145, RoundKey[74]}), .c ({ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1086 ( .a ({new_AGEMA_signal_5150, new_AGEMA_signal_5149, RoundInput[75]}), .b ({new_AGEMA_signal_5152, new_AGEMA_signal_5151, RoundKey[75]}), .c ({ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1087 ( .a ({new_AGEMA_signal_5156, new_AGEMA_signal_5155, RoundInput[76]}), .b ({new_AGEMA_signal_5158, new_AGEMA_signal_5157, RoundKey[76]}), .c ({ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1088 ( .a ({new_AGEMA_signal_5162, new_AGEMA_signal_5161, RoundInput[77]}), .b ({new_AGEMA_signal_5164, new_AGEMA_signal_5163, RoundKey[77]}), .c ({ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1089 ( .a ({new_AGEMA_signal_5168, new_AGEMA_signal_5167, RoundInput[78]}), .b ({new_AGEMA_signal_5170, new_AGEMA_signal_5169, RoundKey[78]}), .c ({ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1090 ( .a ({new_AGEMA_signal_5174, new_AGEMA_signal_5173, RoundInput[79]}), .b ({new_AGEMA_signal_5176, new_AGEMA_signal_5175, RoundKey[79]}), .c ({ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1091 ( .a ({new_AGEMA_signal_5180, new_AGEMA_signal_5179, RoundInput[7]}), .b ({new_AGEMA_signal_5182, new_AGEMA_signal_5181, RoundKey[7]}), .c ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1092 ( .a ({new_AGEMA_signal_5186, new_AGEMA_signal_5185, RoundInput[80]}), .b ({new_AGEMA_signal_5188, new_AGEMA_signal_5187, RoundKey[80]}), .c ({ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1093 ( .a ({new_AGEMA_signal_5192, new_AGEMA_signal_5191, RoundInput[81]}), .b ({new_AGEMA_signal_5194, new_AGEMA_signal_5193, RoundKey[81]}), .c ({ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1094 ( .a ({new_AGEMA_signal_5198, new_AGEMA_signal_5197, RoundInput[82]}), .b ({new_AGEMA_signal_5200, new_AGEMA_signal_5199, RoundKey[82]}), .c ({ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1095 ( .a ({new_AGEMA_signal_5204, new_AGEMA_signal_5203, RoundInput[83]}), .b ({new_AGEMA_signal_5206, new_AGEMA_signal_5205, RoundKey[83]}), .c ({ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1096 ( .a ({new_AGEMA_signal_5210, new_AGEMA_signal_5209, RoundInput[84]}), .b ({new_AGEMA_signal_5212, new_AGEMA_signal_5211, RoundKey[84]}), .c ({ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1097 ( .a ({new_AGEMA_signal_5216, new_AGEMA_signal_5215, RoundInput[85]}), .b ({new_AGEMA_signal_5218, new_AGEMA_signal_5217, RoundKey[85]}), .c ({ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1098 ( .a ({new_AGEMA_signal_5222, new_AGEMA_signal_5221, RoundInput[86]}), .b ({new_AGEMA_signal_5224, new_AGEMA_signal_5223, RoundKey[86]}), .c ({ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1099 ( .a ({new_AGEMA_signal_5228, new_AGEMA_signal_5227, RoundInput[87]}), .b ({new_AGEMA_signal_5230, new_AGEMA_signal_5229, RoundKey[87]}), .c ({ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1100 ( .a ({new_AGEMA_signal_5234, new_AGEMA_signal_5233, RoundInput[88]}), .b ({new_AGEMA_signal_5236, new_AGEMA_signal_5235, RoundKey[88]}), .c ({ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1101 ( .a ({new_AGEMA_signal_5240, new_AGEMA_signal_5239, RoundInput[89]}), .b ({new_AGEMA_signal_5242, new_AGEMA_signal_5241, RoundKey[89]}), .c ({ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1102 ( .a ({new_AGEMA_signal_5246, new_AGEMA_signal_5245, RoundInput[8]}), .b ({new_AGEMA_signal_5248, new_AGEMA_signal_5247, RoundKey[8]}), .c ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1103 ( .a ({new_AGEMA_signal_5252, new_AGEMA_signal_5251, RoundInput[90]}), .b ({new_AGEMA_signal_5254, new_AGEMA_signal_5253, RoundKey[90]}), .c ({ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1104 ( .a ({new_AGEMA_signal_5258, new_AGEMA_signal_5257, RoundInput[91]}), .b ({new_AGEMA_signal_5260, new_AGEMA_signal_5259, RoundKey[91]}), .c ({ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1105 ( .a ({new_AGEMA_signal_5264, new_AGEMA_signal_5263, RoundInput[92]}), .b ({new_AGEMA_signal_5266, new_AGEMA_signal_5265, RoundKey[92]}), .c ({ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1106 ( .a ({new_AGEMA_signal_5270, new_AGEMA_signal_5269, RoundInput[93]}), .b ({new_AGEMA_signal_5272, new_AGEMA_signal_5271, RoundKey[93]}), .c ({ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1107 ( .a ({new_AGEMA_signal_5276, new_AGEMA_signal_5275, RoundInput[94]}), .b ({new_AGEMA_signal_5278, new_AGEMA_signal_5277, RoundKey[94]}), .c ({ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1108 ( .a ({new_AGEMA_signal_5282, new_AGEMA_signal_5281, RoundInput[95]}), .b ({new_AGEMA_signal_5284, new_AGEMA_signal_5283, RoundKey[95]}), .c ({ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1109 ( .a ({new_AGEMA_signal_5288, new_AGEMA_signal_5287, RoundInput[96]}), .b ({new_AGEMA_signal_5290, new_AGEMA_signal_5289, RoundKey[96]}), .c ({ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1110 ( .a ({new_AGEMA_signal_5294, new_AGEMA_signal_5293, RoundInput[97]}), .b ({new_AGEMA_signal_5296, new_AGEMA_signal_5295, RoundKey[97]}), .c ({ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1111 ( .a ({new_AGEMA_signal_5300, new_AGEMA_signal_5299, RoundInput[98]}), .b ({new_AGEMA_signal_5302, new_AGEMA_signal_5301, RoundKey[98]}), .c ({ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1112 ( .a ({new_AGEMA_signal_5306, new_AGEMA_signal_5305, RoundInput[99]}), .b ({new_AGEMA_signal_5308, new_AGEMA_signal_5307, RoundKey[99]}), .c ({ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U1113 ( .a ({new_AGEMA_signal_5312, new_AGEMA_signal_5311, RoundInput[9]}), .b ({new_AGEMA_signal_5314, new_AGEMA_signal_5313, RoundKey[9]}), .c ({ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    NAND2_X1 U1114 ( .A1 (RoundCounter[3]), .A2 (n333), .ZN (n334) ) ;
    NOR2_X1 U1115 ( .A1 (RoundCounter[0]), .A2 (n334), .ZN (done) ) ;
    INV_X1 U1116 ( .A (n335), .ZN (n336) ) ;
    NAND2_X1 U1117 ( .A1 (RoundCounter[2]), .A2 (RoundCounter[1]), .ZN (n338) ) ;
    NOR2_X1 U1118 ( .A1 (n336), .A2 (n338), .ZN (n283) ) ;
    INV_X1 U1119 ( .A (n337), .ZN (n339) ) ;
    NOR2_X1 U1120 ( .A1 (n339), .A2 (n338), .ZN (n285) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T1_U1 ( .a ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .c ({new_AGEMA_signal_5398, new_AGEMA_signal_5397, SubBytesIns_Inst_Sbox_0_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T2_U1 ( .a ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, SubBytesIns_Inst_Sbox_0_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T3_U1 ( .a ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_5402, new_AGEMA_signal_5401, SubBytesIns_Inst_Sbox_0_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T4_U1 ( .a ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_5404, new_AGEMA_signal_5403, SubBytesIns_Inst_Sbox_0_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T5_U1 ( .a ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .b ({ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_5406, new_AGEMA_signal_5405, SubBytesIns_Inst_Sbox_0_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T6_U1 ( .a ({new_AGEMA_signal_5398, new_AGEMA_signal_5397, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5406, new_AGEMA_signal_5405, SubBytesIns_Inst_Sbox_0_T5}), .c ({new_AGEMA_signal_5782, new_AGEMA_signal_5781, SubBytesIns_Inst_Sbox_0_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T7_U1 ( .a ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .c ({new_AGEMA_signal_5408, new_AGEMA_signal_5407, SubBytesIns_Inst_Sbox_0_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T8_U1 ( .a ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_5782, new_AGEMA_signal_5781, SubBytesIns_Inst_Sbox_0_T6}), .c ({new_AGEMA_signal_6142, new_AGEMA_signal_6141, SubBytesIns_Inst_Sbox_0_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T9_U1 ( .a ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_5408, new_AGEMA_signal_5407, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_5784, new_AGEMA_signal_5783, SubBytesIns_Inst_Sbox_0_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T10_U1 ( .a ({new_AGEMA_signal_5782, new_AGEMA_signal_5781, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_5408, new_AGEMA_signal_5407, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_6144, new_AGEMA_signal_6143, SubBytesIns_Inst_Sbox_0_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T11_U1 ( .a ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_5410, new_AGEMA_signal_5409, SubBytesIns_Inst_Sbox_0_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T12_U1 ( .a ({ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .b ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_5412, new_AGEMA_signal_5411, SubBytesIns_Inst_Sbox_0_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T13_U1 ( .a ({new_AGEMA_signal_5402, new_AGEMA_signal_5401, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5404, new_AGEMA_signal_5403, SubBytesIns_Inst_Sbox_0_T4}), .c ({new_AGEMA_signal_5786, new_AGEMA_signal_5785, SubBytesIns_Inst_Sbox_0_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T14_U1 ( .a ({new_AGEMA_signal_5782, new_AGEMA_signal_5781, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_5410, new_AGEMA_signal_5409, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_6146, new_AGEMA_signal_6145, SubBytesIns_Inst_Sbox_0_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T15_U1 ( .a ({new_AGEMA_signal_5406, new_AGEMA_signal_5405, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_5410, new_AGEMA_signal_5409, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_5788, new_AGEMA_signal_5787, SubBytesIns_Inst_Sbox_0_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T16_U1 ( .a ({new_AGEMA_signal_5406, new_AGEMA_signal_5405, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_5412, new_AGEMA_signal_5411, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_5790, new_AGEMA_signal_5789, SubBytesIns_Inst_Sbox_0_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T17_U1 ( .a ({new_AGEMA_signal_5784, new_AGEMA_signal_5783, SubBytesIns_Inst_Sbox_0_T9}), .b ({new_AGEMA_signal_5790, new_AGEMA_signal_5789, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_6148, new_AGEMA_signal_6147, SubBytesIns_Inst_Sbox_0_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T18_U1 ( .a ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_5414, new_AGEMA_signal_5413, SubBytesIns_Inst_Sbox_0_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T19_U1 ( .a ({new_AGEMA_signal_5408, new_AGEMA_signal_5407, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_5414, new_AGEMA_signal_5413, SubBytesIns_Inst_Sbox_0_T18}), .c ({new_AGEMA_signal_5792, new_AGEMA_signal_5791, SubBytesIns_Inst_Sbox_0_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T20_U1 ( .a ({new_AGEMA_signal_5398, new_AGEMA_signal_5397, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5792, new_AGEMA_signal_5791, SubBytesIns_Inst_Sbox_0_T19}), .c ({new_AGEMA_signal_6150, new_AGEMA_signal_6149, SubBytesIns_Inst_Sbox_0_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T21_U1 ( .a ({ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .b ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_5416, new_AGEMA_signal_5415, SubBytesIns_Inst_Sbox_0_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T22_U1 ( .a ({new_AGEMA_signal_5408, new_AGEMA_signal_5407, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_5416, new_AGEMA_signal_5415, SubBytesIns_Inst_Sbox_0_T21}), .c ({new_AGEMA_signal_5794, new_AGEMA_signal_5793, SubBytesIns_Inst_Sbox_0_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T23_U1 ( .a ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_5794, new_AGEMA_signal_5793, SubBytesIns_Inst_Sbox_0_T22}), .c ({new_AGEMA_signal_6152, new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_0_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T24_U1 ( .a ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6144, new_AGEMA_signal_6143, SubBytesIns_Inst_Sbox_0_T10}), .c ({new_AGEMA_signal_6630, new_AGEMA_signal_6629, SubBytesIns_Inst_Sbox_0_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T25_U1 ( .a ({new_AGEMA_signal_6150, new_AGEMA_signal_6149, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_6148, new_AGEMA_signal_6147, SubBytesIns_Inst_Sbox_0_T17}), .c ({new_AGEMA_signal_6632, new_AGEMA_signal_6631, SubBytesIns_Inst_Sbox_0_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T26_U1 ( .a ({new_AGEMA_signal_5402, new_AGEMA_signal_5401, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5790, new_AGEMA_signal_5789, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_6154, new_AGEMA_signal_6153, SubBytesIns_Inst_Sbox_0_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T27_U1 ( .a ({new_AGEMA_signal_5398, new_AGEMA_signal_5397, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5412, new_AGEMA_signal_5411, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_5796, new_AGEMA_signal_5795, SubBytesIns_Inst_Sbox_0_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T1_U1 ( .a ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .c ({new_AGEMA_signal_5418, new_AGEMA_signal_5417, SubBytesIns_Inst_Sbox_1_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T2_U1 ( .a ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_5420, new_AGEMA_signal_5419, SubBytesIns_Inst_Sbox_1_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T3_U1 ( .a ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .c ({new_AGEMA_signal_5422, new_AGEMA_signal_5421, SubBytesIns_Inst_Sbox_1_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T4_U1 ( .a ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_5424, new_AGEMA_signal_5423, SubBytesIns_Inst_Sbox_1_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T5_U1 ( .a ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .b ({ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .c ({new_AGEMA_signal_5426, new_AGEMA_signal_5425, SubBytesIns_Inst_Sbox_1_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T6_U1 ( .a ({new_AGEMA_signal_5418, new_AGEMA_signal_5417, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5426, new_AGEMA_signal_5425, SubBytesIns_Inst_Sbox_1_T5}), .c ({new_AGEMA_signal_5798, new_AGEMA_signal_5797, SubBytesIns_Inst_Sbox_1_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T7_U1 ( .a ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .c ({new_AGEMA_signal_5428, new_AGEMA_signal_5427, SubBytesIns_Inst_Sbox_1_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T8_U1 ( .a ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_5798, new_AGEMA_signal_5797, SubBytesIns_Inst_Sbox_1_T6}), .c ({new_AGEMA_signal_6168, new_AGEMA_signal_6167, SubBytesIns_Inst_Sbox_1_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T9_U1 ( .a ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_5428, new_AGEMA_signal_5427, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_5800, new_AGEMA_signal_5799, SubBytesIns_Inst_Sbox_1_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T10_U1 ( .a ({new_AGEMA_signal_5798, new_AGEMA_signal_5797, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_5428, new_AGEMA_signal_5427, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_6170, new_AGEMA_signal_6169, SubBytesIns_Inst_Sbox_1_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T11_U1 ( .a ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_5430, new_AGEMA_signal_5429, SubBytesIns_Inst_Sbox_1_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T12_U1 ( .a ({ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .b ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_5432, new_AGEMA_signal_5431, SubBytesIns_Inst_Sbox_1_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T13_U1 ( .a ({new_AGEMA_signal_5422, new_AGEMA_signal_5421, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5424, new_AGEMA_signal_5423, SubBytesIns_Inst_Sbox_1_T4}), .c ({new_AGEMA_signal_5802, new_AGEMA_signal_5801, SubBytesIns_Inst_Sbox_1_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T14_U1 ( .a ({new_AGEMA_signal_5798, new_AGEMA_signal_5797, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_5430, new_AGEMA_signal_5429, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_6172, new_AGEMA_signal_6171, SubBytesIns_Inst_Sbox_1_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T15_U1 ( .a ({new_AGEMA_signal_5426, new_AGEMA_signal_5425, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_5430, new_AGEMA_signal_5429, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_5804, new_AGEMA_signal_5803, SubBytesIns_Inst_Sbox_1_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T16_U1 ( .a ({new_AGEMA_signal_5426, new_AGEMA_signal_5425, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_5432, new_AGEMA_signal_5431, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_5806, new_AGEMA_signal_5805, SubBytesIns_Inst_Sbox_1_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T17_U1 ( .a ({new_AGEMA_signal_5800, new_AGEMA_signal_5799, SubBytesIns_Inst_Sbox_1_T9}), .b ({new_AGEMA_signal_5806, new_AGEMA_signal_5805, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_6174, new_AGEMA_signal_6173, SubBytesIns_Inst_Sbox_1_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T18_U1 ( .a ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .c ({new_AGEMA_signal_5434, new_AGEMA_signal_5433, SubBytesIns_Inst_Sbox_1_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T19_U1 ( .a ({new_AGEMA_signal_5428, new_AGEMA_signal_5427, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_5434, new_AGEMA_signal_5433, SubBytesIns_Inst_Sbox_1_T18}), .c ({new_AGEMA_signal_5808, new_AGEMA_signal_5807, SubBytesIns_Inst_Sbox_1_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T20_U1 ( .a ({new_AGEMA_signal_5418, new_AGEMA_signal_5417, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5808, new_AGEMA_signal_5807, SubBytesIns_Inst_Sbox_1_T19}), .c ({new_AGEMA_signal_6176, new_AGEMA_signal_6175, SubBytesIns_Inst_Sbox_1_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T21_U1 ( .a ({ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .b ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .c ({new_AGEMA_signal_5436, new_AGEMA_signal_5435, SubBytesIns_Inst_Sbox_1_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T22_U1 ( .a ({new_AGEMA_signal_5428, new_AGEMA_signal_5427, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_5436, new_AGEMA_signal_5435, SubBytesIns_Inst_Sbox_1_T21}), .c ({new_AGEMA_signal_5810, new_AGEMA_signal_5809, SubBytesIns_Inst_Sbox_1_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T23_U1 ( .a ({new_AGEMA_signal_5420, new_AGEMA_signal_5419, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_5810, new_AGEMA_signal_5809, SubBytesIns_Inst_Sbox_1_T22}), .c ({new_AGEMA_signal_6178, new_AGEMA_signal_6177, SubBytesIns_Inst_Sbox_1_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T24_U1 ( .a ({new_AGEMA_signal_5420, new_AGEMA_signal_5419, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6170, new_AGEMA_signal_6169, SubBytesIns_Inst_Sbox_1_T10}), .c ({new_AGEMA_signal_6648, new_AGEMA_signal_6647, SubBytesIns_Inst_Sbox_1_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T25_U1 ( .a ({new_AGEMA_signal_6176, new_AGEMA_signal_6175, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_6174, new_AGEMA_signal_6173, SubBytesIns_Inst_Sbox_1_T17}), .c ({new_AGEMA_signal_6650, new_AGEMA_signal_6649, SubBytesIns_Inst_Sbox_1_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T26_U1 ( .a ({new_AGEMA_signal_5422, new_AGEMA_signal_5421, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5806, new_AGEMA_signal_5805, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_6180, new_AGEMA_signal_6179, SubBytesIns_Inst_Sbox_1_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T27_U1 ( .a ({new_AGEMA_signal_5418, new_AGEMA_signal_5417, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5432, new_AGEMA_signal_5431, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_5812, new_AGEMA_signal_5811, SubBytesIns_Inst_Sbox_1_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T1_U1 ( .a ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .c ({new_AGEMA_signal_5438, new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_2_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T2_U1 ( .a ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_5440, new_AGEMA_signal_5439, SubBytesIns_Inst_Sbox_2_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T3_U1 ( .a ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_5442, new_AGEMA_signal_5441, SubBytesIns_Inst_Sbox_2_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T4_U1 ( .a ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_5444, new_AGEMA_signal_5443, SubBytesIns_Inst_Sbox_2_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T5_U1 ( .a ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .b ({ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_5446, new_AGEMA_signal_5445, SubBytesIns_Inst_Sbox_2_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T6_U1 ( .a ({new_AGEMA_signal_5438, new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5446, new_AGEMA_signal_5445, SubBytesIns_Inst_Sbox_2_T5}), .c ({new_AGEMA_signal_5814, new_AGEMA_signal_5813, SubBytesIns_Inst_Sbox_2_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T7_U1 ( .a ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .c ({new_AGEMA_signal_5448, new_AGEMA_signal_5447, SubBytesIns_Inst_Sbox_2_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T8_U1 ( .a ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_5814, new_AGEMA_signal_5813, SubBytesIns_Inst_Sbox_2_T6}), .c ({new_AGEMA_signal_6194, new_AGEMA_signal_6193, SubBytesIns_Inst_Sbox_2_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T9_U1 ( .a ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_5448, new_AGEMA_signal_5447, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_5816, new_AGEMA_signal_5815, SubBytesIns_Inst_Sbox_2_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T10_U1 ( .a ({new_AGEMA_signal_5814, new_AGEMA_signal_5813, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_5448, new_AGEMA_signal_5447, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_6196, new_AGEMA_signal_6195, SubBytesIns_Inst_Sbox_2_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T11_U1 ( .a ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_5450, new_AGEMA_signal_5449, SubBytesIns_Inst_Sbox_2_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T12_U1 ( .a ({ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .b ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_5452, new_AGEMA_signal_5451, SubBytesIns_Inst_Sbox_2_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T13_U1 ( .a ({new_AGEMA_signal_5442, new_AGEMA_signal_5441, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5444, new_AGEMA_signal_5443, SubBytesIns_Inst_Sbox_2_T4}), .c ({new_AGEMA_signal_5818, new_AGEMA_signal_5817, SubBytesIns_Inst_Sbox_2_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T14_U1 ( .a ({new_AGEMA_signal_5814, new_AGEMA_signal_5813, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_5450, new_AGEMA_signal_5449, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_6198, new_AGEMA_signal_6197, SubBytesIns_Inst_Sbox_2_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T15_U1 ( .a ({new_AGEMA_signal_5446, new_AGEMA_signal_5445, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_5450, new_AGEMA_signal_5449, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_5820, new_AGEMA_signal_5819, SubBytesIns_Inst_Sbox_2_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T16_U1 ( .a ({new_AGEMA_signal_5446, new_AGEMA_signal_5445, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_5452, new_AGEMA_signal_5451, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_2_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T17_U1 ( .a ({new_AGEMA_signal_5816, new_AGEMA_signal_5815, SubBytesIns_Inst_Sbox_2_T9}), .b ({new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_6200, new_AGEMA_signal_6199, SubBytesIns_Inst_Sbox_2_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T18_U1 ( .a ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_5454, new_AGEMA_signal_5453, SubBytesIns_Inst_Sbox_2_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T19_U1 ( .a ({new_AGEMA_signal_5448, new_AGEMA_signal_5447, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5454, new_AGEMA_signal_5453, SubBytesIns_Inst_Sbox_2_T18}), .c ({new_AGEMA_signal_5824, new_AGEMA_signal_5823, SubBytesIns_Inst_Sbox_2_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T20_U1 ( .a ({new_AGEMA_signal_5438, new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5824, new_AGEMA_signal_5823, SubBytesIns_Inst_Sbox_2_T19}), .c ({new_AGEMA_signal_6202, new_AGEMA_signal_6201, SubBytesIns_Inst_Sbox_2_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T21_U1 ( .a ({ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .b ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_5456, new_AGEMA_signal_5455, SubBytesIns_Inst_Sbox_2_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T22_U1 ( .a ({new_AGEMA_signal_5448, new_AGEMA_signal_5447, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5456, new_AGEMA_signal_5455, SubBytesIns_Inst_Sbox_2_T21}), .c ({new_AGEMA_signal_5826, new_AGEMA_signal_5825, SubBytesIns_Inst_Sbox_2_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T23_U1 ( .a ({new_AGEMA_signal_5440, new_AGEMA_signal_5439, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_5826, new_AGEMA_signal_5825, SubBytesIns_Inst_Sbox_2_T22}), .c ({new_AGEMA_signal_6204, new_AGEMA_signal_6203, SubBytesIns_Inst_Sbox_2_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T24_U1 ( .a ({new_AGEMA_signal_5440, new_AGEMA_signal_5439, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_6196, new_AGEMA_signal_6195, SubBytesIns_Inst_Sbox_2_T10}), .c ({new_AGEMA_signal_6666, new_AGEMA_signal_6665, SubBytesIns_Inst_Sbox_2_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T25_U1 ( .a ({new_AGEMA_signal_6202, new_AGEMA_signal_6201, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_6200, new_AGEMA_signal_6199, SubBytesIns_Inst_Sbox_2_T17}), .c ({new_AGEMA_signal_6668, new_AGEMA_signal_6667, SubBytesIns_Inst_Sbox_2_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T26_U1 ( .a ({new_AGEMA_signal_5442, new_AGEMA_signal_5441, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_6206, new_AGEMA_signal_6205, SubBytesIns_Inst_Sbox_2_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T27_U1 ( .a ({new_AGEMA_signal_5438, new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5452, new_AGEMA_signal_5451, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_5828, new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_2_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T1_U1 ( .a ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_5458, new_AGEMA_signal_5457, SubBytesIns_Inst_Sbox_3_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T2_U1 ( .a ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5460, new_AGEMA_signal_5459, SubBytesIns_Inst_Sbox_3_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T3_U1 ( .a ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_5462, new_AGEMA_signal_5461, SubBytesIns_Inst_Sbox_3_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T4_U1 ( .a ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5464, new_AGEMA_signal_5463, SubBytesIns_Inst_Sbox_3_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T5_U1 ( .a ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .b ({ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_5466, new_AGEMA_signal_5465, SubBytesIns_Inst_Sbox_3_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T6_U1 ( .a ({new_AGEMA_signal_5458, new_AGEMA_signal_5457, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5466, new_AGEMA_signal_5465, SubBytesIns_Inst_Sbox_3_T5}), .c ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, SubBytesIns_Inst_Sbox_3_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T7_U1 ( .a ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_5468, new_AGEMA_signal_5467, SubBytesIns_Inst_Sbox_3_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T8_U1 ( .a ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, SubBytesIns_Inst_Sbox_3_T6}), .c ({new_AGEMA_signal_6220, new_AGEMA_signal_6219, SubBytesIns_Inst_Sbox_3_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T9_U1 ( .a ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_5468, new_AGEMA_signal_5467, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_5832, new_AGEMA_signal_5831, SubBytesIns_Inst_Sbox_3_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T10_U1 ( .a ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5468, new_AGEMA_signal_5467, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_6222, new_AGEMA_signal_6221, SubBytesIns_Inst_Sbox_3_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T11_U1 ( .a ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5470, new_AGEMA_signal_5469, SubBytesIns_Inst_Sbox_3_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T12_U1 ( .a ({ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5472, new_AGEMA_signal_5471, SubBytesIns_Inst_Sbox_3_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T13_U1 ( .a ({new_AGEMA_signal_5462, new_AGEMA_signal_5461, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5464, new_AGEMA_signal_5463, SubBytesIns_Inst_Sbox_3_T4}), .c ({new_AGEMA_signal_5834, new_AGEMA_signal_5833, SubBytesIns_Inst_Sbox_3_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T14_U1 ( .a ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5470, new_AGEMA_signal_5469, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_6224, new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_3_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T15_U1 ( .a ({new_AGEMA_signal_5466, new_AGEMA_signal_5465, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5470, new_AGEMA_signal_5469, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_5836, new_AGEMA_signal_5835, SubBytesIns_Inst_Sbox_3_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T16_U1 ( .a ({new_AGEMA_signal_5466, new_AGEMA_signal_5465, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5472, new_AGEMA_signal_5471, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, SubBytesIns_Inst_Sbox_3_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T17_U1 ( .a ({new_AGEMA_signal_5832, new_AGEMA_signal_5831, SubBytesIns_Inst_Sbox_3_T9}), .b ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_6226, new_AGEMA_signal_6225, SubBytesIns_Inst_Sbox_3_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T18_U1 ( .a ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_5474, new_AGEMA_signal_5473, SubBytesIns_Inst_Sbox_3_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T19_U1 ( .a ({new_AGEMA_signal_5468, new_AGEMA_signal_5467, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5474, new_AGEMA_signal_5473, SubBytesIns_Inst_Sbox_3_T18}), .c ({new_AGEMA_signal_5840, new_AGEMA_signal_5839, SubBytesIns_Inst_Sbox_3_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T20_U1 ( .a ({new_AGEMA_signal_5458, new_AGEMA_signal_5457, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5840, new_AGEMA_signal_5839, SubBytesIns_Inst_Sbox_3_T19}), .c ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, SubBytesIns_Inst_Sbox_3_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T21_U1 ( .a ({ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .b ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_5476, new_AGEMA_signal_5475, SubBytesIns_Inst_Sbox_3_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T22_U1 ( .a ({new_AGEMA_signal_5468, new_AGEMA_signal_5467, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5476, new_AGEMA_signal_5475, SubBytesIns_Inst_Sbox_3_T21}), .c ({new_AGEMA_signal_5842, new_AGEMA_signal_5841, SubBytesIns_Inst_Sbox_3_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T23_U1 ( .a ({new_AGEMA_signal_5460, new_AGEMA_signal_5459, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_5842, new_AGEMA_signal_5841, SubBytesIns_Inst_Sbox_3_T22}), .c ({new_AGEMA_signal_6230, new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_3_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T24_U1 ( .a ({new_AGEMA_signal_5460, new_AGEMA_signal_5459, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_6222, new_AGEMA_signal_6221, SubBytesIns_Inst_Sbox_3_T10}), .c ({new_AGEMA_signal_6684, new_AGEMA_signal_6683, SubBytesIns_Inst_Sbox_3_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T25_U1 ( .a ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_6226, new_AGEMA_signal_6225, SubBytesIns_Inst_Sbox_3_T17}), .c ({new_AGEMA_signal_6686, new_AGEMA_signal_6685, SubBytesIns_Inst_Sbox_3_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T26_U1 ( .a ({new_AGEMA_signal_5462, new_AGEMA_signal_5461, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_6232, new_AGEMA_signal_6231, SubBytesIns_Inst_Sbox_3_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T27_U1 ( .a ({new_AGEMA_signal_5458, new_AGEMA_signal_5457, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5472, new_AGEMA_signal_5471, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_5844, new_AGEMA_signal_5843, SubBytesIns_Inst_Sbox_3_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T1_U1 ( .a ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .c ({new_AGEMA_signal_5478, new_AGEMA_signal_5477, SubBytesIns_Inst_Sbox_4_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T2_U1 ( .a ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5480, new_AGEMA_signal_5479, SubBytesIns_Inst_Sbox_4_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T3_U1 ( .a ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_5482, new_AGEMA_signal_5481, SubBytesIns_Inst_Sbox_4_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T4_U1 ( .a ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5484, new_AGEMA_signal_5483, SubBytesIns_Inst_Sbox_4_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T5_U1 ( .a ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .b ({ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_5486, new_AGEMA_signal_5485, SubBytesIns_Inst_Sbox_4_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T6_U1 ( .a ({new_AGEMA_signal_5478, new_AGEMA_signal_5477, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5486, new_AGEMA_signal_5485, SubBytesIns_Inst_Sbox_4_T5}), .c ({new_AGEMA_signal_5846, new_AGEMA_signal_5845, SubBytesIns_Inst_Sbox_4_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T7_U1 ( .a ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .c ({new_AGEMA_signal_5488, new_AGEMA_signal_5487, SubBytesIns_Inst_Sbox_4_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T8_U1 ( .a ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_5846, new_AGEMA_signal_5845, SubBytesIns_Inst_Sbox_4_T6}), .c ({new_AGEMA_signal_6246, new_AGEMA_signal_6245, SubBytesIns_Inst_Sbox_4_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T9_U1 ( .a ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_5488, new_AGEMA_signal_5487, SubBytesIns_Inst_Sbox_4_T7}), .c ({new_AGEMA_signal_5848, new_AGEMA_signal_5847, SubBytesIns_Inst_Sbox_4_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T10_U1 ( .a ({new_AGEMA_signal_5846, new_AGEMA_signal_5845, SubBytesIns_Inst_Sbox_4_T6}), .b ({new_AGEMA_signal_5488, new_AGEMA_signal_5487, SubBytesIns_Inst_Sbox_4_T7}), .c ({new_AGEMA_signal_6248, new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_4_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T11_U1 ( .a ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5490, new_AGEMA_signal_5489, SubBytesIns_Inst_Sbox_4_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T12_U1 ( .a ({ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .b ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5492, new_AGEMA_signal_5491, SubBytesIns_Inst_Sbox_4_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T13_U1 ( .a ({new_AGEMA_signal_5482, new_AGEMA_signal_5481, SubBytesIns_Inst_Sbox_4_T3}), .b ({new_AGEMA_signal_5484, new_AGEMA_signal_5483, SubBytesIns_Inst_Sbox_4_T4}), .c ({new_AGEMA_signal_5850, new_AGEMA_signal_5849, SubBytesIns_Inst_Sbox_4_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T14_U1 ( .a ({new_AGEMA_signal_5846, new_AGEMA_signal_5845, SubBytesIns_Inst_Sbox_4_T6}), .b ({new_AGEMA_signal_5490, new_AGEMA_signal_5489, SubBytesIns_Inst_Sbox_4_T11}), .c ({new_AGEMA_signal_6250, new_AGEMA_signal_6249, SubBytesIns_Inst_Sbox_4_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T15_U1 ( .a ({new_AGEMA_signal_5486, new_AGEMA_signal_5485, SubBytesIns_Inst_Sbox_4_T5}), .b ({new_AGEMA_signal_5490, new_AGEMA_signal_5489, SubBytesIns_Inst_Sbox_4_T11}), .c ({new_AGEMA_signal_5852, new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_4_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T16_U1 ( .a ({new_AGEMA_signal_5486, new_AGEMA_signal_5485, SubBytesIns_Inst_Sbox_4_T5}), .b ({new_AGEMA_signal_5492, new_AGEMA_signal_5491, SubBytesIns_Inst_Sbox_4_T12}), .c ({new_AGEMA_signal_5854, new_AGEMA_signal_5853, SubBytesIns_Inst_Sbox_4_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T17_U1 ( .a ({new_AGEMA_signal_5848, new_AGEMA_signal_5847, SubBytesIns_Inst_Sbox_4_T9}), .b ({new_AGEMA_signal_5854, new_AGEMA_signal_5853, SubBytesIns_Inst_Sbox_4_T16}), .c ({new_AGEMA_signal_6252, new_AGEMA_signal_6251, SubBytesIns_Inst_Sbox_4_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T18_U1 ( .a ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_5494, new_AGEMA_signal_5493, SubBytesIns_Inst_Sbox_4_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T19_U1 ( .a ({new_AGEMA_signal_5488, new_AGEMA_signal_5487, SubBytesIns_Inst_Sbox_4_T7}), .b ({new_AGEMA_signal_5494, new_AGEMA_signal_5493, SubBytesIns_Inst_Sbox_4_T18}), .c ({new_AGEMA_signal_5856, new_AGEMA_signal_5855, SubBytesIns_Inst_Sbox_4_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T20_U1 ( .a ({new_AGEMA_signal_5478, new_AGEMA_signal_5477, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5856, new_AGEMA_signal_5855, SubBytesIns_Inst_Sbox_4_T19}), .c ({new_AGEMA_signal_6254, new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_4_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T21_U1 ( .a ({ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .b ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_5496, new_AGEMA_signal_5495, SubBytesIns_Inst_Sbox_4_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T22_U1 ( .a ({new_AGEMA_signal_5488, new_AGEMA_signal_5487, SubBytesIns_Inst_Sbox_4_T7}), .b ({new_AGEMA_signal_5496, new_AGEMA_signal_5495, SubBytesIns_Inst_Sbox_4_T21}), .c ({new_AGEMA_signal_5858, new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_4_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T23_U1 ( .a ({new_AGEMA_signal_5480, new_AGEMA_signal_5479, SubBytesIns_Inst_Sbox_4_T2}), .b ({new_AGEMA_signal_5858, new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_4_T22}), .c ({new_AGEMA_signal_6256, new_AGEMA_signal_6255, SubBytesIns_Inst_Sbox_4_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T24_U1 ( .a ({new_AGEMA_signal_5480, new_AGEMA_signal_5479, SubBytesIns_Inst_Sbox_4_T2}), .b ({new_AGEMA_signal_6248, new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_4_T10}), .c ({new_AGEMA_signal_6702, new_AGEMA_signal_6701, SubBytesIns_Inst_Sbox_4_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T25_U1 ( .a ({new_AGEMA_signal_6254, new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_4_T20}), .b ({new_AGEMA_signal_6252, new_AGEMA_signal_6251, SubBytesIns_Inst_Sbox_4_T17}), .c ({new_AGEMA_signal_6704, new_AGEMA_signal_6703, SubBytesIns_Inst_Sbox_4_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T26_U1 ( .a ({new_AGEMA_signal_5482, new_AGEMA_signal_5481, SubBytesIns_Inst_Sbox_4_T3}), .b ({new_AGEMA_signal_5854, new_AGEMA_signal_5853, SubBytesIns_Inst_Sbox_4_T16}), .c ({new_AGEMA_signal_6258, new_AGEMA_signal_6257, SubBytesIns_Inst_Sbox_4_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T27_U1 ( .a ({new_AGEMA_signal_5478, new_AGEMA_signal_5477, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5492, new_AGEMA_signal_5491, SubBytesIns_Inst_Sbox_4_T12}), .c ({new_AGEMA_signal_5860, new_AGEMA_signal_5859, SubBytesIns_Inst_Sbox_4_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T1_U1 ( .a ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .c ({new_AGEMA_signal_5498, new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_5_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T2_U1 ( .a ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5500, new_AGEMA_signal_5499, SubBytesIns_Inst_Sbox_5_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T3_U1 ( .a ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_5502, new_AGEMA_signal_5501, SubBytesIns_Inst_Sbox_5_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T4_U1 ( .a ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5504, new_AGEMA_signal_5503, SubBytesIns_Inst_Sbox_5_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T5_U1 ( .a ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .b ({ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_5506, new_AGEMA_signal_5505, SubBytesIns_Inst_Sbox_5_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T6_U1 ( .a ({new_AGEMA_signal_5498, new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5506, new_AGEMA_signal_5505, SubBytesIns_Inst_Sbox_5_T5}), .c ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, SubBytesIns_Inst_Sbox_5_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T7_U1 ( .a ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .c ({new_AGEMA_signal_5508, new_AGEMA_signal_5507, SubBytesIns_Inst_Sbox_5_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T8_U1 ( .a ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, SubBytesIns_Inst_Sbox_5_T6}), .c ({new_AGEMA_signal_6272, new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_5_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T9_U1 ( .a ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_5508, new_AGEMA_signal_5507, SubBytesIns_Inst_Sbox_5_T7}), .c ({new_AGEMA_signal_5864, new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_5_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T10_U1 ( .a ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, SubBytesIns_Inst_Sbox_5_T6}), .b ({new_AGEMA_signal_5508, new_AGEMA_signal_5507, SubBytesIns_Inst_Sbox_5_T7}), .c ({new_AGEMA_signal_6274, new_AGEMA_signal_6273, SubBytesIns_Inst_Sbox_5_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T11_U1 ( .a ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5510, new_AGEMA_signal_5509, SubBytesIns_Inst_Sbox_5_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T12_U1 ( .a ({ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .b ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5512, new_AGEMA_signal_5511, SubBytesIns_Inst_Sbox_5_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T13_U1 ( .a ({new_AGEMA_signal_5502, new_AGEMA_signal_5501, SubBytesIns_Inst_Sbox_5_T3}), .b ({new_AGEMA_signal_5504, new_AGEMA_signal_5503, SubBytesIns_Inst_Sbox_5_T4}), .c ({new_AGEMA_signal_5866, new_AGEMA_signal_5865, SubBytesIns_Inst_Sbox_5_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T14_U1 ( .a ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, SubBytesIns_Inst_Sbox_5_T6}), .b ({new_AGEMA_signal_5510, new_AGEMA_signal_5509, SubBytesIns_Inst_Sbox_5_T11}), .c ({new_AGEMA_signal_6276, new_AGEMA_signal_6275, SubBytesIns_Inst_Sbox_5_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T15_U1 ( .a ({new_AGEMA_signal_5506, new_AGEMA_signal_5505, SubBytesIns_Inst_Sbox_5_T5}), .b ({new_AGEMA_signal_5510, new_AGEMA_signal_5509, SubBytesIns_Inst_Sbox_5_T11}), .c ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, SubBytesIns_Inst_Sbox_5_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T16_U1 ( .a ({new_AGEMA_signal_5506, new_AGEMA_signal_5505, SubBytesIns_Inst_Sbox_5_T5}), .b ({new_AGEMA_signal_5512, new_AGEMA_signal_5511, SubBytesIns_Inst_Sbox_5_T12}), .c ({new_AGEMA_signal_5870, new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_5_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T17_U1 ( .a ({new_AGEMA_signal_5864, new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_5_T9}), .b ({new_AGEMA_signal_5870, new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_5_T16}), .c ({new_AGEMA_signal_6278, new_AGEMA_signal_6277, SubBytesIns_Inst_Sbox_5_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T18_U1 ( .a ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_5514, new_AGEMA_signal_5513, SubBytesIns_Inst_Sbox_5_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T19_U1 ( .a ({new_AGEMA_signal_5508, new_AGEMA_signal_5507, SubBytesIns_Inst_Sbox_5_T7}), .b ({new_AGEMA_signal_5514, new_AGEMA_signal_5513, SubBytesIns_Inst_Sbox_5_T18}), .c ({new_AGEMA_signal_5872, new_AGEMA_signal_5871, SubBytesIns_Inst_Sbox_5_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T20_U1 ( .a ({new_AGEMA_signal_5498, new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5872, new_AGEMA_signal_5871, SubBytesIns_Inst_Sbox_5_T19}), .c ({new_AGEMA_signal_6280, new_AGEMA_signal_6279, SubBytesIns_Inst_Sbox_5_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T21_U1 ( .a ({ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .b ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_5516, new_AGEMA_signal_5515, SubBytesIns_Inst_Sbox_5_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T22_U1 ( .a ({new_AGEMA_signal_5508, new_AGEMA_signal_5507, SubBytesIns_Inst_Sbox_5_T7}), .b ({new_AGEMA_signal_5516, new_AGEMA_signal_5515, SubBytesIns_Inst_Sbox_5_T21}), .c ({new_AGEMA_signal_5874, new_AGEMA_signal_5873, SubBytesIns_Inst_Sbox_5_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T23_U1 ( .a ({new_AGEMA_signal_5500, new_AGEMA_signal_5499, SubBytesIns_Inst_Sbox_5_T2}), .b ({new_AGEMA_signal_5874, new_AGEMA_signal_5873, SubBytesIns_Inst_Sbox_5_T22}), .c ({new_AGEMA_signal_6282, new_AGEMA_signal_6281, SubBytesIns_Inst_Sbox_5_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T24_U1 ( .a ({new_AGEMA_signal_5500, new_AGEMA_signal_5499, SubBytesIns_Inst_Sbox_5_T2}), .b ({new_AGEMA_signal_6274, new_AGEMA_signal_6273, SubBytesIns_Inst_Sbox_5_T10}), .c ({new_AGEMA_signal_6720, new_AGEMA_signal_6719, SubBytesIns_Inst_Sbox_5_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T25_U1 ( .a ({new_AGEMA_signal_6280, new_AGEMA_signal_6279, SubBytesIns_Inst_Sbox_5_T20}), .b ({new_AGEMA_signal_6278, new_AGEMA_signal_6277, SubBytesIns_Inst_Sbox_5_T17}), .c ({new_AGEMA_signal_6722, new_AGEMA_signal_6721, SubBytesIns_Inst_Sbox_5_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T26_U1 ( .a ({new_AGEMA_signal_5502, new_AGEMA_signal_5501, SubBytesIns_Inst_Sbox_5_T3}), .b ({new_AGEMA_signal_5870, new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_5_T16}), .c ({new_AGEMA_signal_6284, new_AGEMA_signal_6283, SubBytesIns_Inst_Sbox_5_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T27_U1 ( .a ({new_AGEMA_signal_5498, new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5512, new_AGEMA_signal_5511, SubBytesIns_Inst_Sbox_5_T12}), .c ({new_AGEMA_signal_5876, new_AGEMA_signal_5875, SubBytesIns_Inst_Sbox_5_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T1_U1 ( .a ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .c ({new_AGEMA_signal_5518, new_AGEMA_signal_5517, SubBytesIns_Inst_Sbox_6_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T2_U1 ( .a ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_5520, new_AGEMA_signal_5519, SubBytesIns_Inst_Sbox_6_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T3_U1 ( .a ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_5522, new_AGEMA_signal_5521, SubBytesIns_Inst_Sbox_6_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T4_U1 ( .a ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_5524, new_AGEMA_signal_5523, SubBytesIns_Inst_Sbox_6_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T5_U1 ( .a ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .b ({ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_5526, new_AGEMA_signal_5525, SubBytesIns_Inst_Sbox_6_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T6_U1 ( .a ({new_AGEMA_signal_5518, new_AGEMA_signal_5517, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_5526, new_AGEMA_signal_5525, SubBytesIns_Inst_Sbox_6_T5}), .c ({new_AGEMA_signal_5878, new_AGEMA_signal_5877, SubBytesIns_Inst_Sbox_6_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T7_U1 ( .a ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .c ({new_AGEMA_signal_5528, new_AGEMA_signal_5527, SubBytesIns_Inst_Sbox_6_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T8_U1 ( .a ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_5878, new_AGEMA_signal_5877, SubBytesIns_Inst_Sbox_6_T6}), .c ({new_AGEMA_signal_6298, new_AGEMA_signal_6297, SubBytesIns_Inst_Sbox_6_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T9_U1 ( .a ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_5528, new_AGEMA_signal_5527, SubBytesIns_Inst_Sbox_6_T7}), .c ({new_AGEMA_signal_5880, new_AGEMA_signal_5879, SubBytesIns_Inst_Sbox_6_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T10_U1 ( .a ({new_AGEMA_signal_5878, new_AGEMA_signal_5877, SubBytesIns_Inst_Sbox_6_T6}), .b ({new_AGEMA_signal_5528, new_AGEMA_signal_5527, SubBytesIns_Inst_Sbox_6_T7}), .c ({new_AGEMA_signal_6300, new_AGEMA_signal_6299, SubBytesIns_Inst_Sbox_6_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T11_U1 ( .a ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_5530, new_AGEMA_signal_5529, SubBytesIns_Inst_Sbox_6_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T12_U1 ( .a ({ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .b ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_5532, new_AGEMA_signal_5531, SubBytesIns_Inst_Sbox_6_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T13_U1 ( .a ({new_AGEMA_signal_5522, new_AGEMA_signal_5521, SubBytesIns_Inst_Sbox_6_T3}), .b ({new_AGEMA_signal_5524, new_AGEMA_signal_5523, SubBytesIns_Inst_Sbox_6_T4}), .c ({new_AGEMA_signal_5882, new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_6_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T14_U1 ( .a ({new_AGEMA_signal_5878, new_AGEMA_signal_5877, SubBytesIns_Inst_Sbox_6_T6}), .b ({new_AGEMA_signal_5530, new_AGEMA_signal_5529, SubBytesIns_Inst_Sbox_6_T11}), .c ({new_AGEMA_signal_6302, new_AGEMA_signal_6301, SubBytesIns_Inst_Sbox_6_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T15_U1 ( .a ({new_AGEMA_signal_5526, new_AGEMA_signal_5525, SubBytesIns_Inst_Sbox_6_T5}), .b ({new_AGEMA_signal_5530, new_AGEMA_signal_5529, SubBytesIns_Inst_Sbox_6_T11}), .c ({new_AGEMA_signal_5884, new_AGEMA_signal_5883, SubBytesIns_Inst_Sbox_6_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T16_U1 ( .a ({new_AGEMA_signal_5526, new_AGEMA_signal_5525, SubBytesIns_Inst_Sbox_6_T5}), .b ({new_AGEMA_signal_5532, new_AGEMA_signal_5531, SubBytesIns_Inst_Sbox_6_T12}), .c ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, SubBytesIns_Inst_Sbox_6_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T17_U1 ( .a ({new_AGEMA_signal_5880, new_AGEMA_signal_5879, SubBytesIns_Inst_Sbox_6_T9}), .b ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, SubBytesIns_Inst_Sbox_6_T16}), .c ({new_AGEMA_signal_6304, new_AGEMA_signal_6303, SubBytesIns_Inst_Sbox_6_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T18_U1 ( .a ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_5534, new_AGEMA_signal_5533, SubBytesIns_Inst_Sbox_6_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T19_U1 ( .a ({new_AGEMA_signal_5528, new_AGEMA_signal_5527, SubBytesIns_Inst_Sbox_6_T7}), .b ({new_AGEMA_signal_5534, new_AGEMA_signal_5533, SubBytesIns_Inst_Sbox_6_T18}), .c ({new_AGEMA_signal_5888, new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_6_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T20_U1 ( .a ({new_AGEMA_signal_5518, new_AGEMA_signal_5517, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_5888, new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_6_T19}), .c ({new_AGEMA_signal_6306, new_AGEMA_signal_6305, SubBytesIns_Inst_Sbox_6_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T21_U1 ( .a ({ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .b ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_5536, new_AGEMA_signal_5535, SubBytesIns_Inst_Sbox_6_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T22_U1 ( .a ({new_AGEMA_signal_5528, new_AGEMA_signal_5527, SubBytesIns_Inst_Sbox_6_T7}), .b ({new_AGEMA_signal_5536, new_AGEMA_signal_5535, SubBytesIns_Inst_Sbox_6_T21}), .c ({new_AGEMA_signal_5890, new_AGEMA_signal_5889, SubBytesIns_Inst_Sbox_6_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T23_U1 ( .a ({new_AGEMA_signal_5520, new_AGEMA_signal_5519, SubBytesIns_Inst_Sbox_6_T2}), .b ({new_AGEMA_signal_5890, new_AGEMA_signal_5889, SubBytesIns_Inst_Sbox_6_T22}), .c ({new_AGEMA_signal_6308, new_AGEMA_signal_6307, SubBytesIns_Inst_Sbox_6_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T24_U1 ( .a ({new_AGEMA_signal_5520, new_AGEMA_signal_5519, SubBytesIns_Inst_Sbox_6_T2}), .b ({new_AGEMA_signal_6300, new_AGEMA_signal_6299, SubBytesIns_Inst_Sbox_6_T10}), .c ({new_AGEMA_signal_6738, new_AGEMA_signal_6737, SubBytesIns_Inst_Sbox_6_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T25_U1 ( .a ({new_AGEMA_signal_6306, new_AGEMA_signal_6305, SubBytesIns_Inst_Sbox_6_T20}), .b ({new_AGEMA_signal_6304, new_AGEMA_signal_6303, SubBytesIns_Inst_Sbox_6_T17}), .c ({new_AGEMA_signal_6740, new_AGEMA_signal_6739, SubBytesIns_Inst_Sbox_6_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T26_U1 ( .a ({new_AGEMA_signal_5522, new_AGEMA_signal_5521, SubBytesIns_Inst_Sbox_6_T3}), .b ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, SubBytesIns_Inst_Sbox_6_T16}), .c ({new_AGEMA_signal_6310, new_AGEMA_signal_6309, SubBytesIns_Inst_Sbox_6_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T27_U1 ( .a ({new_AGEMA_signal_5518, new_AGEMA_signal_5517, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_5532, new_AGEMA_signal_5531, SubBytesIns_Inst_Sbox_6_T12}), .c ({new_AGEMA_signal_5892, new_AGEMA_signal_5891, SubBytesIns_Inst_Sbox_6_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T1_U1 ( .a ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_5538, new_AGEMA_signal_5537, SubBytesIns_Inst_Sbox_7_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T2_U1 ( .a ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_5540, new_AGEMA_signal_5539, SubBytesIns_Inst_Sbox_7_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T3_U1 ( .a ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_5542, new_AGEMA_signal_5541, SubBytesIns_Inst_Sbox_7_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T4_U1 ( .a ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_5544, new_AGEMA_signal_5543, SubBytesIns_Inst_Sbox_7_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T5_U1 ( .a ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .b ({ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_5546, new_AGEMA_signal_5545, SubBytesIns_Inst_Sbox_7_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T6_U1 ( .a ({new_AGEMA_signal_5538, new_AGEMA_signal_5537, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_5546, new_AGEMA_signal_5545, SubBytesIns_Inst_Sbox_7_T5}), .c ({new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_7_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T7_U1 ( .a ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_5548, new_AGEMA_signal_5547, SubBytesIns_Inst_Sbox_7_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T8_U1 ( .a ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_7_T6}), .c ({new_AGEMA_signal_6324, new_AGEMA_signal_6323, SubBytesIns_Inst_Sbox_7_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T9_U1 ( .a ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_5548, new_AGEMA_signal_5547, SubBytesIns_Inst_Sbox_7_T7}), .c ({new_AGEMA_signal_5896, new_AGEMA_signal_5895, SubBytesIns_Inst_Sbox_7_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T10_U1 ( .a ({new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_7_T6}), .b ({new_AGEMA_signal_5548, new_AGEMA_signal_5547, SubBytesIns_Inst_Sbox_7_T7}), .c ({new_AGEMA_signal_6326, new_AGEMA_signal_6325, SubBytesIns_Inst_Sbox_7_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T11_U1 ( .a ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_5550, new_AGEMA_signal_5549, SubBytesIns_Inst_Sbox_7_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T12_U1 ( .a ({ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_5552, new_AGEMA_signal_5551, SubBytesIns_Inst_Sbox_7_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T13_U1 ( .a ({new_AGEMA_signal_5542, new_AGEMA_signal_5541, SubBytesIns_Inst_Sbox_7_T3}), .b ({new_AGEMA_signal_5544, new_AGEMA_signal_5543, SubBytesIns_Inst_Sbox_7_T4}), .c ({new_AGEMA_signal_5898, new_AGEMA_signal_5897, SubBytesIns_Inst_Sbox_7_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T14_U1 ( .a ({new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_7_T6}), .b ({new_AGEMA_signal_5550, new_AGEMA_signal_5549, SubBytesIns_Inst_Sbox_7_T11}), .c ({new_AGEMA_signal_6328, new_AGEMA_signal_6327, SubBytesIns_Inst_Sbox_7_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T15_U1 ( .a ({new_AGEMA_signal_5546, new_AGEMA_signal_5545, SubBytesIns_Inst_Sbox_7_T5}), .b ({new_AGEMA_signal_5550, new_AGEMA_signal_5549, SubBytesIns_Inst_Sbox_7_T11}), .c ({new_AGEMA_signal_5900, new_AGEMA_signal_5899, SubBytesIns_Inst_Sbox_7_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T16_U1 ( .a ({new_AGEMA_signal_5546, new_AGEMA_signal_5545, SubBytesIns_Inst_Sbox_7_T5}), .b ({new_AGEMA_signal_5552, new_AGEMA_signal_5551, SubBytesIns_Inst_Sbox_7_T12}), .c ({new_AGEMA_signal_5902, new_AGEMA_signal_5901, SubBytesIns_Inst_Sbox_7_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T17_U1 ( .a ({new_AGEMA_signal_5896, new_AGEMA_signal_5895, SubBytesIns_Inst_Sbox_7_T9}), .b ({new_AGEMA_signal_5902, new_AGEMA_signal_5901, SubBytesIns_Inst_Sbox_7_T16}), .c ({new_AGEMA_signal_6330, new_AGEMA_signal_6329, SubBytesIns_Inst_Sbox_7_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T18_U1 ( .a ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_5554, new_AGEMA_signal_5553, SubBytesIns_Inst_Sbox_7_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T19_U1 ( .a ({new_AGEMA_signal_5548, new_AGEMA_signal_5547, SubBytesIns_Inst_Sbox_7_T7}), .b ({new_AGEMA_signal_5554, new_AGEMA_signal_5553, SubBytesIns_Inst_Sbox_7_T18}), .c ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, SubBytesIns_Inst_Sbox_7_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T20_U1 ( .a ({new_AGEMA_signal_5538, new_AGEMA_signal_5537, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, SubBytesIns_Inst_Sbox_7_T19}), .c ({new_AGEMA_signal_6332, new_AGEMA_signal_6331, SubBytesIns_Inst_Sbox_7_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T21_U1 ( .a ({ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .b ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_5556, new_AGEMA_signal_5555, SubBytesIns_Inst_Sbox_7_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T22_U1 ( .a ({new_AGEMA_signal_5548, new_AGEMA_signal_5547, SubBytesIns_Inst_Sbox_7_T7}), .b ({new_AGEMA_signal_5556, new_AGEMA_signal_5555, SubBytesIns_Inst_Sbox_7_T21}), .c ({new_AGEMA_signal_5906, new_AGEMA_signal_5905, SubBytesIns_Inst_Sbox_7_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T23_U1 ( .a ({new_AGEMA_signal_5540, new_AGEMA_signal_5539, SubBytesIns_Inst_Sbox_7_T2}), .b ({new_AGEMA_signal_5906, new_AGEMA_signal_5905, SubBytesIns_Inst_Sbox_7_T22}), .c ({new_AGEMA_signal_6334, new_AGEMA_signal_6333, SubBytesIns_Inst_Sbox_7_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T24_U1 ( .a ({new_AGEMA_signal_5540, new_AGEMA_signal_5539, SubBytesIns_Inst_Sbox_7_T2}), .b ({new_AGEMA_signal_6326, new_AGEMA_signal_6325, SubBytesIns_Inst_Sbox_7_T10}), .c ({new_AGEMA_signal_6756, new_AGEMA_signal_6755, SubBytesIns_Inst_Sbox_7_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T25_U1 ( .a ({new_AGEMA_signal_6332, new_AGEMA_signal_6331, SubBytesIns_Inst_Sbox_7_T20}), .b ({new_AGEMA_signal_6330, new_AGEMA_signal_6329, SubBytesIns_Inst_Sbox_7_T17}), .c ({new_AGEMA_signal_6758, new_AGEMA_signal_6757, SubBytesIns_Inst_Sbox_7_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T26_U1 ( .a ({new_AGEMA_signal_5542, new_AGEMA_signal_5541, SubBytesIns_Inst_Sbox_7_T3}), .b ({new_AGEMA_signal_5902, new_AGEMA_signal_5901, SubBytesIns_Inst_Sbox_7_T16}), .c ({new_AGEMA_signal_6336, new_AGEMA_signal_6335, SubBytesIns_Inst_Sbox_7_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T27_U1 ( .a ({new_AGEMA_signal_5538, new_AGEMA_signal_5537, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_5552, new_AGEMA_signal_5551, SubBytesIns_Inst_Sbox_7_T12}), .c ({new_AGEMA_signal_5908, new_AGEMA_signal_5907, SubBytesIns_Inst_Sbox_7_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T1_U1 ( .a ({ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .b ({ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .c ({new_AGEMA_signal_5558, new_AGEMA_signal_5557, SubBytesIns_Inst_Sbox_8_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T2_U1 ( .a ({ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .b ({ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_5560, new_AGEMA_signal_5559, SubBytesIns_Inst_Sbox_8_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T3_U1 ( .a ({ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .b ({ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_5562, new_AGEMA_signal_5561, SubBytesIns_Inst_Sbox_8_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T4_U1 ( .a ({ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .b ({ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_5564, new_AGEMA_signal_5563, SubBytesIns_Inst_Sbox_8_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T5_U1 ( .a ({ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}), .b ({ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_5566, new_AGEMA_signal_5565, SubBytesIns_Inst_Sbox_8_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T6_U1 ( .a ({new_AGEMA_signal_5558, new_AGEMA_signal_5557, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_5566, new_AGEMA_signal_5565, SubBytesIns_Inst_Sbox_8_T5}), .c ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, SubBytesIns_Inst_Sbox_8_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T7_U1 ( .a ({ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}), .b ({ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}), .c ({new_AGEMA_signal_5568, new_AGEMA_signal_5567, SubBytesIns_Inst_Sbox_8_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T8_U1 ( .a ({ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .b ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, SubBytesIns_Inst_Sbox_8_T6}), .c ({new_AGEMA_signal_6350, new_AGEMA_signal_6349, SubBytesIns_Inst_Sbox_8_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T9_U1 ( .a ({ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .b ({new_AGEMA_signal_5568, new_AGEMA_signal_5567, SubBytesIns_Inst_Sbox_8_T7}), .c ({new_AGEMA_signal_5912, new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_8_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T10_U1 ( .a ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, SubBytesIns_Inst_Sbox_8_T6}), .b ({new_AGEMA_signal_5568, new_AGEMA_signal_5567, SubBytesIns_Inst_Sbox_8_T7}), .c ({new_AGEMA_signal_6352, new_AGEMA_signal_6351, SubBytesIns_Inst_Sbox_8_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T11_U1 ( .a ({ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}), .b ({ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_5570, new_AGEMA_signal_5569, SubBytesIns_Inst_Sbox_8_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T12_U1 ( .a ({ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}), .b ({ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_5572, new_AGEMA_signal_5571, SubBytesIns_Inst_Sbox_8_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T13_U1 ( .a ({new_AGEMA_signal_5562, new_AGEMA_signal_5561, SubBytesIns_Inst_Sbox_8_T3}), .b ({new_AGEMA_signal_5564, new_AGEMA_signal_5563, SubBytesIns_Inst_Sbox_8_T4}), .c ({new_AGEMA_signal_5914, new_AGEMA_signal_5913, SubBytesIns_Inst_Sbox_8_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T14_U1 ( .a ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, SubBytesIns_Inst_Sbox_8_T6}), .b ({new_AGEMA_signal_5570, new_AGEMA_signal_5569, SubBytesIns_Inst_Sbox_8_T11}), .c ({new_AGEMA_signal_6354, new_AGEMA_signal_6353, SubBytesIns_Inst_Sbox_8_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T15_U1 ( .a ({new_AGEMA_signal_5566, new_AGEMA_signal_5565, SubBytesIns_Inst_Sbox_8_T5}), .b ({new_AGEMA_signal_5570, new_AGEMA_signal_5569, SubBytesIns_Inst_Sbox_8_T11}), .c ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, SubBytesIns_Inst_Sbox_8_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T16_U1 ( .a ({new_AGEMA_signal_5566, new_AGEMA_signal_5565, SubBytesIns_Inst_Sbox_8_T5}), .b ({new_AGEMA_signal_5572, new_AGEMA_signal_5571, SubBytesIns_Inst_Sbox_8_T12}), .c ({new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesIns_Inst_Sbox_8_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T17_U1 ( .a ({new_AGEMA_signal_5912, new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_8_T9}), .b ({new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesIns_Inst_Sbox_8_T16}), .c ({new_AGEMA_signal_6356, new_AGEMA_signal_6355, SubBytesIns_Inst_Sbox_8_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T18_U1 ( .a ({ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .b ({ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_5574, new_AGEMA_signal_5573, SubBytesIns_Inst_Sbox_8_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T19_U1 ( .a ({new_AGEMA_signal_5568, new_AGEMA_signal_5567, SubBytesIns_Inst_Sbox_8_T7}), .b ({new_AGEMA_signal_5574, new_AGEMA_signal_5573, SubBytesIns_Inst_Sbox_8_T18}), .c ({new_AGEMA_signal_5920, new_AGEMA_signal_5919, SubBytesIns_Inst_Sbox_8_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T20_U1 ( .a ({new_AGEMA_signal_5558, new_AGEMA_signal_5557, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_5920, new_AGEMA_signal_5919, SubBytesIns_Inst_Sbox_8_T19}), .c ({new_AGEMA_signal_6358, new_AGEMA_signal_6357, SubBytesIns_Inst_Sbox_8_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T21_U1 ( .a ({ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .b ({ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_5576, new_AGEMA_signal_5575, SubBytesIns_Inst_Sbox_8_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T22_U1 ( .a ({new_AGEMA_signal_5568, new_AGEMA_signal_5567, SubBytesIns_Inst_Sbox_8_T7}), .b ({new_AGEMA_signal_5576, new_AGEMA_signal_5575, SubBytesIns_Inst_Sbox_8_T21}), .c ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, SubBytesIns_Inst_Sbox_8_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T23_U1 ( .a ({new_AGEMA_signal_5560, new_AGEMA_signal_5559, SubBytesIns_Inst_Sbox_8_T2}), .b ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, SubBytesIns_Inst_Sbox_8_T22}), .c ({new_AGEMA_signal_6360, new_AGEMA_signal_6359, SubBytesIns_Inst_Sbox_8_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T24_U1 ( .a ({new_AGEMA_signal_5560, new_AGEMA_signal_5559, SubBytesIns_Inst_Sbox_8_T2}), .b ({new_AGEMA_signal_6352, new_AGEMA_signal_6351, SubBytesIns_Inst_Sbox_8_T10}), .c ({new_AGEMA_signal_6774, new_AGEMA_signal_6773, SubBytesIns_Inst_Sbox_8_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T25_U1 ( .a ({new_AGEMA_signal_6358, new_AGEMA_signal_6357, SubBytesIns_Inst_Sbox_8_T20}), .b ({new_AGEMA_signal_6356, new_AGEMA_signal_6355, SubBytesIns_Inst_Sbox_8_T17}), .c ({new_AGEMA_signal_6776, new_AGEMA_signal_6775, SubBytesIns_Inst_Sbox_8_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T26_U1 ( .a ({new_AGEMA_signal_5562, new_AGEMA_signal_5561, SubBytesIns_Inst_Sbox_8_T3}), .b ({new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesIns_Inst_Sbox_8_T16}), .c ({new_AGEMA_signal_6362, new_AGEMA_signal_6361, SubBytesIns_Inst_Sbox_8_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T27_U1 ( .a ({new_AGEMA_signal_5558, new_AGEMA_signal_5557, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_5572, new_AGEMA_signal_5571, SubBytesIns_Inst_Sbox_8_T12}), .c ({new_AGEMA_signal_5924, new_AGEMA_signal_5923, SubBytesIns_Inst_Sbox_8_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T1_U1 ( .a ({ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .b ({ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .c ({new_AGEMA_signal_5578, new_AGEMA_signal_5577, SubBytesIns_Inst_Sbox_9_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T2_U1 ( .a ({ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .b ({ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_5580, new_AGEMA_signal_5579, SubBytesIns_Inst_Sbox_9_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T3_U1 ( .a ({ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .b ({ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_5582, new_AGEMA_signal_5581, SubBytesIns_Inst_Sbox_9_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T4_U1 ( .a ({ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .b ({ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_5584, new_AGEMA_signal_5583, SubBytesIns_Inst_Sbox_9_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T5_U1 ( .a ({ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}), .b ({ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_5586, new_AGEMA_signal_5585, SubBytesIns_Inst_Sbox_9_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T6_U1 ( .a ({new_AGEMA_signal_5578, new_AGEMA_signal_5577, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_5586, new_AGEMA_signal_5585, SubBytesIns_Inst_Sbox_9_T5}), .c ({new_AGEMA_signal_5926, new_AGEMA_signal_5925, SubBytesIns_Inst_Sbox_9_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T7_U1 ( .a ({ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}), .b ({ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}), .c ({new_AGEMA_signal_5588, new_AGEMA_signal_5587, SubBytesIns_Inst_Sbox_9_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T8_U1 ( .a ({ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .b ({new_AGEMA_signal_5926, new_AGEMA_signal_5925, SubBytesIns_Inst_Sbox_9_T6}), .c ({new_AGEMA_signal_6376, new_AGEMA_signal_6375, SubBytesIns_Inst_Sbox_9_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T9_U1 ( .a ({ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .b ({new_AGEMA_signal_5588, new_AGEMA_signal_5587, SubBytesIns_Inst_Sbox_9_T7}), .c ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, SubBytesIns_Inst_Sbox_9_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T10_U1 ( .a ({new_AGEMA_signal_5926, new_AGEMA_signal_5925, SubBytesIns_Inst_Sbox_9_T6}), .b ({new_AGEMA_signal_5588, new_AGEMA_signal_5587, SubBytesIns_Inst_Sbox_9_T7}), .c ({new_AGEMA_signal_6378, new_AGEMA_signal_6377, SubBytesIns_Inst_Sbox_9_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T11_U1 ( .a ({ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}), .b ({ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_5590, new_AGEMA_signal_5589, SubBytesIns_Inst_Sbox_9_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T12_U1 ( .a ({ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}), .b ({ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_5592, new_AGEMA_signal_5591, SubBytesIns_Inst_Sbox_9_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T13_U1 ( .a ({new_AGEMA_signal_5582, new_AGEMA_signal_5581, SubBytesIns_Inst_Sbox_9_T3}), .b ({new_AGEMA_signal_5584, new_AGEMA_signal_5583, SubBytesIns_Inst_Sbox_9_T4}), .c ({new_AGEMA_signal_5930, new_AGEMA_signal_5929, SubBytesIns_Inst_Sbox_9_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T14_U1 ( .a ({new_AGEMA_signal_5926, new_AGEMA_signal_5925, SubBytesIns_Inst_Sbox_9_T6}), .b ({new_AGEMA_signal_5590, new_AGEMA_signal_5589, SubBytesIns_Inst_Sbox_9_T11}), .c ({new_AGEMA_signal_6380, new_AGEMA_signal_6379, SubBytesIns_Inst_Sbox_9_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T15_U1 ( .a ({new_AGEMA_signal_5586, new_AGEMA_signal_5585, SubBytesIns_Inst_Sbox_9_T5}), .b ({new_AGEMA_signal_5590, new_AGEMA_signal_5589, SubBytesIns_Inst_Sbox_9_T11}), .c ({new_AGEMA_signal_5932, new_AGEMA_signal_5931, SubBytesIns_Inst_Sbox_9_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T16_U1 ( .a ({new_AGEMA_signal_5586, new_AGEMA_signal_5585, SubBytesIns_Inst_Sbox_9_T5}), .b ({new_AGEMA_signal_5592, new_AGEMA_signal_5591, SubBytesIns_Inst_Sbox_9_T12}), .c ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, SubBytesIns_Inst_Sbox_9_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T17_U1 ( .a ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, SubBytesIns_Inst_Sbox_9_T9}), .b ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, SubBytesIns_Inst_Sbox_9_T16}), .c ({new_AGEMA_signal_6382, new_AGEMA_signal_6381, SubBytesIns_Inst_Sbox_9_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T18_U1 ( .a ({ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .b ({ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_5594, new_AGEMA_signal_5593, SubBytesIns_Inst_Sbox_9_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T19_U1 ( .a ({new_AGEMA_signal_5588, new_AGEMA_signal_5587, SubBytesIns_Inst_Sbox_9_T7}), .b ({new_AGEMA_signal_5594, new_AGEMA_signal_5593, SubBytesIns_Inst_Sbox_9_T18}), .c ({new_AGEMA_signal_5936, new_AGEMA_signal_5935, SubBytesIns_Inst_Sbox_9_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T20_U1 ( .a ({new_AGEMA_signal_5578, new_AGEMA_signal_5577, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_5936, new_AGEMA_signal_5935, SubBytesIns_Inst_Sbox_9_T19}), .c ({new_AGEMA_signal_6384, new_AGEMA_signal_6383, SubBytesIns_Inst_Sbox_9_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T21_U1 ( .a ({ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .b ({ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_5596, new_AGEMA_signal_5595, SubBytesIns_Inst_Sbox_9_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T22_U1 ( .a ({new_AGEMA_signal_5588, new_AGEMA_signal_5587, SubBytesIns_Inst_Sbox_9_T7}), .b ({new_AGEMA_signal_5596, new_AGEMA_signal_5595, SubBytesIns_Inst_Sbox_9_T21}), .c ({new_AGEMA_signal_5938, new_AGEMA_signal_5937, SubBytesIns_Inst_Sbox_9_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T23_U1 ( .a ({new_AGEMA_signal_5580, new_AGEMA_signal_5579, SubBytesIns_Inst_Sbox_9_T2}), .b ({new_AGEMA_signal_5938, new_AGEMA_signal_5937, SubBytesIns_Inst_Sbox_9_T22}), .c ({new_AGEMA_signal_6386, new_AGEMA_signal_6385, SubBytesIns_Inst_Sbox_9_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T24_U1 ( .a ({new_AGEMA_signal_5580, new_AGEMA_signal_5579, SubBytesIns_Inst_Sbox_9_T2}), .b ({new_AGEMA_signal_6378, new_AGEMA_signal_6377, SubBytesIns_Inst_Sbox_9_T10}), .c ({new_AGEMA_signal_6792, new_AGEMA_signal_6791, SubBytesIns_Inst_Sbox_9_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T25_U1 ( .a ({new_AGEMA_signal_6384, new_AGEMA_signal_6383, SubBytesIns_Inst_Sbox_9_T20}), .b ({new_AGEMA_signal_6382, new_AGEMA_signal_6381, SubBytesIns_Inst_Sbox_9_T17}), .c ({new_AGEMA_signal_6794, new_AGEMA_signal_6793, SubBytesIns_Inst_Sbox_9_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T26_U1 ( .a ({new_AGEMA_signal_5582, new_AGEMA_signal_5581, SubBytesIns_Inst_Sbox_9_T3}), .b ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, SubBytesIns_Inst_Sbox_9_T16}), .c ({new_AGEMA_signal_6388, new_AGEMA_signal_6387, SubBytesIns_Inst_Sbox_9_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T27_U1 ( .a ({new_AGEMA_signal_5578, new_AGEMA_signal_5577, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_5592, new_AGEMA_signal_5591, SubBytesIns_Inst_Sbox_9_T12}), .c ({new_AGEMA_signal_5940, new_AGEMA_signal_5939, SubBytesIns_Inst_Sbox_9_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T1_U1 ( .a ({ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .b ({ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .c ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, SubBytesIns_Inst_Sbox_10_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T2_U1 ( .a ({ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .b ({ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_5600, new_AGEMA_signal_5599, SubBytesIns_Inst_Sbox_10_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T3_U1 ( .a ({ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .b ({ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_5602, new_AGEMA_signal_5601, SubBytesIns_Inst_Sbox_10_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T4_U1 ( .a ({ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .b ({ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_5604, new_AGEMA_signal_5603, SubBytesIns_Inst_Sbox_10_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T5_U1 ( .a ({ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}), .b ({ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_5606, new_AGEMA_signal_5605, SubBytesIns_Inst_Sbox_10_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T6_U1 ( .a ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_5606, new_AGEMA_signal_5605, SubBytesIns_Inst_Sbox_10_T5}), .c ({new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_10_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T7_U1 ( .a ({ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}), .b ({ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}), .c ({new_AGEMA_signal_5608, new_AGEMA_signal_5607, SubBytesIns_Inst_Sbox_10_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T8_U1 ( .a ({ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .b ({new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_10_T6}), .c ({new_AGEMA_signal_6402, new_AGEMA_signal_6401, SubBytesIns_Inst_Sbox_10_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T9_U1 ( .a ({ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .b ({new_AGEMA_signal_5608, new_AGEMA_signal_5607, SubBytesIns_Inst_Sbox_10_T7}), .c ({new_AGEMA_signal_5944, new_AGEMA_signal_5943, SubBytesIns_Inst_Sbox_10_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T10_U1 ( .a ({new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_10_T6}), .b ({new_AGEMA_signal_5608, new_AGEMA_signal_5607, SubBytesIns_Inst_Sbox_10_T7}), .c ({new_AGEMA_signal_6404, new_AGEMA_signal_6403, SubBytesIns_Inst_Sbox_10_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T11_U1 ( .a ({ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}), .b ({ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_5610, new_AGEMA_signal_5609, SubBytesIns_Inst_Sbox_10_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T12_U1 ( .a ({ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}), .b ({ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_5612, new_AGEMA_signal_5611, SubBytesIns_Inst_Sbox_10_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T13_U1 ( .a ({new_AGEMA_signal_5602, new_AGEMA_signal_5601, SubBytesIns_Inst_Sbox_10_T3}), .b ({new_AGEMA_signal_5604, new_AGEMA_signal_5603, SubBytesIns_Inst_Sbox_10_T4}), .c ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, SubBytesIns_Inst_Sbox_10_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T14_U1 ( .a ({new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_10_T6}), .b ({new_AGEMA_signal_5610, new_AGEMA_signal_5609, SubBytesIns_Inst_Sbox_10_T11}), .c ({new_AGEMA_signal_6406, new_AGEMA_signal_6405, SubBytesIns_Inst_Sbox_10_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T15_U1 ( .a ({new_AGEMA_signal_5606, new_AGEMA_signal_5605, SubBytesIns_Inst_Sbox_10_T5}), .b ({new_AGEMA_signal_5610, new_AGEMA_signal_5609, SubBytesIns_Inst_Sbox_10_T11}), .c ({new_AGEMA_signal_5948, new_AGEMA_signal_5947, SubBytesIns_Inst_Sbox_10_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T16_U1 ( .a ({new_AGEMA_signal_5606, new_AGEMA_signal_5605, SubBytesIns_Inst_Sbox_10_T5}), .b ({new_AGEMA_signal_5612, new_AGEMA_signal_5611, SubBytesIns_Inst_Sbox_10_T12}), .c ({new_AGEMA_signal_5950, new_AGEMA_signal_5949, SubBytesIns_Inst_Sbox_10_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T17_U1 ( .a ({new_AGEMA_signal_5944, new_AGEMA_signal_5943, SubBytesIns_Inst_Sbox_10_T9}), .b ({new_AGEMA_signal_5950, new_AGEMA_signal_5949, SubBytesIns_Inst_Sbox_10_T16}), .c ({new_AGEMA_signal_6408, new_AGEMA_signal_6407, SubBytesIns_Inst_Sbox_10_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T18_U1 ( .a ({ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .b ({ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_5614, new_AGEMA_signal_5613, SubBytesIns_Inst_Sbox_10_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T19_U1 ( .a ({new_AGEMA_signal_5608, new_AGEMA_signal_5607, SubBytesIns_Inst_Sbox_10_T7}), .b ({new_AGEMA_signal_5614, new_AGEMA_signal_5613, SubBytesIns_Inst_Sbox_10_T18}), .c ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, SubBytesIns_Inst_Sbox_10_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T20_U1 ( .a ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, SubBytesIns_Inst_Sbox_10_T19}), .c ({new_AGEMA_signal_6410, new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_10_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T21_U1 ( .a ({ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .b ({ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_5616, new_AGEMA_signal_5615, SubBytesIns_Inst_Sbox_10_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T22_U1 ( .a ({new_AGEMA_signal_5608, new_AGEMA_signal_5607, SubBytesIns_Inst_Sbox_10_T7}), .b ({new_AGEMA_signal_5616, new_AGEMA_signal_5615, SubBytesIns_Inst_Sbox_10_T21}), .c ({new_AGEMA_signal_5954, new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_10_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T23_U1 ( .a ({new_AGEMA_signal_5600, new_AGEMA_signal_5599, SubBytesIns_Inst_Sbox_10_T2}), .b ({new_AGEMA_signal_5954, new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_10_T22}), .c ({new_AGEMA_signal_6412, new_AGEMA_signal_6411, SubBytesIns_Inst_Sbox_10_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T24_U1 ( .a ({new_AGEMA_signal_5600, new_AGEMA_signal_5599, SubBytesIns_Inst_Sbox_10_T2}), .b ({new_AGEMA_signal_6404, new_AGEMA_signal_6403, SubBytesIns_Inst_Sbox_10_T10}), .c ({new_AGEMA_signal_6810, new_AGEMA_signal_6809, SubBytesIns_Inst_Sbox_10_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T25_U1 ( .a ({new_AGEMA_signal_6410, new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_10_T20}), .b ({new_AGEMA_signal_6408, new_AGEMA_signal_6407, SubBytesIns_Inst_Sbox_10_T17}), .c ({new_AGEMA_signal_6812, new_AGEMA_signal_6811, SubBytesIns_Inst_Sbox_10_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T26_U1 ( .a ({new_AGEMA_signal_5602, new_AGEMA_signal_5601, SubBytesIns_Inst_Sbox_10_T3}), .b ({new_AGEMA_signal_5950, new_AGEMA_signal_5949, SubBytesIns_Inst_Sbox_10_T16}), .c ({new_AGEMA_signal_6414, new_AGEMA_signal_6413, SubBytesIns_Inst_Sbox_10_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T27_U1 ( .a ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_5612, new_AGEMA_signal_5611, SubBytesIns_Inst_Sbox_10_T12}), .c ({new_AGEMA_signal_5956, new_AGEMA_signal_5955, SubBytesIns_Inst_Sbox_10_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T1_U1 ( .a ({ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_5618, new_AGEMA_signal_5617, SubBytesIns_Inst_Sbox_11_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T2_U1 ( .a ({ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_5620, new_AGEMA_signal_5619, SubBytesIns_Inst_Sbox_11_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T3_U1 ( .a ({ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_5622, new_AGEMA_signal_5621, SubBytesIns_Inst_Sbox_11_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T4_U1 ( .a ({ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_5624, new_AGEMA_signal_5623, SubBytesIns_Inst_Sbox_11_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T5_U1 ( .a ({ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}), .b ({ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_5626, new_AGEMA_signal_5625, SubBytesIns_Inst_Sbox_11_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T6_U1 ( .a ({new_AGEMA_signal_5618, new_AGEMA_signal_5617, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_5626, new_AGEMA_signal_5625, SubBytesIns_Inst_Sbox_11_T5}), .c ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, SubBytesIns_Inst_Sbox_11_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T7_U1 ( .a ({ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_5628, new_AGEMA_signal_5627, SubBytesIns_Inst_Sbox_11_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T8_U1 ( .a ({ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .b ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, SubBytesIns_Inst_Sbox_11_T6}), .c ({new_AGEMA_signal_6428, new_AGEMA_signal_6427, SubBytesIns_Inst_Sbox_11_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T9_U1 ( .a ({ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .b ({new_AGEMA_signal_5628, new_AGEMA_signal_5627, SubBytesIns_Inst_Sbox_11_T7}), .c ({new_AGEMA_signal_5960, new_AGEMA_signal_5959, SubBytesIns_Inst_Sbox_11_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T10_U1 ( .a ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, SubBytesIns_Inst_Sbox_11_T6}), .b ({new_AGEMA_signal_5628, new_AGEMA_signal_5627, SubBytesIns_Inst_Sbox_11_T7}), .c ({new_AGEMA_signal_6430, new_AGEMA_signal_6429, SubBytesIns_Inst_Sbox_11_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T11_U1 ( .a ({ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_5630, new_AGEMA_signal_5629, SubBytesIns_Inst_Sbox_11_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T12_U1 ( .a ({ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_5632, new_AGEMA_signal_5631, SubBytesIns_Inst_Sbox_11_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T13_U1 ( .a ({new_AGEMA_signal_5622, new_AGEMA_signal_5621, SubBytesIns_Inst_Sbox_11_T3}), .b ({new_AGEMA_signal_5624, new_AGEMA_signal_5623, SubBytesIns_Inst_Sbox_11_T4}), .c ({new_AGEMA_signal_5962, new_AGEMA_signal_5961, SubBytesIns_Inst_Sbox_11_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T14_U1 ( .a ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, SubBytesIns_Inst_Sbox_11_T6}), .b ({new_AGEMA_signal_5630, new_AGEMA_signal_5629, SubBytesIns_Inst_Sbox_11_T11}), .c ({new_AGEMA_signal_6432, new_AGEMA_signal_6431, SubBytesIns_Inst_Sbox_11_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T15_U1 ( .a ({new_AGEMA_signal_5626, new_AGEMA_signal_5625, SubBytesIns_Inst_Sbox_11_T5}), .b ({new_AGEMA_signal_5630, new_AGEMA_signal_5629, SubBytesIns_Inst_Sbox_11_T11}), .c ({new_AGEMA_signal_5964, new_AGEMA_signal_5963, SubBytesIns_Inst_Sbox_11_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T16_U1 ( .a ({new_AGEMA_signal_5626, new_AGEMA_signal_5625, SubBytesIns_Inst_Sbox_11_T5}), .b ({new_AGEMA_signal_5632, new_AGEMA_signal_5631, SubBytesIns_Inst_Sbox_11_T12}), .c ({new_AGEMA_signal_5966, new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_11_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T17_U1 ( .a ({new_AGEMA_signal_5960, new_AGEMA_signal_5959, SubBytesIns_Inst_Sbox_11_T9}), .b ({new_AGEMA_signal_5966, new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_11_T16}), .c ({new_AGEMA_signal_6434, new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_11_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T18_U1 ( .a ({ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_5634, new_AGEMA_signal_5633, SubBytesIns_Inst_Sbox_11_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T19_U1 ( .a ({new_AGEMA_signal_5628, new_AGEMA_signal_5627, SubBytesIns_Inst_Sbox_11_T7}), .b ({new_AGEMA_signal_5634, new_AGEMA_signal_5633, SubBytesIns_Inst_Sbox_11_T18}), .c ({new_AGEMA_signal_5968, new_AGEMA_signal_5967, SubBytesIns_Inst_Sbox_11_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T20_U1 ( .a ({new_AGEMA_signal_5618, new_AGEMA_signal_5617, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_5968, new_AGEMA_signal_5967, SubBytesIns_Inst_Sbox_11_T19}), .c ({new_AGEMA_signal_6436, new_AGEMA_signal_6435, SubBytesIns_Inst_Sbox_11_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T21_U1 ( .a ({ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .b ({ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_5636, new_AGEMA_signal_5635, SubBytesIns_Inst_Sbox_11_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T22_U1 ( .a ({new_AGEMA_signal_5628, new_AGEMA_signal_5627, SubBytesIns_Inst_Sbox_11_T7}), .b ({new_AGEMA_signal_5636, new_AGEMA_signal_5635, SubBytesIns_Inst_Sbox_11_T21}), .c ({new_AGEMA_signal_5970, new_AGEMA_signal_5969, SubBytesIns_Inst_Sbox_11_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T23_U1 ( .a ({new_AGEMA_signal_5620, new_AGEMA_signal_5619, SubBytesIns_Inst_Sbox_11_T2}), .b ({new_AGEMA_signal_5970, new_AGEMA_signal_5969, SubBytesIns_Inst_Sbox_11_T22}), .c ({new_AGEMA_signal_6438, new_AGEMA_signal_6437, SubBytesIns_Inst_Sbox_11_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T24_U1 ( .a ({new_AGEMA_signal_5620, new_AGEMA_signal_5619, SubBytesIns_Inst_Sbox_11_T2}), .b ({new_AGEMA_signal_6430, new_AGEMA_signal_6429, SubBytesIns_Inst_Sbox_11_T10}), .c ({new_AGEMA_signal_6828, new_AGEMA_signal_6827, SubBytesIns_Inst_Sbox_11_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T25_U1 ( .a ({new_AGEMA_signal_6436, new_AGEMA_signal_6435, SubBytesIns_Inst_Sbox_11_T20}), .b ({new_AGEMA_signal_6434, new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_11_T17}), .c ({new_AGEMA_signal_6830, new_AGEMA_signal_6829, SubBytesIns_Inst_Sbox_11_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T26_U1 ( .a ({new_AGEMA_signal_5622, new_AGEMA_signal_5621, SubBytesIns_Inst_Sbox_11_T3}), .b ({new_AGEMA_signal_5966, new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_11_T16}), .c ({new_AGEMA_signal_6440, new_AGEMA_signal_6439, SubBytesIns_Inst_Sbox_11_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T27_U1 ( .a ({new_AGEMA_signal_5618, new_AGEMA_signal_5617, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_5632, new_AGEMA_signal_5631, SubBytesIns_Inst_Sbox_11_T12}), .c ({new_AGEMA_signal_5972, new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_11_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T1_U1 ( .a ({ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .c ({new_AGEMA_signal_5638, new_AGEMA_signal_5637, SubBytesIns_Inst_Sbox_12_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T2_U1 ( .a ({ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_5640, new_AGEMA_signal_5639, SubBytesIns_Inst_Sbox_12_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T3_U1 ( .a ({ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_5642, new_AGEMA_signal_5641, SubBytesIns_Inst_Sbox_12_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T4_U1 ( .a ({ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .b ({ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_5644, new_AGEMA_signal_5643, SubBytesIns_Inst_Sbox_12_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T5_U1 ( .a ({ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}), .b ({ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_5646, new_AGEMA_signal_5645, SubBytesIns_Inst_Sbox_12_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T6_U1 ( .a ({new_AGEMA_signal_5638, new_AGEMA_signal_5637, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_5646, new_AGEMA_signal_5645, SubBytesIns_Inst_Sbox_12_T5}), .c ({new_AGEMA_signal_5974, new_AGEMA_signal_5973, SubBytesIns_Inst_Sbox_12_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T7_U1 ( .a ({ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}), .b ({ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}), .c ({new_AGEMA_signal_5648, new_AGEMA_signal_5647, SubBytesIns_Inst_Sbox_12_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T8_U1 ( .a ({ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .b ({new_AGEMA_signal_5974, new_AGEMA_signal_5973, SubBytesIns_Inst_Sbox_12_T6}), .c ({new_AGEMA_signal_6454, new_AGEMA_signal_6453, SubBytesIns_Inst_Sbox_12_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T9_U1 ( .a ({ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .b ({new_AGEMA_signal_5648, new_AGEMA_signal_5647, SubBytesIns_Inst_Sbox_12_T7}), .c ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, SubBytesIns_Inst_Sbox_12_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T10_U1 ( .a ({new_AGEMA_signal_5974, new_AGEMA_signal_5973, SubBytesIns_Inst_Sbox_12_T6}), .b ({new_AGEMA_signal_5648, new_AGEMA_signal_5647, SubBytesIns_Inst_Sbox_12_T7}), .c ({new_AGEMA_signal_6456, new_AGEMA_signal_6455, SubBytesIns_Inst_Sbox_12_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T11_U1 ( .a ({ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}), .b ({ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_5650, new_AGEMA_signal_5649, SubBytesIns_Inst_Sbox_12_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T12_U1 ( .a ({ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}), .b ({ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_5652, new_AGEMA_signal_5651, SubBytesIns_Inst_Sbox_12_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T13_U1 ( .a ({new_AGEMA_signal_5642, new_AGEMA_signal_5641, SubBytesIns_Inst_Sbox_12_T3}), .b ({new_AGEMA_signal_5644, new_AGEMA_signal_5643, SubBytesIns_Inst_Sbox_12_T4}), .c ({new_AGEMA_signal_5978, new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_12_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T14_U1 ( .a ({new_AGEMA_signal_5974, new_AGEMA_signal_5973, SubBytesIns_Inst_Sbox_12_T6}), .b ({new_AGEMA_signal_5650, new_AGEMA_signal_5649, SubBytesIns_Inst_Sbox_12_T11}), .c ({new_AGEMA_signal_6458, new_AGEMA_signal_6457, SubBytesIns_Inst_Sbox_12_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T15_U1 ( .a ({new_AGEMA_signal_5646, new_AGEMA_signal_5645, SubBytesIns_Inst_Sbox_12_T5}), .b ({new_AGEMA_signal_5650, new_AGEMA_signal_5649, SubBytesIns_Inst_Sbox_12_T11}), .c ({new_AGEMA_signal_5980, new_AGEMA_signal_5979, SubBytesIns_Inst_Sbox_12_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T16_U1 ( .a ({new_AGEMA_signal_5646, new_AGEMA_signal_5645, SubBytesIns_Inst_Sbox_12_T5}), .b ({new_AGEMA_signal_5652, new_AGEMA_signal_5651, SubBytesIns_Inst_Sbox_12_T12}), .c ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, SubBytesIns_Inst_Sbox_12_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T17_U1 ( .a ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, SubBytesIns_Inst_Sbox_12_T9}), .b ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, SubBytesIns_Inst_Sbox_12_T16}), .c ({new_AGEMA_signal_6460, new_AGEMA_signal_6459, SubBytesIns_Inst_Sbox_12_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T18_U1 ( .a ({ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .b ({ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_5654, new_AGEMA_signal_5653, SubBytesIns_Inst_Sbox_12_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T19_U1 ( .a ({new_AGEMA_signal_5648, new_AGEMA_signal_5647, SubBytesIns_Inst_Sbox_12_T7}), .b ({new_AGEMA_signal_5654, new_AGEMA_signal_5653, SubBytesIns_Inst_Sbox_12_T18}), .c ({new_AGEMA_signal_5984, new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_12_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T20_U1 ( .a ({new_AGEMA_signal_5638, new_AGEMA_signal_5637, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_5984, new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_12_T19}), .c ({new_AGEMA_signal_6462, new_AGEMA_signal_6461, SubBytesIns_Inst_Sbox_12_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T21_U1 ( .a ({ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .b ({ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_5656, new_AGEMA_signal_5655, SubBytesIns_Inst_Sbox_12_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T22_U1 ( .a ({new_AGEMA_signal_5648, new_AGEMA_signal_5647, SubBytesIns_Inst_Sbox_12_T7}), .b ({new_AGEMA_signal_5656, new_AGEMA_signal_5655, SubBytesIns_Inst_Sbox_12_T21}), .c ({new_AGEMA_signal_5986, new_AGEMA_signal_5985, SubBytesIns_Inst_Sbox_12_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T23_U1 ( .a ({new_AGEMA_signal_5640, new_AGEMA_signal_5639, SubBytesIns_Inst_Sbox_12_T2}), .b ({new_AGEMA_signal_5986, new_AGEMA_signal_5985, SubBytesIns_Inst_Sbox_12_T22}), .c ({new_AGEMA_signal_6464, new_AGEMA_signal_6463, SubBytesIns_Inst_Sbox_12_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T24_U1 ( .a ({new_AGEMA_signal_5640, new_AGEMA_signal_5639, SubBytesIns_Inst_Sbox_12_T2}), .b ({new_AGEMA_signal_6456, new_AGEMA_signal_6455, SubBytesIns_Inst_Sbox_12_T10}), .c ({new_AGEMA_signal_6846, new_AGEMA_signal_6845, SubBytesIns_Inst_Sbox_12_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T25_U1 ( .a ({new_AGEMA_signal_6462, new_AGEMA_signal_6461, SubBytesIns_Inst_Sbox_12_T20}), .b ({new_AGEMA_signal_6460, new_AGEMA_signal_6459, SubBytesIns_Inst_Sbox_12_T17}), .c ({new_AGEMA_signal_6848, new_AGEMA_signal_6847, SubBytesIns_Inst_Sbox_12_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T26_U1 ( .a ({new_AGEMA_signal_5642, new_AGEMA_signal_5641, SubBytesIns_Inst_Sbox_12_T3}), .b ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, SubBytesIns_Inst_Sbox_12_T16}), .c ({new_AGEMA_signal_6466, new_AGEMA_signal_6465, SubBytesIns_Inst_Sbox_12_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T27_U1 ( .a ({new_AGEMA_signal_5638, new_AGEMA_signal_5637, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_5652, new_AGEMA_signal_5651, SubBytesIns_Inst_Sbox_12_T12}), .c ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, SubBytesIns_Inst_Sbox_12_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T1_U1 ( .a ({ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .b ({ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .c ({new_AGEMA_signal_5658, new_AGEMA_signal_5657, SubBytesIns_Inst_Sbox_13_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T2_U1 ( .a ({ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .b ({ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_5660, new_AGEMA_signal_5659, SubBytesIns_Inst_Sbox_13_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T3_U1 ( .a ({ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .b ({ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_5662, new_AGEMA_signal_5661, SubBytesIns_Inst_Sbox_13_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T4_U1 ( .a ({ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .b ({ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_5664, new_AGEMA_signal_5663, SubBytesIns_Inst_Sbox_13_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T5_U1 ( .a ({ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}), .b ({ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_5666, new_AGEMA_signal_5665, SubBytesIns_Inst_Sbox_13_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T6_U1 ( .a ({new_AGEMA_signal_5658, new_AGEMA_signal_5657, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_5666, new_AGEMA_signal_5665, SubBytesIns_Inst_Sbox_13_T5}), .c ({new_AGEMA_signal_5990, new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_13_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T7_U1 ( .a ({ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}), .b ({ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}), .c ({new_AGEMA_signal_5668, new_AGEMA_signal_5667, SubBytesIns_Inst_Sbox_13_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T8_U1 ( .a ({ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .b ({new_AGEMA_signal_5990, new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_13_T6}), .c ({new_AGEMA_signal_6480, new_AGEMA_signal_6479, SubBytesIns_Inst_Sbox_13_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T9_U1 ( .a ({ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .b ({new_AGEMA_signal_5668, new_AGEMA_signal_5667, SubBytesIns_Inst_Sbox_13_T7}), .c ({new_AGEMA_signal_5992, new_AGEMA_signal_5991, SubBytesIns_Inst_Sbox_13_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T10_U1 ( .a ({new_AGEMA_signal_5990, new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_13_T6}), .b ({new_AGEMA_signal_5668, new_AGEMA_signal_5667, SubBytesIns_Inst_Sbox_13_T7}), .c ({new_AGEMA_signal_6482, new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_13_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T11_U1 ( .a ({ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}), .b ({ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_5670, new_AGEMA_signal_5669, SubBytesIns_Inst_Sbox_13_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T12_U1 ( .a ({ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}), .b ({ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_5672, new_AGEMA_signal_5671, SubBytesIns_Inst_Sbox_13_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T13_U1 ( .a ({new_AGEMA_signal_5662, new_AGEMA_signal_5661, SubBytesIns_Inst_Sbox_13_T3}), .b ({new_AGEMA_signal_5664, new_AGEMA_signal_5663, SubBytesIns_Inst_Sbox_13_T4}), .c ({new_AGEMA_signal_5994, new_AGEMA_signal_5993, SubBytesIns_Inst_Sbox_13_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T14_U1 ( .a ({new_AGEMA_signal_5990, new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_13_T6}), .b ({new_AGEMA_signal_5670, new_AGEMA_signal_5669, SubBytesIns_Inst_Sbox_13_T11}), .c ({new_AGEMA_signal_6484, new_AGEMA_signal_6483, SubBytesIns_Inst_Sbox_13_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T15_U1 ( .a ({new_AGEMA_signal_5666, new_AGEMA_signal_5665, SubBytesIns_Inst_Sbox_13_T5}), .b ({new_AGEMA_signal_5670, new_AGEMA_signal_5669, SubBytesIns_Inst_Sbox_13_T11}), .c ({new_AGEMA_signal_5996, new_AGEMA_signal_5995, SubBytesIns_Inst_Sbox_13_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T16_U1 ( .a ({new_AGEMA_signal_5666, new_AGEMA_signal_5665, SubBytesIns_Inst_Sbox_13_T5}), .b ({new_AGEMA_signal_5672, new_AGEMA_signal_5671, SubBytesIns_Inst_Sbox_13_T12}), .c ({new_AGEMA_signal_5998, new_AGEMA_signal_5997, SubBytesIns_Inst_Sbox_13_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T17_U1 ( .a ({new_AGEMA_signal_5992, new_AGEMA_signal_5991, SubBytesIns_Inst_Sbox_13_T9}), .b ({new_AGEMA_signal_5998, new_AGEMA_signal_5997, SubBytesIns_Inst_Sbox_13_T16}), .c ({new_AGEMA_signal_6486, new_AGEMA_signal_6485, SubBytesIns_Inst_Sbox_13_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T18_U1 ( .a ({ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .b ({ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_5674, new_AGEMA_signal_5673, SubBytesIns_Inst_Sbox_13_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T19_U1 ( .a ({new_AGEMA_signal_5668, new_AGEMA_signal_5667, SubBytesIns_Inst_Sbox_13_T7}), .b ({new_AGEMA_signal_5674, new_AGEMA_signal_5673, SubBytesIns_Inst_Sbox_13_T18}), .c ({new_AGEMA_signal_6000, new_AGEMA_signal_5999, SubBytesIns_Inst_Sbox_13_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T20_U1 ( .a ({new_AGEMA_signal_5658, new_AGEMA_signal_5657, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_6000, new_AGEMA_signal_5999, SubBytesIns_Inst_Sbox_13_T19}), .c ({new_AGEMA_signal_6488, new_AGEMA_signal_6487, SubBytesIns_Inst_Sbox_13_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T21_U1 ( .a ({ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .b ({ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_5676, new_AGEMA_signal_5675, SubBytesIns_Inst_Sbox_13_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T22_U1 ( .a ({new_AGEMA_signal_5668, new_AGEMA_signal_5667, SubBytesIns_Inst_Sbox_13_T7}), .b ({new_AGEMA_signal_5676, new_AGEMA_signal_5675, SubBytesIns_Inst_Sbox_13_T21}), .c ({new_AGEMA_signal_6002, new_AGEMA_signal_6001, SubBytesIns_Inst_Sbox_13_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T23_U1 ( .a ({new_AGEMA_signal_5660, new_AGEMA_signal_5659, SubBytesIns_Inst_Sbox_13_T2}), .b ({new_AGEMA_signal_6002, new_AGEMA_signal_6001, SubBytesIns_Inst_Sbox_13_T22}), .c ({new_AGEMA_signal_6490, new_AGEMA_signal_6489, SubBytesIns_Inst_Sbox_13_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T24_U1 ( .a ({new_AGEMA_signal_5660, new_AGEMA_signal_5659, SubBytesIns_Inst_Sbox_13_T2}), .b ({new_AGEMA_signal_6482, new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_13_T10}), .c ({new_AGEMA_signal_6864, new_AGEMA_signal_6863, SubBytesIns_Inst_Sbox_13_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T25_U1 ( .a ({new_AGEMA_signal_6488, new_AGEMA_signal_6487, SubBytesIns_Inst_Sbox_13_T20}), .b ({new_AGEMA_signal_6486, new_AGEMA_signal_6485, SubBytesIns_Inst_Sbox_13_T17}), .c ({new_AGEMA_signal_6866, new_AGEMA_signal_6865, SubBytesIns_Inst_Sbox_13_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T26_U1 ( .a ({new_AGEMA_signal_5662, new_AGEMA_signal_5661, SubBytesIns_Inst_Sbox_13_T3}), .b ({new_AGEMA_signal_5998, new_AGEMA_signal_5997, SubBytesIns_Inst_Sbox_13_T16}), .c ({new_AGEMA_signal_6492, new_AGEMA_signal_6491, SubBytesIns_Inst_Sbox_13_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T27_U1 ( .a ({new_AGEMA_signal_5658, new_AGEMA_signal_5657, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_5672, new_AGEMA_signal_5671, SubBytesIns_Inst_Sbox_13_T12}), .c ({new_AGEMA_signal_6004, new_AGEMA_signal_6003, SubBytesIns_Inst_Sbox_13_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T1_U1 ( .a ({ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .b ({ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .c ({new_AGEMA_signal_5678, new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_14_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T2_U1 ( .a ({ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .b ({ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_5680, new_AGEMA_signal_5679, SubBytesIns_Inst_Sbox_14_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T3_U1 ( .a ({ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .b ({ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_5682, new_AGEMA_signal_5681, SubBytesIns_Inst_Sbox_14_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T4_U1 ( .a ({ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .b ({ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_5684, new_AGEMA_signal_5683, SubBytesIns_Inst_Sbox_14_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T5_U1 ( .a ({ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}), .b ({ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_5686, new_AGEMA_signal_5685, SubBytesIns_Inst_Sbox_14_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T6_U1 ( .a ({new_AGEMA_signal_5678, new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_5686, new_AGEMA_signal_5685, SubBytesIns_Inst_Sbox_14_T5}), .c ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, SubBytesIns_Inst_Sbox_14_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T7_U1 ( .a ({ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}), .b ({ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}), .c ({new_AGEMA_signal_5688, new_AGEMA_signal_5687, SubBytesIns_Inst_Sbox_14_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T8_U1 ( .a ({ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .b ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, SubBytesIns_Inst_Sbox_14_T6}), .c ({new_AGEMA_signal_6506, new_AGEMA_signal_6505, SubBytesIns_Inst_Sbox_14_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T9_U1 ( .a ({ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .b ({new_AGEMA_signal_5688, new_AGEMA_signal_5687, SubBytesIns_Inst_Sbox_14_T7}), .c ({new_AGEMA_signal_6008, new_AGEMA_signal_6007, SubBytesIns_Inst_Sbox_14_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T10_U1 ( .a ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, SubBytesIns_Inst_Sbox_14_T6}), .b ({new_AGEMA_signal_5688, new_AGEMA_signal_5687, SubBytesIns_Inst_Sbox_14_T7}), .c ({new_AGEMA_signal_6508, new_AGEMA_signal_6507, SubBytesIns_Inst_Sbox_14_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T11_U1 ( .a ({ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}), .b ({ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_5690, new_AGEMA_signal_5689, SubBytesIns_Inst_Sbox_14_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T12_U1 ( .a ({ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}), .b ({ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_5692, new_AGEMA_signal_5691, SubBytesIns_Inst_Sbox_14_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T13_U1 ( .a ({new_AGEMA_signal_5682, new_AGEMA_signal_5681, SubBytesIns_Inst_Sbox_14_T3}), .b ({new_AGEMA_signal_5684, new_AGEMA_signal_5683, SubBytesIns_Inst_Sbox_14_T4}), .c ({new_AGEMA_signal_6010, new_AGEMA_signal_6009, SubBytesIns_Inst_Sbox_14_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T14_U1 ( .a ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, SubBytesIns_Inst_Sbox_14_T6}), .b ({new_AGEMA_signal_5690, new_AGEMA_signal_5689, SubBytesIns_Inst_Sbox_14_T11}), .c ({new_AGEMA_signal_6510, new_AGEMA_signal_6509, SubBytesIns_Inst_Sbox_14_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T15_U1 ( .a ({new_AGEMA_signal_5686, new_AGEMA_signal_5685, SubBytesIns_Inst_Sbox_14_T5}), .b ({new_AGEMA_signal_5690, new_AGEMA_signal_5689, SubBytesIns_Inst_Sbox_14_T11}), .c ({new_AGEMA_signal_6012, new_AGEMA_signal_6011, SubBytesIns_Inst_Sbox_14_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T16_U1 ( .a ({new_AGEMA_signal_5686, new_AGEMA_signal_5685, SubBytesIns_Inst_Sbox_14_T5}), .b ({new_AGEMA_signal_5692, new_AGEMA_signal_5691, SubBytesIns_Inst_Sbox_14_T12}), .c ({new_AGEMA_signal_6014, new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_14_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T17_U1 ( .a ({new_AGEMA_signal_6008, new_AGEMA_signal_6007, SubBytesIns_Inst_Sbox_14_T9}), .b ({new_AGEMA_signal_6014, new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_14_T16}), .c ({new_AGEMA_signal_6512, new_AGEMA_signal_6511, SubBytesIns_Inst_Sbox_14_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T18_U1 ( .a ({ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .b ({ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_5694, new_AGEMA_signal_5693, SubBytesIns_Inst_Sbox_14_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T19_U1 ( .a ({new_AGEMA_signal_5688, new_AGEMA_signal_5687, SubBytesIns_Inst_Sbox_14_T7}), .b ({new_AGEMA_signal_5694, new_AGEMA_signal_5693, SubBytesIns_Inst_Sbox_14_T18}), .c ({new_AGEMA_signal_6016, new_AGEMA_signal_6015, SubBytesIns_Inst_Sbox_14_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T20_U1 ( .a ({new_AGEMA_signal_5678, new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_6016, new_AGEMA_signal_6015, SubBytesIns_Inst_Sbox_14_T19}), .c ({new_AGEMA_signal_6514, new_AGEMA_signal_6513, SubBytesIns_Inst_Sbox_14_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T21_U1 ( .a ({ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .b ({ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_5696, new_AGEMA_signal_5695, SubBytesIns_Inst_Sbox_14_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T22_U1 ( .a ({new_AGEMA_signal_5688, new_AGEMA_signal_5687, SubBytesIns_Inst_Sbox_14_T7}), .b ({new_AGEMA_signal_5696, new_AGEMA_signal_5695, SubBytesIns_Inst_Sbox_14_T21}), .c ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, SubBytesIns_Inst_Sbox_14_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T23_U1 ( .a ({new_AGEMA_signal_5680, new_AGEMA_signal_5679, SubBytesIns_Inst_Sbox_14_T2}), .b ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, SubBytesIns_Inst_Sbox_14_T22}), .c ({new_AGEMA_signal_6516, new_AGEMA_signal_6515, SubBytesIns_Inst_Sbox_14_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T24_U1 ( .a ({new_AGEMA_signal_5680, new_AGEMA_signal_5679, SubBytesIns_Inst_Sbox_14_T2}), .b ({new_AGEMA_signal_6508, new_AGEMA_signal_6507, SubBytesIns_Inst_Sbox_14_T10}), .c ({new_AGEMA_signal_6882, new_AGEMA_signal_6881, SubBytesIns_Inst_Sbox_14_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T25_U1 ( .a ({new_AGEMA_signal_6514, new_AGEMA_signal_6513, SubBytesIns_Inst_Sbox_14_T20}), .b ({new_AGEMA_signal_6512, new_AGEMA_signal_6511, SubBytesIns_Inst_Sbox_14_T17}), .c ({new_AGEMA_signal_6884, new_AGEMA_signal_6883, SubBytesIns_Inst_Sbox_14_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T26_U1 ( .a ({new_AGEMA_signal_5682, new_AGEMA_signal_5681, SubBytesIns_Inst_Sbox_14_T3}), .b ({new_AGEMA_signal_6014, new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_14_T16}), .c ({new_AGEMA_signal_6518, new_AGEMA_signal_6517, SubBytesIns_Inst_Sbox_14_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T27_U1 ( .a ({new_AGEMA_signal_5678, new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_5692, new_AGEMA_signal_5691, SubBytesIns_Inst_Sbox_14_T12}), .c ({new_AGEMA_signal_6020, new_AGEMA_signal_6019, SubBytesIns_Inst_Sbox_14_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T1_U1 ( .a ({ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_5698, new_AGEMA_signal_5697, SubBytesIns_Inst_Sbox_15_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T2_U1 ( .a ({ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_5700, new_AGEMA_signal_5699, SubBytesIns_Inst_Sbox_15_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T3_U1 ( .a ({ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_5702, new_AGEMA_signal_5701, SubBytesIns_Inst_Sbox_15_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T4_U1 ( .a ({ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_5704, new_AGEMA_signal_5703, SubBytesIns_Inst_Sbox_15_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T5_U1 ( .a ({ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}), .b ({ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, SubBytesIns_Inst_Sbox_15_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T6_U1 ( .a ({new_AGEMA_signal_5698, new_AGEMA_signal_5697, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, SubBytesIns_Inst_Sbox_15_T5}), .c ({new_AGEMA_signal_6022, new_AGEMA_signal_6021, SubBytesIns_Inst_Sbox_15_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T7_U1 ( .a ({ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_5708, new_AGEMA_signal_5707, SubBytesIns_Inst_Sbox_15_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T8_U1 ( .a ({ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_6022, new_AGEMA_signal_6021, SubBytesIns_Inst_Sbox_15_T6}), .c ({new_AGEMA_signal_6532, new_AGEMA_signal_6531, SubBytesIns_Inst_Sbox_15_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T9_U1 ( .a ({ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_5708, new_AGEMA_signal_5707, SubBytesIns_Inst_Sbox_15_T7}), .c ({new_AGEMA_signal_6024, new_AGEMA_signal_6023, SubBytesIns_Inst_Sbox_15_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T10_U1 ( .a ({new_AGEMA_signal_6022, new_AGEMA_signal_6021, SubBytesIns_Inst_Sbox_15_T6}), .b ({new_AGEMA_signal_5708, new_AGEMA_signal_5707, SubBytesIns_Inst_Sbox_15_T7}), .c ({new_AGEMA_signal_6534, new_AGEMA_signal_6533, SubBytesIns_Inst_Sbox_15_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T11_U1 ( .a ({ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_5710, new_AGEMA_signal_5709, SubBytesIns_Inst_Sbox_15_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T12_U1 ( .a ({ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_5712, new_AGEMA_signal_5711, SubBytesIns_Inst_Sbox_15_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T13_U1 ( .a ({new_AGEMA_signal_5702, new_AGEMA_signal_5701, SubBytesIns_Inst_Sbox_15_T3}), .b ({new_AGEMA_signal_5704, new_AGEMA_signal_5703, SubBytesIns_Inst_Sbox_15_T4}), .c ({new_AGEMA_signal_6026, new_AGEMA_signal_6025, SubBytesIns_Inst_Sbox_15_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T14_U1 ( .a ({new_AGEMA_signal_6022, new_AGEMA_signal_6021, SubBytesIns_Inst_Sbox_15_T6}), .b ({new_AGEMA_signal_5710, new_AGEMA_signal_5709, SubBytesIns_Inst_Sbox_15_T11}), .c ({new_AGEMA_signal_6536, new_AGEMA_signal_6535, SubBytesIns_Inst_Sbox_15_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T15_U1 ( .a ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, SubBytesIns_Inst_Sbox_15_T5}), .b ({new_AGEMA_signal_5710, new_AGEMA_signal_5709, SubBytesIns_Inst_Sbox_15_T11}), .c ({new_AGEMA_signal_6028, new_AGEMA_signal_6027, SubBytesIns_Inst_Sbox_15_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T16_U1 ( .a ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, SubBytesIns_Inst_Sbox_15_T5}), .b ({new_AGEMA_signal_5712, new_AGEMA_signal_5711, SubBytesIns_Inst_Sbox_15_T12}), .c ({new_AGEMA_signal_6030, new_AGEMA_signal_6029, SubBytesIns_Inst_Sbox_15_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T17_U1 ( .a ({new_AGEMA_signal_6024, new_AGEMA_signal_6023, SubBytesIns_Inst_Sbox_15_T9}), .b ({new_AGEMA_signal_6030, new_AGEMA_signal_6029, SubBytesIns_Inst_Sbox_15_T16}), .c ({new_AGEMA_signal_6538, new_AGEMA_signal_6537, SubBytesIns_Inst_Sbox_15_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T18_U1 ( .a ({ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_5714, new_AGEMA_signal_5713, SubBytesIns_Inst_Sbox_15_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T19_U1 ( .a ({new_AGEMA_signal_5708, new_AGEMA_signal_5707, SubBytesIns_Inst_Sbox_15_T7}), .b ({new_AGEMA_signal_5714, new_AGEMA_signal_5713, SubBytesIns_Inst_Sbox_15_T18}), .c ({new_AGEMA_signal_6032, new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_15_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T20_U1 ( .a ({new_AGEMA_signal_5698, new_AGEMA_signal_5697, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_6032, new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_15_T19}), .c ({new_AGEMA_signal_6540, new_AGEMA_signal_6539, SubBytesIns_Inst_Sbox_15_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T21_U1 ( .a ({ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .b ({ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_5716, new_AGEMA_signal_5715, SubBytesIns_Inst_Sbox_15_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T22_U1 ( .a ({new_AGEMA_signal_5708, new_AGEMA_signal_5707, SubBytesIns_Inst_Sbox_15_T7}), .b ({new_AGEMA_signal_5716, new_AGEMA_signal_5715, SubBytesIns_Inst_Sbox_15_T21}), .c ({new_AGEMA_signal_6034, new_AGEMA_signal_6033, SubBytesIns_Inst_Sbox_15_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T23_U1 ( .a ({new_AGEMA_signal_5700, new_AGEMA_signal_5699, SubBytesIns_Inst_Sbox_15_T2}), .b ({new_AGEMA_signal_6034, new_AGEMA_signal_6033, SubBytesIns_Inst_Sbox_15_T22}), .c ({new_AGEMA_signal_6542, new_AGEMA_signal_6541, SubBytesIns_Inst_Sbox_15_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T24_U1 ( .a ({new_AGEMA_signal_5700, new_AGEMA_signal_5699, SubBytesIns_Inst_Sbox_15_T2}), .b ({new_AGEMA_signal_6534, new_AGEMA_signal_6533, SubBytesIns_Inst_Sbox_15_T10}), .c ({new_AGEMA_signal_6900, new_AGEMA_signal_6899, SubBytesIns_Inst_Sbox_15_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T25_U1 ( .a ({new_AGEMA_signal_6540, new_AGEMA_signal_6539, SubBytesIns_Inst_Sbox_15_T20}), .b ({new_AGEMA_signal_6538, new_AGEMA_signal_6537, SubBytesIns_Inst_Sbox_15_T17}), .c ({new_AGEMA_signal_6902, new_AGEMA_signal_6901, SubBytesIns_Inst_Sbox_15_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T26_U1 ( .a ({new_AGEMA_signal_5702, new_AGEMA_signal_5701, SubBytesIns_Inst_Sbox_15_T3}), .b ({new_AGEMA_signal_6030, new_AGEMA_signal_6029, SubBytesIns_Inst_Sbox_15_T16}), .c ({new_AGEMA_signal_6544, new_AGEMA_signal_6543, SubBytesIns_Inst_Sbox_15_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T27_U1 ( .a ({new_AGEMA_signal_5698, new_AGEMA_signal_5697, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_5712, new_AGEMA_signal_5711, SubBytesIns_Inst_Sbox_15_T12}), .c ({new_AGEMA_signal_6036, new_AGEMA_signal_6035, SubBytesIns_Inst_Sbox_15_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T1_U1 ( .a ({new_AGEMA_signal_4810, new_AGEMA_signal_4809, RoundKey[23]}), .b ({new_AGEMA_signal_4792, new_AGEMA_signal_4791, RoundKey[20]}), .c ({new_AGEMA_signal_5318, new_AGEMA_signal_5317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T2_U1 ( .a ({new_AGEMA_signal_4810, new_AGEMA_signal_4809, RoundKey[23]}), .b ({new_AGEMA_signal_4774, new_AGEMA_signal_4773, RoundKey[18]}), .c ({new_AGEMA_signal_5320, new_AGEMA_signal_5319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T3_U1 ( .a ({new_AGEMA_signal_4810, new_AGEMA_signal_4809, RoundKey[23]}), .b ({new_AGEMA_signal_4768, new_AGEMA_signal_4767, RoundKey[17]}), .c ({new_AGEMA_signal_5322, new_AGEMA_signal_5321, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T4_U1 ( .a ({new_AGEMA_signal_4792, new_AGEMA_signal_4791, RoundKey[20]}), .b ({new_AGEMA_signal_4774, new_AGEMA_signal_4773, RoundKey[18]}), .c ({new_AGEMA_signal_5324, new_AGEMA_signal_5323, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T5_U1 ( .a ({new_AGEMA_signal_4780, new_AGEMA_signal_4779, RoundKey[19]}), .b ({new_AGEMA_signal_4768, new_AGEMA_signal_4767, RoundKey[17]}), .c ({new_AGEMA_signal_5326, new_AGEMA_signal_5325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T6_U1 ( .a ({new_AGEMA_signal_5318, new_AGEMA_signal_5317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5326, new_AGEMA_signal_5325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}), .c ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T7_U1 ( .a ({new_AGEMA_signal_4804, new_AGEMA_signal_4803, RoundKey[22]}), .b ({new_AGEMA_signal_4798, new_AGEMA_signal_4797, RoundKey[21]}), .c ({new_AGEMA_signal_5328, new_AGEMA_signal_5327, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T8_U1 ( .a ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, RoundKey[16]}), .b ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .c ({new_AGEMA_signal_6038, new_AGEMA_signal_6037, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T9_U1 ( .a ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, RoundKey[16]}), .b ({new_AGEMA_signal_5328, new_AGEMA_signal_5327, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_5720, new_AGEMA_signal_5719, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T10_U1 ( .a ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_5328, new_AGEMA_signal_5327, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_6040, new_AGEMA_signal_6039, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T11_U1 ( .a ({new_AGEMA_signal_4804, new_AGEMA_signal_4803, RoundKey[22]}), .b ({new_AGEMA_signal_4774, new_AGEMA_signal_4773, RoundKey[18]}), .c ({new_AGEMA_signal_5330, new_AGEMA_signal_5329, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T12_U1 ( .a ({new_AGEMA_signal_4798, new_AGEMA_signal_4797, RoundKey[21]}), .b ({new_AGEMA_signal_4774, new_AGEMA_signal_4773, RoundKey[18]}), .c ({new_AGEMA_signal_5332, new_AGEMA_signal_5331, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T13_U1 ( .a ({new_AGEMA_signal_5322, new_AGEMA_signal_5321, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5324, new_AGEMA_signal_5323, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}), .c ({new_AGEMA_signal_5722, new_AGEMA_signal_5721, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T14_U1 ( .a ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_5330, new_AGEMA_signal_5329, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_6042, new_AGEMA_signal_6041, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T15_U1 ( .a ({new_AGEMA_signal_5326, new_AGEMA_signal_5325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_5330, new_AGEMA_signal_5329, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_5724, new_AGEMA_signal_5723, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T16_U1 ( .a ({new_AGEMA_signal_5326, new_AGEMA_signal_5325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_5332, new_AGEMA_signal_5331, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_5726, new_AGEMA_signal_5725, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T17_U1 ( .a ({new_AGEMA_signal_5720, new_AGEMA_signal_5719, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}), .b ({new_AGEMA_signal_5726, new_AGEMA_signal_5725, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_6044, new_AGEMA_signal_6043, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T18_U1 ( .a ({new_AGEMA_signal_4792, new_AGEMA_signal_4791, RoundKey[20]}), .b ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, RoundKey[16]}), .c ({new_AGEMA_signal_5334, new_AGEMA_signal_5333, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T19_U1 ( .a ({new_AGEMA_signal_5328, new_AGEMA_signal_5327, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_5334, new_AGEMA_signal_5333, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18}), .c ({new_AGEMA_signal_5728, new_AGEMA_signal_5727, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T20_U1 ( .a ({new_AGEMA_signal_5318, new_AGEMA_signal_5317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5728, new_AGEMA_signal_5727, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}), .c ({new_AGEMA_signal_6046, new_AGEMA_signal_6045, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T21_U1 ( .a ({new_AGEMA_signal_4768, new_AGEMA_signal_4767, RoundKey[17]}), .b ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, RoundKey[16]}), .c ({new_AGEMA_signal_5336, new_AGEMA_signal_5335, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T22_U1 ( .a ({new_AGEMA_signal_5328, new_AGEMA_signal_5327, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_5336, new_AGEMA_signal_5335, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21}), .c ({new_AGEMA_signal_5730, new_AGEMA_signal_5729, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T23_U1 ( .a ({new_AGEMA_signal_5320, new_AGEMA_signal_5319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_5730, new_AGEMA_signal_5729, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}), .c ({new_AGEMA_signal_6048, new_AGEMA_signal_6047, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T24_U1 ( .a ({new_AGEMA_signal_5320, new_AGEMA_signal_5319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6040, new_AGEMA_signal_6039, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}), .c ({new_AGEMA_signal_6558, new_AGEMA_signal_6557, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T25_U1 ( .a ({new_AGEMA_signal_6046, new_AGEMA_signal_6045, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_6044, new_AGEMA_signal_6043, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}), .c ({new_AGEMA_signal_6560, new_AGEMA_signal_6559, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T26_U1 ( .a ({new_AGEMA_signal_5322, new_AGEMA_signal_5321, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5726, new_AGEMA_signal_5725, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_6050, new_AGEMA_signal_6049, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T27_U1 ( .a ({new_AGEMA_signal_5318, new_AGEMA_signal_5317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5332, new_AGEMA_signal_5331, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_5732, new_AGEMA_signal_5731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T1_U1 ( .a ({new_AGEMA_signal_4756, new_AGEMA_signal_4755, RoundKey[15]}), .b ({new_AGEMA_signal_4738, new_AGEMA_signal_4737, RoundKey[12]}), .c ({new_AGEMA_signal_5338, new_AGEMA_signal_5337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T2_U1 ( .a ({new_AGEMA_signal_4756, new_AGEMA_signal_4755, RoundKey[15]}), .b ({new_AGEMA_signal_4618, new_AGEMA_signal_4617, RoundKey[10]}), .c ({new_AGEMA_signal_5340, new_AGEMA_signal_5339, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T3_U1 ( .a ({new_AGEMA_signal_4756, new_AGEMA_signal_4755, RoundKey[15]}), .b ({new_AGEMA_signal_5314, new_AGEMA_signal_5313, RoundKey[9]}), .c ({new_AGEMA_signal_5342, new_AGEMA_signal_5341, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T4_U1 ( .a ({new_AGEMA_signal_4738, new_AGEMA_signal_4737, RoundKey[12]}), .b ({new_AGEMA_signal_4618, new_AGEMA_signal_4617, RoundKey[10]}), .c ({new_AGEMA_signal_5344, new_AGEMA_signal_5343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T5_U1 ( .a ({new_AGEMA_signal_4684, new_AGEMA_signal_4683, RoundKey[11]}), .b ({new_AGEMA_signal_5314, new_AGEMA_signal_5313, RoundKey[9]}), .c ({new_AGEMA_signal_5346, new_AGEMA_signal_5345, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T6_U1 ( .a ({new_AGEMA_signal_5338, new_AGEMA_signal_5337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5346, new_AGEMA_signal_5345, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}), .c ({new_AGEMA_signal_5734, new_AGEMA_signal_5733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T7_U1 ( .a ({new_AGEMA_signal_4750, new_AGEMA_signal_4749, RoundKey[14]}), .b ({new_AGEMA_signal_4744, new_AGEMA_signal_4743, RoundKey[13]}), .c ({new_AGEMA_signal_5348, new_AGEMA_signal_5347, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T8_U1 ( .a ({new_AGEMA_signal_5248, new_AGEMA_signal_5247, RoundKey[8]}), .b ({new_AGEMA_signal_5734, new_AGEMA_signal_5733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .c ({new_AGEMA_signal_6064, new_AGEMA_signal_6063, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T9_U1 ( .a ({new_AGEMA_signal_5248, new_AGEMA_signal_5247, RoundKey[8]}), .b ({new_AGEMA_signal_5348, new_AGEMA_signal_5347, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_5736, new_AGEMA_signal_5735, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T10_U1 ( .a ({new_AGEMA_signal_5734, new_AGEMA_signal_5733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_5348, new_AGEMA_signal_5347, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_6066, new_AGEMA_signal_6065, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T11_U1 ( .a ({new_AGEMA_signal_4750, new_AGEMA_signal_4749, RoundKey[14]}), .b ({new_AGEMA_signal_4618, new_AGEMA_signal_4617, RoundKey[10]}), .c ({new_AGEMA_signal_5350, new_AGEMA_signal_5349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T12_U1 ( .a ({new_AGEMA_signal_4744, new_AGEMA_signal_4743, RoundKey[13]}), .b ({new_AGEMA_signal_4618, new_AGEMA_signal_4617, RoundKey[10]}), .c ({new_AGEMA_signal_5352, new_AGEMA_signal_5351, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T13_U1 ( .a ({new_AGEMA_signal_5342, new_AGEMA_signal_5341, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5344, new_AGEMA_signal_5343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}), .c ({new_AGEMA_signal_5738, new_AGEMA_signal_5737, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T14_U1 ( .a ({new_AGEMA_signal_5734, new_AGEMA_signal_5733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_5350, new_AGEMA_signal_5349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_6068, new_AGEMA_signal_6067, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T15_U1 ( .a ({new_AGEMA_signal_5346, new_AGEMA_signal_5345, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_5350, new_AGEMA_signal_5349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_5740, new_AGEMA_signal_5739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T16_U1 ( .a ({new_AGEMA_signal_5346, new_AGEMA_signal_5345, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_5352, new_AGEMA_signal_5351, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T17_U1 ( .a ({new_AGEMA_signal_5736, new_AGEMA_signal_5735, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}), .b ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_6070, new_AGEMA_signal_6069, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T18_U1 ( .a ({new_AGEMA_signal_4738, new_AGEMA_signal_4737, RoundKey[12]}), .b ({new_AGEMA_signal_5248, new_AGEMA_signal_5247, RoundKey[8]}), .c ({new_AGEMA_signal_5354, new_AGEMA_signal_5353, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T19_U1 ( .a ({new_AGEMA_signal_5348, new_AGEMA_signal_5347, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_5354, new_AGEMA_signal_5353, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18}), .c ({new_AGEMA_signal_5744, new_AGEMA_signal_5743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T20_U1 ( .a ({new_AGEMA_signal_5338, new_AGEMA_signal_5337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5744, new_AGEMA_signal_5743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}), .c ({new_AGEMA_signal_6072, new_AGEMA_signal_6071, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T21_U1 ( .a ({new_AGEMA_signal_5314, new_AGEMA_signal_5313, RoundKey[9]}), .b ({new_AGEMA_signal_5248, new_AGEMA_signal_5247, RoundKey[8]}), .c ({new_AGEMA_signal_5356, new_AGEMA_signal_5355, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T22_U1 ( .a ({new_AGEMA_signal_5348, new_AGEMA_signal_5347, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_5356, new_AGEMA_signal_5355, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21}), .c ({new_AGEMA_signal_5746, new_AGEMA_signal_5745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T23_U1 ( .a ({new_AGEMA_signal_5340, new_AGEMA_signal_5339, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_5746, new_AGEMA_signal_5745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}), .c ({new_AGEMA_signal_6074, new_AGEMA_signal_6073, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T24_U1 ( .a ({new_AGEMA_signal_5340, new_AGEMA_signal_5339, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6066, new_AGEMA_signal_6065, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}), .c ({new_AGEMA_signal_6576, new_AGEMA_signal_6575, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T25_U1 ( .a ({new_AGEMA_signal_6072, new_AGEMA_signal_6071, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_6070, new_AGEMA_signal_6069, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}), .c ({new_AGEMA_signal_6578, new_AGEMA_signal_6577, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T26_U1 ( .a ({new_AGEMA_signal_5342, new_AGEMA_signal_5341, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_6076, new_AGEMA_signal_6075, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T27_U1 ( .a ({new_AGEMA_signal_5338, new_AGEMA_signal_5337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5352, new_AGEMA_signal_5351, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T1_U1 ( .a ({new_AGEMA_signal_5182, new_AGEMA_signal_5181, RoundKey[7]}), .b ({new_AGEMA_signal_4984, new_AGEMA_signal_4983, RoundKey[4]}), .c ({new_AGEMA_signal_5358, new_AGEMA_signal_5357, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T2_U1 ( .a ({new_AGEMA_signal_5182, new_AGEMA_signal_5181, RoundKey[7]}), .b ({new_AGEMA_signal_4852, new_AGEMA_signal_4851, RoundKey[2]}), .c ({new_AGEMA_signal_5360, new_AGEMA_signal_5359, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T3_U1 ( .a ({new_AGEMA_signal_5182, new_AGEMA_signal_5181, RoundKey[7]}), .b ({new_AGEMA_signal_4786, new_AGEMA_signal_4785, RoundKey[1]}), .c ({new_AGEMA_signal_5362, new_AGEMA_signal_5361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T4_U1 ( .a ({new_AGEMA_signal_4984, new_AGEMA_signal_4983, RoundKey[4]}), .b ({new_AGEMA_signal_4852, new_AGEMA_signal_4851, RoundKey[2]}), .c ({new_AGEMA_signal_5364, new_AGEMA_signal_5363, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T5_U1 ( .a ({new_AGEMA_signal_4918, new_AGEMA_signal_4917, RoundKey[3]}), .b ({new_AGEMA_signal_4786, new_AGEMA_signal_4785, RoundKey[1]}), .c ({new_AGEMA_signal_5366, new_AGEMA_signal_5365, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T6_U1 ( .a ({new_AGEMA_signal_5358, new_AGEMA_signal_5357, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5366, new_AGEMA_signal_5365, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}), .c ({new_AGEMA_signal_5750, new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T7_U1 ( .a ({new_AGEMA_signal_5116, new_AGEMA_signal_5115, RoundKey[6]}), .b ({new_AGEMA_signal_5050, new_AGEMA_signal_5049, RoundKey[5]}), .c ({new_AGEMA_signal_5368, new_AGEMA_signal_5367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T8_U1 ( .a ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, RoundKey[0]}), .b ({new_AGEMA_signal_5750, new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .c ({new_AGEMA_signal_6090, new_AGEMA_signal_6089, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T9_U1 ( .a ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, RoundKey[0]}), .b ({new_AGEMA_signal_5368, new_AGEMA_signal_5367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_5752, new_AGEMA_signal_5751, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T10_U1 ( .a ({new_AGEMA_signal_5750, new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_5368, new_AGEMA_signal_5367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_6092, new_AGEMA_signal_6091, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T11_U1 ( .a ({new_AGEMA_signal_5116, new_AGEMA_signal_5115, RoundKey[6]}), .b ({new_AGEMA_signal_4852, new_AGEMA_signal_4851, RoundKey[2]}), .c ({new_AGEMA_signal_5370, new_AGEMA_signal_5369, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T12_U1 ( .a ({new_AGEMA_signal_5050, new_AGEMA_signal_5049, RoundKey[5]}), .b ({new_AGEMA_signal_4852, new_AGEMA_signal_4851, RoundKey[2]}), .c ({new_AGEMA_signal_5372, new_AGEMA_signal_5371, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T13_U1 ( .a ({new_AGEMA_signal_5362, new_AGEMA_signal_5361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5364, new_AGEMA_signal_5363, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}), .c ({new_AGEMA_signal_5754, new_AGEMA_signal_5753, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T14_U1 ( .a ({new_AGEMA_signal_5750, new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_5370, new_AGEMA_signal_5369, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_6094, new_AGEMA_signal_6093, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T15_U1 ( .a ({new_AGEMA_signal_5366, new_AGEMA_signal_5365, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_5370, new_AGEMA_signal_5369, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_5756, new_AGEMA_signal_5755, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T16_U1 ( .a ({new_AGEMA_signal_5366, new_AGEMA_signal_5365, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_5372, new_AGEMA_signal_5371, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_5758, new_AGEMA_signal_5757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T17_U1 ( .a ({new_AGEMA_signal_5752, new_AGEMA_signal_5751, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}), .b ({new_AGEMA_signal_5758, new_AGEMA_signal_5757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_6096, new_AGEMA_signal_6095, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T18_U1 ( .a ({new_AGEMA_signal_4984, new_AGEMA_signal_4983, RoundKey[4]}), .b ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, RoundKey[0]}), .c ({new_AGEMA_signal_5374, new_AGEMA_signal_5373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T19_U1 ( .a ({new_AGEMA_signal_5368, new_AGEMA_signal_5367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5374, new_AGEMA_signal_5373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18}), .c ({new_AGEMA_signal_5760, new_AGEMA_signal_5759, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T20_U1 ( .a ({new_AGEMA_signal_5358, new_AGEMA_signal_5357, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5760, new_AGEMA_signal_5759, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}), .c ({new_AGEMA_signal_6098, new_AGEMA_signal_6097, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T21_U1 ( .a ({new_AGEMA_signal_4786, new_AGEMA_signal_4785, RoundKey[1]}), .b ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, RoundKey[0]}), .c ({new_AGEMA_signal_5376, new_AGEMA_signal_5375, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T22_U1 ( .a ({new_AGEMA_signal_5368, new_AGEMA_signal_5367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5376, new_AGEMA_signal_5375, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21}), .c ({new_AGEMA_signal_5762, new_AGEMA_signal_5761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T23_U1 ( .a ({new_AGEMA_signal_5360, new_AGEMA_signal_5359, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_5762, new_AGEMA_signal_5761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}), .c ({new_AGEMA_signal_6100, new_AGEMA_signal_6099, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T24_U1 ( .a ({new_AGEMA_signal_5360, new_AGEMA_signal_5359, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_6092, new_AGEMA_signal_6091, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}), .c ({new_AGEMA_signal_6594, new_AGEMA_signal_6593, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T25_U1 ( .a ({new_AGEMA_signal_6098, new_AGEMA_signal_6097, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_6096, new_AGEMA_signal_6095, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}), .c ({new_AGEMA_signal_6596, new_AGEMA_signal_6595, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T26_U1 ( .a ({new_AGEMA_signal_5362, new_AGEMA_signal_5361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5758, new_AGEMA_signal_5757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_6102, new_AGEMA_signal_6101, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T27_U1 ( .a ({new_AGEMA_signal_5358, new_AGEMA_signal_5357, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5372, new_AGEMA_signal_5371, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_5764, new_AGEMA_signal_5763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T1_U1 ( .a ({new_AGEMA_signal_4864, new_AGEMA_signal_4863, RoundKey[31]}), .b ({new_AGEMA_signal_4840, new_AGEMA_signal_4839, RoundKey[28]}), .c ({new_AGEMA_signal_5378, new_AGEMA_signal_5377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T2_U1 ( .a ({new_AGEMA_signal_4864, new_AGEMA_signal_4863, RoundKey[31]}), .b ({new_AGEMA_signal_4828, new_AGEMA_signal_4827, RoundKey[26]}), .c ({new_AGEMA_signal_5380, new_AGEMA_signal_5379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T3_U1 ( .a ({new_AGEMA_signal_4864, new_AGEMA_signal_4863, RoundKey[31]}), .b ({new_AGEMA_signal_4822, new_AGEMA_signal_4821, RoundKey[25]}), .c ({new_AGEMA_signal_5382, new_AGEMA_signal_5381, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T4_U1 ( .a ({new_AGEMA_signal_4840, new_AGEMA_signal_4839, RoundKey[28]}), .b ({new_AGEMA_signal_4828, new_AGEMA_signal_4827, RoundKey[26]}), .c ({new_AGEMA_signal_5384, new_AGEMA_signal_5383, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T5_U1 ( .a ({new_AGEMA_signal_4834, new_AGEMA_signal_4833, RoundKey[27]}), .b ({new_AGEMA_signal_4822, new_AGEMA_signal_4821, RoundKey[25]}), .c ({new_AGEMA_signal_5386, new_AGEMA_signal_5385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T6_U1 ( .a ({new_AGEMA_signal_5378, new_AGEMA_signal_5377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5386, new_AGEMA_signal_5385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}), .c ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T7_U1 ( .a ({new_AGEMA_signal_4858, new_AGEMA_signal_4857, RoundKey[30]}), .b ({new_AGEMA_signal_4846, new_AGEMA_signal_4845, RoundKey[29]}), .c ({new_AGEMA_signal_5388, new_AGEMA_signal_5387, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T8_U1 ( .a ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, RoundKey[24]}), .b ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .c ({new_AGEMA_signal_6116, new_AGEMA_signal_6115, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T9_U1 ( .a ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, RoundKey[24]}), .b ({new_AGEMA_signal_5388, new_AGEMA_signal_5387, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_5768, new_AGEMA_signal_5767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T10_U1 ( .a ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5388, new_AGEMA_signal_5387, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_6118, new_AGEMA_signal_6117, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T11_U1 ( .a ({new_AGEMA_signal_4858, new_AGEMA_signal_4857, RoundKey[30]}), .b ({new_AGEMA_signal_4828, new_AGEMA_signal_4827, RoundKey[26]}), .c ({new_AGEMA_signal_5390, new_AGEMA_signal_5389, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T12_U1 ( .a ({new_AGEMA_signal_4846, new_AGEMA_signal_4845, RoundKey[29]}), .b ({new_AGEMA_signal_4828, new_AGEMA_signal_4827, RoundKey[26]}), .c ({new_AGEMA_signal_5392, new_AGEMA_signal_5391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T13_U1 ( .a ({new_AGEMA_signal_5382, new_AGEMA_signal_5381, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5384, new_AGEMA_signal_5383, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}), .c ({new_AGEMA_signal_5770, new_AGEMA_signal_5769, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T14_U1 ( .a ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5390, new_AGEMA_signal_5389, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_6120, new_AGEMA_signal_6119, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T15_U1 ( .a ({new_AGEMA_signal_5386, new_AGEMA_signal_5385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5390, new_AGEMA_signal_5389, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_5772, new_AGEMA_signal_5771, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T16_U1 ( .a ({new_AGEMA_signal_5386, new_AGEMA_signal_5385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5392, new_AGEMA_signal_5391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_5774, new_AGEMA_signal_5773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T17_U1 ( .a ({new_AGEMA_signal_5768, new_AGEMA_signal_5767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}), .b ({new_AGEMA_signal_5774, new_AGEMA_signal_5773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_6122, new_AGEMA_signal_6121, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T18_U1 ( .a ({new_AGEMA_signal_4840, new_AGEMA_signal_4839, RoundKey[28]}), .b ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, RoundKey[24]}), .c ({new_AGEMA_signal_5394, new_AGEMA_signal_5393, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T19_U1 ( .a ({new_AGEMA_signal_5388, new_AGEMA_signal_5387, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5394, new_AGEMA_signal_5393, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18}), .c ({new_AGEMA_signal_5776, new_AGEMA_signal_5775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T20_U1 ( .a ({new_AGEMA_signal_5378, new_AGEMA_signal_5377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5776, new_AGEMA_signal_5775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}), .c ({new_AGEMA_signal_6124, new_AGEMA_signal_6123, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T21_U1 ( .a ({new_AGEMA_signal_4822, new_AGEMA_signal_4821, RoundKey[25]}), .b ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, RoundKey[24]}), .c ({new_AGEMA_signal_5396, new_AGEMA_signal_5395, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T22_U1 ( .a ({new_AGEMA_signal_5388, new_AGEMA_signal_5387, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5396, new_AGEMA_signal_5395, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21}), .c ({new_AGEMA_signal_5778, new_AGEMA_signal_5777, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T23_U1 ( .a ({new_AGEMA_signal_5380, new_AGEMA_signal_5379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_5778, new_AGEMA_signal_5777, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}), .c ({new_AGEMA_signal_6126, new_AGEMA_signal_6125, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T24_U1 ( .a ({new_AGEMA_signal_5380, new_AGEMA_signal_5379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_6118, new_AGEMA_signal_6117, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}), .c ({new_AGEMA_signal_6612, new_AGEMA_signal_6611, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T25_U1 ( .a ({new_AGEMA_signal_6124, new_AGEMA_signal_6123, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_6122, new_AGEMA_signal_6121, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}), .c ({new_AGEMA_signal_6614, new_AGEMA_signal_6613, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T26_U1 ( .a ({new_AGEMA_signal_5382, new_AGEMA_signal_5381, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5774, new_AGEMA_signal_5773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_6128, new_AGEMA_signal_6127, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T27_U1 ( .a ({new_AGEMA_signal_5378, new_AGEMA_signal_5377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5392, new_AGEMA_signal_5391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_5780, new_AGEMA_signal_5779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27}) ) ;
    INV_X1 RoundCounterIns_U14 ( .A (RoundCounterIns_n13), .ZN (RoundCounterIns_n1) ) ;
    MUX2_X1 RoundCounterIns_U13 ( .S (RoundCounterIns_n5), .A (RoundCounterIns_n12), .B (RoundCounterIns_n11), .Z (RoundCounterIns_n13) ) ;
    NOR2_X1 RoundCounterIns_U12 ( .A1 (reset), .A2 (RoundCounterIns_n10), .ZN (RoundCounterIns_N8) ) ;
    XNOR2_X1 RoundCounterIns_U11 ( .A (RoundCounter[0]), .B (RoundCounter[1]), .ZN (RoundCounterIns_n10) ) ;
    MUX2_X1 RoundCounterIns_U10 ( .S (RoundCounter[3]), .A (RoundCounterIns_n9), .B (RoundCounterIns_n8), .Z (RoundCounterIns_N10) ) ;
    NAND2_X1 RoundCounterIns_U9 ( .A1 (RoundCounterIns_n12), .A2 (RoundCounterIns_n7), .ZN (RoundCounterIns_n8) ) ;
    NAND2_X1 RoundCounterIns_U8 ( .A1 (RoundCounterIns_n5), .A2 (RoundCounterIns_n2), .ZN (RoundCounterIns_n7) ) ;
    NOR2_X1 RoundCounterIns_U7 ( .A1 (RoundCounterIns_n4), .A2 (RoundCounterIns_N7), .ZN (RoundCounterIns_n12) ) ;
    NOR2_X1 RoundCounterIns_U6 ( .A1 (RoundCounter[1]), .A2 (reset), .ZN (RoundCounterIns_n4) ) ;
    NOR2_X1 RoundCounterIns_U5 ( .A1 (RoundCounterIns_n5), .A2 (RoundCounterIns_n11), .ZN (RoundCounterIns_n9) ) ;
    NAND2_X1 RoundCounterIns_U4 ( .A1 (RoundCounter[1]), .A2 (RoundCounterIns_n3), .ZN (RoundCounterIns_n11) ) ;
    NOR2_X1 RoundCounterIns_U3 ( .A1 (reset), .A2 (RoundCounterIns_n6), .ZN (RoundCounterIns_n3) ) ;
    NOR2_X1 RoundCounterIns_U2 ( .A1 (reset), .A2 (RoundCounter[0]), .ZN (RoundCounterIns_N7) ) ;
    INV_X1 RoundCounterIns_U1 ( .A (reset), .ZN (RoundCounterIns_n2) ) ;
    INV_X1 RoundCounterIns_count_reg_0__U1 ( .A (RoundCounter[0]), .ZN (RoundCounterIns_n6) ) ;
    INV_X1 RoundCounterIns_count_reg_2__U1 ( .A (RoundCounter[2]), .ZN (RoundCounterIns_n5) ) ;
    ClockGatingController #(9) ClockGatingInst ( .clk (clk), .rst (reset), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M1_U1 ( .a ({new_AGEMA_signal_5786, new_AGEMA_signal_5785, SubBytesIns_Inst_Sbox_0_T13}), .b ({new_AGEMA_signal_5782, new_AGEMA_signal_5781, SubBytesIns_Inst_Sbox_0_T6}), .clk (clk), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_6156, new_AGEMA_signal_6155, SubBytesIns_Inst_Sbox_0_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M2_U1 ( .a ({new_AGEMA_signal_6152, new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_0_T23}), .b ({new_AGEMA_signal_6142, new_AGEMA_signal_6141, SubBytesIns_Inst_Sbox_0_T8}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({new_AGEMA_signal_6634, new_AGEMA_signal_6633, SubBytesIns_Inst_Sbox_0_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M3_U1 ( .a ({new_AGEMA_signal_6146, new_AGEMA_signal_6145, SubBytesIns_Inst_Sbox_0_T14}), .b ({new_AGEMA_signal_6156, new_AGEMA_signal_6155, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_6636, new_AGEMA_signal_6635, SubBytesIns_Inst_Sbox_0_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M4_U1 ( .a ({new_AGEMA_signal_5792, new_AGEMA_signal_5791, SubBytesIns_Inst_Sbox_0_T19}), .b ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .clk (clk), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_6158, new_AGEMA_signal_6157, SubBytesIns_Inst_Sbox_0_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M5_U1 ( .a ({new_AGEMA_signal_6158, new_AGEMA_signal_6157, SubBytesIns_Inst_Sbox_0_M4}), .b ({new_AGEMA_signal_6156, new_AGEMA_signal_6155, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_6638, new_AGEMA_signal_6637, SubBytesIns_Inst_Sbox_0_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M6_U1 ( .a ({new_AGEMA_signal_5402, new_AGEMA_signal_5401, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5790, new_AGEMA_signal_5789, SubBytesIns_Inst_Sbox_0_T16}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({new_AGEMA_signal_6160, new_AGEMA_signal_6159, SubBytesIns_Inst_Sbox_0_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M7_U1 ( .a ({new_AGEMA_signal_5794, new_AGEMA_signal_5793, SubBytesIns_Inst_Sbox_0_T22}), .b ({new_AGEMA_signal_5784, new_AGEMA_signal_5783, SubBytesIns_Inst_Sbox_0_T9}), .clk (clk), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_6162, new_AGEMA_signal_6161, SubBytesIns_Inst_Sbox_0_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M8_U1 ( .a ({new_AGEMA_signal_6154, new_AGEMA_signal_6153, SubBytesIns_Inst_Sbox_0_T26}), .b ({new_AGEMA_signal_6160, new_AGEMA_signal_6159, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_6640, new_AGEMA_signal_6639, SubBytesIns_Inst_Sbox_0_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M9_U1 ( .a ({new_AGEMA_signal_6150, new_AGEMA_signal_6149, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_6148, new_AGEMA_signal_6147, SubBytesIns_Inst_Sbox_0_T17}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({new_AGEMA_signal_6642, new_AGEMA_signal_6641, SubBytesIns_Inst_Sbox_0_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M10_U1 ( .a ({new_AGEMA_signal_6642, new_AGEMA_signal_6641, SubBytesIns_Inst_Sbox_0_M9}), .b ({new_AGEMA_signal_6160, new_AGEMA_signal_6159, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_6958, new_AGEMA_signal_6957, SubBytesIns_Inst_Sbox_0_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M11_U1 ( .a ({new_AGEMA_signal_5398, new_AGEMA_signal_5397, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5788, new_AGEMA_signal_5787, SubBytesIns_Inst_Sbox_0_T15}), .clk (clk), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_6164, new_AGEMA_signal_6163, SubBytesIns_Inst_Sbox_0_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M12_U1 ( .a ({new_AGEMA_signal_5404, new_AGEMA_signal_5403, SubBytesIns_Inst_Sbox_0_T4}), .b ({new_AGEMA_signal_5796, new_AGEMA_signal_5795, SubBytesIns_Inst_Sbox_0_T27}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({new_AGEMA_signal_6166, new_AGEMA_signal_6165, SubBytesIns_Inst_Sbox_0_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M13_U1 ( .a ({new_AGEMA_signal_6166, new_AGEMA_signal_6165, SubBytesIns_Inst_Sbox_0_M12}), .b ({new_AGEMA_signal_6164, new_AGEMA_signal_6163, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_6644, new_AGEMA_signal_6643, SubBytesIns_Inst_Sbox_0_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M14_U1 ( .a ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6144, new_AGEMA_signal_6143, SubBytesIns_Inst_Sbox_0_T10}), .clk (clk), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_6646, new_AGEMA_signal_6645, SubBytesIns_Inst_Sbox_0_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M15_U1 ( .a ({new_AGEMA_signal_6646, new_AGEMA_signal_6645, SubBytesIns_Inst_Sbox_0_M14}), .b ({new_AGEMA_signal_6164, new_AGEMA_signal_6163, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_6960, new_AGEMA_signal_6959, SubBytesIns_Inst_Sbox_0_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M16_U1 ( .a ({new_AGEMA_signal_6636, new_AGEMA_signal_6635, SubBytesIns_Inst_Sbox_0_M3}), .b ({new_AGEMA_signal_6634, new_AGEMA_signal_6633, SubBytesIns_Inst_Sbox_0_M2}), .c ({new_AGEMA_signal_6962, new_AGEMA_signal_6961, SubBytesIns_Inst_Sbox_0_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M17_U1 ( .a ({new_AGEMA_signal_6638, new_AGEMA_signal_6637, SubBytesIns_Inst_Sbox_0_M5}), .b ({new_AGEMA_signal_6630, new_AGEMA_signal_6629, SubBytesIns_Inst_Sbox_0_T24}), .c ({new_AGEMA_signal_6964, new_AGEMA_signal_6963, SubBytesIns_Inst_Sbox_0_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M18_U1 ( .a ({new_AGEMA_signal_6640, new_AGEMA_signal_6639, SubBytesIns_Inst_Sbox_0_M8}), .b ({new_AGEMA_signal_6162, new_AGEMA_signal_6161, SubBytesIns_Inst_Sbox_0_M7}), .c ({new_AGEMA_signal_6966, new_AGEMA_signal_6965, SubBytesIns_Inst_Sbox_0_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M19_U1 ( .a ({new_AGEMA_signal_6958, new_AGEMA_signal_6957, SubBytesIns_Inst_Sbox_0_M10}), .b ({new_AGEMA_signal_6960, new_AGEMA_signal_6959, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_7150, new_AGEMA_signal_7149, SubBytesIns_Inst_Sbox_0_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M20_U1 ( .a ({new_AGEMA_signal_6962, new_AGEMA_signal_6961, SubBytesIns_Inst_Sbox_0_M16}), .b ({new_AGEMA_signal_6644, new_AGEMA_signal_6643, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_7152, new_AGEMA_signal_7151, SubBytesIns_Inst_Sbox_0_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M21_U1 ( .a ({new_AGEMA_signal_6964, new_AGEMA_signal_6963, SubBytesIns_Inst_Sbox_0_M17}), .b ({new_AGEMA_signal_6960, new_AGEMA_signal_6959, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_7154, new_AGEMA_signal_7153, SubBytesIns_Inst_Sbox_0_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M22_U1 ( .a ({new_AGEMA_signal_6966, new_AGEMA_signal_6965, SubBytesIns_Inst_Sbox_0_M18}), .b ({new_AGEMA_signal_6644, new_AGEMA_signal_6643, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_7156, new_AGEMA_signal_7155, SubBytesIns_Inst_Sbox_0_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M23_U1 ( .a ({new_AGEMA_signal_7150, new_AGEMA_signal_7149, SubBytesIns_Inst_Sbox_0_M19}), .b ({new_AGEMA_signal_6632, new_AGEMA_signal_6631, SubBytesIns_Inst_Sbox_0_T25}), .c ({new_AGEMA_signal_7310, new_AGEMA_signal_7309, SubBytesIns_Inst_Sbox_0_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M24_U1 ( .a ({new_AGEMA_signal_7156, new_AGEMA_signal_7155, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_7310, new_AGEMA_signal_7309, SubBytesIns_Inst_Sbox_0_M23}), .c ({new_AGEMA_signal_7478, new_AGEMA_signal_7477, SubBytesIns_Inst_Sbox_0_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M27_U1 ( .a ({new_AGEMA_signal_7152, new_AGEMA_signal_7151, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_7154, new_AGEMA_signal_7153, SubBytesIns_Inst_Sbox_0_M21}), .c ({new_AGEMA_signal_7314, new_AGEMA_signal_7313, SubBytesIns_Inst_Sbox_0_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M1_U1 ( .a ({new_AGEMA_signal_5802, new_AGEMA_signal_5801, SubBytesIns_Inst_Sbox_1_T13}), .b ({new_AGEMA_signal_5798, new_AGEMA_signal_5797, SubBytesIns_Inst_Sbox_1_T6}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({new_AGEMA_signal_6182, new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_1_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M2_U1 ( .a ({new_AGEMA_signal_6178, new_AGEMA_signal_6177, SubBytesIns_Inst_Sbox_1_T23}), .b ({new_AGEMA_signal_6168, new_AGEMA_signal_6167, SubBytesIns_Inst_Sbox_1_T8}), .clk (clk), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_6652, new_AGEMA_signal_6651, SubBytesIns_Inst_Sbox_1_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M3_U1 ( .a ({new_AGEMA_signal_6172, new_AGEMA_signal_6171, SubBytesIns_Inst_Sbox_1_T14}), .b ({new_AGEMA_signal_6182, new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_6654, new_AGEMA_signal_6653, SubBytesIns_Inst_Sbox_1_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M4_U1 ( .a ({new_AGEMA_signal_5808, new_AGEMA_signal_5807, SubBytesIns_Inst_Sbox_1_T19}), .b ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({new_AGEMA_signal_6184, new_AGEMA_signal_6183, SubBytesIns_Inst_Sbox_1_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M5_U1 ( .a ({new_AGEMA_signal_6184, new_AGEMA_signal_6183, SubBytesIns_Inst_Sbox_1_M4}), .b ({new_AGEMA_signal_6182, new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_6656, new_AGEMA_signal_6655, SubBytesIns_Inst_Sbox_1_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M6_U1 ( .a ({new_AGEMA_signal_5422, new_AGEMA_signal_5421, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5806, new_AGEMA_signal_5805, SubBytesIns_Inst_Sbox_1_T16}), .clk (clk), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_6186, new_AGEMA_signal_6185, SubBytesIns_Inst_Sbox_1_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M7_U1 ( .a ({new_AGEMA_signal_5810, new_AGEMA_signal_5809, SubBytesIns_Inst_Sbox_1_T22}), .b ({new_AGEMA_signal_5800, new_AGEMA_signal_5799, SubBytesIns_Inst_Sbox_1_T9}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({new_AGEMA_signal_6188, new_AGEMA_signal_6187, SubBytesIns_Inst_Sbox_1_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M8_U1 ( .a ({new_AGEMA_signal_6180, new_AGEMA_signal_6179, SubBytesIns_Inst_Sbox_1_T26}), .b ({new_AGEMA_signal_6186, new_AGEMA_signal_6185, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_6658, new_AGEMA_signal_6657, SubBytesIns_Inst_Sbox_1_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M9_U1 ( .a ({new_AGEMA_signal_6176, new_AGEMA_signal_6175, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_6174, new_AGEMA_signal_6173, SubBytesIns_Inst_Sbox_1_T17}), .clk (clk), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_6660, new_AGEMA_signal_6659, SubBytesIns_Inst_Sbox_1_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M10_U1 ( .a ({new_AGEMA_signal_6660, new_AGEMA_signal_6659, SubBytesIns_Inst_Sbox_1_M9}), .b ({new_AGEMA_signal_6186, new_AGEMA_signal_6185, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_6968, new_AGEMA_signal_6967, SubBytesIns_Inst_Sbox_1_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M11_U1 ( .a ({new_AGEMA_signal_5418, new_AGEMA_signal_5417, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5804, new_AGEMA_signal_5803, SubBytesIns_Inst_Sbox_1_T15}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({new_AGEMA_signal_6190, new_AGEMA_signal_6189, SubBytesIns_Inst_Sbox_1_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M12_U1 ( .a ({new_AGEMA_signal_5424, new_AGEMA_signal_5423, SubBytesIns_Inst_Sbox_1_T4}), .b ({new_AGEMA_signal_5812, new_AGEMA_signal_5811, SubBytesIns_Inst_Sbox_1_T27}), .clk (clk), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_6192, new_AGEMA_signal_6191, SubBytesIns_Inst_Sbox_1_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M13_U1 ( .a ({new_AGEMA_signal_6192, new_AGEMA_signal_6191, SubBytesIns_Inst_Sbox_1_M12}), .b ({new_AGEMA_signal_6190, new_AGEMA_signal_6189, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_6662, new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_1_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M14_U1 ( .a ({new_AGEMA_signal_5420, new_AGEMA_signal_5419, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6170, new_AGEMA_signal_6169, SubBytesIns_Inst_Sbox_1_T10}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({new_AGEMA_signal_6664, new_AGEMA_signal_6663, SubBytesIns_Inst_Sbox_1_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M15_U1 ( .a ({new_AGEMA_signal_6664, new_AGEMA_signal_6663, SubBytesIns_Inst_Sbox_1_M14}), .b ({new_AGEMA_signal_6190, new_AGEMA_signal_6189, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_6970, new_AGEMA_signal_6969, SubBytesIns_Inst_Sbox_1_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M16_U1 ( .a ({new_AGEMA_signal_6654, new_AGEMA_signal_6653, SubBytesIns_Inst_Sbox_1_M3}), .b ({new_AGEMA_signal_6652, new_AGEMA_signal_6651, SubBytesIns_Inst_Sbox_1_M2}), .c ({new_AGEMA_signal_6972, new_AGEMA_signal_6971, SubBytesIns_Inst_Sbox_1_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M17_U1 ( .a ({new_AGEMA_signal_6656, new_AGEMA_signal_6655, SubBytesIns_Inst_Sbox_1_M5}), .b ({new_AGEMA_signal_6648, new_AGEMA_signal_6647, SubBytesIns_Inst_Sbox_1_T24}), .c ({new_AGEMA_signal_6974, new_AGEMA_signal_6973, SubBytesIns_Inst_Sbox_1_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M18_U1 ( .a ({new_AGEMA_signal_6658, new_AGEMA_signal_6657, SubBytesIns_Inst_Sbox_1_M8}), .b ({new_AGEMA_signal_6188, new_AGEMA_signal_6187, SubBytesIns_Inst_Sbox_1_M7}), .c ({new_AGEMA_signal_6976, new_AGEMA_signal_6975, SubBytesIns_Inst_Sbox_1_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M19_U1 ( .a ({new_AGEMA_signal_6968, new_AGEMA_signal_6967, SubBytesIns_Inst_Sbox_1_M10}), .b ({new_AGEMA_signal_6970, new_AGEMA_signal_6969, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_7158, new_AGEMA_signal_7157, SubBytesIns_Inst_Sbox_1_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M20_U1 ( .a ({new_AGEMA_signal_6972, new_AGEMA_signal_6971, SubBytesIns_Inst_Sbox_1_M16}), .b ({new_AGEMA_signal_6662, new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_7160, new_AGEMA_signal_7159, SubBytesIns_Inst_Sbox_1_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M21_U1 ( .a ({new_AGEMA_signal_6974, new_AGEMA_signal_6973, SubBytesIns_Inst_Sbox_1_M17}), .b ({new_AGEMA_signal_6970, new_AGEMA_signal_6969, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_7162, new_AGEMA_signal_7161, SubBytesIns_Inst_Sbox_1_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M22_U1 ( .a ({new_AGEMA_signal_6976, new_AGEMA_signal_6975, SubBytesIns_Inst_Sbox_1_M18}), .b ({new_AGEMA_signal_6662, new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_7164, new_AGEMA_signal_7163, SubBytesIns_Inst_Sbox_1_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M23_U1 ( .a ({new_AGEMA_signal_7158, new_AGEMA_signal_7157, SubBytesIns_Inst_Sbox_1_M19}), .b ({new_AGEMA_signal_6650, new_AGEMA_signal_6649, SubBytesIns_Inst_Sbox_1_T25}), .c ({new_AGEMA_signal_7318, new_AGEMA_signal_7317, SubBytesIns_Inst_Sbox_1_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M24_U1 ( .a ({new_AGEMA_signal_7164, new_AGEMA_signal_7163, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_7318, new_AGEMA_signal_7317, SubBytesIns_Inst_Sbox_1_M23}), .c ({new_AGEMA_signal_7488, new_AGEMA_signal_7487, SubBytesIns_Inst_Sbox_1_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M27_U1 ( .a ({new_AGEMA_signal_7160, new_AGEMA_signal_7159, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_7162, new_AGEMA_signal_7161, SubBytesIns_Inst_Sbox_1_M21}), .c ({new_AGEMA_signal_7322, new_AGEMA_signal_7321, SubBytesIns_Inst_Sbox_1_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M1_U1 ( .a ({new_AGEMA_signal_5818, new_AGEMA_signal_5817, SubBytesIns_Inst_Sbox_2_T13}), .b ({new_AGEMA_signal_5814, new_AGEMA_signal_5813, SubBytesIns_Inst_Sbox_2_T6}), .clk (clk), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_6208, new_AGEMA_signal_6207, SubBytesIns_Inst_Sbox_2_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M2_U1 ( .a ({new_AGEMA_signal_6204, new_AGEMA_signal_6203, SubBytesIns_Inst_Sbox_2_T23}), .b ({new_AGEMA_signal_6194, new_AGEMA_signal_6193, SubBytesIns_Inst_Sbox_2_T8}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({new_AGEMA_signal_6670, new_AGEMA_signal_6669, SubBytesIns_Inst_Sbox_2_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M3_U1 ( .a ({new_AGEMA_signal_6198, new_AGEMA_signal_6197, SubBytesIns_Inst_Sbox_2_T14}), .b ({new_AGEMA_signal_6208, new_AGEMA_signal_6207, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_6672, new_AGEMA_signal_6671, SubBytesIns_Inst_Sbox_2_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M4_U1 ( .a ({new_AGEMA_signal_5824, new_AGEMA_signal_5823, SubBytesIns_Inst_Sbox_2_T19}), .b ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .clk (clk), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_6210, new_AGEMA_signal_6209, SubBytesIns_Inst_Sbox_2_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M5_U1 ( .a ({new_AGEMA_signal_6210, new_AGEMA_signal_6209, SubBytesIns_Inst_Sbox_2_M4}), .b ({new_AGEMA_signal_6208, new_AGEMA_signal_6207, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_6674, new_AGEMA_signal_6673, SubBytesIns_Inst_Sbox_2_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M6_U1 ( .a ({new_AGEMA_signal_5442, new_AGEMA_signal_5441, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_2_T16}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({new_AGEMA_signal_6212, new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_2_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M7_U1 ( .a ({new_AGEMA_signal_5826, new_AGEMA_signal_5825, SubBytesIns_Inst_Sbox_2_T22}), .b ({new_AGEMA_signal_5816, new_AGEMA_signal_5815, SubBytesIns_Inst_Sbox_2_T9}), .clk (clk), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_6214, new_AGEMA_signal_6213, SubBytesIns_Inst_Sbox_2_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M8_U1 ( .a ({new_AGEMA_signal_6206, new_AGEMA_signal_6205, SubBytesIns_Inst_Sbox_2_T26}), .b ({new_AGEMA_signal_6212, new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_6676, new_AGEMA_signal_6675, SubBytesIns_Inst_Sbox_2_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M9_U1 ( .a ({new_AGEMA_signal_6202, new_AGEMA_signal_6201, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_6200, new_AGEMA_signal_6199, SubBytesIns_Inst_Sbox_2_T17}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({new_AGEMA_signal_6678, new_AGEMA_signal_6677, SubBytesIns_Inst_Sbox_2_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M10_U1 ( .a ({new_AGEMA_signal_6678, new_AGEMA_signal_6677, SubBytesIns_Inst_Sbox_2_M9}), .b ({new_AGEMA_signal_6212, new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_6978, new_AGEMA_signal_6977, SubBytesIns_Inst_Sbox_2_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M11_U1 ( .a ({new_AGEMA_signal_5438, new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5820, new_AGEMA_signal_5819, SubBytesIns_Inst_Sbox_2_T15}), .clk (clk), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_6216, new_AGEMA_signal_6215, SubBytesIns_Inst_Sbox_2_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M12_U1 ( .a ({new_AGEMA_signal_5444, new_AGEMA_signal_5443, SubBytesIns_Inst_Sbox_2_T4}), .b ({new_AGEMA_signal_5828, new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_2_T27}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({new_AGEMA_signal_6218, new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_2_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M13_U1 ( .a ({new_AGEMA_signal_6218, new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_2_M12}), .b ({new_AGEMA_signal_6216, new_AGEMA_signal_6215, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_6680, new_AGEMA_signal_6679, SubBytesIns_Inst_Sbox_2_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M14_U1 ( .a ({new_AGEMA_signal_5440, new_AGEMA_signal_5439, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_6196, new_AGEMA_signal_6195, SubBytesIns_Inst_Sbox_2_T10}), .clk (clk), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_6682, new_AGEMA_signal_6681, SubBytesIns_Inst_Sbox_2_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M15_U1 ( .a ({new_AGEMA_signal_6682, new_AGEMA_signal_6681, SubBytesIns_Inst_Sbox_2_M14}), .b ({new_AGEMA_signal_6216, new_AGEMA_signal_6215, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_6980, new_AGEMA_signal_6979, SubBytesIns_Inst_Sbox_2_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M16_U1 ( .a ({new_AGEMA_signal_6672, new_AGEMA_signal_6671, SubBytesIns_Inst_Sbox_2_M3}), .b ({new_AGEMA_signal_6670, new_AGEMA_signal_6669, SubBytesIns_Inst_Sbox_2_M2}), .c ({new_AGEMA_signal_6982, new_AGEMA_signal_6981, SubBytesIns_Inst_Sbox_2_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M17_U1 ( .a ({new_AGEMA_signal_6674, new_AGEMA_signal_6673, SubBytesIns_Inst_Sbox_2_M5}), .b ({new_AGEMA_signal_6666, new_AGEMA_signal_6665, SubBytesIns_Inst_Sbox_2_T24}), .c ({new_AGEMA_signal_6984, new_AGEMA_signal_6983, SubBytesIns_Inst_Sbox_2_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M18_U1 ( .a ({new_AGEMA_signal_6676, new_AGEMA_signal_6675, SubBytesIns_Inst_Sbox_2_M8}), .b ({new_AGEMA_signal_6214, new_AGEMA_signal_6213, SubBytesIns_Inst_Sbox_2_M7}), .c ({new_AGEMA_signal_6986, new_AGEMA_signal_6985, SubBytesIns_Inst_Sbox_2_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M19_U1 ( .a ({new_AGEMA_signal_6978, new_AGEMA_signal_6977, SubBytesIns_Inst_Sbox_2_M10}), .b ({new_AGEMA_signal_6980, new_AGEMA_signal_6979, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_7166, new_AGEMA_signal_7165, SubBytesIns_Inst_Sbox_2_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M20_U1 ( .a ({new_AGEMA_signal_6982, new_AGEMA_signal_6981, SubBytesIns_Inst_Sbox_2_M16}), .b ({new_AGEMA_signal_6680, new_AGEMA_signal_6679, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_7168, new_AGEMA_signal_7167, SubBytesIns_Inst_Sbox_2_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M21_U1 ( .a ({new_AGEMA_signal_6984, new_AGEMA_signal_6983, SubBytesIns_Inst_Sbox_2_M17}), .b ({new_AGEMA_signal_6980, new_AGEMA_signal_6979, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_7170, new_AGEMA_signal_7169, SubBytesIns_Inst_Sbox_2_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M22_U1 ( .a ({new_AGEMA_signal_6986, new_AGEMA_signal_6985, SubBytesIns_Inst_Sbox_2_M18}), .b ({new_AGEMA_signal_6680, new_AGEMA_signal_6679, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_7172, new_AGEMA_signal_7171, SubBytesIns_Inst_Sbox_2_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M23_U1 ( .a ({new_AGEMA_signal_7166, new_AGEMA_signal_7165, SubBytesIns_Inst_Sbox_2_M19}), .b ({new_AGEMA_signal_6668, new_AGEMA_signal_6667, SubBytesIns_Inst_Sbox_2_T25}), .c ({new_AGEMA_signal_7326, new_AGEMA_signal_7325, SubBytesIns_Inst_Sbox_2_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M24_U1 ( .a ({new_AGEMA_signal_7172, new_AGEMA_signal_7171, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_7326, new_AGEMA_signal_7325, SubBytesIns_Inst_Sbox_2_M23}), .c ({new_AGEMA_signal_7498, new_AGEMA_signal_7497, SubBytesIns_Inst_Sbox_2_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M27_U1 ( .a ({new_AGEMA_signal_7168, new_AGEMA_signal_7167, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_7170, new_AGEMA_signal_7169, SubBytesIns_Inst_Sbox_2_M21}), .c ({new_AGEMA_signal_7330, new_AGEMA_signal_7329, SubBytesIns_Inst_Sbox_2_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M1_U1 ( .a ({new_AGEMA_signal_5834, new_AGEMA_signal_5833, SubBytesIns_Inst_Sbox_3_T13}), .b ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, SubBytesIns_Inst_Sbox_3_T6}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({new_AGEMA_signal_6234, new_AGEMA_signal_6233, SubBytesIns_Inst_Sbox_3_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M2_U1 ( .a ({new_AGEMA_signal_6230, new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_3_T23}), .b ({new_AGEMA_signal_6220, new_AGEMA_signal_6219, SubBytesIns_Inst_Sbox_3_T8}), .clk (clk), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_6688, new_AGEMA_signal_6687, SubBytesIns_Inst_Sbox_3_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M3_U1 ( .a ({new_AGEMA_signal_6224, new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_3_T14}), .b ({new_AGEMA_signal_6234, new_AGEMA_signal_6233, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_6690, new_AGEMA_signal_6689, SubBytesIns_Inst_Sbox_3_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M4_U1 ( .a ({new_AGEMA_signal_5840, new_AGEMA_signal_5839, SubBytesIns_Inst_Sbox_3_T19}), .b ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({new_AGEMA_signal_6236, new_AGEMA_signal_6235, SubBytesIns_Inst_Sbox_3_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M5_U1 ( .a ({new_AGEMA_signal_6236, new_AGEMA_signal_6235, SubBytesIns_Inst_Sbox_3_M4}), .b ({new_AGEMA_signal_6234, new_AGEMA_signal_6233, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_6692, new_AGEMA_signal_6691, SubBytesIns_Inst_Sbox_3_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M6_U1 ( .a ({new_AGEMA_signal_5462, new_AGEMA_signal_5461, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, SubBytesIns_Inst_Sbox_3_T16}), .clk (clk), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_6238, new_AGEMA_signal_6237, SubBytesIns_Inst_Sbox_3_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M7_U1 ( .a ({new_AGEMA_signal_5842, new_AGEMA_signal_5841, SubBytesIns_Inst_Sbox_3_T22}), .b ({new_AGEMA_signal_5832, new_AGEMA_signal_5831, SubBytesIns_Inst_Sbox_3_T9}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({new_AGEMA_signal_6240, new_AGEMA_signal_6239, SubBytesIns_Inst_Sbox_3_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M8_U1 ( .a ({new_AGEMA_signal_6232, new_AGEMA_signal_6231, SubBytesIns_Inst_Sbox_3_T26}), .b ({new_AGEMA_signal_6238, new_AGEMA_signal_6237, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_6694, new_AGEMA_signal_6693, SubBytesIns_Inst_Sbox_3_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M9_U1 ( .a ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_6226, new_AGEMA_signal_6225, SubBytesIns_Inst_Sbox_3_T17}), .clk (clk), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_6696, new_AGEMA_signal_6695, SubBytesIns_Inst_Sbox_3_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M10_U1 ( .a ({new_AGEMA_signal_6696, new_AGEMA_signal_6695, SubBytesIns_Inst_Sbox_3_M9}), .b ({new_AGEMA_signal_6238, new_AGEMA_signal_6237, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_6988, new_AGEMA_signal_6987, SubBytesIns_Inst_Sbox_3_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M11_U1 ( .a ({new_AGEMA_signal_5458, new_AGEMA_signal_5457, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5836, new_AGEMA_signal_5835, SubBytesIns_Inst_Sbox_3_T15}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({new_AGEMA_signal_6242, new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_3_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M12_U1 ( .a ({new_AGEMA_signal_5464, new_AGEMA_signal_5463, SubBytesIns_Inst_Sbox_3_T4}), .b ({new_AGEMA_signal_5844, new_AGEMA_signal_5843, SubBytesIns_Inst_Sbox_3_T27}), .clk (clk), .r ({Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_6244, new_AGEMA_signal_6243, SubBytesIns_Inst_Sbox_3_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M13_U1 ( .a ({new_AGEMA_signal_6244, new_AGEMA_signal_6243, SubBytesIns_Inst_Sbox_3_M12}), .b ({new_AGEMA_signal_6242, new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_6698, new_AGEMA_signal_6697, SubBytesIns_Inst_Sbox_3_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M14_U1 ( .a ({new_AGEMA_signal_5460, new_AGEMA_signal_5459, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_6222, new_AGEMA_signal_6221, SubBytesIns_Inst_Sbox_3_T10}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105]}), .c ({new_AGEMA_signal_6700, new_AGEMA_signal_6699, SubBytesIns_Inst_Sbox_3_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M15_U1 ( .a ({new_AGEMA_signal_6700, new_AGEMA_signal_6699, SubBytesIns_Inst_Sbox_3_M14}), .b ({new_AGEMA_signal_6242, new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_6990, new_AGEMA_signal_6989, SubBytesIns_Inst_Sbox_3_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M16_U1 ( .a ({new_AGEMA_signal_6690, new_AGEMA_signal_6689, SubBytesIns_Inst_Sbox_3_M3}), .b ({new_AGEMA_signal_6688, new_AGEMA_signal_6687, SubBytesIns_Inst_Sbox_3_M2}), .c ({new_AGEMA_signal_6992, new_AGEMA_signal_6991, SubBytesIns_Inst_Sbox_3_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M17_U1 ( .a ({new_AGEMA_signal_6692, new_AGEMA_signal_6691, SubBytesIns_Inst_Sbox_3_M5}), .b ({new_AGEMA_signal_6684, new_AGEMA_signal_6683, SubBytesIns_Inst_Sbox_3_T24}), .c ({new_AGEMA_signal_6994, new_AGEMA_signal_6993, SubBytesIns_Inst_Sbox_3_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M18_U1 ( .a ({new_AGEMA_signal_6694, new_AGEMA_signal_6693, SubBytesIns_Inst_Sbox_3_M8}), .b ({new_AGEMA_signal_6240, new_AGEMA_signal_6239, SubBytesIns_Inst_Sbox_3_M7}), .c ({new_AGEMA_signal_6996, new_AGEMA_signal_6995, SubBytesIns_Inst_Sbox_3_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M19_U1 ( .a ({new_AGEMA_signal_6988, new_AGEMA_signal_6987, SubBytesIns_Inst_Sbox_3_M10}), .b ({new_AGEMA_signal_6990, new_AGEMA_signal_6989, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_7174, new_AGEMA_signal_7173, SubBytesIns_Inst_Sbox_3_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M20_U1 ( .a ({new_AGEMA_signal_6992, new_AGEMA_signal_6991, SubBytesIns_Inst_Sbox_3_M16}), .b ({new_AGEMA_signal_6698, new_AGEMA_signal_6697, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_7176, new_AGEMA_signal_7175, SubBytesIns_Inst_Sbox_3_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M21_U1 ( .a ({new_AGEMA_signal_6994, new_AGEMA_signal_6993, SubBytesIns_Inst_Sbox_3_M17}), .b ({new_AGEMA_signal_6990, new_AGEMA_signal_6989, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_7178, new_AGEMA_signal_7177, SubBytesIns_Inst_Sbox_3_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M22_U1 ( .a ({new_AGEMA_signal_6996, new_AGEMA_signal_6995, SubBytesIns_Inst_Sbox_3_M18}), .b ({new_AGEMA_signal_6698, new_AGEMA_signal_6697, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_7180, new_AGEMA_signal_7179, SubBytesIns_Inst_Sbox_3_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M23_U1 ( .a ({new_AGEMA_signal_7174, new_AGEMA_signal_7173, SubBytesIns_Inst_Sbox_3_M19}), .b ({new_AGEMA_signal_6686, new_AGEMA_signal_6685, SubBytesIns_Inst_Sbox_3_T25}), .c ({new_AGEMA_signal_7334, new_AGEMA_signal_7333, SubBytesIns_Inst_Sbox_3_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M24_U1 ( .a ({new_AGEMA_signal_7180, new_AGEMA_signal_7179, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_7334, new_AGEMA_signal_7333, SubBytesIns_Inst_Sbox_3_M23}), .c ({new_AGEMA_signal_7508, new_AGEMA_signal_7507, SubBytesIns_Inst_Sbox_3_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M27_U1 ( .a ({new_AGEMA_signal_7176, new_AGEMA_signal_7175, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_7178, new_AGEMA_signal_7177, SubBytesIns_Inst_Sbox_3_M21}), .c ({new_AGEMA_signal_7338, new_AGEMA_signal_7337, SubBytesIns_Inst_Sbox_3_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M1_U1 ( .a ({new_AGEMA_signal_5850, new_AGEMA_signal_5849, SubBytesIns_Inst_Sbox_4_T13}), .b ({new_AGEMA_signal_5846, new_AGEMA_signal_5845, SubBytesIns_Inst_Sbox_4_T6}), .clk (clk), .r ({Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_6260, new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_4_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M2_U1 ( .a ({new_AGEMA_signal_6256, new_AGEMA_signal_6255, SubBytesIns_Inst_Sbox_4_T23}), .b ({new_AGEMA_signal_6246, new_AGEMA_signal_6245, SubBytesIns_Inst_Sbox_4_T8}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111]}), .c ({new_AGEMA_signal_6706, new_AGEMA_signal_6705, SubBytesIns_Inst_Sbox_4_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M3_U1 ( .a ({new_AGEMA_signal_6250, new_AGEMA_signal_6249, SubBytesIns_Inst_Sbox_4_T14}), .b ({new_AGEMA_signal_6260, new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_4_M1}), .c ({new_AGEMA_signal_6708, new_AGEMA_signal_6707, SubBytesIns_Inst_Sbox_4_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M4_U1 ( .a ({new_AGEMA_signal_5856, new_AGEMA_signal_5855, SubBytesIns_Inst_Sbox_4_T19}), .b ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .clk (clk), .r ({Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_6262, new_AGEMA_signal_6261, SubBytesIns_Inst_Sbox_4_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M5_U1 ( .a ({new_AGEMA_signal_6262, new_AGEMA_signal_6261, SubBytesIns_Inst_Sbox_4_M4}), .b ({new_AGEMA_signal_6260, new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_4_M1}), .c ({new_AGEMA_signal_6710, new_AGEMA_signal_6709, SubBytesIns_Inst_Sbox_4_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M6_U1 ( .a ({new_AGEMA_signal_5482, new_AGEMA_signal_5481, SubBytesIns_Inst_Sbox_4_T3}), .b ({new_AGEMA_signal_5854, new_AGEMA_signal_5853, SubBytesIns_Inst_Sbox_4_T16}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117]}), .c ({new_AGEMA_signal_6264, new_AGEMA_signal_6263, SubBytesIns_Inst_Sbox_4_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M7_U1 ( .a ({new_AGEMA_signal_5858, new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_4_T22}), .b ({new_AGEMA_signal_5848, new_AGEMA_signal_5847, SubBytesIns_Inst_Sbox_4_T9}), .clk (clk), .r ({Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_6266, new_AGEMA_signal_6265, SubBytesIns_Inst_Sbox_4_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M8_U1 ( .a ({new_AGEMA_signal_6258, new_AGEMA_signal_6257, SubBytesIns_Inst_Sbox_4_T26}), .b ({new_AGEMA_signal_6264, new_AGEMA_signal_6263, SubBytesIns_Inst_Sbox_4_M6}), .c ({new_AGEMA_signal_6712, new_AGEMA_signal_6711, SubBytesIns_Inst_Sbox_4_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M9_U1 ( .a ({new_AGEMA_signal_6254, new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_4_T20}), .b ({new_AGEMA_signal_6252, new_AGEMA_signal_6251, SubBytesIns_Inst_Sbox_4_T17}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123]}), .c ({new_AGEMA_signal_6714, new_AGEMA_signal_6713, SubBytesIns_Inst_Sbox_4_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M10_U1 ( .a ({new_AGEMA_signal_6714, new_AGEMA_signal_6713, SubBytesIns_Inst_Sbox_4_M9}), .b ({new_AGEMA_signal_6264, new_AGEMA_signal_6263, SubBytesIns_Inst_Sbox_4_M6}), .c ({new_AGEMA_signal_6998, new_AGEMA_signal_6997, SubBytesIns_Inst_Sbox_4_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M11_U1 ( .a ({new_AGEMA_signal_5478, new_AGEMA_signal_5477, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5852, new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_4_T15}), .clk (clk), .r ({Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_6268, new_AGEMA_signal_6267, SubBytesIns_Inst_Sbox_4_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M12_U1 ( .a ({new_AGEMA_signal_5484, new_AGEMA_signal_5483, SubBytesIns_Inst_Sbox_4_T4}), .b ({new_AGEMA_signal_5860, new_AGEMA_signal_5859, SubBytesIns_Inst_Sbox_4_T27}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129]}), .c ({new_AGEMA_signal_6270, new_AGEMA_signal_6269, SubBytesIns_Inst_Sbox_4_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M13_U1 ( .a ({new_AGEMA_signal_6270, new_AGEMA_signal_6269, SubBytesIns_Inst_Sbox_4_M12}), .b ({new_AGEMA_signal_6268, new_AGEMA_signal_6267, SubBytesIns_Inst_Sbox_4_M11}), .c ({new_AGEMA_signal_6716, new_AGEMA_signal_6715, SubBytesIns_Inst_Sbox_4_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M14_U1 ( .a ({new_AGEMA_signal_5480, new_AGEMA_signal_5479, SubBytesIns_Inst_Sbox_4_T2}), .b ({new_AGEMA_signal_6248, new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_4_T10}), .clk (clk), .r ({Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_6718, new_AGEMA_signal_6717, SubBytesIns_Inst_Sbox_4_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M15_U1 ( .a ({new_AGEMA_signal_6718, new_AGEMA_signal_6717, SubBytesIns_Inst_Sbox_4_M14}), .b ({new_AGEMA_signal_6268, new_AGEMA_signal_6267, SubBytesIns_Inst_Sbox_4_M11}), .c ({new_AGEMA_signal_7000, new_AGEMA_signal_6999, SubBytesIns_Inst_Sbox_4_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M16_U1 ( .a ({new_AGEMA_signal_6708, new_AGEMA_signal_6707, SubBytesIns_Inst_Sbox_4_M3}), .b ({new_AGEMA_signal_6706, new_AGEMA_signal_6705, SubBytesIns_Inst_Sbox_4_M2}), .c ({new_AGEMA_signal_7002, new_AGEMA_signal_7001, SubBytesIns_Inst_Sbox_4_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M17_U1 ( .a ({new_AGEMA_signal_6710, new_AGEMA_signal_6709, SubBytesIns_Inst_Sbox_4_M5}), .b ({new_AGEMA_signal_6702, new_AGEMA_signal_6701, SubBytesIns_Inst_Sbox_4_T24}), .c ({new_AGEMA_signal_7004, new_AGEMA_signal_7003, SubBytesIns_Inst_Sbox_4_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M18_U1 ( .a ({new_AGEMA_signal_6712, new_AGEMA_signal_6711, SubBytesIns_Inst_Sbox_4_M8}), .b ({new_AGEMA_signal_6266, new_AGEMA_signal_6265, SubBytesIns_Inst_Sbox_4_M7}), .c ({new_AGEMA_signal_7006, new_AGEMA_signal_7005, SubBytesIns_Inst_Sbox_4_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M19_U1 ( .a ({new_AGEMA_signal_6998, new_AGEMA_signal_6997, SubBytesIns_Inst_Sbox_4_M10}), .b ({new_AGEMA_signal_7000, new_AGEMA_signal_6999, SubBytesIns_Inst_Sbox_4_M15}), .c ({new_AGEMA_signal_7182, new_AGEMA_signal_7181, SubBytesIns_Inst_Sbox_4_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M20_U1 ( .a ({new_AGEMA_signal_7002, new_AGEMA_signal_7001, SubBytesIns_Inst_Sbox_4_M16}), .b ({new_AGEMA_signal_6716, new_AGEMA_signal_6715, SubBytesIns_Inst_Sbox_4_M13}), .c ({new_AGEMA_signal_7184, new_AGEMA_signal_7183, SubBytesIns_Inst_Sbox_4_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M21_U1 ( .a ({new_AGEMA_signal_7004, new_AGEMA_signal_7003, SubBytesIns_Inst_Sbox_4_M17}), .b ({new_AGEMA_signal_7000, new_AGEMA_signal_6999, SubBytesIns_Inst_Sbox_4_M15}), .c ({new_AGEMA_signal_7186, new_AGEMA_signal_7185, SubBytesIns_Inst_Sbox_4_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M22_U1 ( .a ({new_AGEMA_signal_7006, new_AGEMA_signal_7005, SubBytesIns_Inst_Sbox_4_M18}), .b ({new_AGEMA_signal_6716, new_AGEMA_signal_6715, SubBytesIns_Inst_Sbox_4_M13}), .c ({new_AGEMA_signal_7188, new_AGEMA_signal_7187, SubBytesIns_Inst_Sbox_4_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M23_U1 ( .a ({new_AGEMA_signal_7182, new_AGEMA_signal_7181, SubBytesIns_Inst_Sbox_4_M19}), .b ({new_AGEMA_signal_6704, new_AGEMA_signal_6703, SubBytesIns_Inst_Sbox_4_T25}), .c ({new_AGEMA_signal_7342, new_AGEMA_signal_7341, SubBytesIns_Inst_Sbox_4_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M24_U1 ( .a ({new_AGEMA_signal_7188, new_AGEMA_signal_7187, SubBytesIns_Inst_Sbox_4_M22}), .b ({new_AGEMA_signal_7342, new_AGEMA_signal_7341, SubBytesIns_Inst_Sbox_4_M23}), .c ({new_AGEMA_signal_7518, new_AGEMA_signal_7517, SubBytesIns_Inst_Sbox_4_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M27_U1 ( .a ({new_AGEMA_signal_7184, new_AGEMA_signal_7183, SubBytesIns_Inst_Sbox_4_M20}), .b ({new_AGEMA_signal_7186, new_AGEMA_signal_7185, SubBytesIns_Inst_Sbox_4_M21}), .c ({new_AGEMA_signal_7346, new_AGEMA_signal_7345, SubBytesIns_Inst_Sbox_4_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M1_U1 ( .a ({new_AGEMA_signal_5866, new_AGEMA_signal_5865, SubBytesIns_Inst_Sbox_5_T13}), .b ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, SubBytesIns_Inst_Sbox_5_T6}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135]}), .c ({new_AGEMA_signal_6286, new_AGEMA_signal_6285, SubBytesIns_Inst_Sbox_5_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M2_U1 ( .a ({new_AGEMA_signal_6282, new_AGEMA_signal_6281, SubBytesIns_Inst_Sbox_5_T23}), .b ({new_AGEMA_signal_6272, new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_5_T8}), .clk (clk), .r ({Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_6724, new_AGEMA_signal_6723, SubBytesIns_Inst_Sbox_5_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M3_U1 ( .a ({new_AGEMA_signal_6276, new_AGEMA_signal_6275, SubBytesIns_Inst_Sbox_5_T14}), .b ({new_AGEMA_signal_6286, new_AGEMA_signal_6285, SubBytesIns_Inst_Sbox_5_M1}), .c ({new_AGEMA_signal_6726, new_AGEMA_signal_6725, SubBytesIns_Inst_Sbox_5_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M4_U1 ( .a ({new_AGEMA_signal_5872, new_AGEMA_signal_5871, SubBytesIns_Inst_Sbox_5_T19}), .b ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141]}), .c ({new_AGEMA_signal_6288, new_AGEMA_signal_6287, SubBytesIns_Inst_Sbox_5_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M5_U1 ( .a ({new_AGEMA_signal_6288, new_AGEMA_signal_6287, SubBytesIns_Inst_Sbox_5_M4}), .b ({new_AGEMA_signal_6286, new_AGEMA_signal_6285, SubBytesIns_Inst_Sbox_5_M1}), .c ({new_AGEMA_signal_6728, new_AGEMA_signal_6727, SubBytesIns_Inst_Sbox_5_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M6_U1 ( .a ({new_AGEMA_signal_5502, new_AGEMA_signal_5501, SubBytesIns_Inst_Sbox_5_T3}), .b ({new_AGEMA_signal_5870, new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_5_T16}), .clk (clk), .r ({Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_6290, new_AGEMA_signal_6289, SubBytesIns_Inst_Sbox_5_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M7_U1 ( .a ({new_AGEMA_signal_5874, new_AGEMA_signal_5873, SubBytesIns_Inst_Sbox_5_T22}), .b ({new_AGEMA_signal_5864, new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_5_T9}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147]}), .c ({new_AGEMA_signal_6292, new_AGEMA_signal_6291, SubBytesIns_Inst_Sbox_5_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M8_U1 ( .a ({new_AGEMA_signal_6284, new_AGEMA_signal_6283, SubBytesIns_Inst_Sbox_5_T26}), .b ({new_AGEMA_signal_6290, new_AGEMA_signal_6289, SubBytesIns_Inst_Sbox_5_M6}), .c ({new_AGEMA_signal_6730, new_AGEMA_signal_6729, SubBytesIns_Inst_Sbox_5_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M9_U1 ( .a ({new_AGEMA_signal_6280, new_AGEMA_signal_6279, SubBytesIns_Inst_Sbox_5_T20}), .b ({new_AGEMA_signal_6278, new_AGEMA_signal_6277, SubBytesIns_Inst_Sbox_5_T17}), .clk (clk), .r ({Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_6732, new_AGEMA_signal_6731, SubBytesIns_Inst_Sbox_5_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M10_U1 ( .a ({new_AGEMA_signal_6732, new_AGEMA_signal_6731, SubBytesIns_Inst_Sbox_5_M9}), .b ({new_AGEMA_signal_6290, new_AGEMA_signal_6289, SubBytesIns_Inst_Sbox_5_M6}), .c ({new_AGEMA_signal_7008, new_AGEMA_signal_7007, SubBytesIns_Inst_Sbox_5_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M11_U1 ( .a ({new_AGEMA_signal_5498, new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, SubBytesIns_Inst_Sbox_5_T15}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153]}), .c ({new_AGEMA_signal_6294, new_AGEMA_signal_6293, SubBytesIns_Inst_Sbox_5_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M12_U1 ( .a ({new_AGEMA_signal_5504, new_AGEMA_signal_5503, SubBytesIns_Inst_Sbox_5_T4}), .b ({new_AGEMA_signal_5876, new_AGEMA_signal_5875, SubBytesIns_Inst_Sbox_5_T27}), .clk (clk), .r ({Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_6296, new_AGEMA_signal_6295, SubBytesIns_Inst_Sbox_5_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M13_U1 ( .a ({new_AGEMA_signal_6296, new_AGEMA_signal_6295, SubBytesIns_Inst_Sbox_5_M12}), .b ({new_AGEMA_signal_6294, new_AGEMA_signal_6293, SubBytesIns_Inst_Sbox_5_M11}), .c ({new_AGEMA_signal_6734, new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_5_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M14_U1 ( .a ({new_AGEMA_signal_5500, new_AGEMA_signal_5499, SubBytesIns_Inst_Sbox_5_T2}), .b ({new_AGEMA_signal_6274, new_AGEMA_signal_6273, SubBytesIns_Inst_Sbox_5_T10}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159]}), .c ({new_AGEMA_signal_6736, new_AGEMA_signal_6735, SubBytesIns_Inst_Sbox_5_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M15_U1 ( .a ({new_AGEMA_signal_6736, new_AGEMA_signal_6735, SubBytesIns_Inst_Sbox_5_M14}), .b ({new_AGEMA_signal_6294, new_AGEMA_signal_6293, SubBytesIns_Inst_Sbox_5_M11}), .c ({new_AGEMA_signal_7010, new_AGEMA_signal_7009, SubBytesIns_Inst_Sbox_5_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M16_U1 ( .a ({new_AGEMA_signal_6726, new_AGEMA_signal_6725, SubBytesIns_Inst_Sbox_5_M3}), .b ({new_AGEMA_signal_6724, new_AGEMA_signal_6723, SubBytesIns_Inst_Sbox_5_M2}), .c ({new_AGEMA_signal_7012, new_AGEMA_signal_7011, SubBytesIns_Inst_Sbox_5_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M17_U1 ( .a ({new_AGEMA_signal_6728, new_AGEMA_signal_6727, SubBytesIns_Inst_Sbox_5_M5}), .b ({new_AGEMA_signal_6720, new_AGEMA_signal_6719, SubBytesIns_Inst_Sbox_5_T24}), .c ({new_AGEMA_signal_7014, new_AGEMA_signal_7013, SubBytesIns_Inst_Sbox_5_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M18_U1 ( .a ({new_AGEMA_signal_6730, new_AGEMA_signal_6729, SubBytesIns_Inst_Sbox_5_M8}), .b ({new_AGEMA_signal_6292, new_AGEMA_signal_6291, SubBytesIns_Inst_Sbox_5_M7}), .c ({new_AGEMA_signal_7016, new_AGEMA_signal_7015, SubBytesIns_Inst_Sbox_5_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M19_U1 ( .a ({new_AGEMA_signal_7008, new_AGEMA_signal_7007, SubBytesIns_Inst_Sbox_5_M10}), .b ({new_AGEMA_signal_7010, new_AGEMA_signal_7009, SubBytesIns_Inst_Sbox_5_M15}), .c ({new_AGEMA_signal_7190, new_AGEMA_signal_7189, SubBytesIns_Inst_Sbox_5_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M20_U1 ( .a ({new_AGEMA_signal_7012, new_AGEMA_signal_7011, SubBytesIns_Inst_Sbox_5_M16}), .b ({new_AGEMA_signal_6734, new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_5_M13}), .c ({new_AGEMA_signal_7192, new_AGEMA_signal_7191, SubBytesIns_Inst_Sbox_5_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M21_U1 ( .a ({new_AGEMA_signal_7014, new_AGEMA_signal_7013, SubBytesIns_Inst_Sbox_5_M17}), .b ({new_AGEMA_signal_7010, new_AGEMA_signal_7009, SubBytesIns_Inst_Sbox_5_M15}), .c ({new_AGEMA_signal_7194, new_AGEMA_signal_7193, SubBytesIns_Inst_Sbox_5_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M22_U1 ( .a ({new_AGEMA_signal_7016, new_AGEMA_signal_7015, SubBytesIns_Inst_Sbox_5_M18}), .b ({new_AGEMA_signal_6734, new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_5_M13}), .c ({new_AGEMA_signal_7196, new_AGEMA_signal_7195, SubBytesIns_Inst_Sbox_5_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M23_U1 ( .a ({new_AGEMA_signal_7190, new_AGEMA_signal_7189, SubBytesIns_Inst_Sbox_5_M19}), .b ({new_AGEMA_signal_6722, new_AGEMA_signal_6721, SubBytesIns_Inst_Sbox_5_T25}), .c ({new_AGEMA_signal_7350, new_AGEMA_signal_7349, SubBytesIns_Inst_Sbox_5_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M24_U1 ( .a ({new_AGEMA_signal_7196, new_AGEMA_signal_7195, SubBytesIns_Inst_Sbox_5_M22}), .b ({new_AGEMA_signal_7350, new_AGEMA_signal_7349, SubBytesIns_Inst_Sbox_5_M23}), .c ({new_AGEMA_signal_7528, new_AGEMA_signal_7527, SubBytesIns_Inst_Sbox_5_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M27_U1 ( .a ({new_AGEMA_signal_7192, new_AGEMA_signal_7191, SubBytesIns_Inst_Sbox_5_M20}), .b ({new_AGEMA_signal_7194, new_AGEMA_signal_7193, SubBytesIns_Inst_Sbox_5_M21}), .c ({new_AGEMA_signal_7354, new_AGEMA_signal_7353, SubBytesIns_Inst_Sbox_5_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M1_U1 ( .a ({new_AGEMA_signal_5882, new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_6_T13}), .b ({new_AGEMA_signal_5878, new_AGEMA_signal_5877, SubBytesIns_Inst_Sbox_6_T6}), .clk (clk), .r ({Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_6312, new_AGEMA_signal_6311, SubBytesIns_Inst_Sbox_6_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M2_U1 ( .a ({new_AGEMA_signal_6308, new_AGEMA_signal_6307, SubBytesIns_Inst_Sbox_6_T23}), .b ({new_AGEMA_signal_6298, new_AGEMA_signal_6297, SubBytesIns_Inst_Sbox_6_T8}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165]}), .c ({new_AGEMA_signal_6742, new_AGEMA_signal_6741, SubBytesIns_Inst_Sbox_6_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M3_U1 ( .a ({new_AGEMA_signal_6302, new_AGEMA_signal_6301, SubBytesIns_Inst_Sbox_6_T14}), .b ({new_AGEMA_signal_6312, new_AGEMA_signal_6311, SubBytesIns_Inst_Sbox_6_M1}), .c ({new_AGEMA_signal_6744, new_AGEMA_signal_6743, SubBytesIns_Inst_Sbox_6_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M4_U1 ( .a ({new_AGEMA_signal_5888, new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_6_T19}), .b ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .clk (clk), .r ({Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_6314, new_AGEMA_signal_6313, SubBytesIns_Inst_Sbox_6_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M5_U1 ( .a ({new_AGEMA_signal_6314, new_AGEMA_signal_6313, SubBytesIns_Inst_Sbox_6_M4}), .b ({new_AGEMA_signal_6312, new_AGEMA_signal_6311, SubBytesIns_Inst_Sbox_6_M1}), .c ({new_AGEMA_signal_6746, new_AGEMA_signal_6745, SubBytesIns_Inst_Sbox_6_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M6_U1 ( .a ({new_AGEMA_signal_5522, new_AGEMA_signal_5521, SubBytesIns_Inst_Sbox_6_T3}), .b ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, SubBytesIns_Inst_Sbox_6_T16}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171]}), .c ({new_AGEMA_signal_6316, new_AGEMA_signal_6315, SubBytesIns_Inst_Sbox_6_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M7_U1 ( .a ({new_AGEMA_signal_5890, new_AGEMA_signal_5889, SubBytesIns_Inst_Sbox_6_T22}), .b ({new_AGEMA_signal_5880, new_AGEMA_signal_5879, SubBytesIns_Inst_Sbox_6_T9}), .clk (clk), .r ({Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_6318, new_AGEMA_signal_6317, SubBytesIns_Inst_Sbox_6_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M8_U1 ( .a ({new_AGEMA_signal_6310, new_AGEMA_signal_6309, SubBytesIns_Inst_Sbox_6_T26}), .b ({new_AGEMA_signal_6316, new_AGEMA_signal_6315, SubBytesIns_Inst_Sbox_6_M6}), .c ({new_AGEMA_signal_6748, new_AGEMA_signal_6747, SubBytesIns_Inst_Sbox_6_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M9_U1 ( .a ({new_AGEMA_signal_6306, new_AGEMA_signal_6305, SubBytesIns_Inst_Sbox_6_T20}), .b ({new_AGEMA_signal_6304, new_AGEMA_signal_6303, SubBytesIns_Inst_Sbox_6_T17}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177]}), .c ({new_AGEMA_signal_6750, new_AGEMA_signal_6749, SubBytesIns_Inst_Sbox_6_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M10_U1 ( .a ({new_AGEMA_signal_6750, new_AGEMA_signal_6749, SubBytesIns_Inst_Sbox_6_M9}), .b ({new_AGEMA_signal_6316, new_AGEMA_signal_6315, SubBytesIns_Inst_Sbox_6_M6}), .c ({new_AGEMA_signal_7018, new_AGEMA_signal_7017, SubBytesIns_Inst_Sbox_6_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M11_U1 ( .a ({new_AGEMA_signal_5518, new_AGEMA_signal_5517, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_5884, new_AGEMA_signal_5883, SubBytesIns_Inst_Sbox_6_T15}), .clk (clk), .r ({Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_6320, new_AGEMA_signal_6319, SubBytesIns_Inst_Sbox_6_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M12_U1 ( .a ({new_AGEMA_signal_5524, new_AGEMA_signal_5523, SubBytesIns_Inst_Sbox_6_T4}), .b ({new_AGEMA_signal_5892, new_AGEMA_signal_5891, SubBytesIns_Inst_Sbox_6_T27}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183]}), .c ({new_AGEMA_signal_6322, new_AGEMA_signal_6321, SubBytesIns_Inst_Sbox_6_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M13_U1 ( .a ({new_AGEMA_signal_6322, new_AGEMA_signal_6321, SubBytesIns_Inst_Sbox_6_M12}), .b ({new_AGEMA_signal_6320, new_AGEMA_signal_6319, SubBytesIns_Inst_Sbox_6_M11}), .c ({new_AGEMA_signal_6752, new_AGEMA_signal_6751, SubBytesIns_Inst_Sbox_6_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M14_U1 ( .a ({new_AGEMA_signal_5520, new_AGEMA_signal_5519, SubBytesIns_Inst_Sbox_6_T2}), .b ({new_AGEMA_signal_6300, new_AGEMA_signal_6299, SubBytesIns_Inst_Sbox_6_T10}), .clk (clk), .r ({Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_6754, new_AGEMA_signal_6753, SubBytesIns_Inst_Sbox_6_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M15_U1 ( .a ({new_AGEMA_signal_6754, new_AGEMA_signal_6753, SubBytesIns_Inst_Sbox_6_M14}), .b ({new_AGEMA_signal_6320, new_AGEMA_signal_6319, SubBytesIns_Inst_Sbox_6_M11}), .c ({new_AGEMA_signal_7020, new_AGEMA_signal_7019, SubBytesIns_Inst_Sbox_6_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M16_U1 ( .a ({new_AGEMA_signal_6744, new_AGEMA_signal_6743, SubBytesIns_Inst_Sbox_6_M3}), .b ({new_AGEMA_signal_6742, new_AGEMA_signal_6741, SubBytesIns_Inst_Sbox_6_M2}), .c ({new_AGEMA_signal_7022, new_AGEMA_signal_7021, SubBytesIns_Inst_Sbox_6_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M17_U1 ( .a ({new_AGEMA_signal_6746, new_AGEMA_signal_6745, SubBytesIns_Inst_Sbox_6_M5}), .b ({new_AGEMA_signal_6738, new_AGEMA_signal_6737, SubBytesIns_Inst_Sbox_6_T24}), .c ({new_AGEMA_signal_7024, new_AGEMA_signal_7023, SubBytesIns_Inst_Sbox_6_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M18_U1 ( .a ({new_AGEMA_signal_6748, new_AGEMA_signal_6747, SubBytesIns_Inst_Sbox_6_M8}), .b ({new_AGEMA_signal_6318, new_AGEMA_signal_6317, SubBytesIns_Inst_Sbox_6_M7}), .c ({new_AGEMA_signal_7026, new_AGEMA_signal_7025, SubBytesIns_Inst_Sbox_6_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M19_U1 ( .a ({new_AGEMA_signal_7018, new_AGEMA_signal_7017, SubBytesIns_Inst_Sbox_6_M10}), .b ({new_AGEMA_signal_7020, new_AGEMA_signal_7019, SubBytesIns_Inst_Sbox_6_M15}), .c ({new_AGEMA_signal_7198, new_AGEMA_signal_7197, SubBytesIns_Inst_Sbox_6_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M20_U1 ( .a ({new_AGEMA_signal_7022, new_AGEMA_signal_7021, SubBytesIns_Inst_Sbox_6_M16}), .b ({new_AGEMA_signal_6752, new_AGEMA_signal_6751, SubBytesIns_Inst_Sbox_6_M13}), .c ({new_AGEMA_signal_7200, new_AGEMA_signal_7199, SubBytesIns_Inst_Sbox_6_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M21_U1 ( .a ({new_AGEMA_signal_7024, new_AGEMA_signal_7023, SubBytesIns_Inst_Sbox_6_M17}), .b ({new_AGEMA_signal_7020, new_AGEMA_signal_7019, SubBytesIns_Inst_Sbox_6_M15}), .c ({new_AGEMA_signal_7202, new_AGEMA_signal_7201, SubBytesIns_Inst_Sbox_6_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M22_U1 ( .a ({new_AGEMA_signal_7026, new_AGEMA_signal_7025, SubBytesIns_Inst_Sbox_6_M18}), .b ({new_AGEMA_signal_6752, new_AGEMA_signal_6751, SubBytesIns_Inst_Sbox_6_M13}), .c ({new_AGEMA_signal_7204, new_AGEMA_signal_7203, SubBytesIns_Inst_Sbox_6_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M23_U1 ( .a ({new_AGEMA_signal_7198, new_AGEMA_signal_7197, SubBytesIns_Inst_Sbox_6_M19}), .b ({new_AGEMA_signal_6740, new_AGEMA_signal_6739, SubBytesIns_Inst_Sbox_6_T25}), .c ({new_AGEMA_signal_7358, new_AGEMA_signal_7357, SubBytesIns_Inst_Sbox_6_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M24_U1 ( .a ({new_AGEMA_signal_7204, new_AGEMA_signal_7203, SubBytesIns_Inst_Sbox_6_M22}), .b ({new_AGEMA_signal_7358, new_AGEMA_signal_7357, SubBytesIns_Inst_Sbox_6_M23}), .c ({new_AGEMA_signal_7538, new_AGEMA_signal_7537, SubBytesIns_Inst_Sbox_6_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M27_U1 ( .a ({new_AGEMA_signal_7200, new_AGEMA_signal_7199, SubBytesIns_Inst_Sbox_6_M20}), .b ({new_AGEMA_signal_7202, new_AGEMA_signal_7201, SubBytesIns_Inst_Sbox_6_M21}), .c ({new_AGEMA_signal_7362, new_AGEMA_signal_7361, SubBytesIns_Inst_Sbox_6_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M1_U1 ( .a ({new_AGEMA_signal_5898, new_AGEMA_signal_5897, SubBytesIns_Inst_Sbox_7_T13}), .b ({new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_7_T6}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189]}), .c ({new_AGEMA_signal_6338, new_AGEMA_signal_6337, SubBytesIns_Inst_Sbox_7_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M2_U1 ( .a ({new_AGEMA_signal_6334, new_AGEMA_signal_6333, SubBytesIns_Inst_Sbox_7_T23}), .b ({new_AGEMA_signal_6324, new_AGEMA_signal_6323, SubBytesIns_Inst_Sbox_7_T8}), .clk (clk), .r ({Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_6760, new_AGEMA_signal_6759, SubBytesIns_Inst_Sbox_7_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M3_U1 ( .a ({new_AGEMA_signal_6328, new_AGEMA_signal_6327, SubBytesIns_Inst_Sbox_7_T14}), .b ({new_AGEMA_signal_6338, new_AGEMA_signal_6337, SubBytesIns_Inst_Sbox_7_M1}), .c ({new_AGEMA_signal_6762, new_AGEMA_signal_6761, SubBytesIns_Inst_Sbox_7_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M4_U1 ( .a ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, SubBytesIns_Inst_Sbox_7_T19}), .b ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195]}), .c ({new_AGEMA_signal_6340, new_AGEMA_signal_6339, SubBytesIns_Inst_Sbox_7_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M5_U1 ( .a ({new_AGEMA_signal_6340, new_AGEMA_signal_6339, SubBytesIns_Inst_Sbox_7_M4}), .b ({new_AGEMA_signal_6338, new_AGEMA_signal_6337, SubBytesIns_Inst_Sbox_7_M1}), .c ({new_AGEMA_signal_6764, new_AGEMA_signal_6763, SubBytesIns_Inst_Sbox_7_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M6_U1 ( .a ({new_AGEMA_signal_5542, new_AGEMA_signal_5541, SubBytesIns_Inst_Sbox_7_T3}), .b ({new_AGEMA_signal_5902, new_AGEMA_signal_5901, SubBytesIns_Inst_Sbox_7_T16}), .clk (clk), .r ({Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_6342, new_AGEMA_signal_6341, SubBytesIns_Inst_Sbox_7_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M7_U1 ( .a ({new_AGEMA_signal_5906, new_AGEMA_signal_5905, SubBytesIns_Inst_Sbox_7_T22}), .b ({new_AGEMA_signal_5896, new_AGEMA_signal_5895, SubBytesIns_Inst_Sbox_7_T9}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201]}), .c ({new_AGEMA_signal_6344, new_AGEMA_signal_6343, SubBytesIns_Inst_Sbox_7_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M8_U1 ( .a ({new_AGEMA_signal_6336, new_AGEMA_signal_6335, SubBytesIns_Inst_Sbox_7_T26}), .b ({new_AGEMA_signal_6342, new_AGEMA_signal_6341, SubBytesIns_Inst_Sbox_7_M6}), .c ({new_AGEMA_signal_6766, new_AGEMA_signal_6765, SubBytesIns_Inst_Sbox_7_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M9_U1 ( .a ({new_AGEMA_signal_6332, new_AGEMA_signal_6331, SubBytesIns_Inst_Sbox_7_T20}), .b ({new_AGEMA_signal_6330, new_AGEMA_signal_6329, SubBytesIns_Inst_Sbox_7_T17}), .clk (clk), .r ({Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_6768, new_AGEMA_signal_6767, SubBytesIns_Inst_Sbox_7_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M10_U1 ( .a ({new_AGEMA_signal_6768, new_AGEMA_signal_6767, SubBytesIns_Inst_Sbox_7_M9}), .b ({new_AGEMA_signal_6342, new_AGEMA_signal_6341, SubBytesIns_Inst_Sbox_7_M6}), .c ({new_AGEMA_signal_7028, new_AGEMA_signal_7027, SubBytesIns_Inst_Sbox_7_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M11_U1 ( .a ({new_AGEMA_signal_5538, new_AGEMA_signal_5537, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_5900, new_AGEMA_signal_5899, SubBytesIns_Inst_Sbox_7_T15}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207]}), .c ({new_AGEMA_signal_6346, new_AGEMA_signal_6345, SubBytesIns_Inst_Sbox_7_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M12_U1 ( .a ({new_AGEMA_signal_5544, new_AGEMA_signal_5543, SubBytesIns_Inst_Sbox_7_T4}), .b ({new_AGEMA_signal_5908, new_AGEMA_signal_5907, SubBytesIns_Inst_Sbox_7_T27}), .clk (clk), .r ({Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_6348, new_AGEMA_signal_6347, SubBytesIns_Inst_Sbox_7_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M13_U1 ( .a ({new_AGEMA_signal_6348, new_AGEMA_signal_6347, SubBytesIns_Inst_Sbox_7_M12}), .b ({new_AGEMA_signal_6346, new_AGEMA_signal_6345, SubBytesIns_Inst_Sbox_7_M11}), .c ({new_AGEMA_signal_6770, new_AGEMA_signal_6769, SubBytesIns_Inst_Sbox_7_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M14_U1 ( .a ({new_AGEMA_signal_5540, new_AGEMA_signal_5539, SubBytesIns_Inst_Sbox_7_T2}), .b ({new_AGEMA_signal_6326, new_AGEMA_signal_6325, SubBytesIns_Inst_Sbox_7_T10}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213]}), .c ({new_AGEMA_signal_6772, new_AGEMA_signal_6771, SubBytesIns_Inst_Sbox_7_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M15_U1 ( .a ({new_AGEMA_signal_6772, new_AGEMA_signal_6771, SubBytesIns_Inst_Sbox_7_M14}), .b ({new_AGEMA_signal_6346, new_AGEMA_signal_6345, SubBytesIns_Inst_Sbox_7_M11}), .c ({new_AGEMA_signal_7030, new_AGEMA_signal_7029, SubBytesIns_Inst_Sbox_7_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M16_U1 ( .a ({new_AGEMA_signal_6762, new_AGEMA_signal_6761, SubBytesIns_Inst_Sbox_7_M3}), .b ({new_AGEMA_signal_6760, new_AGEMA_signal_6759, SubBytesIns_Inst_Sbox_7_M2}), .c ({new_AGEMA_signal_7032, new_AGEMA_signal_7031, SubBytesIns_Inst_Sbox_7_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M17_U1 ( .a ({new_AGEMA_signal_6764, new_AGEMA_signal_6763, SubBytesIns_Inst_Sbox_7_M5}), .b ({new_AGEMA_signal_6756, new_AGEMA_signal_6755, SubBytesIns_Inst_Sbox_7_T24}), .c ({new_AGEMA_signal_7034, new_AGEMA_signal_7033, SubBytesIns_Inst_Sbox_7_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M18_U1 ( .a ({new_AGEMA_signal_6766, new_AGEMA_signal_6765, SubBytesIns_Inst_Sbox_7_M8}), .b ({new_AGEMA_signal_6344, new_AGEMA_signal_6343, SubBytesIns_Inst_Sbox_7_M7}), .c ({new_AGEMA_signal_7036, new_AGEMA_signal_7035, SubBytesIns_Inst_Sbox_7_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M19_U1 ( .a ({new_AGEMA_signal_7028, new_AGEMA_signal_7027, SubBytesIns_Inst_Sbox_7_M10}), .b ({new_AGEMA_signal_7030, new_AGEMA_signal_7029, SubBytesIns_Inst_Sbox_7_M15}), .c ({new_AGEMA_signal_7206, new_AGEMA_signal_7205, SubBytesIns_Inst_Sbox_7_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M20_U1 ( .a ({new_AGEMA_signal_7032, new_AGEMA_signal_7031, SubBytesIns_Inst_Sbox_7_M16}), .b ({new_AGEMA_signal_6770, new_AGEMA_signal_6769, SubBytesIns_Inst_Sbox_7_M13}), .c ({new_AGEMA_signal_7208, new_AGEMA_signal_7207, SubBytesIns_Inst_Sbox_7_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M21_U1 ( .a ({new_AGEMA_signal_7034, new_AGEMA_signal_7033, SubBytesIns_Inst_Sbox_7_M17}), .b ({new_AGEMA_signal_7030, new_AGEMA_signal_7029, SubBytesIns_Inst_Sbox_7_M15}), .c ({new_AGEMA_signal_7210, new_AGEMA_signal_7209, SubBytesIns_Inst_Sbox_7_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M22_U1 ( .a ({new_AGEMA_signal_7036, new_AGEMA_signal_7035, SubBytesIns_Inst_Sbox_7_M18}), .b ({new_AGEMA_signal_6770, new_AGEMA_signal_6769, SubBytesIns_Inst_Sbox_7_M13}), .c ({new_AGEMA_signal_7212, new_AGEMA_signal_7211, SubBytesIns_Inst_Sbox_7_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M23_U1 ( .a ({new_AGEMA_signal_7206, new_AGEMA_signal_7205, SubBytesIns_Inst_Sbox_7_M19}), .b ({new_AGEMA_signal_6758, new_AGEMA_signal_6757, SubBytesIns_Inst_Sbox_7_T25}), .c ({new_AGEMA_signal_7366, new_AGEMA_signal_7365, SubBytesIns_Inst_Sbox_7_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M24_U1 ( .a ({new_AGEMA_signal_7212, new_AGEMA_signal_7211, SubBytesIns_Inst_Sbox_7_M22}), .b ({new_AGEMA_signal_7366, new_AGEMA_signal_7365, SubBytesIns_Inst_Sbox_7_M23}), .c ({new_AGEMA_signal_7548, new_AGEMA_signal_7547, SubBytesIns_Inst_Sbox_7_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M27_U1 ( .a ({new_AGEMA_signal_7208, new_AGEMA_signal_7207, SubBytesIns_Inst_Sbox_7_M20}), .b ({new_AGEMA_signal_7210, new_AGEMA_signal_7209, SubBytesIns_Inst_Sbox_7_M21}), .c ({new_AGEMA_signal_7370, new_AGEMA_signal_7369, SubBytesIns_Inst_Sbox_7_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M1_U1 ( .a ({new_AGEMA_signal_5914, new_AGEMA_signal_5913, SubBytesIns_Inst_Sbox_8_T13}), .b ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, SubBytesIns_Inst_Sbox_8_T6}), .clk (clk), .r ({Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_6364, new_AGEMA_signal_6363, SubBytesIns_Inst_Sbox_8_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M2_U1 ( .a ({new_AGEMA_signal_6360, new_AGEMA_signal_6359, SubBytesIns_Inst_Sbox_8_T23}), .b ({new_AGEMA_signal_6350, new_AGEMA_signal_6349, SubBytesIns_Inst_Sbox_8_T8}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219]}), .c ({new_AGEMA_signal_6778, new_AGEMA_signal_6777, SubBytesIns_Inst_Sbox_8_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M3_U1 ( .a ({new_AGEMA_signal_6354, new_AGEMA_signal_6353, SubBytesIns_Inst_Sbox_8_T14}), .b ({new_AGEMA_signal_6364, new_AGEMA_signal_6363, SubBytesIns_Inst_Sbox_8_M1}), .c ({new_AGEMA_signal_6780, new_AGEMA_signal_6779, SubBytesIns_Inst_Sbox_8_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M4_U1 ( .a ({new_AGEMA_signal_5920, new_AGEMA_signal_5919, SubBytesIns_Inst_Sbox_8_T19}), .b ({ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .clk (clk), .r ({Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_6366, new_AGEMA_signal_6365, SubBytesIns_Inst_Sbox_8_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M5_U1 ( .a ({new_AGEMA_signal_6366, new_AGEMA_signal_6365, SubBytesIns_Inst_Sbox_8_M4}), .b ({new_AGEMA_signal_6364, new_AGEMA_signal_6363, SubBytesIns_Inst_Sbox_8_M1}), .c ({new_AGEMA_signal_6782, new_AGEMA_signal_6781, SubBytesIns_Inst_Sbox_8_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M6_U1 ( .a ({new_AGEMA_signal_5562, new_AGEMA_signal_5561, SubBytesIns_Inst_Sbox_8_T3}), .b ({new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesIns_Inst_Sbox_8_T16}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225]}), .c ({new_AGEMA_signal_6368, new_AGEMA_signal_6367, SubBytesIns_Inst_Sbox_8_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M7_U1 ( .a ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, SubBytesIns_Inst_Sbox_8_T22}), .b ({new_AGEMA_signal_5912, new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_8_T9}), .clk (clk), .r ({Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_6370, new_AGEMA_signal_6369, SubBytesIns_Inst_Sbox_8_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M8_U1 ( .a ({new_AGEMA_signal_6362, new_AGEMA_signal_6361, SubBytesIns_Inst_Sbox_8_T26}), .b ({new_AGEMA_signal_6368, new_AGEMA_signal_6367, SubBytesIns_Inst_Sbox_8_M6}), .c ({new_AGEMA_signal_6784, new_AGEMA_signal_6783, SubBytesIns_Inst_Sbox_8_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M9_U1 ( .a ({new_AGEMA_signal_6358, new_AGEMA_signal_6357, SubBytesIns_Inst_Sbox_8_T20}), .b ({new_AGEMA_signal_6356, new_AGEMA_signal_6355, SubBytesIns_Inst_Sbox_8_T17}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231]}), .c ({new_AGEMA_signal_6786, new_AGEMA_signal_6785, SubBytesIns_Inst_Sbox_8_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M10_U1 ( .a ({new_AGEMA_signal_6786, new_AGEMA_signal_6785, SubBytesIns_Inst_Sbox_8_M9}), .b ({new_AGEMA_signal_6368, new_AGEMA_signal_6367, SubBytesIns_Inst_Sbox_8_M6}), .c ({new_AGEMA_signal_7038, new_AGEMA_signal_7037, SubBytesIns_Inst_Sbox_8_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M11_U1 ( .a ({new_AGEMA_signal_5558, new_AGEMA_signal_5557, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, SubBytesIns_Inst_Sbox_8_T15}), .clk (clk), .r ({Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_6372, new_AGEMA_signal_6371, SubBytesIns_Inst_Sbox_8_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M12_U1 ( .a ({new_AGEMA_signal_5564, new_AGEMA_signal_5563, SubBytesIns_Inst_Sbox_8_T4}), .b ({new_AGEMA_signal_5924, new_AGEMA_signal_5923, SubBytesIns_Inst_Sbox_8_T27}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237]}), .c ({new_AGEMA_signal_6374, new_AGEMA_signal_6373, SubBytesIns_Inst_Sbox_8_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M13_U1 ( .a ({new_AGEMA_signal_6374, new_AGEMA_signal_6373, SubBytesIns_Inst_Sbox_8_M12}), .b ({new_AGEMA_signal_6372, new_AGEMA_signal_6371, SubBytesIns_Inst_Sbox_8_M11}), .c ({new_AGEMA_signal_6788, new_AGEMA_signal_6787, SubBytesIns_Inst_Sbox_8_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M14_U1 ( .a ({new_AGEMA_signal_5560, new_AGEMA_signal_5559, SubBytesIns_Inst_Sbox_8_T2}), .b ({new_AGEMA_signal_6352, new_AGEMA_signal_6351, SubBytesIns_Inst_Sbox_8_T10}), .clk (clk), .r ({Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_6790, new_AGEMA_signal_6789, SubBytesIns_Inst_Sbox_8_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M15_U1 ( .a ({new_AGEMA_signal_6790, new_AGEMA_signal_6789, SubBytesIns_Inst_Sbox_8_M14}), .b ({new_AGEMA_signal_6372, new_AGEMA_signal_6371, SubBytesIns_Inst_Sbox_8_M11}), .c ({new_AGEMA_signal_7040, new_AGEMA_signal_7039, SubBytesIns_Inst_Sbox_8_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M16_U1 ( .a ({new_AGEMA_signal_6780, new_AGEMA_signal_6779, SubBytesIns_Inst_Sbox_8_M3}), .b ({new_AGEMA_signal_6778, new_AGEMA_signal_6777, SubBytesIns_Inst_Sbox_8_M2}), .c ({new_AGEMA_signal_7042, new_AGEMA_signal_7041, SubBytesIns_Inst_Sbox_8_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M17_U1 ( .a ({new_AGEMA_signal_6782, new_AGEMA_signal_6781, SubBytesIns_Inst_Sbox_8_M5}), .b ({new_AGEMA_signal_6774, new_AGEMA_signal_6773, SubBytesIns_Inst_Sbox_8_T24}), .c ({new_AGEMA_signal_7044, new_AGEMA_signal_7043, SubBytesIns_Inst_Sbox_8_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M18_U1 ( .a ({new_AGEMA_signal_6784, new_AGEMA_signal_6783, SubBytesIns_Inst_Sbox_8_M8}), .b ({new_AGEMA_signal_6370, new_AGEMA_signal_6369, SubBytesIns_Inst_Sbox_8_M7}), .c ({new_AGEMA_signal_7046, new_AGEMA_signal_7045, SubBytesIns_Inst_Sbox_8_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M19_U1 ( .a ({new_AGEMA_signal_7038, new_AGEMA_signal_7037, SubBytesIns_Inst_Sbox_8_M10}), .b ({new_AGEMA_signal_7040, new_AGEMA_signal_7039, SubBytesIns_Inst_Sbox_8_M15}), .c ({new_AGEMA_signal_7214, new_AGEMA_signal_7213, SubBytesIns_Inst_Sbox_8_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M20_U1 ( .a ({new_AGEMA_signal_7042, new_AGEMA_signal_7041, SubBytesIns_Inst_Sbox_8_M16}), .b ({new_AGEMA_signal_6788, new_AGEMA_signal_6787, SubBytesIns_Inst_Sbox_8_M13}), .c ({new_AGEMA_signal_7216, new_AGEMA_signal_7215, SubBytesIns_Inst_Sbox_8_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M21_U1 ( .a ({new_AGEMA_signal_7044, new_AGEMA_signal_7043, SubBytesIns_Inst_Sbox_8_M17}), .b ({new_AGEMA_signal_7040, new_AGEMA_signal_7039, SubBytesIns_Inst_Sbox_8_M15}), .c ({new_AGEMA_signal_7218, new_AGEMA_signal_7217, SubBytesIns_Inst_Sbox_8_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M22_U1 ( .a ({new_AGEMA_signal_7046, new_AGEMA_signal_7045, SubBytesIns_Inst_Sbox_8_M18}), .b ({new_AGEMA_signal_6788, new_AGEMA_signal_6787, SubBytesIns_Inst_Sbox_8_M13}), .c ({new_AGEMA_signal_7220, new_AGEMA_signal_7219, SubBytesIns_Inst_Sbox_8_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M23_U1 ( .a ({new_AGEMA_signal_7214, new_AGEMA_signal_7213, SubBytesIns_Inst_Sbox_8_M19}), .b ({new_AGEMA_signal_6776, new_AGEMA_signal_6775, SubBytesIns_Inst_Sbox_8_T25}), .c ({new_AGEMA_signal_7374, new_AGEMA_signal_7373, SubBytesIns_Inst_Sbox_8_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M24_U1 ( .a ({new_AGEMA_signal_7220, new_AGEMA_signal_7219, SubBytesIns_Inst_Sbox_8_M22}), .b ({new_AGEMA_signal_7374, new_AGEMA_signal_7373, SubBytesIns_Inst_Sbox_8_M23}), .c ({new_AGEMA_signal_7558, new_AGEMA_signal_7557, SubBytesIns_Inst_Sbox_8_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M27_U1 ( .a ({new_AGEMA_signal_7216, new_AGEMA_signal_7215, SubBytesIns_Inst_Sbox_8_M20}), .b ({new_AGEMA_signal_7218, new_AGEMA_signal_7217, SubBytesIns_Inst_Sbox_8_M21}), .c ({new_AGEMA_signal_7378, new_AGEMA_signal_7377, SubBytesIns_Inst_Sbox_8_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M1_U1 ( .a ({new_AGEMA_signal_5930, new_AGEMA_signal_5929, SubBytesIns_Inst_Sbox_9_T13}), .b ({new_AGEMA_signal_5926, new_AGEMA_signal_5925, SubBytesIns_Inst_Sbox_9_T6}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243]}), .c ({new_AGEMA_signal_6390, new_AGEMA_signal_6389, SubBytesIns_Inst_Sbox_9_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M2_U1 ( .a ({new_AGEMA_signal_6386, new_AGEMA_signal_6385, SubBytesIns_Inst_Sbox_9_T23}), .b ({new_AGEMA_signal_6376, new_AGEMA_signal_6375, SubBytesIns_Inst_Sbox_9_T8}), .clk (clk), .r ({Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_6796, new_AGEMA_signal_6795, SubBytesIns_Inst_Sbox_9_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M3_U1 ( .a ({new_AGEMA_signal_6380, new_AGEMA_signal_6379, SubBytesIns_Inst_Sbox_9_T14}), .b ({new_AGEMA_signal_6390, new_AGEMA_signal_6389, SubBytesIns_Inst_Sbox_9_M1}), .c ({new_AGEMA_signal_6798, new_AGEMA_signal_6797, SubBytesIns_Inst_Sbox_9_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M4_U1 ( .a ({new_AGEMA_signal_5936, new_AGEMA_signal_5935, SubBytesIns_Inst_Sbox_9_T19}), .b ({ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249]}), .c ({new_AGEMA_signal_6392, new_AGEMA_signal_6391, SubBytesIns_Inst_Sbox_9_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M5_U1 ( .a ({new_AGEMA_signal_6392, new_AGEMA_signal_6391, SubBytesIns_Inst_Sbox_9_M4}), .b ({new_AGEMA_signal_6390, new_AGEMA_signal_6389, SubBytesIns_Inst_Sbox_9_M1}), .c ({new_AGEMA_signal_6800, new_AGEMA_signal_6799, SubBytesIns_Inst_Sbox_9_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M6_U1 ( .a ({new_AGEMA_signal_5582, new_AGEMA_signal_5581, SubBytesIns_Inst_Sbox_9_T3}), .b ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, SubBytesIns_Inst_Sbox_9_T16}), .clk (clk), .r ({Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_6394, new_AGEMA_signal_6393, SubBytesIns_Inst_Sbox_9_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M7_U1 ( .a ({new_AGEMA_signal_5938, new_AGEMA_signal_5937, SubBytesIns_Inst_Sbox_9_T22}), .b ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, SubBytesIns_Inst_Sbox_9_T9}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255]}), .c ({new_AGEMA_signal_6396, new_AGEMA_signal_6395, SubBytesIns_Inst_Sbox_9_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M8_U1 ( .a ({new_AGEMA_signal_6388, new_AGEMA_signal_6387, SubBytesIns_Inst_Sbox_9_T26}), .b ({new_AGEMA_signal_6394, new_AGEMA_signal_6393, SubBytesIns_Inst_Sbox_9_M6}), .c ({new_AGEMA_signal_6802, new_AGEMA_signal_6801, SubBytesIns_Inst_Sbox_9_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M9_U1 ( .a ({new_AGEMA_signal_6384, new_AGEMA_signal_6383, SubBytesIns_Inst_Sbox_9_T20}), .b ({new_AGEMA_signal_6382, new_AGEMA_signal_6381, SubBytesIns_Inst_Sbox_9_T17}), .clk (clk), .r ({Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_6804, new_AGEMA_signal_6803, SubBytesIns_Inst_Sbox_9_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M10_U1 ( .a ({new_AGEMA_signal_6804, new_AGEMA_signal_6803, SubBytesIns_Inst_Sbox_9_M9}), .b ({new_AGEMA_signal_6394, new_AGEMA_signal_6393, SubBytesIns_Inst_Sbox_9_M6}), .c ({new_AGEMA_signal_7048, new_AGEMA_signal_7047, SubBytesIns_Inst_Sbox_9_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M11_U1 ( .a ({new_AGEMA_signal_5578, new_AGEMA_signal_5577, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_5932, new_AGEMA_signal_5931, SubBytesIns_Inst_Sbox_9_T15}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261]}), .c ({new_AGEMA_signal_6398, new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_9_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M12_U1 ( .a ({new_AGEMA_signal_5584, new_AGEMA_signal_5583, SubBytesIns_Inst_Sbox_9_T4}), .b ({new_AGEMA_signal_5940, new_AGEMA_signal_5939, SubBytesIns_Inst_Sbox_9_T27}), .clk (clk), .r ({Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_6400, new_AGEMA_signal_6399, SubBytesIns_Inst_Sbox_9_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M13_U1 ( .a ({new_AGEMA_signal_6400, new_AGEMA_signal_6399, SubBytesIns_Inst_Sbox_9_M12}), .b ({new_AGEMA_signal_6398, new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_9_M11}), .c ({new_AGEMA_signal_6806, new_AGEMA_signal_6805, SubBytesIns_Inst_Sbox_9_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M14_U1 ( .a ({new_AGEMA_signal_5580, new_AGEMA_signal_5579, SubBytesIns_Inst_Sbox_9_T2}), .b ({new_AGEMA_signal_6378, new_AGEMA_signal_6377, SubBytesIns_Inst_Sbox_9_T10}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267]}), .c ({new_AGEMA_signal_6808, new_AGEMA_signal_6807, SubBytesIns_Inst_Sbox_9_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M15_U1 ( .a ({new_AGEMA_signal_6808, new_AGEMA_signal_6807, SubBytesIns_Inst_Sbox_9_M14}), .b ({new_AGEMA_signal_6398, new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_9_M11}), .c ({new_AGEMA_signal_7050, new_AGEMA_signal_7049, SubBytesIns_Inst_Sbox_9_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M16_U1 ( .a ({new_AGEMA_signal_6798, new_AGEMA_signal_6797, SubBytesIns_Inst_Sbox_9_M3}), .b ({new_AGEMA_signal_6796, new_AGEMA_signal_6795, SubBytesIns_Inst_Sbox_9_M2}), .c ({new_AGEMA_signal_7052, new_AGEMA_signal_7051, SubBytesIns_Inst_Sbox_9_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M17_U1 ( .a ({new_AGEMA_signal_6800, new_AGEMA_signal_6799, SubBytesIns_Inst_Sbox_9_M5}), .b ({new_AGEMA_signal_6792, new_AGEMA_signal_6791, SubBytesIns_Inst_Sbox_9_T24}), .c ({new_AGEMA_signal_7054, new_AGEMA_signal_7053, SubBytesIns_Inst_Sbox_9_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M18_U1 ( .a ({new_AGEMA_signal_6802, new_AGEMA_signal_6801, SubBytesIns_Inst_Sbox_9_M8}), .b ({new_AGEMA_signal_6396, new_AGEMA_signal_6395, SubBytesIns_Inst_Sbox_9_M7}), .c ({new_AGEMA_signal_7056, new_AGEMA_signal_7055, SubBytesIns_Inst_Sbox_9_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M19_U1 ( .a ({new_AGEMA_signal_7048, new_AGEMA_signal_7047, SubBytesIns_Inst_Sbox_9_M10}), .b ({new_AGEMA_signal_7050, new_AGEMA_signal_7049, SubBytesIns_Inst_Sbox_9_M15}), .c ({new_AGEMA_signal_7222, new_AGEMA_signal_7221, SubBytesIns_Inst_Sbox_9_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M20_U1 ( .a ({new_AGEMA_signal_7052, new_AGEMA_signal_7051, SubBytesIns_Inst_Sbox_9_M16}), .b ({new_AGEMA_signal_6806, new_AGEMA_signal_6805, SubBytesIns_Inst_Sbox_9_M13}), .c ({new_AGEMA_signal_7224, new_AGEMA_signal_7223, SubBytesIns_Inst_Sbox_9_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M21_U1 ( .a ({new_AGEMA_signal_7054, new_AGEMA_signal_7053, SubBytesIns_Inst_Sbox_9_M17}), .b ({new_AGEMA_signal_7050, new_AGEMA_signal_7049, SubBytesIns_Inst_Sbox_9_M15}), .c ({new_AGEMA_signal_7226, new_AGEMA_signal_7225, SubBytesIns_Inst_Sbox_9_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M22_U1 ( .a ({new_AGEMA_signal_7056, new_AGEMA_signal_7055, SubBytesIns_Inst_Sbox_9_M18}), .b ({new_AGEMA_signal_6806, new_AGEMA_signal_6805, SubBytesIns_Inst_Sbox_9_M13}), .c ({new_AGEMA_signal_7228, new_AGEMA_signal_7227, SubBytesIns_Inst_Sbox_9_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M23_U1 ( .a ({new_AGEMA_signal_7222, new_AGEMA_signal_7221, SubBytesIns_Inst_Sbox_9_M19}), .b ({new_AGEMA_signal_6794, new_AGEMA_signal_6793, SubBytesIns_Inst_Sbox_9_T25}), .c ({new_AGEMA_signal_7382, new_AGEMA_signal_7381, SubBytesIns_Inst_Sbox_9_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M24_U1 ( .a ({new_AGEMA_signal_7228, new_AGEMA_signal_7227, SubBytesIns_Inst_Sbox_9_M22}), .b ({new_AGEMA_signal_7382, new_AGEMA_signal_7381, SubBytesIns_Inst_Sbox_9_M23}), .c ({new_AGEMA_signal_7568, new_AGEMA_signal_7567, SubBytesIns_Inst_Sbox_9_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M27_U1 ( .a ({new_AGEMA_signal_7224, new_AGEMA_signal_7223, SubBytesIns_Inst_Sbox_9_M20}), .b ({new_AGEMA_signal_7226, new_AGEMA_signal_7225, SubBytesIns_Inst_Sbox_9_M21}), .c ({new_AGEMA_signal_7386, new_AGEMA_signal_7385, SubBytesIns_Inst_Sbox_9_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M1_U1 ( .a ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, SubBytesIns_Inst_Sbox_10_T13}), .b ({new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_10_T6}), .clk (clk), .r ({Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_6416, new_AGEMA_signal_6415, SubBytesIns_Inst_Sbox_10_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M2_U1 ( .a ({new_AGEMA_signal_6412, new_AGEMA_signal_6411, SubBytesIns_Inst_Sbox_10_T23}), .b ({new_AGEMA_signal_6402, new_AGEMA_signal_6401, SubBytesIns_Inst_Sbox_10_T8}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273]}), .c ({new_AGEMA_signal_6814, new_AGEMA_signal_6813, SubBytesIns_Inst_Sbox_10_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M3_U1 ( .a ({new_AGEMA_signal_6406, new_AGEMA_signal_6405, SubBytesIns_Inst_Sbox_10_T14}), .b ({new_AGEMA_signal_6416, new_AGEMA_signal_6415, SubBytesIns_Inst_Sbox_10_M1}), .c ({new_AGEMA_signal_6816, new_AGEMA_signal_6815, SubBytesIns_Inst_Sbox_10_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M4_U1 ( .a ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, SubBytesIns_Inst_Sbox_10_T19}), .b ({ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .clk (clk), .r ({Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_6418, new_AGEMA_signal_6417, SubBytesIns_Inst_Sbox_10_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M5_U1 ( .a ({new_AGEMA_signal_6418, new_AGEMA_signal_6417, SubBytesIns_Inst_Sbox_10_M4}), .b ({new_AGEMA_signal_6416, new_AGEMA_signal_6415, SubBytesIns_Inst_Sbox_10_M1}), .c ({new_AGEMA_signal_6818, new_AGEMA_signal_6817, SubBytesIns_Inst_Sbox_10_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M6_U1 ( .a ({new_AGEMA_signal_5602, new_AGEMA_signal_5601, SubBytesIns_Inst_Sbox_10_T3}), .b ({new_AGEMA_signal_5950, new_AGEMA_signal_5949, SubBytesIns_Inst_Sbox_10_T16}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279]}), .c ({new_AGEMA_signal_6420, new_AGEMA_signal_6419, SubBytesIns_Inst_Sbox_10_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M7_U1 ( .a ({new_AGEMA_signal_5954, new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_10_T22}), .b ({new_AGEMA_signal_5944, new_AGEMA_signal_5943, SubBytesIns_Inst_Sbox_10_T9}), .clk (clk), .r ({Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_6422, new_AGEMA_signal_6421, SubBytesIns_Inst_Sbox_10_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M8_U1 ( .a ({new_AGEMA_signal_6414, new_AGEMA_signal_6413, SubBytesIns_Inst_Sbox_10_T26}), .b ({new_AGEMA_signal_6420, new_AGEMA_signal_6419, SubBytesIns_Inst_Sbox_10_M6}), .c ({new_AGEMA_signal_6820, new_AGEMA_signal_6819, SubBytesIns_Inst_Sbox_10_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M9_U1 ( .a ({new_AGEMA_signal_6410, new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_10_T20}), .b ({new_AGEMA_signal_6408, new_AGEMA_signal_6407, SubBytesIns_Inst_Sbox_10_T17}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285]}), .c ({new_AGEMA_signal_6822, new_AGEMA_signal_6821, SubBytesIns_Inst_Sbox_10_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M10_U1 ( .a ({new_AGEMA_signal_6822, new_AGEMA_signal_6821, SubBytesIns_Inst_Sbox_10_M9}), .b ({new_AGEMA_signal_6420, new_AGEMA_signal_6419, SubBytesIns_Inst_Sbox_10_M6}), .c ({new_AGEMA_signal_7058, new_AGEMA_signal_7057, SubBytesIns_Inst_Sbox_10_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M11_U1 ( .a ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_5948, new_AGEMA_signal_5947, SubBytesIns_Inst_Sbox_10_T15}), .clk (clk), .r ({Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_6424, new_AGEMA_signal_6423, SubBytesIns_Inst_Sbox_10_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M12_U1 ( .a ({new_AGEMA_signal_5604, new_AGEMA_signal_5603, SubBytesIns_Inst_Sbox_10_T4}), .b ({new_AGEMA_signal_5956, new_AGEMA_signal_5955, SubBytesIns_Inst_Sbox_10_T27}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291]}), .c ({new_AGEMA_signal_6426, new_AGEMA_signal_6425, SubBytesIns_Inst_Sbox_10_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M13_U1 ( .a ({new_AGEMA_signal_6426, new_AGEMA_signal_6425, SubBytesIns_Inst_Sbox_10_M12}), .b ({new_AGEMA_signal_6424, new_AGEMA_signal_6423, SubBytesIns_Inst_Sbox_10_M11}), .c ({new_AGEMA_signal_6824, new_AGEMA_signal_6823, SubBytesIns_Inst_Sbox_10_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M14_U1 ( .a ({new_AGEMA_signal_5600, new_AGEMA_signal_5599, SubBytesIns_Inst_Sbox_10_T2}), .b ({new_AGEMA_signal_6404, new_AGEMA_signal_6403, SubBytesIns_Inst_Sbox_10_T10}), .clk (clk), .r ({Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_6826, new_AGEMA_signal_6825, SubBytesIns_Inst_Sbox_10_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M15_U1 ( .a ({new_AGEMA_signal_6826, new_AGEMA_signal_6825, SubBytesIns_Inst_Sbox_10_M14}), .b ({new_AGEMA_signal_6424, new_AGEMA_signal_6423, SubBytesIns_Inst_Sbox_10_M11}), .c ({new_AGEMA_signal_7060, new_AGEMA_signal_7059, SubBytesIns_Inst_Sbox_10_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M16_U1 ( .a ({new_AGEMA_signal_6816, new_AGEMA_signal_6815, SubBytesIns_Inst_Sbox_10_M3}), .b ({new_AGEMA_signal_6814, new_AGEMA_signal_6813, SubBytesIns_Inst_Sbox_10_M2}), .c ({new_AGEMA_signal_7062, new_AGEMA_signal_7061, SubBytesIns_Inst_Sbox_10_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M17_U1 ( .a ({new_AGEMA_signal_6818, new_AGEMA_signal_6817, SubBytesIns_Inst_Sbox_10_M5}), .b ({new_AGEMA_signal_6810, new_AGEMA_signal_6809, SubBytesIns_Inst_Sbox_10_T24}), .c ({new_AGEMA_signal_7064, new_AGEMA_signal_7063, SubBytesIns_Inst_Sbox_10_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M18_U1 ( .a ({new_AGEMA_signal_6820, new_AGEMA_signal_6819, SubBytesIns_Inst_Sbox_10_M8}), .b ({new_AGEMA_signal_6422, new_AGEMA_signal_6421, SubBytesIns_Inst_Sbox_10_M7}), .c ({new_AGEMA_signal_7066, new_AGEMA_signal_7065, SubBytesIns_Inst_Sbox_10_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M19_U1 ( .a ({new_AGEMA_signal_7058, new_AGEMA_signal_7057, SubBytesIns_Inst_Sbox_10_M10}), .b ({new_AGEMA_signal_7060, new_AGEMA_signal_7059, SubBytesIns_Inst_Sbox_10_M15}), .c ({new_AGEMA_signal_7230, new_AGEMA_signal_7229, SubBytesIns_Inst_Sbox_10_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M20_U1 ( .a ({new_AGEMA_signal_7062, new_AGEMA_signal_7061, SubBytesIns_Inst_Sbox_10_M16}), .b ({new_AGEMA_signal_6824, new_AGEMA_signal_6823, SubBytesIns_Inst_Sbox_10_M13}), .c ({new_AGEMA_signal_7232, new_AGEMA_signal_7231, SubBytesIns_Inst_Sbox_10_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M21_U1 ( .a ({new_AGEMA_signal_7064, new_AGEMA_signal_7063, SubBytesIns_Inst_Sbox_10_M17}), .b ({new_AGEMA_signal_7060, new_AGEMA_signal_7059, SubBytesIns_Inst_Sbox_10_M15}), .c ({new_AGEMA_signal_7234, new_AGEMA_signal_7233, SubBytesIns_Inst_Sbox_10_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M22_U1 ( .a ({new_AGEMA_signal_7066, new_AGEMA_signal_7065, SubBytesIns_Inst_Sbox_10_M18}), .b ({new_AGEMA_signal_6824, new_AGEMA_signal_6823, SubBytesIns_Inst_Sbox_10_M13}), .c ({new_AGEMA_signal_7236, new_AGEMA_signal_7235, SubBytesIns_Inst_Sbox_10_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M23_U1 ( .a ({new_AGEMA_signal_7230, new_AGEMA_signal_7229, SubBytesIns_Inst_Sbox_10_M19}), .b ({new_AGEMA_signal_6812, new_AGEMA_signal_6811, SubBytesIns_Inst_Sbox_10_T25}), .c ({new_AGEMA_signal_7390, new_AGEMA_signal_7389, SubBytesIns_Inst_Sbox_10_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M24_U1 ( .a ({new_AGEMA_signal_7236, new_AGEMA_signal_7235, SubBytesIns_Inst_Sbox_10_M22}), .b ({new_AGEMA_signal_7390, new_AGEMA_signal_7389, SubBytesIns_Inst_Sbox_10_M23}), .c ({new_AGEMA_signal_7578, new_AGEMA_signal_7577, SubBytesIns_Inst_Sbox_10_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M27_U1 ( .a ({new_AGEMA_signal_7232, new_AGEMA_signal_7231, SubBytesIns_Inst_Sbox_10_M20}), .b ({new_AGEMA_signal_7234, new_AGEMA_signal_7233, SubBytesIns_Inst_Sbox_10_M21}), .c ({new_AGEMA_signal_7394, new_AGEMA_signal_7393, SubBytesIns_Inst_Sbox_10_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M1_U1 ( .a ({new_AGEMA_signal_5962, new_AGEMA_signal_5961, SubBytesIns_Inst_Sbox_11_T13}), .b ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, SubBytesIns_Inst_Sbox_11_T6}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297]}), .c ({new_AGEMA_signal_6442, new_AGEMA_signal_6441, SubBytesIns_Inst_Sbox_11_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M2_U1 ( .a ({new_AGEMA_signal_6438, new_AGEMA_signal_6437, SubBytesIns_Inst_Sbox_11_T23}), .b ({new_AGEMA_signal_6428, new_AGEMA_signal_6427, SubBytesIns_Inst_Sbox_11_T8}), .clk (clk), .r ({Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_6832, new_AGEMA_signal_6831, SubBytesIns_Inst_Sbox_11_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M3_U1 ( .a ({new_AGEMA_signal_6432, new_AGEMA_signal_6431, SubBytesIns_Inst_Sbox_11_T14}), .b ({new_AGEMA_signal_6442, new_AGEMA_signal_6441, SubBytesIns_Inst_Sbox_11_M1}), .c ({new_AGEMA_signal_6834, new_AGEMA_signal_6833, SubBytesIns_Inst_Sbox_11_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M4_U1 ( .a ({new_AGEMA_signal_5968, new_AGEMA_signal_5967, SubBytesIns_Inst_Sbox_11_T19}), .b ({ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303]}), .c ({new_AGEMA_signal_6444, new_AGEMA_signal_6443, SubBytesIns_Inst_Sbox_11_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M5_U1 ( .a ({new_AGEMA_signal_6444, new_AGEMA_signal_6443, SubBytesIns_Inst_Sbox_11_M4}), .b ({new_AGEMA_signal_6442, new_AGEMA_signal_6441, SubBytesIns_Inst_Sbox_11_M1}), .c ({new_AGEMA_signal_6836, new_AGEMA_signal_6835, SubBytesIns_Inst_Sbox_11_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M6_U1 ( .a ({new_AGEMA_signal_5622, new_AGEMA_signal_5621, SubBytesIns_Inst_Sbox_11_T3}), .b ({new_AGEMA_signal_5966, new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_11_T16}), .clk (clk), .r ({Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_6446, new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_11_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M7_U1 ( .a ({new_AGEMA_signal_5970, new_AGEMA_signal_5969, SubBytesIns_Inst_Sbox_11_T22}), .b ({new_AGEMA_signal_5960, new_AGEMA_signal_5959, SubBytesIns_Inst_Sbox_11_T9}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309]}), .c ({new_AGEMA_signal_6448, new_AGEMA_signal_6447, SubBytesIns_Inst_Sbox_11_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M8_U1 ( .a ({new_AGEMA_signal_6440, new_AGEMA_signal_6439, SubBytesIns_Inst_Sbox_11_T26}), .b ({new_AGEMA_signal_6446, new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_11_M6}), .c ({new_AGEMA_signal_6838, new_AGEMA_signal_6837, SubBytesIns_Inst_Sbox_11_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M9_U1 ( .a ({new_AGEMA_signal_6436, new_AGEMA_signal_6435, SubBytesIns_Inst_Sbox_11_T20}), .b ({new_AGEMA_signal_6434, new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_11_T17}), .clk (clk), .r ({Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_6840, new_AGEMA_signal_6839, SubBytesIns_Inst_Sbox_11_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M10_U1 ( .a ({new_AGEMA_signal_6840, new_AGEMA_signal_6839, SubBytesIns_Inst_Sbox_11_M9}), .b ({new_AGEMA_signal_6446, new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_11_M6}), .c ({new_AGEMA_signal_7068, new_AGEMA_signal_7067, SubBytesIns_Inst_Sbox_11_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M11_U1 ( .a ({new_AGEMA_signal_5618, new_AGEMA_signal_5617, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_5964, new_AGEMA_signal_5963, SubBytesIns_Inst_Sbox_11_T15}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315]}), .c ({new_AGEMA_signal_6450, new_AGEMA_signal_6449, SubBytesIns_Inst_Sbox_11_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M12_U1 ( .a ({new_AGEMA_signal_5624, new_AGEMA_signal_5623, SubBytesIns_Inst_Sbox_11_T4}), .b ({new_AGEMA_signal_5972, new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_11_T27}), .clk (clk), .r ({Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_6452, new_AGEMA_signal_6451, SubBytesIns_Inst_Sbox_11_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M13_U1 ( .a ({new_AGEMA_signal_6452, new_AGEMA_signal_6451, SubBytesIns_Inst_Sbox_11_M12}), .b ({new_AGEMA_signal_6450, new_AGEMA_signal_6449, SubBytesIns_Inst_Sbox_11_M11}), .c ({new_AGEMA_signal_6842, new_AGEMA_signal_6841, SubBytesIns_Inst_Sbox_11_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M14_U1 ( .a ({new_AGEMA_signal_5620, new_AGEMA_signal_5619, SubBytesIns_Inst_Sbox_11_T2}), .b ({new_AGEMA_signal_6430, new_AGEMA_signal_6429, SubBytesIns_Inst_Sbox_11_T10}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321]}), .c ({new_AGEMA_signal_6844, new_AGEMA_signal_6843, SubBytesIns_Inst_Sbox_11_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M15_U1 ( .a ({new_AGEMA_signal_6844, new_AGEMA_signal_6843, SubBytesIns_Inst_Sbox_11_M14}), .b ({new_AGEMA_signal_6450, new_AGEMA_signal_6449, SubBytesIns_Inst_Sbox_11_M11}), .c ({new_AGEMA_signal_7070, new_AGEMA_signal_7069, SubBytesIns_Inst_Sbox_11_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M16_U1 ( .a ({new_AGEMA_signal_6834, new_AGEMA_signal_6833, SubBytesIns_Inst_Sbox_11_M3}), .b ({new_AGEMA_signal_6832, new_AGEMA_signal_6831, SubBytesIns_Inst_Sbox_11_M2}), .c ({new_AGEMA_signal_7072, new_AGEMA_signal_7071, SubBytesIns_Inst_Sbox_11_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M17_U1 ( .a ({new_AGEMA_signal_6836, new_AGEMA_signal_6835, SubBytesIns_Inst_Sbox_11_M5}), .b ({new_AGEMA_signal_6828, new_AGEMA_signal_6827, SubBytesIns_Inst_Sbox_11_T24}), .c ({new_AGEMA_signal_7074, new_AGEMA_signal_7073, SubBytesIns_Inst_Sbox_11_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M18_U1 ( .a ({new_AGEMA_signal_6838, new_AGEMA_signal_6837, SubBytesIns_Inst_Sbox_11_M8}), .b ({new_AGEMA_signal_6448, new_AGEMA_signal_6447, SubBytesIns_Inst_Sbox_11_M7}), .c ({new_AGEMA_signal_7076, new_AGEMA_signal_7075, SubBytesIns_Inst_Sbox_11_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M19_U1 ( .a ({new_AGEMA_signal_7068, new_AGEMA_signal_7067, SubBytesIns_Inst_Sbox_11_M10}), .b ({new_AGEMA_signal_7070, new_AGEMA_signal_7069, SubBytesIns_Inst_Sbox_11_M15}), .c ({new_AGEMA_signal_7238, new_AGEMA_signal_7237, SubBytesIns_Inst_Sbox_11_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M20_U1 ( .a ({new_AGEMA_signal_7072, new_AGEMA_signal_7071, SubBytesIns_Inst_Sbox_11_M16}), .b ({new_AGEMA_signal_6842, new_AGEMA_signal_6841, SubBytesIns_Inst_Sbox_11_M13}), .c ({new_AGEMA_signal_7240, new_AGEMA_signal_7239, SubBytesIns_Inst_Sbox_11_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M21_U1 ( .a ({new_AGEMA_signal_7074, new_AGEMA_signal_7073, SubBytesIns_Inst_Sbox_11_M17}), .b ({new_AGEMA_signal_7070, new_AGEMA_signal_7069, SubBytesIns_Inst_Sbox_11_M15}), .c ({new_AGEMA_signal_7242, new_AGEMA_signal_7241, SubBytesIns_Inst_Sbox_11_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M22_U1 ( .a ({new_AGEMA_signal_7076, new_AGEMA_signal_7075, SubBytesIns_Inst_Sbox_11_M18}), .b ({new_AGEMA_signal_6842, new_AGEMA_signal_6841, SubBytesIns_Inst_Sbox_11_M13}), .c ({new_AGEMA_signal_7244, new_AGEMA_signal_7243, SubBytesIns_Inst_Sbox_11_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M23_U1 ( .a ({new_AGEMA_signal_7238, new_AGEMA_signal_7237, SubBytesIns_Inst_Sbox_11_M19}), .b ({new_AGEMA_signal_6830, new_AGEMA_signal_6829, SubBytesIns_Inst_Sbox_11_T25}), .c ({new_AGEMA_signal_7398, new_AGEMA_signal_7397, SubBytesIns_Inst_Sbox_11_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M24_U1 ( .a ({new_AGEMA_signal_7244, new_AGEMA_signal_7243, SubBytesIns_Inst_Sbox_11_M22}), .b ({new_AGEMA_signal_7398, new_AGEMA_signal_7397, SubBytesIns_Inst_Sbox_11_M23}), .c ({new_AGEMA_signal_7588, new_AGEMA_signal_7587, SubBytesIns_Inst_Sbox_11_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M27_U1 ( .a ({new_AGEMA_signal_7240, new_AGEMA_signal_7239, SubBytesIns_Inst_Sbox_11_M20}), .b ({new_AGEMA_signal_7242, new_AGEMA_signal_7241, SubBytesIns_Inst_Sbox_11_M21}), .c ({new_AGEMA_signal_7402, new_AGEMA_signal_7401, SubBytesIns_Inst_Sbox_11_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M1_U1 ( .a ({new_AGEMA_signal_5978, new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_12_T13}), .b ({new_AGEMA_signal_5974, new_AGEMA_signal_5973, SubBytesIns_Inst_Sbox_12_T6}), .clk (clk), .r ({Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_6468, new_AGEMA_signal_6467, SubBytesIns_Inst_Sbox_12_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M2_U1 ( .a ({new_AGEMA_signal_6464, new_AGEMA_signal_6463, SubBytesIns_Inst_Sbox_12_T23}), .b ({new_AGEMA_signal_6454, new_AGEMA_signal_6453, SubBytesIns_Inst_Sbox_12_T8}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327]}), .c ({new_AGEMA_signal_6850, new_AGEMA_signal_6849, SubBytesIns_Inst_Sbox_12_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M3_U1 ( .a ({new_AGEMA_signal_6458, new_AGEMA_signal_6457, SubBytesIns_Inst_Sbox_12_T14}), .b ({new_AGEMA_signal_6468, new_AGEMA_signal_6467, SubBytesIns_Inst_Sbox_12_M1}), .c ({new_AGEMA_signal_6852, new_AGEMA_signal_6851, SubBytesIns_Inst_Sbox_12_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M4_U1 ( .a ({new_AGEMA_signal_5984, new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_12_T19}), .b ({ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .clk (clk), .r ({Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_6470, new_AGEMA_signal_6469, SubBytesIns_Inst_Sbox_12_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M5_U1 ( .a ({new_AGEMA_signal_6470, new_AGEMA_signal_6469, SubBytesIns_Inst_Sbox_12_M4}), .b ({new_AGEMA_signal_6468, new_AGEMA_signal_6467, SubBytesIns_Inst_Sbox_12_M1}), .c ({new_AGEMA_signal_6854, new_AGEMA_signal_6853, SubBytesIns_Inst_Sbox_12_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M6_U1 ( .a ({new_AGEMA_signal_5642, new_AGEMA_signal_5641, SubBytesIns_Inst_Sbox_12_T3}), .b ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, SubBytesIns_Inst_Sbox_12_T16}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333]}), .c ({new_AGEMA_signal_6472, new_AGEMA_signal_6471, SubBytesIns_Inst_Sbox_12_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M7_U1 ( .a ({new_AGEMA_signal_5986, new_AGEMA_signal_5985, SubBytesIns_Inst_Sbox_12_T22}), .b ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, SubBytesIns_Inst_Sbox_12_T9}), .clk (clk), .r ({Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_6474, new_AGEMA_signal_6473, SubBytesIns_Inst_Sbox_12_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M8_U1 ( .a ({new_AGEMA_signal_6466, new_AGEMA_signal_6465, SubBytesIns_Inst_Sbox_12_T26}), .b ({new_AGEMA_signal_6472, new_AGEMA_signal_6471, SubBytesIns_Inst_Sbox_12_M6}), .c ({new_AGEMA_signal_6856, new_AGEMA_signal_6855, SubBytesIns_Inst_Sbox_12_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M9_U1 ( .a ({new_AGEMA_signal_6462, new_AGEMA_signal_6461, SubBytesIns_Inst_Sbox_12_T20}), .b ({new_AGEMA_signal_6460, new_AGEMA_signal_6459, SubBytesIns_Inst_Sbox_12_T17}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339]}), .c ({new_AGEMA_signal_6858, new_AGEMA_signal_6857, SubBytesIns_Inst_Sbox_12_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M10_U1 ( .a ({new_AGEMA_signal_6858, new_AGEMA_signal_6857, SubBytesIns_Inst_Sbox_12_M9}), .b ({new_AGEMA_signal_6472, new_AGEMA_signal_6471, SubBytesIns_Inst_Sbox_12_M6}), .c ({new_AGEMA_signal_7078, new_AGEMA_signal_7077, SubBytesIns_Inst_Sbox_12_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M11_U1 ( .a ({new_AGEMA_signal_5638, new_AGEMA_signal_5637, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_5980, new_AGEMA_signal_5979, SubBytesIns_Inst_Sbox_12_T15}), .clk (clk), .r ({Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_6476, new_AGEMA_signal_6475, SubBytesIns_Inst_Sbox_12_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M12_U1 ( .a ({new_AGEMA_signal_5644, new_AGEMA_signal_5643, SubBytesIns_Inst_Sbox_12_T4}), .b ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, SubBytesIns_Inst_Sbox_12_T27}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345]}), .c ({new_AGEMA_signal_6478, new_AGEMA_signal_6477, SubBytesIns_Inst_Sbox_12_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M13_U1 ( .a ({new_AGEMA_signal_6478, new_AGEMA_signal_6477, SubBytesIns_Inst_Sbox_12_M12}), .b ({new_AGEMA_signal_6476, new_AGEMA_signal_6475, SubBytesIns_Inst_Sbox_12_M11}), .c ({new_AGEMA_signal_6860, new_AGEMA_signal_6859, SubBytesIns_Inst_Sbox_12_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M14_U1 ( .a ({new_AGEMA_signal_5640, new_AGEMA_signal_5639, SubBytesIns_Inst_Sbox_12_T2}), .b ({new_AGEMA_signal_6456, new_AGEMA_signal_6455, SubBytesIns_Inst_Sbox_12_T10}), .clk (clk), .r ({Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_6862, new_AGEMA_signal_6861, SubBytesIns_Inst_Sbox_12_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M15_U1 ( .a ({new_AGEMA_signal_6862, new_AGEMA_signal_6861, SubBytesIns_Inst_Sbox_12_M14}), .b ({new_AGEMA_signal_6476, new_AGEMA_signal_6475, SubBytesIns_Inst_Sbox_12_M11}), .c ({new_AGEMA_signal_7080, new_AGEMA_signal_7079, SubBytesIns_Inst_Sbox_12_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M16_U1 ( .a ({new_AGEMA_signal_6852, new_AGEMA_signal_6851, SubBytesIns_Inst_Sbox_12_M3}), .b ({new_AGEMA_signal_6850, new_AGEMA_signal_6849, SubBytesIns_Inst_Sbox_12_M2}), .c ({new_AGEMA_signal_7082, new_AGEMA_signal_7081, SubBytesIns_Inst_Sbox_12_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M17_U1 ( .a ({new_AGEMA_signal_6854, new_AGEMA_signal_6853, SubBytesIns_Inst_Sbox_12_M5}), .b ({new_AGEMA_signal_6846, new_AGEMA_signal_6845, SubBytesIns_Inst_Sbox_12_T24}), .c ({new_AGEMA_signal_7084, new_AGEMA_signal_7083, SubBytesIns_Inst_Sbox_12_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M18_U1 ( .a ({new_AGEMA_signal_6856, new_AGEMA_signal_6855, SubBytesIns_Inst_Sbox_12_M8}), .b ({new_AGEMA_signal_6474, new_AGEMA_signal_6473, SubBytesIns_Inst_Sbox_12_M7}), .c ({new_AGEMA_signal_7086, new_AGEMA_signal_7085, SubBytesIns_Inst_Sbox_12_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M19_U1 ( .a ({new_AGEMA_signal_7078, new_AGEMA_signal_7077, SubBytesIns_Inst_Sbox_12_M10}), .b ({new_AGEMA_signal_7080, new_AGEMA_signal_7079, SubBytesIns_Inst_Sbox_12_M15}), .c ({new_AGEMA_signal_7246, new_AGEMA_signal_7245, SubBytesIns_Inst_Sbox_12_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M20_U1 ( .a ({new_AGEMA_signal_7082, new_AGEMA_signal_7081, SubBytesIns_Inst_Sbox_12_M16}), .b ({new_AGEMA_signal_6860, new_AGEMA_signal_6859, SubBytesIns_Inst_Sbox_12_M13}), .c ({new_AGEMA_signal_7248, new_AGEMA_signal_7247, SubBytesIns_Inst_Sbox_12_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M21_U1 ( .a ({new_AGEMA_signal_7084, new_AGEMA_signal_7083, SubBytesIns_Inst_Sbox_12_M17}), .b ({new_AGEMA_signal_7080, new_AGEMA_signal_7079, SubBytesIns_Inst_Sbox_12_M15}), .c ({new_AGEMA_signal_7250, new_AGEMA_signal_7249, SubBytesIns_Inst_Sbox_12_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M22_U1 ( .a ({new_AGEMA_signal_7086, new_AGEMA_signal_7085, SubBytesIns_Inst_Sbox_12_M18}), .b ({new_AGEMA_signal_6860, new_AGEMA_signal_6859, SubBytesIns_Inst_Sbox_12_M13}), .c ({new_AGEMA_signal_7252, new_AGEMA_signal_7251, SubBytesIns_Inst_Sbox_12_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M23_U1 ( .a ({new_AGEMA_signal_7246, new_AGEMA_signal_7245, SubBytesIns_Inst_Sbox_12_M19}), .b ({new_AGEMA_signal_6848, new_AGEMA_signal_6847, SubBytesIns_Inst_Sbox_12_T25}), .c ({new_AGEMA_signal_7406, new_AGEMA_signal_7405, SubBytesIns_Inst_Sbox_12_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M24_U1 ( .a ({new_AGEMA_signal_7252, new_AGEMA_signal_7251, SubBytesIns_Inst_Sbox_12_M22}), .b ({new_AGEMA_signal_7406, new_AGEMA_signal_7405, SubBytesIns_Inst_Sbox_12_M23}), .c ({new_AGEMA_signal_7598, new_AGEMA_signal_7597, SubBytesIns_Inst_Sbox_12_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M27_U1 ( .a ({new_AGEMA_signal_7248, new_AGEMA_signal_7247, SubBytesIns_Inst_Sbox_12_M20}), .b ({new_AGEMA_signal_7250, new_AGEMA_signal_7249, SubBytesIns_Inst_Sbox_12_M21}), .c ({new_AGEMA_signal_7410, new_AGEMA_signal_7409, SubBytesIns_Inst_Sbox_12_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M1_U1 ( .a ({new_AGEMA_signal_5994, new_AGEMA_signal_5993, SubBytesIns_Inst_Sbox_13_T13}), .b ({new_AGEMA_signal_5990, new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_13_T6}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351]}), .c ({new_AGEMA_signal_6494, new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_13_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M2_U1 ( .a ({new_AGEMA_signal_6490, new_AGEMA_signal_6489, SubBytesIns_Inst_Sbox_13_T23}), .b ({new_AGEMA_signal_6480, new_AGEMA_signal_6479, SubBytesIns_Inst_Sbox_13_T8}), .clk (clk), .r ({Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_6868, new_AGEMA_signal_6867, SubBytesIns_Inst_Sbox_13_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M3_U1 ( .a ({new_AGEMA_signal_6484, new_AGEMA_signal_6483, SubBytesIns_Inst_Sbox_13_T14}), .b ({new_AGEMA_signal_6494, new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_13_M1}), .c ({new_AGEMA_signal_6870, new_AGEMA_signal_6869, SubBytesIns_Inst_Sbox_13_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M4_U1 ( .a ({new_AGEMA_signal_6000, new_AGEMA_signal_5999, SubBytesIns_Inst_Sbox_13_T19}), .b ({ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357]}), .c ({new_AGEMA_signal_6496, new_AGEMA_signal_6495, SubBytesIns_Inst_Sbox_13_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M5_U1 ( .a ({new_AGEMA_signal_6496, new_AGEMA_signal_6495, SubBytesIns_Inst_Sbox_13_M4}), .b ({new_AGEMA_signal_6494, new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_13_M1}), .c ({new_AGEMA_signal_6872, new_AGEMA_signal_6871, SubBytesIns_Inst_Sbox_13_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M6_U1 ( .a ({new_AGEMA_signal_5662, new_AGEMA_signal_5661, SubBytesIns_Inst_Sbox_13_T3}), .b ({new_AGEMA_signal_5998, new_AGEMA_signal_5997, SubBytesIns_Inst_Sbox_13_T16}), .clk (clk), .r ({Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_6498, new_AGEMA_signal_6497, SubBytesIns_Inst_Sbox_13_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M7_U1 ( .a ({new_AGEMA_signal_6002, new_AGEMA_signal_6001, SubBytesIns_Inst_Sbox_13_T22}), .b ({new_AGEMA_signal_5992, new_AGEMA_signal_5991, SubBytesIns_Inst_Sbox_13_T9}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363]}), .c ({new_AGEMA_signal_6500, new_AGEMA_signal_6499, SubBytesIns_Inst_Sbox_13_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M8_U1 ( .a ({new_AGEMA_signal_6492, new_AGEMA_signal_6491, SubBytesIns_Inst_Sbox_13_T26}), .b ({new_AGEMA_signal_6498, new_AGEMA_signal_6497, SubBytesIns_Inst_Sbox_13_M6}), .c ({new_AGEMA_signal_6874, new_AGEMA_signal_6873, SubBytesIns_Inst_Sbox_13_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M9_U1 ( .a ({new_AGEMA_signal_6488, new_AGEMA_signal_6487, SubBytesIns_Inst_Sbox_13_T20}), .b ({new_AGEMA_signal_6486, new_AGEMA_signal_6485, SubBytesIns_Inst_Sbox_13_T17}), .clk (clk), .r ({Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_6876, new_AGEMA_signal_6875, SubBytesIns_Inst_Sbox_13_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M10_U1 ( .a ({new_AGEMA_signal_6876, new_AGEMA_signal_6875, SubBytesIns_Inst_Sbox_13_M9}), .b ({new_AGEMA_signal_6498, new_AGEMA_signal_6497, SubBytesIns_Inst_Sbox_13_M6}), .c ({new_AGEMA_signal_7088, new_AGEMA_signal_7087, SubBytesIns_Inst_Sbox_13_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M11_U1 ( .a ({new_AGEMA_signal_5658, new_AGEMA_signal_5657, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_5996, new_AGEMA_signal_5995, SubBytesIns_Inst_Sbox_13_T15}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369]}), .c ({new_AGEMA_signal_6502, new_AGEMA_signal_6501, SubBytesIns_Inst_Sbox_13_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M12_U1 ( .a ({new_AGEMA_signal_5664, new_AGEMA_signal_5663, SubBytesIns_Inst_Sbox_13_T4}), .b ({new_AGEMA_signal_6004, new_AGEMA_signal_6003, SubBytesIns_Inst_Sbox_13_T27}), .clk (clk), .r ({Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_6504, new_AGEMA_signal_6503, SubBytesIns_Inst_Sbox_13_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M13_U1 ( .a ({new_AGEMA_signal_6504, new_AGEMA_signal_6503, SubBytesIns_Inst_Sbox_13_M12}), .b ({new_AGEMA_signal_6502, new_AGEMA_signal_6501, SubBytesIns_Inst_Sbox_13_M11}), .c ({new_AGEMA_signal_6878, new_AGEMA_signal_6877, SubBytesIns_Inst_Sbox_13_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M14_U1 ( .a ({new_AGEMA_signal_5660, new_AGEMA_signal_5659, SubBytesIns_Inst_Sbox_13_T2}), .b ({new_AGEMA_signal_6482, new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_13_T10}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375]}), .c ({new_AGEMA_signal_6880, new_AGEMA_signal_6879, SubBytesIns_Inst_Sbox_13_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M15_U1 ( .a ({new_AGEMA_signal_6880, new_AGEMA_signal_6879, SubBytesIns_Inst_Sbox_13_M14}), .b ({new_AGEMA_signal_6502, new_AGEMA_signal_6501, SubBytesIns_Inst_Sbox_13_M11}), .c ({new_AGEMA_signal_7090, new_AGEMA_signal_7089, SubBytesIns_Inst_Sbox_13_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M16_U1 ( .a ({new_AGEMA_signal_6870, new_AGEMA_signal_6869, SubBytesIns_Inst_Sbox_13_M3}), .b ({new_AGEMA_signal_6868, new_AGEMA_signal_6867, SubBytesIns_Inst_Sbox_13_M2}), .c ({new_AGEMA_signal_7092, new_AGEMA_signal_7091, SubBytesIns_Inst_Sbox_13_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M17_U1 ( .a ({new_AGEMA_signal_6872, new_AGEMA_signal_6871, SubBytesIns_Inst_Sbox_13_M5}), .b ({new_AGEMA_signal_6864, new_AGEMA_signal_6863, SubBytesIns_Inst_Sbox_13_T24}), .c ({new_AGEMA_signal_7094, new_AGEMA_signal_7093, SubBytesIns_Inst_Sbox_13_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M18_U1 ( .a ({new_AGEMA_signal_6874, new_AGEMA_signal_6873, SubBytesIns_Inst_Sbox_13_M8}), .b ({new_AGEMA_signal_6500, new_AGEMA_signal_6499, SubBytesIns_Inst_Sbox_13_M7}), .c ({new_AGEMA_signal_7096, new_AGEMA_signal_7095, SubBytesIns_Inst_Sbox_13_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M19_U1 ( .a ({new_AGEMA_signal_7088, new_AGEMA_signal_7087, SubBytesIns_Inst_Sbox_13_M10}), .b ({new_AGEMA_signal_7090, new_AGEMA_signal_7089, SubBytesIns_Inst_Sbox_13_M15}), .c ({new_AGEMA_signal_7254, new_AGEMA_signal_7253, SubBytesIns_Inst_Sbox_13_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M20_U1 ( .a ({new_AGEMA_signal_7092, new_AGEMA_signal_7091, SubBytesIns_Inst_Sbox_13_M16}), .b ({new_AGEMA_signal_6878, new_AGEMA_signal_6877, SubBytesIns_Inst_Sbox_13_M13}), .c ({new_AGEMA_signal_7256, new_AGEMA_signal_7255, SubBytesIns_Inst_Sbox_13_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M21_U1 ( .a ({new_AGEMA_signal_7094, new_AGEMA_signal_7093, SubBytesIns_Inst_Sbox_13_M17}), .b ({new_AGEMA_signal_7090, new_AGEMA_signal_7089, SubBytesIns_Inst_Sbox_13_M15}), .c ({new_AGEMA_signal_7258, new_AGEMA_signal_7257, SubBytesIns_Inst_Sbox_13_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M22_U1 ( .a ({new_AGEMA_signal_7096, new_AGEMA_signal_7095, SubBytesIns_Inst_Sbox_13_M18}), .b ({new_AGEMA_signal_6878, new_AGEMA_signal_6877, SubBytesIns_Inst_Sbox_13_M13}), .c ({new_AGEMA_signal_7260, new_AGEMA_signal_7259, SubBytesIns_Inst_Sbox_13_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M23_U1 ( .a ({new_AGEMA_signal_7254, new_AGEMA_signal_7253, SubBytesIns_Inst_Sbox_13_M19}), .b ({new_AGEMA_signal_6866, new_AGEMA_signal_6865, SubBytesIns_Inst_Sbox_13_T25}), .c ({new_AGEMA_signal_7414, new_AGEMA_signal_7413, SubBytesIns_Inst_Sbox_13_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M24_U1 ( .a ({new_AGEMA_signal_7260, new_AGEMA_signal_7259, SubBytesIns_Inst_Sbox_13_M22}), .b ({new_AGEMA_signal_7414, new_AGEMA_signal_7413, SubBytesIns_Inst_Sbox_13_M23}), .c ({new_AGEMA_signal_7608, new_AGEMA_signal_7607, SubBytesIns_Inst_Sbox_13_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M27_U1 ( .a ({new_AGEMA_signal_7256, new_AGEMA_signal_7255, SubBytesIns_Inst_Sbox_13_M20}), .b ({new_AGEMA_signal_7258, new_AGEMA_signal_7257, SubBytesIns_Inst_Sbox_13_M21}), .c ({new_AGEMA_signal_7418, new_AGEMA_signal_7417, SubBytesIns_Inst_Sbox_13_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M1_U1 ( .a ({new_AGEMA_signal_6010, new_AGEMA_signal_6009, SubBytesIns_Inst_Sbox_14_T13}), .b ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, SubBytesIns_Inst_Sbox_14_T6}), .clk (clk), .r ({Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_6520, new_AGEMA_signal_6519, SubBytesIns_Inst_Sbox_14_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M2_U1 ( .a ({new_AGEMA_signal_6516, new_AGEMA_signal_6515, SubBytesIns_Inst_Sbox_14_T23}), .b ({new_AGEMA_signal_6506, new_AGEMA_signal_6505, SubBytesIns_Inst_Sbox_14_T8}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381]}), .c ({new_AGEMA_signal_6886, new_AGEMA_signal_6885, SubBytesIns_Inst_Sbox_14_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M3_U1 ( .a ({new_AGEMA_signal_6510, new_AGEMA_signal_6509, SubBytesIns_Inst_Sbox_14_T14}), .b ({new_AGEMA_signal_6520, new_AGEMA_signal_6519, SubBytesIns_Inst_Sbox_14_M1}), .c ({new_AGEMA_signal_6888, new_AGEMA_signal_6887, SubBytesIns_Inst_Sbox_14_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M4_U1 ( .a ({new_AGEMA_signal_6016, new_AGEMA_signal_6015, SubBytesIns_Inst_Sbox_14_T19}), .b ({ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .clk (clk), .r ({Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_6522, new_AGEMA_signal_6521, SubBytesIns_Inst_Sbox_14_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M5_U1 ( .a ({new_AGEMA_signal_6522, new_AGEMA_signal_6521, SubBytesIns_Inst_Sbox_14_M4}), .b ({new_AGEMA_signal_6520, new_AGEMA_signal_6519, SubBytesIns_Inst_Sbox_14_M1}), .c ({new_AGEMA_signal_6890, new_AGEMA_signal_6889, SubBytesIns_Inst_Sbox_14_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M6_U1 ( .a ({new_AGEMA_signal_5682, new_AGEMA_signal_5681, SubBytesIns_Inst_Sbox_14_T3}), .b ({new_AGEMA_signal_6014, new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_14_T16}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387]}), .c ({new_AGEMA_signal_6524, new_AGEMA_signal_6523, SubBytesIns_Inst_Sbox_14_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M7_U1 ( .a ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, SubBytesIns_Inst_Sbox_14_T22}), .b ({new_AGEMA_signal_6008, new_AGEMA_signal_6007, SubBytesIns_Inst_Sbox_14_T9}), .clk (clk), .r ({Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_6526, new_AGEMA_signal_6525, SubBytesIns_Inst_Sbox_14_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M8_U1 ( .a ({new_AGEMA_signal_6518, new_AGEMA_signal_6517, SubBytesIns_Inst_Sbox_14_T26}), .b ({new_AGEMA_signal_6524, new_AGEMA_signal_6523, SubBytesIns_Inst_Sbox_14_M6}), .c ({new_AGEMA_signal_6892, new_AGEMA_signal_6891, SubBytesIns_Inst_Sbox_14_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M9_U1 ( .a ({new_AGEMA_signal_6514, new_AGEMA_signal_6513, SubBytesIns_Inst_Sbox_14_T20}), .b ({new_AGEMA_signal_6512, new_AGEMA_signal_6511, SubBytesIns_Inst_Sbox_14_T17}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393]}), .c ({new_AGEMA_signal_6894, new_AGEMA_signal_6893, SubBytesIns_Inst_Sbox_14_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M10_U1 ( .a ({new_AGEMA_signal_6894, new_AGEMA_signal_6893, SubBytesIns_Inst_Sbox_14_M9}), .b ({new_AGEMA_signal_6524, new_AGEMA_signal_6523, SubBytesIns_Inst_Sbox_14_M6}), .c ({new_AGEMA_signal_7098, new_AGEMA_signal_7097, SubBytesIns_Inst_Sbox_14_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M11_U1 ( .a ({new_AGEMA_signal_5678, new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_6012, new_AGEMA_signal_6011, SubBytesIns_Inst_Sbox_14_T15}), .clk (clk), .r ({Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_6528, new_AGEMA_signal_6527, SubBytesIns_Inst_Sbox_14_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M12_U1 ( .a ({new_AGEMA_signal_5684, new_AGEMA_signal_5683, SubBytesIns_Inst_Sbox_14_T4}), .b ({new_AGEMA_signal_6020, new_AGEMA_signal_6019, SubBytesIns_Inst_Sbox_14_T27}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399]}), .c ({new_AGEMA_signal_6530, new_AGEMA_signal_6529, SubBytesIns_Inst_Sbox_14_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M13_U1 ( .a ({new_AGEMA_signal_6530, new_AGEMA_signal_6529, SubBytesIns_Inst_Sbox_14_M12}), .b ({new_AGEMA_signal_6528, new_AGEMA_signal_6527, SubBytesIns_Inst_Sbox_14_M11}), .c ({new_AGEMA_signal_6896, new_AGEMA_signal_6895, SubBytesIns_Inst_Sbox_14_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M14_U1 ( .a ({new_AGEMA_signal_5680, new_AGEMA_signal_5679, SubBytesIns_Inst_Sbox_14_T2}), .b ({new_AGEMA_signal_6508, new_AGEMA_signal_6507, SubBytesIns_Inst_Sbox_14_T10}), .clk (clk), .r ({Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_6898, new_AGEMA_signal_6897, SubBytesIns_Inst_Sbox_14_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M15_U1 ( .a ({new_AGEMA_signal_6898, new_AGEMA_signal_6897, SubBytesIns_Inst_Sbox_14_M14}), .b ({new_AGEMA_signal_6528, new_AGEMA_signal_6527, SubBytesIns_Inst_Sbox_14_M11}), .c ({new_AGEMA_signal_7100, new_AGEMA_signal_7099, SubBytesIns_Inst_Sbox_14_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M16_U1 ( .a ({new_AGEMA_signal_6888, new_AGEMA_signal_6887, SubBytesIns_Inst_Sbox_14_M3}), .b ({new_AGEMA_signal_6886, new_AGEMA_signal_6885, SubBytesIns_Inst_Sbox_14_M2}), .c ({new_AGEMA_signal_7102, new_AGEMA_signal_7101, SubBytesIns_Inst_Sbox_14_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M17_U1 ( .a ({new_AGEMA_signal_6890, new_AGEMA_signal_6889, SubBytesIns_Inst_Sbox_14_M5}), .b ({new_AGEMA_signal_6882, new_AGEMA_signal_6881, SubBytesIns_Inst_Sbox_14_T24}), .c ({new_AGEMA_signal_7104, new_AGEMA_signal_7103, SubBytesIns_Inst_Sbox_14_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M18_U1 ( .a ({new_AGEMA_signal_6892, new_AGEMA_signal_6891, SubBytesIns_Inst_Sbox_14_M8}), .b ({new_AGEMA_signal_6526, new_AGEMA_signal_6525, SubBytesIns_Inst_Sbox_14_M7}), .c ({new_AGEMA_signal_7106, new_AGEMA_signal_7105, SubBytesIns_Inst_Sbox_14_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M19_U1 ( .a ({new_AGEMA_signal_7098, new_AGEMA_signal_7097, SubBytesIns_Inst_Sbox_14_M10}), .b ({new_AGEMA_signal_7100, new_AGEMA_signal_7099, SubBytesIns_Inst_Sbox_14_M15}), .c ({new_AGEMA_signal_7262, new_AGEMA_signal_7261, SubBytesIns_Inst_Sbox_14_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M20_U1 ( .a ({new_AGEMA_signal_7102, new_AGEMA_signal_7101, SubBytesIns_Inst_Sbox_14_M16}), .b ({new_AGEMA_signal_6896, new_AGEMA_signal_6895, SubBytesIns_Inst_Sbox_14_M13}), .c ({new_AGEMA_signal_7264, new_AGEMA_signal_7263, SubBytesIns_Inst_Sbox_14_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M21_U1 ( .a ({new_AGEMA_signal_7104, new_AGEMA_signal_7103, SubBytesIns_Inst_Sbox_14_M17}), .b ({new_AGEMA_signal_7100, new_AGEMA_signal_7099, SubBytesIns_Inst_Sbox_14_M15}), .c ({new_AGEMA_signal_7266, new_AGEMA_signal_7265, SubBytesIns_Inst_Sbox_14_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M22_U1 ( .a ({new_AGEMA_signal_7106, new_AGEMA_signal_7105, SubBytesIns_Inst_Sbox_14_M18}), .b ({new_AGEMA_signal_6896, new_AGEMA_signal_6895, SubBytesIns_Inst_Sbox_14_M13}), .c ({new_AGEMA_signal_7268, new_AGEMA_signal_7267, SubBytesIns_Inst_Sbox_14_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M23_U1 ( .a ({new_AGEMA_signal_7262, new_AGEMA_signal_7261, SubBytesIns_Inst_Sbox_14_M19}), .b ({new_AGEMA_signal_6884, new_AGEMA_signal_6883, SubBytesIns_Inst_Sbox_14_T25}), .c ({new_AGEMA_signal_7422, new_AGEMA_signal_7421, SubBytesIns_Inst_Sbox_14_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M24_U1 ( .a ({new_AGEMA_signal_7268, new_AGEMA_signal_7267, SubBytesIns_Inst_Sbox_14_M22}), .b ({new_AGEMA_signal_7422, new_AGEMA_signal_7421, SubBytesIns_Inst_Sbox_14_M23}), .c ({new_AGEMA_signal_7618, new_AGEMA_signal_7617, SubBytesIns_Inst_Sbox_14_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M27_U1 ( .a ({new_AGEMA_signal_7264, new_AGEMA_signal_7263, SubBytesIns_Inst_Sbox_14_M20}), .b ({new_AGEMA_signal_7266, new_AGEMA_signal_7265, SubBytesIns_Inst_Sbox_14_M21}), .c ({new_AGEMA_signal_7426, new_AGEMA_signal_7425, SubBytesIns_Inst_Sbox_14_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M1_U1 ( .a ({new_AGEMA_signal_6026, new_AGEMA_signal_6025, SubBytesIns_Inst_Sbox_15_T13}), .b ({new_AGEMA_signal_6022, new_AGEMA_signal_6021, SubBytesIns_Inst_Sbox_15_T6}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405]}), .c ({new_AGEMA_signal_6546, new_AGEMA_signal_6545, SubBytesIns_Inst_Sbox_15_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M2_U1 ( .a ({new_AGEMA_signal_6542, new_AGEMA_signal_6541, SubBytesIns_Inst_Sbox_15_T23}), .b ({new_AGEMA_signal_6532, new_AGEMA_signal_6531, SubBytesIns_Inst_Sbox_15_T8}), .clk (clk), .r ({Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_6904, new_AGEMA_signal_6903, SubBytesIns_Inst_Sbox_15_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M3_U1 ( .a ({new_AGEMA_signal_6536, new_AGEMA_signal_6535, SubBytesIns_Inst_Sbox_15_T14}), .b ({new_AGEMA_signal_6546, new_AGEMA_signal_6545, SubBytesIns_Inst_Sbox_15_M1}), .c ({new_AGEMA_signal_6906, new_AGEMA_signal_6905, SubBytesIns_Inst_Sbox_15_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M4_U1 ( .a ({new_AGEMA_signal_6032, new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_15_T19}), .b ({ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411]}), .c ({new_AGEMA_signal_6548, new_AGEMA_signal_6547, SubBytesIns_Inst_Sbox_15_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M5_U1 ( .a ({new_AGEMA_signal_6548, new_AGEMA_signal_6547, SubBytesIns_Inst_Sbox_15_M4}), .b ({new_AGEMA_signal_6546, new_AGEMA_signal_6545, SubBytesIns_Inst_Sbox_15_M1}), .c ({new_AGEMA_signal_6908, new_AGEMA_signal_6907, SubBytesIns_Inst_Sbox_15_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M6_U1 ( .a ({new_AGEMA_signal_5702, new_AGEMA_signal_5701, SubBytesIns_Inst_Sbox_15_T3}), .b ({new_AGEMA_signal_6030, new_AGEMA_signal_6029, SubBytesIns_Inst_Sbox_15_T16}), .clk (clk), .r ({Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_6550, new_AGEMA_signal_6549, SubBytesIns_Inst_Sbox_15_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M7_U1 ( .a ({new_AGEMA_signal_6034, new_AGEMA_signal_6033, SubBytesIns_Inst_Sbox_15_T22}), .b ({new_AGEMA_signal_6024, new_AGEMA_signal_6023, SubBytesIns_Inst_Sbox_15_T9}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417]}), .c ({new_AGEMA_signal_6552, new_AGEMA_signal_6551, SubBytesIns_Inst_Sbox_15_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M8_U1 ( .a ({new_AGEMA_signal_6544, new_AGEMA_signal_6543, SubBytesIns_Inst_Sbox_15_T26}), .b ({new_AGEMA_signal_6550, new_AGEMA_signal_6549, SubBytesIns_Inst_Sbox_15_M6}), .c ({new_AGEMA_signal_6910, new_AGEMA_signal_6909, SubBytesIns_Inst_Sbox_15_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M9_U1 ( .a ({new_AGEMA_signal_6540, new_AGEMA_signal_6539, SubBytesIns_Inst_Sbox_15_T20}), .b ({new_AGEMA_signal_6538, new_AGEMA_signal_6537, SubBytesIns_Inst_Sbox_15_T17}), .clk (clk), .r ({Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_6912, new_AGEMA_signal_6911, SubBytesIns_Inst_Sbox_15_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M10_U1 ( .a ({new_AGEMA_signal_6912, new_AGEMA_signal_6911, SubBytesIns_Inst_Sbox_15_M9}), .b ({new_AGEMA_signal_6550, new_AGEMA_signal_6549, SubBytesIns_Inst_Sbox_15_M6}), .c ({new_AGEMA_signal_7108, new_AGEMA_signal_7107, SubBytesIns_Inst_Sbox_15_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M11_U1 ( .a ({new_AGEMA_signal_5698, new_AGEMA_signal_5697, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_6028, new_AGEMA_signal_6027, SubBytesIns_Inst_Sbox_15_T15}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423]}), .c ({new_AGEMA_signal_6554, new_AGEMA_signal_6553, SubBytesIns_Inst_Sbox_15_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M12_U1 ( .a ({new_AGEMA_signal_5704, new_AGEMA_signal_5703, SubBytesIns_Inst_Sbox_15_T4}), .b ({new_AGEMA_signal_6036, new_AGEMA_signal_6035, SubBytesIns_Inst_Sbox_15_T27}), .clk (clk), .r ({Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_6556, new_AGEMA_signal_6555, SubBytesIns_Inst_Sbox_15_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M13_U1 ( .a ({new_AGEMA_signal_6556, new_AGEMA_signal_6555, SubBytesIns_Inst_Sbox_15_M12}), .b ({new_AGEMA_signal_6554, new_AGEMA_signal_6553, SubBytesIns_Inst_Sbox_15_M11}), .c ({new_AGEMA_signal_6914, new_AGEMA_signal_6913, SubBytesIns_Inst_Sbox_15_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M14_U1 ( .a ({new_AGEMA_signal_5700, new_AGEMA_signal_5699, SubBytesIns_Inst_Sbox_15_T2}), .b ({new_AGEMA_signal_6534, new_AGEMA_signal_6533, SubBytesIns_Inst_Sbox_15_T10}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429]}), .c ({new_AGEMA_signal_6916, new_AGEMA_signal_6915, SubBytesIns_Inst_Sbox_15_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M15_U1 ( .a ({new_AGEMA_signal_6916, new_AGEMA_signal_6915, SubBytesIns_Inst_Sbox_15_M14}), .b ({new_AGEMA_signal_6554, new_AGEMA_signal_6553, SubBytesIns_Inst_Sbox_15_M11}), .c ({new_AGEMA_signal_7110, new_AGEMA_signal_7109, SubBytesIns_Inst_Sbox_15_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M16_U1 ( .a ({new_AGEMA_signal_6906, new_AGEMA_signal_6905, SubBytesIns_Inst_Sbox_15_M3}), .b ({new_AGEMA_signal_6904, new_AGEMA_signal_6903, SubBytesIns_Inst_Sbox_15_M2}), .c ({new_AGEMA_signal_7112, new_AGEMA_signal_7111, SubBytesIns_Inst_Sbox_15_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M17_U1 ( .a ({new_AGEMA_signal_6908, new_AGEMA_signal_6907, SubBytesIns_Inst_Sbox_15_M5}), .b ({new_AGEMA_signal_6900, new_AGEMA_signal_6899, SubBytesIns_Inst_Sbox_15_T24}), .c ({new_AGEMA_signal_7114, new_AGEMA_signal_7113, SubBytesIns_Inst_Sbox_15_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M18_U1 ( .a ({new_AGEMA_signal_6910, new_AGEMA_signal_6909, SubBytesIns_Inst_Sbox_15_M8}), .b ({new_AGEMA_signal_6552, new_AGEMA_signal_6551, SubBytesIns_Inst_Sbox_15_M7}), .c ({new_AGEMA_signal_7116, new_AGEMA_signal_7115, SubBytesIns_Inst_Sbox_15_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M19_U1 ( .a ({new_AGEMA_signal_7108, new_AGEMA_signal_7107, SubBytesIns_Inst_Sbox_15_M10}), .b ({new_AGEMA_signal_7110, new_AGEMA_signal_7109, SubBytesIns_Inst_Sbox_15_M15}), .c ({new_AGEMA_signal_7270, new_AGEMA_signal_7269, SubBytesIns_Inst_Sbox_15_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M20_U1 ( .a ({new_AGEMA_signal_7112, new_AGEMA_signal_7111, SubBytesIns_Inst_Sbox_15_M16}), .b ({new_AGEMA_signal_6914, new_AGEMA_signal_6913, SubBytesIns_Inst_Sbox_15_M13}), .c ({new_AGEMA_signal_7272, new_AGEMA_signal_7271, SubBytesIns_Inst_Sbox_15_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M21_U1 ( .a ({new_AGEMA_signal_7114, new_AGEMA_signal_7113, SubBytesIns_Inst_Sbox_15_M17}), .b ({new_AGEMA_signal_7110, new_AGEMA_signal_7109, SubBytesIns_Inst_Sbox_15_M15}), .c ({new_AGEMA_signal_7274, new_AGEMA_signal_7273, SubBytesIns_Inst_Sbox_15_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M22_U1 ( .a ({new_AGEMA_signal_7116, new_AGEMA_signal_7115, SubBytesIns_Inst_Sbox_15_M18}), .b ({new_AGEMA_signal_6914, new_AGEMA_signal_6913, SubBytesIns_Inst_Sbox_15_M13}), .c ({new_AGEMA_signal_7276, new_AGEMA_signal_7275, SubBytesIns_Inst_Sbox_15_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M23_U1 ( .a ({new_AGEMA_signal_7270, new_AGEMA_signal_7269, SubBytesIns_Inst_Sbox_15_M19}), .b ({new_AGEMA_signal_6902, new_AGEMA_signal_6901, SubBytesIns_Inst_Sbox_15_T25}), .c ({new_AGEMA_signal_7430, new_AGEMA_signal_7429, SubBytesIns_Inst_Sbox_15_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M24_U1 ( .a ({new_AGEMA_signal_7276, new_AGEMA_signal_7275, SubBytesIns_Inst_Sbox_15_M22}), .b ({new_AGEMA_signal_7430, new_AGEMA_signal_7429, SubBytesIns_Inst_Sbox_15_M23}), .c ({new_AGEMA_signal_7628, new_AGEMA_signal_7627, SubBytesIns_Inst_Sbox_15_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M27_U1 ( .a ({new_AGEMA_signal_7272, new_AGEMA_signal_7271, SubBytesIns_Inst_Sbox_15_M20}), .b ({new_AGEMA_signal_7274, new_AGEMA_signal_7273, SubBytesIns_Inst_Sbox_15_M21}), .c ({new_AGEMA_signal_7434, new_AGEMA_signal_7433, SubBytesIns_Inst_Sbox_15_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M1_U1 ( .a ({new_AGEMA_signal_5722, new_AGEMA_signal_5721, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13}), .b ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .clk (clk), .r ({Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_6052, new_AGEMA_signal_6051, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M2_U1 ( .a ({new_AGEMA_signal_6048, new_AGEMA_signal_6047, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23}), .b ({new_AGEMA_signal_6038, new_AGEMA_signal_6037, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435]}), .c ({new_AGEMA_signal_6562, new_AGEMA_signal_6561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M3_U1 ( .a ({new_AGEMA_signal_6042, new_AGEMA_signal_6041, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14}), .b ({new_AGEMA_signal_6052, new_AGEMA_signal_6051, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_6564, new_AGEMA_signal_6563, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M4_U1 ( .a ({new_AGEMA_signal_5728, new_AGEMA_signal_5727, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}), .b ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, RoundKey[16]}), .clk (clk), .r ({Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_6054, new_AGEMA_signal_6053, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M5_U1 ( .a ({new_AGEMA_signal_6054, new_AGEMA_signal_6053, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4}), .b ({new_AGEMA_signal_6052, new_AGEMA_signal_6051, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_6566, new_AGEMA_signal_6565, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M6_U1 ( .a ({new_AGEMA_signal_5322, new_AGEMA_signal_5321, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5726, new_AGEMA_signal_5725, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441]}), .c ({new_AGEMA_signal_6056, new_AGEMA_signal_6055, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M7_U1 ( .a ({new_AGEMA_signal_5730, new_AGEMA_signal_5729, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}), .b ({new_AGEMA_signal_5720, new_AGEMA_signal_5719, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}), .clk (clk), .r ({Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_6058, new_AGEMA_signal_6057, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M8_U1 ( .a ({new_AGEMA_signal_6050, new_AGEMA_signal_6049, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26}), .b ({new_AGEMA_signal_6056, new_AGEMA_signal_6055, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_6568, new_AGEMA_signal_6567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M9_U1 ( .a ({new_AGEMA_signal_6046, new_AGEMA_signal_6045, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_6044, new_AGEMA_signal_6043, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447]}), .c ({new_AGEMA_signal_6570, new_AGEMA_signal_6569, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M10_U1 ( .a ({new_AGEMA_signal_6570, new_AGEMA_signal_6569, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9}), .b ({new_AGEMA_signal_6056, new_AGEMA_signal_6055, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_6918, new_AGEMA_signal_6917, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M11_U1 ( .a ({new_AGEMA_signal_5318, new_AGEMA_signal_5317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5724, new_AGEMA_signal_5723, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15}), .clk (clk), .r ({Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_6060, new_AGEMA_signal_6059, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M12_U1 ( .a ({new_AGEMA_signal_5324, new_AGEMA_signal_5323, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}), .b ({new_AGEMA_signal_5732, new_AGEMA_signal_5731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453]}), .c ({new_AGEMA_signal_6062, new_AGEMA_signal_6061, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M13_U1 ( .a ({new_AGEMA_signal_6062, new_AGEMA_signal_6061, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12}), .b ({new_AGEMA_signal_6060, new_AGEMA_signal_6059, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_6572, new_AGEMA_signal_6571, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M14_U1 ( .a ({new_AGEMA_signal_5320, new_AGEMA_signal_5319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6040, new_AGEMA_signal_6039, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}), .clk (clk), .r ({Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_6574, new_AGEMA_signal_6573, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M15_U1 ( .a ({new_AGEMA_signal_6574, new_AGEMA_signal_6573, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14}), .b ({new_AGEMA_signal_6060, new_AGEMA_signal_6059, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_6920, new_AGEMA_signal_6919, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M16_U1 ( .a ({new_AGEMA_signal_6564, new_AGEMA_signal_6563, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3}), .b ({new_AGEMA_signal_6562, new_AGEMA_signal_6561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2}), .c ({new_AGEMA_signal_6922, new_AGEMA_signal_6921, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M17_U1 ( .a ({new_AGEMA_signal_6566, new_AGEMA_signal_6565, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5}), .b ({new_AGEMA_signal_6558, new_AGEMA_signal_6557, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24}), .c ({new_AGEMA_signal_6924, new_AGEMA_signal_6923, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M18_U1 ( .a ({new_AGEMA_signal_6568, new_AGEMA_signal_6567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8}), .b ({new_AGEMA_signal_6058, new_AGEMA_signal_6057, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7}), .c ({new_AGEMA_signal_6926, new_AGEMA_signal_6925, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M19_U1 ( .a ({new_AGEMA_signal_6918, new_AGEMA_signal_6917, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10}), .b ({new_AGEMA_signal_6920, new_AGEMA_signal_6919, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_7118, new_AGEMA_signal_7117, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M20_U1 ( .a ({new_AGEMA_signal_6922, new_AGEMA_signal_6921, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16}), .b ({new_AGEMA_signal_6572, new_AGEMA_signal_6571, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_7120, new_AGEMA_signal_7119, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M21_U1 ( .a ({new_AGEMA_signal_6924, new_AGEMA_signal_6923, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17}), .b ({new_AGEMA_signal_6920, new_AGEMA_signal_6919, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_7122, new_AGEMA_signal_7121, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M22_U1 ( .a ({new_AGEMA_signal_6926, new_AGEMA_signal_6925, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18}), .b ({new_AGEMA_signal_6572, new_AGEMA_signal_6571, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_7124, new_AGEMA_signal_7123, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M23_U1 ( .a ({new_AGEMA_signal_7118, new_AGEMA_signal_7117, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19}), .b ({new_AGEMA_signal_6560, new_AGEMA_signal_6559, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25}), .c ({new_AGEMA_signal_7278, new_AGEMA_signal_7277, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M24_U1 ( .a ({new_AGEMA_signal_7124, new_AGEMA_signal_7123, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_7278, new_AGEMA_signal_7277, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}), .c ({new_AGEMA_signal_7438, new_AGEMA_signal_7437, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M27_U1 ( .a ({new_AGEMA_signal_7120, new_AGEMA_signal_7119, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_7122, new_AGEMA_signal_7121, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}), .c ({new_AGEMA_signal_7282, new_AGEMA_signal_7281, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M1_U1 ( .a ({new_AGEMA_signal_5738, new_AGEMA_signal_5737, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13}), .b ({new_AGEMA_signal_5734, new_AGEMA_signal_5733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459]}), .c ({new_AGEMA_signal_6078, new_AGEMA_signal_6077, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M2_U1 ( .a ({new_AGEMA_signal_6074, new_AGEMA_signal_6073, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23}), .b ({new_AGEMA_signal_6064, new_AGEMA_signal_6063, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8}), .clk (clk), .r ({Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_6580, new_AGEMA_signal_6579, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M3_U1 ( .a ({new_AGEMA_signal_6068, new_AGEMA_signal_6067, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14}), .b ({new_AGEMA_signal_6078, new_AGEMA_signal_6077, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_6582, new_AGEMA_signal_6581, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M4_U1 ( .a ({new_AGEMA_signal_5744, new_AGEMA_signal_5743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}), .b ({new_AGEMA_signal_5248, new_AGEMA_signal_5247, RoundKey[8]}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465]}), .c ({new_AGEMA_signal_6080, new_AGEMA_signal_6079, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M5_U1 ( .a ({new_AGEMA_signal_6080, new_AGEMA_signal_6079, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4}), .b ({new_AGEMA_signal_6078, new_AGEMA_signal_6077, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_6584, new_AGEMA_signal_6583, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M6_U1 ( .a ({new_AGEMA_signal_5342, new_AGEMA_signal_5341, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .clk (clk), .r ({Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_6082, new_AGEMA_signal_6081, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M7_U1 ( .a ({new_AGEMA_signal_5746, new_AGEMA_signal_5745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}), .b ({new_AGEMA_signal_5736, new_AGEMA_signal_5735, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471]}), .c ({new_AGEMA_signal_6084, new_AGEMA_signal_6083, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M8_U1 ( .a ({new_AGEMA_signal_6076, new_AGEMA_signal_6075, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26}), .b ({new_AGEMA_signal_6082, new_AGEMA_signal_6081, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_6586, new_AGEMA_signal_6585, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M9_U1 ( .a ({new_AGEMA_signal_6072, new_AGEMA_signal_6071, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_6070, new_AGEMA_signal_6069, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}), .clk (clk), .r ({Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_6588, new_AGEMA_signal_6587, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M10_U1 ( .a ({new_AGEMA_signal_6588, new_AGEMA_signal_6587, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9}), .b ({new_AGEMA_signal_6082, new_AGEMA_signal_6081, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_6928, new_AGEMA_signal_6927, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M11_U1 ( .a ({new_AGEMA_signal_5338, new_AGEMA_signal_5337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5740, new_AGEMA_signal_5739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477]}), .c ({new_AGEMA_signal_6086, new_AGEMA_signal_6085, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M12_U1 ( .a ({new_AGEMA_signal_5344, new_AGEMA_signal_5343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}), .b ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27}), .clk (clk), .r ({Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_6088, new_AGEMA_signal_6087, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M13_U1 ( .a ({new_AGEMA_signal_6088, new_AGEMA_signal_6087, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12}), .b ({new_AGEMA_signal_6086, new_AGEMA_signal_6085, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_6590, new_AGEMA_signal_6589, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M14_U1 ( .a ({new_AGEMA_signal_5340, new_AGEMA_signal_5339, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6066, new_AGEMA_signal_6065, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483]}), .c ({new_AGEMA_signal_6592, new_AGEMA_signal_6591, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M15_U1 ( .a ({new_AGEMA_signal_6592, new_AGEMA_signal_6591, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14}), .b ({new_AGEMA_signal_6086, new_AGEMA_signal_6085, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_6930, new_AGEMA_signal_6929, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M16_U1 ( .a ({new_AGEMA_signal_6582, new_AGEMA_signal_6581, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3}), .b ({new_AGEMA_signal_6580, new_AGEMA_signal_6579, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2}), .c ({new_AGEMA_signal_6932, new_AGEMA_signal_6931, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M17_U1 ( .a ({new_AGEMA_signal_6584, new_AGEMA_signal_6583, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5}), .b ({new_AGEMA_signal_6576, new_AGEMA_signal_6575, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24}), .c ({new_AGEMA_signal_6934, new_AGEMA_signal_6933, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M18_U1 ( .a ({new_AGEMA_signal_6586, new_AGEMA_signal_6585, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8}), .b ({new_AGEMA_signal_6084, new_AGEMA_signal_6083, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7}), .c ({new_AGEMA_signal_6936, new_AGEMA_signal_6935, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M19_U1 ( .a ({new_AGEMA_signal_6928, new_AGEMA_signal_6927, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10}), .b ({new_AGEMA_signal_6930, new_AGEMA_signal_6929, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_7126, new_AGEMA_signal_7125, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M20_U1 ( .a ({new_AGEMA_signal_6932, new_AGEMA_signal_6931, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16}), .b ({new_AGEMA_signal_6590, new_AGEMA_signal_6589, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_7128, new_AGEMA_signal_7127, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M21_U1 ( .a ({new_AGEMA_signal_6934, new_AGEMA_signal_6933, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17}), .b ({new_AGEMA_signal_6930, new_AGEMA_signal_6929, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_7130, new_AGEMA_signal_7129, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M22_U1 ( .a ({new_AGEMA_signal_6936, new_AGEMA_signal_6935, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18}), .b ({new_AGEMA_signal_6590, new_AGEMA_signal_6589, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_7132, new_AGEMA_signal_7131, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M23_U1 ( .a ({new_AGEMA_signal_7126, new_AGEMA_signal_7125, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19}), .b ({new_AGEMA_signal_6578, new_AGEMA_signal_6577, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25}), .c ({new_AGEMA_signal_7286, new_AGEMA_signal_7285, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M24_U1 ( .a ({new_AGEMA_signal_7132, new_AGEMA_signal_7131, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_7286, new_AGEMA_signal_7285, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}), .c ({new_AGEMA_signal_7448, new_AGEMA_signal_7447, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M27_U1 ( .a ({new_AGEMA_signal_7128, new_AGEMA_signal_7127, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_7130, new_AGEMA_signal_7129, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}), .c ({new_AGEMA_signal_7290, new_AGEMA_signal_7289, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M1_U1 ( .a ({new_AGEMA_signal_5754, new_AGEMA_signal_5753, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13}), .b ({new_AGEMA_signal_5750, new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .clk (clk), .r ({Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_6104, new_AGEMA_signal_6103, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M2_U1 ( .a ({new_AGEMA_signal_6100, new_AGEMA_signal_6099, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23}), .b ({new_AGEMA_signal_6090, new_AGEMA_signal_6089, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489]}), .c ({new_AGEMA_signal_6598, new_AGEMA_signal_6597, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M3_U1 ( .a ({new_AGEMA_signal_6094, new_AGEMA_signal_6093, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14}), .b ({new_AGEMA_signal_6104, new_AGEMA_signal_6103, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_6600, new_AGEMA_signal_6599, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M4_U1 ( .a ({new_AGEMA_signal_5760, new_AGEMA_signal_5759, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}), .b ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, RoundKey[0]}), .clk (clk), .r ({Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_6106, new_AGEMA_signal_6105, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M5_U1 ( .a ({new_AGEMA_signal_6106, new_AGEMA_signal_6105, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4}), .b ({new_AGEMA_signal_6104, new_AGEMA_signal_6103, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_6602, new_AGEMA_signal_6601, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M6_U1 ( .a ({new_AGEMA_signal_5362, new_AGEMA_signal_5361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5758, new_AGEMA_signal_5757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495]}), .c ({new_AGEMA_signal_6108, new_AGEMA_signal_6107, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M7_U1 ( .a ({new_AGEMA_signal_5762, new_AGEMA_signal_5761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}), .b ({new_AGEMA_signal_5752, new_AGEMA_signal_5751, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}), .clk (clk), .r ({Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_6110, new_AGEMA_signal_6109, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M8_U1 ( .a ({new_AGEMA_signal_6102, new_AGEMA_signal_6101, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26}), .b ({new_AGEMA_signal_6108, new_AGEMA_signal_6107, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_6604, new_AGEMA_signal_6603, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M9_U1 ( .a ({new_AGEMA_signal_6098, new_AGEMA_signal_6097, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_6096, new_AGEMA_signal_6095, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501]}), .c ({new_AGEMA_signal_6606, new_AGEMA_signal_6605, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M10_U1 ( .a ({new_AGEMA_signal_6606, new_AGEMA_signal_6605, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9}), .b ({new_AGEMA_signal_6108, new_AGEMA_signal_6107, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_6938, new_AGEMA_signal_6937, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M11_U1 ( .a ({new_AGEMA_signal_5358, new_AGEMA_signal_5357, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5756, new_AGEMA_signal_5755, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15}), .clk (clk), .r ({Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_6112, new_AGEMA_signal_6111, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M12_U1 ( .a ({new_AGEMA_signal_5364, new_AGEMA_signal_5363, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}), .b ({new_AGEMA_signal_5764, new_AGEMA_signal_5763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507]}), .c ({new_AGEMA_signal_6114, new_AGEMA_signal_6113, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M13_U1 ( .a ({new_AGEMA_signal_6114, new_AGEMA_signal_6113, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12}), .b ({new_AGEMA_signal_6112, new_AGEMA_signal_6111, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_6608, new_AGEMA_signal_6607, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M14_U1 ( .a ({new_AGEMA_signal_5360, new_AGEMA_signal_5359, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_6092, new_AGEMA_signal_6091, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}), .clk (clk), .r ({Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_6610, new_AGEMA_signal_6609, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M15_U1 ( .a ({new_AGEMA_signal_6610, new_AGEMA_signal_6609, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14}), .b ({new_AGEMA_signal_6112, new_AGEMA_signal_6111, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_6940, new_AGEMA_signal_6939, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M16_U1 ( .a ({new_AGEMA_signal_6600, new_AGEMA_signal_6599, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3}), .b ({new_AGEMA_signal_6598, new_AGEMA_signal_6597, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2}), .c ({new_AGEMA_signal_6942, new_AGEMA_signal_6941, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M17_U1 ( .a ({new_AGEMA_signal_6602, new_AGEMA_signal_6601, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5}), .b ({new_AGEMA_signal_6594, new_AGEMA_signal_6593, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24}), .c ({new_AGEMA_signal_6944, new_AGEMA_signal_6943, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M18_U1 ( .a ({new_AGEMA_signal_6604, new_AGEMA_signal_6603, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8}), .b ({new_AGEMA_signal_6110, new_AGEMA_signal_6109, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7}), .c ({new_AGEMA_signal_6946, new_AGEMA_signal_6945, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M19_U1 ( .a ({new_AGEMA_signal_6938, new_AGEMA_signal_6937, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10}), .b ({new_AGEMA_signal_6940, new_AGEMA_signal_6939, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_7134, new_AGEMA_signal_7133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M20_U1 ( .a ({new_AGEMA_signal_6942, new_AGEMA_signal_6941, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16}), .b ({new_AGEMA_signal_6608, new_AGEMA_signal_6607, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_7136, new_AGEMA_signal_7135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M21_U1 ( .a ({new_AGEMA_signal_6944, new_AGEMA_signal_6943, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17}), .b ({new_AGEMA_signal_6940, new_AGEMA_signal_6939, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_7138, new_AGEMA_signal_7137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M22_U1 ( .a ({new_AGEMA_signal_6946, new_AGEMA_signal_6945, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18}), .b ({new_AGEMA_signal_6608, new_AGEMA_signal_6607, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_7140, new_AGEMA_signal_7139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M23_U1 ( .a ({new_AGEMA_signal_7134, new_AGEMA_signal_7133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19}), .b ({new_AGEMA_signal_6596, new_AGEMA_signal_6595, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25}), .c ({new_AGEMA_signal_7294, new_AGEMA_signal_7293, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M24_U1 ( .a ({new_AGEMA_signal_7140, new_AGEMA_signal_7139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_7294, new_AGEMA_signal_7293, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}), .c ({new_AGEMA_signal_7458, new_AGEMA_signal_7457, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M27_U1 ( .a ({new_AGEMA_signal_7136, new_AGEMA_signal_7135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_7138, new_AGEMA_signal_7137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}), .c ({new_AGEMA_signal_7298, new_AGEMA_signal_7297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M1_U1 ( .a ({new_AGEMA_signal_5770, new_AGEMA_signal_5769, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13}), .b ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513]}), .c ({new_AGEMA_signal_6130, new_AGEMA_signal_6129, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M2_U1 ( .a ({new_AGEMA_signal_6126, new_AGEMA_signal_6125, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23}), .b ({new_AGEMA_signal_6116, new_AGEMA_signal_6115, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8}), .clk (clk), .r ({Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_6616, new_AGEMA_signal_6615, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M3_U1 ( .a ({new_AGEMA_signal_6120, new_AGEMA_signal_6119, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14}), .b ({new_AGEMA_signal_6130, new_AGEMA_signal_6129, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_6618, new_AGEMA_signal_6617, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M4_U1 ( .a ({new_AGEMA_signal_5776, new_AGEMA_signal_5775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}), .b ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, RoundKey[24]}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519]}), .c ({new_AGEMA_signal_6132, new_AGEMA_signal_6131, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M5_U1 ( .a ({new_AGEMA_signal_6132, new_AGEMA_signal_6131, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4}), .b ({new_AGEMA_signal_6130, new_AGEMA_signal_6129, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_6620, new_AGEMA_signal_6619, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M6_U1 ( .a ({new_AGEMA_signal_5382, new_AGEMA_signal_5381, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5774, new_AGEMA_signal_5773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .clk (clk), .r ({Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_6134, new_AGEMA_signal_6133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M7_U1 ( .a ({new_AGEMA_signal_5778, new_AGEMA_signal_5777, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}), .b ({new_AGEMA_signal_5768, new_AGEMA_signal_5767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525]}), .c ({new_AGEMA_signal_6136, new_AGEMA_signal_6135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M8_U1 ( .a ({new_AGEMA_signal_6128, new_AGEMA_signal_6127, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26}), .b ({new_AGEMA_signal_6134, new_AGEMA_signal_6133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_6622, new_AGEMA_signal_6621, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M9_U1 ( .a ({new_AGEMA_signal_6124, new_AGEMA_signal_6123, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_6122, new_AGEMA_signal_6121, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}), .clk (clk), .r ({Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_6624, new_AGEMA_signal_6623, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M10_U1 ( .a ({new_AGEMA_signal_6624, new_AGEMA_signal_6623, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9}), .b ({new_AGEMA_signal_6134, new_AGEMA_signal_6133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_6948, new_AGEMA_signal_6947, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M11_U1 ( .a ({new_AGEMA_signal_5378, new_AGEMA_signal_5377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5772, new_AGEMA_signal_5771, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531]}), .c ({new_AGEMA_signal_6138, new_AGEMA_signal_6137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M12_U1 ( .a ({new_AGEMA_signal_5384, new_AGEMA_signal_5383, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}), .b ({new_AGEMA_signal_5780, new_AGEMA_signal_5779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27}), .clk (clk), .r ({Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_6140, new_AGEMA_signal_6139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M13_U1 ( .a ({new_AGEMA_signal_6140, new_AGEMA_signal_6139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12}), .b ({new_AGEMA_signal_6138, new_AGEMA_signal_6137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_6626, new_AGEMA_signal_6625, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M14_U1 ( .a ({new_AGEMA_signal_5380, new_AGEMA_signal_5379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_6118, new_AGEMA_signal_6117, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537]}), .c ({new_AGEMA_signal_6628, new_AGEMA_signal_6627, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M15_U1 ( .a ({new_AGEMA_signal_6628, new_AGEMA_signal_6627, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14}), .b ({new_AGEMA_signal_6138, new_AGEMA_signal_6137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_6950, new_AGEMA_signal_6949, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M16_U1 ( .a ({new_AGEMA_signal_6618, new_AGEMA_signal_6617, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3}), .b ({new_AGEMA_signal_6616, new_AGEMA_signal_6615, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2}), .c ({new_AGEMA_signal_6952, new_AGEMA_signal_6951, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M17_U1 ( .a ({new_AGEMA_signal_6620, new_AGEMA_signal_6619, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5}), .b ({new_AGEMA_signal_6612, new_AGEMA_signal_6611, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24}), .c ({new_AGEMA_signal_6954, new_AGEMA_signal_6953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M18_U1 ( .a ({new_AGEMA_signal_6622, new_AGEMA_signal_6621, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8}), .b ({new_AGEMA_signal_6136, new_AGEMA_signal_6135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7}), .c ({new_AGEMA_signal_6956, new_AGEMA_signal_6955, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M19_U1 ( .a ({new_AGEMA_signal_6948, new_AGEMA_signal_6947, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10}), .b ({new_AGEMA_signal_6950, new_AGEMA_signal_6949, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_7142, new_AGEMA_signal_7141, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M20_U1 ( .a ({new_AGEMA_signal_6952, new_AGEMA_signal_6951, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16}), .b ({new_AGEMA_signal_6626, new_AGEMA_signal_6625, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_7144, new_AGEMA_signal_7143, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M21_U1 ( .a ({new_AGEMA_signal_6954, new_AGEMA_signal_6953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17}), .b ({new_AGEMA_signal_6950, new_AGEMA_signal_6949, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_7146, new_AGEMA_signal_7145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M22_U1 ( .a ({new_AGEMA_signal_6956, new_AGEMA_signal_6955, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18}), .b ({new_AGEMA_signal_6626, new_AGEMA_signal_6625, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_7148, new_AGEMA_signal_7147, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M23_U1 ( .a ({new_AGEMA_signal_7142, new_AGEMA_signal_7141, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19}), .b ({new_AGEMA_signal_6614, new_AGEMA_signal_6613, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25}), .c ({new_AGEMA_signal_7302, new_AGEMA_signal_7301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M24_U1 ( .a ({new_AGEMA_signal_7148, new_AGEMA_signal_7147, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_7302, new_AGEMA_signal_7301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}), .c ({new_AGEMA_signal_7468, new_AGEMA_signal_7467, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M27_U1 ( .a ({new_AGEMA_signal_7144, new_AGEMA_signal_7143, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_7146, new_AGEMA_signal_7145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}), .c ({new_AGEMA_signal_7306, new_AGEMA_signal_7305, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M25_U1 ( .a ({new_AGEMA_signal_7156, new_AGEMA_signal_7155, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_7152, new_AGEMA_signal_7151, SubBytesIns_Inst_Sbox_0_M20}), .clk (clk), .r ({Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_7312, new_AGEMA_signal_7311, SubBytesIns_Inst_Sbox_0_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M26_U1 ( .a ({new_AGEMA_signal_7154, new_AGEMA_signal_7153, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_7312, new_AGEMA_signal_7311, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_7480, new_AGEMA_signal_7479, SubBytesIns_Inst_Sbox_0_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M28_U1 ( .a ({new_AGEMA_signal_7310, new_AGEMA_signal_7309, SubBytesIns_Inst_Sbox_0_M23}), .b ({new_AGEMA_signal_7312, new_AGEMA_signal_7311, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_7482, new_AGEMA_signal_7481, SubBytesIns_Inst_Sbox_0_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M31_U1 ( .a ({new_AGEMA_signal_7152, new_AGEMA_signal_7151, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_7310, new_AGEMA_signal_7309, SubBytesIns_Inst_Sbox_0_M23}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543]}), .c ({new_AGEMA_signal_7484, new_AGEMA_signal_7483, SubBytesIns_Inst_Sbox_0_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M33_U1 ( .a ({new_AGEMA_signal_7314, new_AGEMA_signal_7313, SubBytesIns_Inst_Sbox_0_M27}), .b ({new_AGEMA_signal_7312, new_AGEMA_signal_7311, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_7486, new_AGEMA_signal_7485, SubBytesIns_Inst_Sbox_0_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M34_U1 ( .a ({new_AGEMA_signal_7154, new_AGEMA_signal_7153, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_7156, new_AGEMA_signal_7155, SubBytesIns_Inst_Sbox_0_M22}), .clk (clk), .r ({Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_7316, new_AGEMA_signal_7315, SubBytesIns_Inst_Sbox_0_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M36_U1 ( .a ({new_AGEMA_signal_7478, new_AGEMA_signal_7477, SubBytesIns_Inst_Sbox_0_M24}), .b ({new_AGEMA_signal_7312, new_AGEMA_signal_7311, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_7686, new_AGEMA_signal_7685, SubBytesIns_Inst_Sbox_0_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M25_U1 ( .a ({new_AGEMA_signal_7164, new_AGEMA_signal_7163, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_7160, new_AGEMA_signal_7159, SubBytesIns_Inst_Sbox_1_M20}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549]}), .c ({new_AGEMA_signal_7320, new_AGEMA_signal_7319, SubBytesIns_Inst_Sbox_1_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M26_U1 ( .a ({new_AGEMA_signal_7162, new_AGEMA_signal_7161, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_7320, new_AGEMA_signal_7319, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_7490, new_AGEMA_signal_7489, SubBytesIns_Inst_Sbox_1_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M28_U1 ( .a ({new_AGEMA_signal_7318, new_AGEMA_signal_7317, SubBytesIns_Inst_Sbox_1_M23}), .b ({new_AGEMA_signal_7320, new_AGEMA_signal_7319, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_7492, new_AGEMA_signal_7491, SubBytesIns_Inst_Sbox_1_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M31_U1 ( .a ({new_AGEMA_signal_7160, new_AGEMA_signal_7159, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_7318, new_AGEMA_signal_7317, SubBytesIns_Inst_Sbox_1_M23}), .clk (clk), .r ({Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_7494, new_AGEMA_signal_7493, SubBytesIns_Inst_Sbox_1_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M33_U1 ( .a ({new_AGEMA_signal_7322, new_AGEMA_signal_7321, SubBytesIns_Inst_Sbox_1_M27}), .b ({new_AGEMA_signal_7320, new_AGEMA_signal_7319, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_7496, new_AGEMA_signal_7495, SubBytesIns_Inst_Sbox_1_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M34_U1 ( .a ({new_AGEMA_signal_7162, new_AGEMA_signal_7161, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_7164, new_AGEMA_signal_7163, SubBytesIns_Inst_Sbox_1_M22}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555]}), .c ({new_AGEMA_signal_7324, new_AGEMA_signal_7323, SubBytesIns_Inst_Sbox_1_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M36_U1 ( .a ({new_AGEMA_signal_7488, new_AGEMA_signal_7487, SubBytesIns_Inst_Sbox_1_M24}), .b ({new_AGEMA_signal_7320, new_AGEMA_signal_7319, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_7696, new_AGEMA_signal_7695, SubBytesIns_Inst_Sbox_1_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M25_U1 ( .a ({new_AGEMA_signal_7172, new_AGEMA_signal_7171, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_7168, new_AGEMA_signal_7167, SubBytesIns_Inst_Sbox_2_M20}), .clk (clk), .r ({Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_7328, new_AGEMA_signal_7327, SubBytesIns_Inst_Sbox_2_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M26_U1 ( .a ({new_AGEMA_signal_7170, new_AGEMA_signal_7169, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_7328, new_AGEMA_signal_7327, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_7500, new_AGEMA_signal_7499, SubBytesIns_Inst_Sbox_2_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M28_U1 ( .a ({new_AGEMA_signal_7326, new_AGEMA_signal_7325, SubBytesIns_Inst_Sbox_2_M23}), .b ({new_AGEMA_signal_7328, new_AGEMA_signal_7327, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_7502, new_AGEMA_signal_7501, SubBytesIns_Inst_Sbox_2_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M31_U1 ( .a ({new_AGEMA_signal_7168, new_AGEMA_signal_7167, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_7326, new_AGEMA_signal_7325, SubBytesIns_Inst_Sbox_2_M23}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561]}), .c ({new_AGEMA_signal_7504, new_AGEMA_signal_7503, SubBytesIns_Inst_Sbox_2_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M33_U1 ( .a ({new_AGEMA_signal_7330, new_AGEMA_signal_7329, SubBytesIns_Inst_Sbox_2_M27}), .b ({new_AGEMA_signal_7328, new_AGEMA_signal_7327, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_7506, new_AGEMA_signal_7505, SubBytesIns_Inst_Sbox_2_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M34_U1 ( .a ({new_AGEMA_signal_7170, new_AGEMA_signal_7169, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_7172, new_AGEMA_signal_7171, SubBytesIns_Inst_Sbox_2_M22}), .clk (clk), .r ({Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_7332, new_AGEMA_signal_7331, SubBytesIns_Inst_Sbox_2_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M36_U1 ( .a ({new_AGEMA_signal_7498, new_AGEMA_signal_7497, SubBytesIns_Inst_Sbox_2_M24}), .b ({new_AGEMA_signal_7328, new_AGEMA_signal_7327, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_7706, new_AGEMA_signal_7705, SubBytesIns_Inst_Sbox_2_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M25_U1 ( .a ({new_AGEMA_signal_7180, new_AGEMA_signal_7179, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_7176, new_AGEMA_signal_7175, SubBytesIns_Inst_Sbox_3_M20}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567]}), .c ({new_AGEMA_signal_7336, new_AGEMA_signal_7335, SubBytesIns_Inst_Sbox_3_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M26_U1 ( .a ({new_AGEMA_signal_7178, new_AGEMA_signal_7177, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_7336, new_AGEMA_signal_7335, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_7510, new_AGEMA_signal_7509, SubBytesIns_Inst_Sbox_3_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M28_U1 ( .a ({new_AGEMA_signal_7334, new_AGEMA_signal_7333, SubBytesIns_Inst_Sbox_3_M23}), .b ({new_AGEMA_signal_7336, new_AGEMA_signal_7335, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_7512, new_AGEMA_signal_7511, SubBytesIns_Inst_Sbox_3_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M31_U1 ( .a ({new_AGEMA_signal_7176, new_AGEMA_signal_7175, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_7334, new_AGEMA_signal_7333, SubBytesIns_Inst_Sbox_3_M23}), .clk (clk), .r ({Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_7514, new_AGEMA_signal_7513, SubBytesIns_Inst_Sbox_3_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M33_U1 ( .a ({new_AGEMA_signal_7338, new_AGEMA_signal_7337, SubBytesIns_Inst_Sbox_3_M27}), .b ({new_AGEMA_signal_7336, new_AGEMA_signal_7335, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_7516, new_AGEMA_signal_7515, SubBytesIns_Inst_Sbox_3_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M34_U1 ( .a ({new_AGEMA_signal_7178, new_AGEMA_signal_7177, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_7180, new_AGEMA_signal_7179, SubBytesIns_Inst_Sbox_3_M22}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573]}), .c ({new_AGEMA_signal_7340, new_AGEMA_signal_7339, SubBytesIns_Inst_Sbox_3_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M36_U1 ( .a ({new_AGEMA_signal_7508, new_AGEMA_signal_7507, SubBytesIns_Inst_Sbox_3_M24}), .b ({new_AGEMA_signal_7336, new_AGEMA_signal_7335, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_7716, new_AGEMA_signal_7715, SubBytesIns_Inst_Sbox_3_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M25_U1 ( .a ({new_AGEMA_signal_7188, new_AGEMA_signal_7187, SubBytesIns_Inst_Sbox_4_M22}), .b ({new_AGEMA_signal_7184, new_AGEMA_signal_7183, SubBytesIns_Inst_Sbox_4_M20}), .clk (clk), .r ({Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_7344, new_AGEMA_signal_7343, SubBytesIns_Inst_Sbox_4_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M26_U1 ( .a ({new_AGEMA_signal_7186, new_AGEMA_signal_7185, SubBytesIns_Inst_Sbox_4_M21}), .b ({new_AGEMA_signal_7344, new_AGEMA_signal_7343, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_7520, new_AGEMA_signal_7519, SubBytesIns_Inst_Sbox_4_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M28_U1 ( .a ({new_AGEMA_signal_7342, new_AGEMA_signal_7341, SubBytesIns_Inst_Sbox_4_M23}), .b ({new_AGEMA_signal_7344, new_AGEMA_signal_7343, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_7522, new_AGEMA_signal_7521, SubBytesIns_Inst_Sbox_4_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M31_U1 ( .a ({new_AGEMA_signal_7184, new_AGEMA_signal_7183, SubBytesIns_Inst_Sbox_4_M20}), .b ({new_AGEMA_signal_7342, new_AGEMA_signal_7341, SubBytesIns_Inst_Sbox_4_M23}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579]}), .c ({new_AGEMA_signal_7524, new_AGEMA_signal_7523, SubBytesIns_Inst_Sbox_4_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M33_U1 ( .a ({new_AGEMA_signal_7346, new_AGEMA_signal_7345, SubBytesIns_Inst_Sbox_4_M27}), .b ({new_AGEMA_signal_7344, new_AGEMA_signal_7343, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_7526, new_AGEMA_signal_7525, SubBytesIns_Inst_Sbox_4_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M34_U1 ( .a ({new_AGEMA_signal_7186, new_AGEMA_signal_7185, SubBytesIns_Inst_Sbox_4_M21}), .b ({new_AGEMA_signal_7188, new_AGEMA_signal_7187, SubBytesIns_Inst_Sbox_4_M22}), .clk (clk), .r ({Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_7348, new_AGEMA_signal_7347, SubBytesIns_Inst_Sbox_4_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M36_U1 ( .a ({new_AGEMA_signal_7518, new_AGEMA_signal_7517, SubBytesIns_Inst_Sbox_4_M24}), .b ({new_AGEMA_signal_7344, new_AGEMA_signal_7343, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_7726, new_AGEMA_signal_7725, SubBytesIns_Inst_Sbox_4_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M25_U1 ( .a ({new_AGEMA_signal_7196, new_AGEMA_signal_7195, SubBytesIns_Inst_Sbox_5_M22}), .b ({new_AGEMA_signal_7192, new_AGEMA_signal_7191, SubBytesIns_Inst_Sbox_5_M20}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585]}), .c ({new_AGEMA_signal_7352, new_AGEMA_signal_7351, SubBytesIns_Inst_Sbox_5_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M26_U1 ( .a ({new_AGEMA_signal_7194, new_AGEMA_signal_7193, SubBytesIns_Inst_Sbox_5_M21}), .b ({new_AGEMA_signal_7352, new_AGEMA_signal_7351, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_7530, new_AGEMA_signal_7529, SubBytesIns_Inst_Sbox_5_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M28_U1 ( .a ({new_AGEMA_signal_7350, new_AGEMA_signal_7349, SubBytesIns_Inst_Sbox_5_M23}), .b ({new_AGEMA_signal_7352, new_AGEMA_signal_7351, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_7532, new_AGEMA_signal_7531, SubBytesIns_Inst_Sbox_5_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M31_U1 ( .a ({new_AGEMA_signal_7192, new_AGEMA_signal_7191, SubBytesIns_Inst_Sbox_5_M20}), .b ({new_AGEMA_signal_7350, new_AGEMA_signal_7349, SubBytesIns_Inst_Sbox_5_M23}), .clk (clk), .r ({Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_7534, new_AGEMA_signal_7533, SubBytesIns_Inst_Sbox_5_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M33_U1 ( .a ({new_AGEMA_signal_7354, new_AGEMA_signal_7353, SubBytesIns_Inst_Sbox_5_M27}), .b ({new_AGEMA_signal_7352, new_AGEMA_signal_7351, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_7536, new_AGEMA_signal_7535, SubBytesIns_Inst_Sbox_5_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M34_U1 ( .a ({new_AGEMA_signal_7194, new_AGEMA_signal_7193, SubBytesIns_Inst_Sbox_5_M21}), .b ({new_AGEMA_signal_7196, new_AGEMA_signal_7195, SubBytesIns_Inst_Sbox_5_M22}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591]}), .c ({new_AGEMA_signal_7356, new_AGEMA_signal_7355, SubBytesIns_Inst_Sbox_5_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M36_U1 ( .a ({new_AGEMA_signal_7528, new_AGEMA_signal_7527, SubBytesIns_Inst_Sbox_5_M24}), .b ({new_AGEMA_signal_7352, new_AGEMA_signal_7351, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_7736, new_AGEMA_signal_7735, SubBytesIns_Inst_Sbox_5_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M25_U1 ( .a ({new_AGEMA_signal_7204, new_AGEMA_signal_7203, SubBytesIns_Inst_Sbox_6_M22}), .b ({new_AGEMA_signal_7200, new_AGEMA_signal_7199, SubBytesIns_Inst_Sbox_6_M20}), .clk (clk), .r ({Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_7360, new_AGEMA_signal_7359, SubBytesIns_Inst_Sbox_6_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M26_U1 ( .a ({new_AGEMA_signal_7202, new_AGEMA_signal_7201, SubBytesIns_Inst_Sbox_6_M21}), .b ({new_AGEMA_signal_7360, new_AGEMA_signal_7359, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_7540, new_AGEMA_signal_7539, SubBytesIns_Inst_Sbox_6_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M28_U1 ( .a ({new_AGEMA_signal_7358, new_AGEMA_signal_7357, SubBytesIns_Inst_Sbox_6_M23}), .b ({new_AGEMA_signal_7360, new_AGEMA_signal_7359, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_7542, new_AGEMA_signal_7541, SubBytesIns_Inst_Sbox_6_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M31_U1 ( .a ({new_AGEMA_signal_7200, new_AGEMA_signal_7199, SubBytesIns_Inst_Sbox_6_M20}), .b ({new_AGEMA_signal_7358, new_AGEMA_signal_7357, SubBytesIns_Inst_Sbox_6_M23}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597]}), .c ({new_AGEMA_signal_7544, new_AGEMA_signal_7543, SubBytesIns_Inst_Sbox_6_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M33_U1 ( .a ({new_AGEMA_signal_7362, new_AGEMA_signal_7361, SubBytesIns_Inst_Sbox_6_M27}), .b ({new_AGEMA_signal_7360, new_AGEMA_signal_7359, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_7546, new_AGEMA_signal_7545, SubBytesIns_Inst_Sbox_6_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M34_U1 ( .a ({new_AGEMA_signal_7202, new_AGEMA_signal_7201, SubBytesIns_Inst_Sbox_6_M21}), .b ({new_AGEMA_signal_7204, new_AGEMA_signal_7203, SubBytesIns_Inst_Sbox_6_M22}), .clk (clk), .r ({Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_7364, new_AGEMA_signal_7363, SubBytesIns_Inst_Sbox_6_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M36_U1 ( .a ({new_AGEMA_signal_7538, new_AGEMA_signal_7537, SubBytesIns_Inst_Sbox_6_M24}), .b ({new_AGEMA_signal_7360, new_AGEMA_signal_7359, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_7746, new_AGEMA_signal_7745, SubBytesIns_Inst_Sbox_6_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M25_U1 ( .a ({new_AGEMA_signal_7212, new_AGEMA_signal_7211, SubBytesIns_Inst_Sbox_7_M22}), .b ({new_AGEMA_signal_7208, new_AGEMA_signal_7207, SubBytesIns_Inst_Sbox_7_M20}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603]}), .c ({new_AGEMA_signal_7368, new_AGEMA_signal_7367, SubBytesIns_Inst_Sbox_7_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M26_U1 ( .a ({new_AGEMA_signal_7210, new_AGEMA_signal_7209, SubBytesIns_Inst_Sbox_7_M21}), .b ({new_AGEMA_signal_7368, new_AGEMA_signal_7367, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_7550, new_AGEMA_signal_7549, SubBytesIns_Inst_Sbox_7_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M28_U1 ( .a ({new_AGEMA_signal_7366, new_AGEMA_signal_7365, SubBytesIns_Inst_Sbox_7_M23}), .b ({new_AGEMA_signal_7368, new_AGEMA_signal_7367, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_7552, new_AGEMA_signal_7551, SubBytesIns_Inst_Sbox_7_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M31_U1 ( .a ({new_AGEMA_signal_7208, new_AGEMA_signal_7207, SubBytesIns_Inst_Sbox_7_M20}), .b ({new_AGEMA_signal_7366, new_AGEMA_signal_7365, SubBytesIns_Inst_Sbox_7_M23}), .clk (clk), .r ({Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_7554, new_AGEMA_signal_7553, SubBytesIns_Inst_Sbox_7_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M33_U1 ( .a ({new_AGEMA_signal_7370, new_AGEMA_signal_7369, SubBytesIns_Inst_Sbox_7_M27}), .b ({new_AGEMA_signal_7368, new_AGEMA_signal_7367, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_7556, new_AGEMA_signal_7555, SubBytesIns_Inst_Sbox_7_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M34_U1 ( .a ({new_AGEMA_signal_7210, new_AGEMA_signal_7209, SubBytesIns_Inst_Sbox_7_M21}), .b ({new_AGEMA_signal_7212, new_AGEMA_signal_7211, SubBytesIns_Inst_Sbox_7_M22}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609]}), .c ({new_AGEMA_signal_7372, new_AGEMA_signal_7371, SubBytesIns_Inst_Sbox_7_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M36_U1 ( .a ({new_AGEMA_signal_7548, new_AGEMA_signal_7547, SubBytesIns_Inst_Sbox_7_M24}), .b ({new_AGEMA_signal_7368, new_AGEMA_signal_7367, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_7756, new_AGEMA_signal_7755, SubBytesIns_Inst_Sbox_7_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M25_U1 ( .a ({new_AGEMA_signal_7220, new_AGEMA_signal_7219, SubBytesIns_Inst_Sbox_8_M22}), .b ({new_AGEMA_signal_7216, new_AGEMA_signal_7215, SubBytesIns_Inst_Sbox_8_M20}), .clk (clk), .r ({Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_7376, new_AGEMA_signal_7375, SubBytesIns_Inst_Sbox_8_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M26_U1 ( .a ({new_AGEMA_signal_7218, new_AGEMA_signal_7217, SubBytesIns_Inst_Sbox_8_M21}), .b ({new_AGEMA_signal_7376, new_AGEMA_signal_7375, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_7560, new_AGEMA_signal_7559, SubBytesIns_Inst_Sbox_8_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M28_U1 ( .a ({new_AGEMA_signal_7374, new_AGEMA_signal_7373, SubBytesIns_Inst_Sbox_8_M23}), .b ({new_AGEMA_signal_7376, new_AGEMA_signal_7375, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_7562, new_AGEMA_signal_7561, SubBytesIns_Inst_Sbox_8_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M31_U1 ( .a ({new_AGEMA_signal_7216, new_AGEMA_signal_7215, SubBytesIns_Inst_Sbox_8_M20}), .b ({new_AGEMA_signal_7374, new_AGEMA_signal_7373, SubBytesIns_Inst_Sbox_8_M23}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615]}), .c ({new_AGEMA_signal_7564, new_AGEMA_signal_7563, SubBytesIns_Inst_Sbox_8_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M33_U1 ( .a ({new_AGEMA_signal_7378, new_AGEMA_signal_7377, SubBytesIns_Inst_Sbox_8_M27}), .b ({new_AGEMA_signal_7376, new_AGEMA_signal_7375, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_7566, new_AGEMA_signal_7565, SubBytesIns_Inst_Sbox_8_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M34_U1 ( .a ({new_AGEMA_signal_7218, new_AGEMA_signal_7217, SubBytesIns_Inst_Sbox_8_M21}), .b ({new_AGEMA_signal_7220, new_AGEMA_signal_7219, SubBytesIns_Inst_Sbox_8_M22}), .clk (clk), .r ({Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_7380, new_AGEMA_signal_7379, SubBytesIns_Inst_Sbox_8_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M36_U1 ( .a ({new_AGEMA_signal_7558, new_AGEMA_signal_7557, SubBytesIns_Inst_Sbox_8_M24}), .b ({new_AGEMA_signal_7376, new_AGEMA_signal_7375, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_7766, new_AGEMA_signal_7765, SubBytesIns_Inst_Sbox_8_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M25_U1 ( .a ({new_AGEMA_signal_7228, new_AGEMA_signal_7227, SubBytesIns_Inst_Sbox_9_M22}), .b ({new_AGEMA_signal_7224, new_AGEMA_signal_7223, SubBytesIns_Inst_Sbox_9_M20}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621]}), .c ({new_AGEMA_signal_7384, new_AGEMA_signal_7383, SubBytesIns_Inst_Sbox_9_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M26_U1 ( .a ({new_AGEMA_signal_7226, new_AGEMA_signal_7225, SubBytesIns_Inst_Sbox_9_M21}), .b ({new_AGEMA_signal_7384, new_AGEMA_signal_7383, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_7570, new_AGEMA_signal_7569, SubBytesIns_Inst_Sbox_9_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M28_U1 ( .a ({new_AGEMA_signal_7382, new_AGEMA_signal_7381, SubBytesIns_Inst_Sbox_9_M23}), .b ({new_AGEMA_signal_7384, new_AGEMA_signal_7383, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_7572, new_AGEMA_signal_7571, SubBytesIns_Inst_Sbox_9_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M31_U1 ( .a ({new_AGEMA_signal_7224, new_AGEMA_signal_7223, SubBytesIns_Inst_Sbox_9_M20}), .b ({new_AGEMA_signal_7382, new_AGEMA_signal_7381, SubBytesIns_Inst_Sbox_9_M23}), .clk (clk), .r ({Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_7574, new_AGEMA_signal_7573, SubBytesIns_Inst_Sbox_9_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M33_U1 ( .a ({new_AGEMA_signal_7386, new_AGEMA_signal_7385, SubBytesIns_Inst_Sbox_9_M27}), .b ({new_AGEMA_signal_7384, new_AGEMA_signal_7383, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_7576, new_AGEMA_signal_7575, SubBytesIns_Inst_Sbox_9_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M34_U1 ( .a ({new_AGEMA_signal_7226, new_AGEMA_signal_7225, SubBytesIns_Inst_Sbox_9_M21}), .b ({new_AGEMA_signal_7228, new_AGEMA_signal_7227, SubBytesIns_Inst_Sbox_9_M22}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627]}), .c ({new_AGEMA_signal_7388, new_AGEMA_signal_7387, SubBytesIns_Inst_Sbox_9_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M36_U1 ( .a ({new_AGEMA_signal_7568, new_AGEMA_signal_7567, SubBytesIns_Inst_Sbox_9_M24}), .b ({new_AGEMA_signal_7384, new_AGEMA_signal_7383, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_7776, new_AGEMA_signal_7775, SubBytesIns_Inst_Sbox_9_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M25_U1 ( .a ({new_AGEMA_signal_7236, new_AGEMA_signal_7235, SubBytesIns_Inst_Sbox_10_M22}), .b ({new_AGEMA_signal_7232, new_AGEMA_signal_7231, SubBytesIns_Inst_Sbox_10_M20}), .clk (clk), .r ({Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_7392, new_AGEMA_signal_7391, SubBytesIns_Inst_Sbox_10_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M26_U1 ( .a ({new_AGEMA_signal_7234, new_AGEMA_signal_7233, SubBytesIns_Inst_Sbox_10_M21}), .b ({new_AGEMA_signal_7392, new_AGEMA_signal_7391, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_7580, new_AGEMA_signal_7579, SubBytesIns_Inst_Sbox_10_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M28_U1 ( .a ({new_AGEMA_signal_7390, new_AGEMA_signal_7389, SubBytesIns_Inst_Sbox_10_M23}), .b ({new_AGEMA_signal_7392, new_AGEMA_signal_7391, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_7582, new_AGEMA_signal_7581, SubBytesIns_Inst_Sbox_10_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M31_U1 ( .a ({new_AGEMA_signal_7232, new_AGEMA_signal_7231, SubBytesIns_Inst_Sbox_10_M20}), .b ({new_AGEMA_signal_7390, new_AGEMA_signal_7389, SubBytesIns_Inst_Sbox_10_M23}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633]}), .c ({new_AGEMA_signal_7584, new_AGEMA_signal_7583, SubBytesIns_Inst_Sbox_10_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M33_U1 ( .a ({new_AGEMA_signal_7394, new_AGEMA_signal_7393, SubBytesIns_Inst_Sbox_10_M27}), .b ({new_AGEMA_signal_7392, new_AGEMA_signal_7391, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_7586, new_AGEMA_signal_7585, SubBytesIns_Inst_Sbox_10_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M34_U1 ( .a ({new_AGEMA_signal_7234, new_AGEMA_signal_7233, SubBytesIns_Inst_Sbox_10_M21}), .b ({new_AGEMA_signal_7236, new_AGEMA_signal_7235, SubBytesIns_Inst_Sbox_10_M22}), .clk (clk), .r ({Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_7396, new_AGEMA_signal_7395, SubBytesIns_Inst_Sbox_10_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M36_U1 ( .a ({new_AGEMA_signal_7578, new_AGEMA_signal_7577, SubBytesIns_Inst_Sbox_10_M24}), .b ({new_AGEMA_signal_7392, new_AGEMA_signal_7391, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_7786, new_AGEMA_signal_7785, SubBytesIns_Inst_Sbox_10_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M25_U1 ( .a ({new_AGEMA_signal_7244, new_AGEMA_signal_7243, SubBytesIns_Inst_Sbox_11_M22}), .b ({new_AGEMA_signal_7240, new_AGEMA_signal_7239, SubBytesIns_Inst_Sbox_11_M20}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639]}), .c ({new_AGEMA_signal_7400, new_AGEMA_signal_7399, SubBytesIns_Inst_Sbox_11_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M26_U1 ( .a ({new_AGEMA_signal_7242, new_AGEMA_signal_7241, SubBytesIns_Inst_Sbox_11_M21}), .b ({new_AGEMA_signal_7400, new_AGEMA_signal_7399, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_7590, new_AGEMA_signal_7589, SubBytesIns_Inst_Sbox_11_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M28_U1 ( .a ({new_AGEMA_signal_7398, new_AGEMA_signal_7397, SubBytesIns_Inst_Sbox_11_M23}), .b ({new_AGEMA_signal_7400, new_AGEMA_signal_7399, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_7592, new_AGEMA_signal_7591, SubBytesIns_Inst_Sbox_11_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M31_U1 ( .a ({new_AGEMA_signal_7240, new_AGEMA_signal_7239, SubBytesIns_Inst_Sbox_11_M20}), .b ({new_AGEMA_signal_7398, new_AGEMA_signal_7397, SubBytesIns_Inst_Sbox_11_M23}), .clk (clk), .r ({Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_7594, new_AGEMA_signal_7593, SubBytesIns_Inst_Sbox_11_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M33_U1 ( .a ({new_AGEMA_signal_7402, new_AGEMA_signal_7401, SubBytesIns_Inst_Sbox_11_M27}), .b ({new_AGEMA_signal_7400, new_AGEMA_signal_7399, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_7596, new_AGEMA_signal_7595, SubBytesIns_Inst_Sbox_11_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M34_U1 ( .a ({new_AGEMA_signal_7242, new_AGEMA_signal_7241, SubBytesIns_Inst_Sbox_11_M21}), .b ({new_AGEMA_signal_7244, new_AGEMA_signal_7243, SubBytesIns_Inst_Sbox_11_M22}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645]}), .c ({new_AGEMA_signal_7404, new_AGEMA_signal_7403, SubBytesIns_Inst_Sbox_11_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M36_U1 ( .a ({new_AGEMA_signal_7588, new_AGEMA_signal_7587, SubBytesIns_Inst_Sbox_11_M24}), .b ({new_AGEMA_signal_7400, new_AGEMA_signal_7399, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_7796, new_AGEMA_signal_7795, SubBytesIns_Inst_Sbox_11_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M25_U1 ( .a ({new_AGEMA_signal_7252, new_AGEMA_signal_7251, SubBytesIns_Inst_Sbox_12_M22}), .b ({new_AGEMA_signal_7248, new_AGEMA_signal_7247, SubBytesIns_Inst_Sbox_12_M20}), .clk (clk), .r ({Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_7408, new_AGEMA_signal_7407, SubBytesIns_Inst_Sbox_12_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M26_U1 ( .a ({new_AGEMA_signal_7250, new_AGEMA_signal_7249, SubBytesIns_Inst_Sbox_12_M21}), .b ({new_AGEMA_signal_7408, new_AGEMA_signal_7407, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_7600, new_AGEMA_signal_7599, SubBytesIns_Inst_Sbox_12_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M28_U1 ( .a ({new_AGEMA_signal_7406, new_AGEMA_signal_7405, SubBytesIns_Inst_Sbox_12_M23}), .b ({new_AGEMA_signal_7408, new_AGEMA_signal_7407, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_7602, new_AGEMA_signal_7601, SubBytesIns_Inst_Sbox_12_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M31_U1 ( .a ({new_AGEMA_signal_7248, new_AGEMA_signal_7247, SubBytesIns_Inst_Sbox_12_M20}), .b ({new_AGEMA_signal_7406, new_AGEMA_signal_7405, SubBytesIns_Inst_Sbox_12_M23}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651]}), .c ({new_AGEMA_signal_7604, new_AGEMA_signal_7603, SubBytesIns_Inst_Sbox_12_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M33_U1 ( .a ({new_AGEMA_signal_7410, new_AGEMA_signal_7409, SubBytesIns_Inst_Sbox_12_M27}), .b ({new_AGEMA_signal_7408, new_AGEMA_signal_7407, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_7606, new_AGEMA_signal_7605, SubBytesIns_Inst_Sbox_12_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M34_U1 ( .a ({new_AGEMA_signal_7250, new_AGEMA_signal_7249, SubBytesIns_Inst_Sbox_12_M21}), .b ({new_AGEMA_signal_7252, new_AGEMA_signal_7251, SubBytesIns_Inst_Sbox_12_M22}), .clk (clk), .r ({Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_7412, new_AGEMA_signal_7411, SubBytesIns_Inst_Sbox_12_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M36_U1 ( .a ({new_AGEMA_signal_7598, new_AGEMA_signal_7597, SubBytesIns_Inst_Sbox_12_M24}), .b ({new_AGEMA_signal_7408, new_AGEMA_signal_7407, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_7806, new_AGEMA_signal_7805, SubBytesIns_Inst_Sbox_12_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M25_U1 ( .a ({new_AGEMA_signal_7260, new_AGEMA_signal_7259, SubBytesIns_Inst_Sbox_13_M22}), .b ({new_AGEMA_signal_7256, new_AGEMA_signal_7255, SubBytesIns_Inst_Sbox_13_M20}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657]}), .c ({new_AGEMA_signal_7416, new_AGEMA_signal_7415, SubBytesIns_Inst_Sbox_13_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M26_U1 ( .a ({new_AGEMA_signal_7258, new_AGEMA_signal_7257, SubBytesIns_Inst_Sbox_13_M21}), .b ({new_AGEMA_signal_7416, new_AGEMA_signal_7415, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_7610, new_AGEMA_signal_7609, SubBytesIns_Inst_Sbox_13_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M28_U1 ( .a ({new_AGEMA_signal_7414, new_AGEMA_signal_7413, SubBytesIns_Inst_Sbox_13_M23}), .b ({new_AGEMA_signal_7416, new_AGEMA_signal_7415, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_7612, new_AGEMA_signal_7611, SubBytesIns_Inst_Sbox_13_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M31_U1 ( .a ({new_AGEMA_signal_7256, new_AGEMA_signal_7255, SubBytesIns_Inst_Sbox_13_M20}), .b ({new_AGEMA_signal_7414, new_AGEMA_signal_7413, SubBytesIns_Inst_Sbox_13_M23}), .clk (clk), .r ({Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_7614, new_AGEMA_signal_7613, SubBytesIns_Inst_Sbox_13_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M33_U1 ( .a ({new_AGEMA_signal_7418, new_AGEMA_signal_7417, SubBytesIns_Inst_Sbox_13_M27}), .b ({new_AGEMA_signal_7416, new_AGEMA_signal_7415, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_7616, new_AGEMA_signal_7615, SubBytesIns_Inst_Sbox_13_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M34_U1 ( .a ({new_AGEMA_signal_7258, new_AGEMA_signal_7257, SubBytesIns_Inst_Sbox_13_M21}), .b ({new_AGEMA_signal_7260, new_AGEMA_signal_7259, SubBytesIns_Inst_Sbox_13_M22}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663]}), .c ({new_AGEMA_signal_7420, new_AGEMA_signal_7419, SubBytesIns_Inst_Sbox_13_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M36_U1 ( .a ({new_AGEMA_signal_7608, new_AGEMA_signal_7607, SubBytesIns_Inst_Sbox_13_M24}), .b ({new_AGEMA_signal_7416, new_AGEMA_signal_7415, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_7816, new_AGEMA_signal_7815, SubBytesIns_Inst_Sbox_13_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M25_U1 ( .a ({new_AGEMA_signal_7268, new_AGEMA_signal_7267, SubBytesIns_Inst_Sbox_14_M22}), .b ({new_AGEMA_signal_7264, new_AGEMA_signal_7263, SubBytesIns_Inst_Sbox_14_M20}), .clk (clk), .r ({Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_7424, new_AGEMA_signal_7423, SubBytesIns_Inst_Sbox_14_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M26_U1 ( .a ({new_AGEMA_signal_7266, new_AGEMA_signal_7265, SubBytesIns_Inst_Sbox_14_M21}), .b ({new_AGEMA_signal_7424, new_AGEMA_signal_7423, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_7620, new_AGEMA_signal_7619, SubBytesIns_Inst_Sbox_14_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M28_U1 ( .a ({new_AGEMA_signal_7422, new_AGEMA_signal_7421, SubBytesIns_Inst_Sbox_14_M23}), .b ({new_AGEMA_signal_7424, new_AGEMA_signal_7423, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_7622, new_AGEMA_signal_7621, SubBytesIns_Inst_Sbox_14_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M31_U1 ( .a ({new_AGEMA_signal_7264, new_AGEMA_signal_7263, SubBytesIns_Inst_Sbox_14_M20}), .b ({new_AGEMA_signal_7422, new_AGEMA_signal_7421, SubBytesIns_Inst_Sbox_14_M23}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669]}), .c ({new_AGEMA_signal_7624, new_AGEMA_signal_7623, SubBytesIns_Inst_Sbox_14_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M33_U1 ( .a ({new_AGEMA_signal_7426, new_AGEMA_signal_7425, SubBytesIns_Inst_Sbox_14_M27}), .b ({new_AGEMA_signal_7424, new_AGEMA_signal_7423, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_7626, new_AGEMA_signal_7625, SubBytesIns_Inst_Sbox_14_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M34_U1 ( .a ({new_AGEMA_signal_7266, new_AGEMA_signal_7265, SubBytesIns_Inst_Sbox_14_M21}), .b ({new_AGEMA_signal_7268, new_AGEMA_signal_7267, SubBytesIns_Inst_Sbox_14_M22}), .clk (clk), .r ({Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_7428, new_AGEMA_signal_7427, SubBytesIns_Inst_Sbox_14_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M36_U1 ( .a ({new_AGEMA_signal_7618, new_AGEMA_signal_7617, SubBytesIns_Inst_Sbox_14_M24}), .b ({new_AGEMA_signal_7424, new_AGEMA_signal_7423, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_7826, new_AGEMA_signal_7825, SubBytesIns_Inst_Sbox_14_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M25_U1 ( .a ({new_AGEMA_signal_7276, new_AGEMA_signal_7275, SubBytesIns_Inst_Sbox_15_M22}), .b ({new_AGEMA_signal_7272, new_AGEMA_signal_7271, SubBytesIns_Inst_Sbox_15_M20}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675]}), .c ({new_AGEMA_signal_7432, new_AGEMA_signal_7431, SubBytesIns_Inst_Sbox_15_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M26_U1 ( .a ({new_AGEMA_signal_7274, new_AGEMA_signal_7273, SubBytesIns_Inst_Sbox_15_M21}), .b ({new_AGEMA_signal_7432, new_AGEMA_signal_7431, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_7630, new_AGEMA_signal_7629, SubBytesIns_Inst_Sbox_15_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M28_U1 ( .a ({new_AGEMA_signal_7430, new_AGEMA_signal_7429, SubBytesIns_Inst_Sbox_15_M23}), .b ({new_AGEMA_signal_7432, new_AGEMA_signal_7431, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_7632, new_AGEMA_signal_7631, SubBytesIns_Inst_Sbox_15_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M31_U1 ( .a ({new_AGEMA_signal_7272, new_AGEMA_signal_7271, SubBytesIns_Inst_Sbox_15_M20}), .b ({new_AGEMA_signal_7430, new_AGEMA_signal_7429, SubBytesIns_Inst_Sbox_15_M23}), .clk (clk), .r ({Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_7634, new_AGEMA_signal_7633, SubBytesIns_Inst_Sbox_15_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M33_U1 ( .a ({new_AGEMA_signal_7434, new_AGEMA_signal_7433, SubBytesIns_Inst_Sbox_15_M27}), .b ({new_AGEMA_signal_7432, new_AGEMA_signal_7431, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_7636, new_AGEMA_signal_7635, SubBytesIns_Inst_Sbox_15_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M34_U1 ( .a ({new_AGEMA_signal_7274, new_AGEMA_signal_7273, SubBytesIns_Inst_Sbox_15_M21}), .b ({new_AGEMA_signal_7276, new_AGEMA_signal_7275, SubBytesIns_Inst_Sbox_15_M22}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681]}), .c ({new_AGEMA_signal_7436, new_AGEMA_signal_7435, SubBytesIns_Inst_Sbox_15_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M36_U1 ( .a ({new_AGEMA_signal_7628, new_AGEMA_signal_7627, SubBytesIns_Inst_Sbox_15_M24}), .b ({new_AGEMA_signal_7432, new_AGEMA_signal_7431, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_7836, new_AGEMA_signal_7835, SubBytesIns_Inst_Sbox_15_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M25_U1 ( .a ({new_AGEMA_signal_7124, new_AGEMA_signal_7123, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_7120, new_AGEMA_signal_7119, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}), .clk (clk), .r ({Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_7280, new_AGEMA_signal_7279, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M26_U1 ( .a ({new_AGEMA_signal_7122, new_AGEMA_signal_7121, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_7280, new_AGEMA_signal_7279, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_7440, new_AGEMA_signal_7439, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M28_U1 ( .a ({new_AGEMA_signal_7278, new_AGEMA_signal_7277, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}), .b ({new_AGEMA_signal_7280, new_AGEMA_signal_7279, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_7442, new_AGEMA_signal_7441, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M31_U1 ( .a ({new_AGEMA_signal_7120, new_AGEMA_signal_7119, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_7278, new_AGEMA_signal_7277, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687]}), .c ({new_AGEMA_signal_7444, new_AGEMA_signal_7443, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M33_U1 ( .a ({new_AGEMA_signal_7282, new_AGEMA_signal_7281, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27}), .b ({new_AGEMA_signal_7280, new_AGEMA_signal_7279, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_7446, new_AGEMA_signal_7445, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M34_U1 ( .a ({new_AGEMA_signal_7122, new_AGEMA_signal_7121, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_7124, new_AGEMA_signal_7123, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}), .clk (clk), .r ({Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_7284, new_AGEMA_signal_7283, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M36_U1 ( .a ({new_AGEMA_signal_7438, new_AGEMA_signal_7437, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24}), .b ({new_AGEMA_signal_7280, new_AGEMA_signal_7279, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_7646, new_AGEMA_signal_7645, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M25_U1 ( .a ({new_AGEMA_signal_7132, new_AGEMA_signal_7131, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_7128, new_AGEMA_signal_7127, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693]}), .c ({new_AGEMA_signal_7288, new_AGEMA_signal_7287, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M26_U1 ( .a ({new_AGEMA_signal_7130, new_AGEMA_signal_7129, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_7288, new_AGEMA_signal_7287, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_7450, new_AGEMA_signal_7449, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M28_U1 ( .a ({new_AGEMA_signal_7286, new_AGEMA_signal_7285, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}), .b ({new_AGEMA_signal_7288, new_AGEMA_signal_7287, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_7452, new_AGEMA_signal_7451, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M31_U1 ( .a ({new_AGEMA_signal_7128, new_AGEMA_signal_7127, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_7286, new_AGEMA_signal_7285, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}), .clk (clk), .r ({Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_7454, new_AGEMA_signal_7453, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M33_U1 ( .a ({new_AGEMA_signal_7290, new_AGEMA_signal_7289, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27}), .b ({new_AGEMA_signal_7288, new_AGEMA_signal_7287, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_7456, new_AGEMA_signal_7455, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M34_U1 ( .a ({new_AGEMA_signal_7130, new_AGEMA_signal_7129, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_7132, new_AGEMA_signal_7131, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699]}), .c ({new_AGEMA_signal_7292, new_AGEMA_signal_7291, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M36_U1 ( .a ({new_AGEMA_signal_7448, new_AGEMA_signal_7447, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24}), .b ({new_AGEMA_signal_7288, new_AGEMA_signal_7287, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_7656, new_AGEMA_signal_7655, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M25_U1 ( .a ({new_AGEMA_signal_7140, new_AGEMA_signal_7139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_7136, new_AGEMA_signal_7135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}), .clk (clk), .r ({Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_7296, new_AGEMA_signal_7295, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M26_U1 ( .a ({new_AGEMA_signal_7138, new_AGEMA_signal_7137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_7296, new_AGEMA_signal_7295, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_7460, new_AGEMA_signal_7459, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M28_U1 ( .a ({new_AGEMA_signal_7294, new_AGEMA_signal_7293, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}), .b ({new_AGEMA_signal_7296, new_AGEMA_signal_7295, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_7462, new_AGEMA_signal_7461, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M31_U1 ( .a ({new_AGEMA_signal_7136, new_AGEMA_signal_7135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_7294, new_AGEMA_signal_7293, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705]}), .c ({new_AGEMA_signal_7464, new_AGEMA_signal_7463, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M33_U1 ( .a ({new_AGEMA_signal_7298, new_AGEMA_signal_7297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27}), .b ({new_AGEMA_signal_7296, new_AGEMA_signal_7295, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_7466, new_AGEMA_signal_7465, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M34_U1 ( .a ({new_AGEMA_signal_7138, new_AGEMA_signal_7137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_7140, new_AGEMA_signal_7139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}), .clk (clk), .r ({Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_7300, new_AGEMA_signal_7299, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M36_U1 ( .a ({new_AGEMA_signal_7458, new_AGEMA_signal_7457, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24}), .b ({new_AGEMA_signal_7296, new_AGEMA_signal_7295, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_7666, new_AGEMA_signal_7665, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M25_U1 ( .a ({new_AGEMA_signal_7148, new_AGEMA_signal_7147, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_7144, new_AGEMA_signal_7143, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711]}), .c ({new_AGEMA_signal_7304, new_AGEMA_signal_7303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M26_U1 ( .a ({new_AGEMA_signal_7146, new_AGEMA_signal_7145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_7304, new_AGEMA_signal_7303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_7470, new_AGEMA_signal_7469, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M28_U1 ( .a ({new_AGEMA_signal_7302, new_AGEMA_signal_7301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}), .b ({new_AGEMA_signal_7304, new_AGEMA_signal_7303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_7472, new_AGEMA_signal_7471, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M31_U1 ( .a ({new_AGEMA_signal_7144, new_AGEMA_signal_7143, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_7302, new_AGEMA_signal_7301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}), .clk (clk), .r ({Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_7474, new_AGEMA_signal_7473, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M33_U1 ( .a ({new_AGEMA_signal_7306, new_AGEMA_signal_7305, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27}), .b ({new_AGEMA_signal_7304, new_AGEMA_signal_7303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_7476, new_AGEMA_signal_7475, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M34_U1 ( .a ({new_AGEMA_signal_7146, new_AGEMA_signal_7145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_7148, new_AGEMA_signal_7147, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717]}), .c ({new_AGEMA_signal_7308, new_AGEMA_signal_7307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M36_U1 ( .a ({new_AGEMA_signal_7468, new_AGEMA_signal_7467, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24}), .b ({new_AGEMA_signal_7304, new_AGEMA_signal_7303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_7676, new_AGEMA_signal_7675, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M29_U1 ( .a ({new_AGEMA_signal_7482, new_AGEMA_signal_7481, SubBytesIns_Inst_Sbox_0_M28}), .b ({new_AGEMA_signal_7314, new_AGEMA_signal_7313, SubBytesIns_Inst_Sbox_0_M27}), .clk (clk), .r ({Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_7678, new_AGEMA_signal_7677, SubBytesIns_Inst_Sbox_0_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M30_U1 ( .a ({new_AGEMA_signal_7480, new_AGEMA_signal_7479, SubBytesIns_Inst_Sbox_0_M26}), .b ({new_AGEMA_signal_7478, new_AGEMA_signal_7477, SubBytesIns_Inst_Sbox_0_M24}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723]}), .c ({new_AGEMA_signal_7680, new_AGEMA_signal_7679, SubBytesIns_Inst_Sbox_0_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M32_U1 ( .a ({new_AGEMA_signal_7314, new_AGEMA_signal_7313, SubBytesIns_Inst_Sbox_0_M27}), .b ({new_AGEMA_signal_7484, new_AGEMA_signal_7483, SubBytesIns_Inst_Sbox_0_M31}), .clk (clk), .r ({Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_7682, new_AGEMA_signal_7681, SubBytesIns_Inst_Sbox_0_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M35_U1 ( .a ({new_AGEMA_signal_7478, new_AGEMA_signal_7477, SubBytesIns_Inst_Sbox_0_M24}), .b ({new_AGEMA_signal_7316, new_AGEMA_signal_7315, SubBytesIns_Inst_Sbox_0_M34}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729]}), .c ({new_AGEMA_signal_7684, new_AGEMA_signal_7683, SubBytesIns_Inst_Sbox_0_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M37_U1 ( .a ({new_AGEMA_signal_7154, new_AGEMA_signal_7153, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_7678, new_AGEMA_signal_7677, SubBytesIns_Inst_Sbox_0_M29}), .c ({new_AGEMA_signal_7870, new_AGEMA_signal_7869, SubBytesIns_Inst_Sbox_0_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M38_U1 ( .a ({new_AGEMA_signal_7682, new_AGEMA_signal_7681, SubBytesIns_Inst_Sbox_0_M32}), .b ({new_AGEMA_signal_7486, new_AGEMA_signal_7485, SubBytesIns_Inst_Sbox_0_M33}), .c ({new_AGEMA_signal_7872, new_AGEMA_signal_7871, SubBytesIns_Inst_Sbox_0_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M39_U1 ( .a ({new_AGEMA_signal_7310, new_AGEMA_signal_7309, SubBytesIns_Inst_Sbox_0_M23}), .b ({new_AGEMA_signal_7680, new_AGEMA_signal_7679, SubBytesIns_Inst_Sbox_0_M30}), .c ({new_AGEMA_signal_7874, new_AGEMA_signal_7873, SubBytesIns_Inst_Sbox_0_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M40_U1 ( .a ({new_AGEMA_signal_7684, new_AGEMA_signal_7683, SubBytesIns_Inst_Sbox_0_M35}), .b ({new_AGEMA_signal_7686, new_AGEMA_signal_7685, SubBytesIns_Inst_Sbox_0_M36}), .c ({new_AGEMA_signal_7876, new_AGEMA_signal_7875, SubBytesIns_Inst_Sbox_0_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M41_U1 ( .a ({new_AGEMA_signal_7872, new_AGEMA_signal_7871, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_7876, new_AGEMA_signal_7875, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_8094, new_AGEMA_signal_8093, SubBytesIns_Inst_Sbox_0_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M42_U1 ( .a ({new_AGEMA_signal_7870, new_AGEMA_signal_7869, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_7874, new_AGEMA_signal_7873, SubBytesIns_Inst_Sbox_0_M39}), .c ({new_AGEMA_signal_8096, new_AGEMA_signal_8095, SubBytesIns_Inst_Sbox_0_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M43_U1 ( .a ({new_AGEMA_signal_7870, new_AGEMA_signal_7869, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_7872, new_AGEMA_signal_7871, SubBytesIns_Inst_Sbox_0_M38}), .c ({new_AGEMA_signal_8098, new_AGEMA_signal_8097, SubBytesIns_Inst_Sbox_0_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M44_U1 ( .a ({new_AGEMA_signal_7874, new_AGEMA_signal_7873, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_7876, new_AGEMA_signal_7875, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_8100, new_AGEMA_signal_8099, SubBytesIns_Inst_Sbox_0_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M45_U1 ( .a ({new_AGEMA_signal_8096, new_AGEMA_signal_8095, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_8094, new_AGEMA_signal_8093, SubBytesIns_Inst_Sbox_0_M41}), .c ({new_AGEMA_signal_8574, new_AGEMA_signal_8573, SubBytesIns_Inst_Sbox_0_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M29_U1 ( .a ({new_AGEMA_signal_7492, new_AGEMA_signal_7491, SubBytesIns_Inst_Sbox_1_M28}), .b ({new_AGEMA_signal_7322, new_AGEMA_signal_7321, SubBytesIns_Inst_Sbox_1_M27}), .clk (clk), .r ({Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_7688, new_AGEMA_signal_7687, SubBytesIns_Inst_Sbox_1_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M30_U1 ( .a ({new_AGEMA_signal_7490, new_AGEMA_signal_7489, SubBytesIns_Inst_Sbox_1_M26}), .b ({new_AGEMA_signal_7488, new_AGEMA_signal_7487, SubBytesIns_Inst_Sbox_1_M24}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735]}), .c ({new_AGEMA_signal_7690, new_AGEMA_signal_7689, SubBytesIns_Inst_Sbox_1_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M32_U1 ( .a ({new_AGEMA_signal_7322, new_AGEMA_signal_7321, SubBytesIns_Inst_Sbox_1_M27}), .b ({new_AGEMA_signal_7494, new_AGEMA_signal_7493, SubBytesIns_Inst_Sbox_1_M31}), .clk (clk), .r ({Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_7692, new_AGEMA_signal_7691, SubBytesIns_Inst_Sbox_1_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M35_U1 ( .a ({new_AGEMA_signal_7488, new_AGEMA_signal_7487, SubBytesIns_Inst_Sbox_1_M24}), .b ({new_AGEMA_signal_7324, new_AGEMA_signal_7323, SubBytesIns_Inst_Sbox_1_M34}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741]}), .c ({new_AGEMA_signal_7694, new_AGEMA_signal_7693, SubBytesIns_Inst_Sbox_1_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M37_U1 ( .a ({new_AGEMA_signal_7162, new_AGEMA_signal_7161, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_7688, new_AGEMA_signal_7687, SubBytesIns_Inst_Sbox_1_M29}), .c ({new_AGEMA_signal_7878, new_AGEMA_signal_7877, SubBytesIns_Inst_Sbox_1_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M38_U1 ( .a ({new_AGEMA_signal_7692, new_AGEMA_signal_7691, SubBytesIns_Inst_Sbox_1_M32}), .b ({new_AGEMA_signal_7496, new_AGEMA_signal_7495, SubBytesIns_Inst_Sbox_1_M33}), .c ({new_AGEMA_signal_7880, new_AGEMA_signal_7879, SubBytesIns_Inst_Sbox_1_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M39_U1 ( .a ({new_AGEMA_signal_7318, new_AGEMA_signal_7317, SubBytesIns_Inst_Sbox_1_M23}), .b ({new_AGEMA_signal_7690, new_AGEMA_signal_7689, SubBytesIns_Inst_Sbox_1_M30}), .c ({new_AGEMA_signal_7882, new_AGEMA_signal_7881, SubBytesIns_Inst_Sbox_1_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M40_U1 ( .a ({new_AGEMA_signal_7694, new_AGEMA_signal_7693, SubBytesIns_Inst_Sbox_1_M35}), .b ({new_AGEMA_signal_7696, new_AGEMA_signal_7695, SubBytesIns_Inst_Sbox_1_M36}), .c ({new_AGEMA_signal_7884, new_AGEMA_signal_7883, SubBytesIns_Inst_Sbox_1_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M41_U1 ( .a ({new_AGEMA_signal_7880, new_AGEMA_signal_7879, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_7884, new_AGEMA_signal_7883, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_8118, new_AGEMA_signal_8117, SubBytesIns_Inst_Sbox_1_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M42_U1 ( .a ({new_AGEMA_signal_7878, new_AGEMA_signal_7877, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_7882, new_AGEMA_signal_7881, SubBytesIns_Inst_Sbox_1_M39}), .c ({new_AGEMA_signal_8120, new_AGEMA_signal_8119, SubBytesIns_Inst_Sbox_1_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M43_U1 ( .a ({new_AGEMA_signal_7878, new_AGEMA_signal_7877, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_7880, new_AGEMA_signal_7879, SubBytesIns_Inst_Sbox_1_M38}), .c ({new_AGEMA_signal_8122, new_AGEMA_signal_8121, SubBytesIns_Inst_Sbox_1_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M44_U1 ( .a ({new_AGEMA_signal_7882, new_AGEMA_signal_7881, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_7884, new_AGEMA_signal_7883, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_8124, new_AGEMA_signal_8123, SubBytesIns_Inst_Sbox_1_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M45_U1 ( .a ({new_AGEMA_signal_8120, new_AGEMA_signal_8119, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_8118, new_AGEMA_signal_8117, SubBytesIns_Inst_Sbox_1_M41}), .c ({new_AGEMA_signal_8598, new_AGEMA_signal_8597, SubBytesIns_Inst_Sbox_1_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M29_U1 ( .a ({new_AGEMA_signal_7502, new_AGEMA_signal_7501, SubBytesIns_Inst_Sbox_2_M28}), .b ({new_AGEMA_signal_7330, new_AGEMA_signal_7329, SubBytesIns_Inst_Sbox_2_M27}), .clk (clk), .r ({Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_7698, new_AGEMA_signal_7697, SubBytesIns_Inst_Sbox_2_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M30_U1 ( .a ({new_AGEMA_signal_7500, new_AGEMA_signal_7499, SubBytesIns_Inst_Sbox_2_M26}), .b ({new_AGEMA_signal_7498, new_AGEMA_signal_7497, SubBytesIns_Inst_Sbox_2_M24}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747]}), .c ({new_AGEMA_signal_7700, new_AGEMA_signal_7699, SubBytesIns_Inst_Sbox_2_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M32_U1 ( .a ({new_AGEMA_signal_7330, new_AGEMA_signal_7329, SubBytesIns_Inst_Sbox_2_M27}), .b ({new_AGEMA_signal_7504, new_AGEMA_signal_7503, SubBytesIns_Inst_Sbox_2_M31}), .clk (clk), .r ({Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_7702, new_AGEMA_signal_7701, SubBytesIns_Inst_Sbox_2_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M35_U1 ( .a ({new_AGEMA_signal_7498, new_AGEMA_signal_7497, SubBytesIns_Inst_Sbox_2_M24}), .b ({new_AGEMA_signal_7332, new_AGEMA_signal_7331, SubBytesIns_Inst_Sbox_2_M34}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753]}), .c ({new_AGEMA_signal_7704, new_AGEMA_signal_7703, SubBytesIns_Inst_Sbox_2_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M37_U1 ( .a ({new_AGEMA_signal_7170, new_AGEMA_signal_7169, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_7698, new_AGEMA_signal_7697, SubBytesIns_Inst_Sbox_2_M29}), .c ({new_AGEMA_signal_7886, new_AGEMA_signal_7885, SubBytesIns_Inst_Sbox_2_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M38_U1 ( .a ({new_AGEMA_signal_7702, new_AGEMA_signal_7701, SubBytesIns_Inst_Sbox_2_M32}), .b ({new_AGEMA_signal_7506, new_AGEMA_signal_7505, SubBytesIns_Inst_Sbox_2_M33}), .c ({new_AGEMA_signal_7888, new_AGEMA_signal_7887, SubBytesIns_Inst_Sbox_2_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M39_U1 ( .a ({new_AGEMA_signal_7326, new_AGEMA_signal_7325, SubBytesIns_Inst_Sbox_2_M23}), .b ({new_AGEMA_signal_7700, new_AGEMA_signal_7699, SubBytesIns_Inst_Sbox_2_M30}), .c ({new_AGEMA_signal_7890, new_AGEMA_signal_7889, SubBytesIns_Inst_Sbox_2_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M40_U1 ( .a ({new_AGEMA_signal_7704, new_AGEMA_signal_7703, SubBytesIns_Inst_Sbox_2_M35}), .b ({new_AGEMA_signal_7706, new_AGEMA_signal_7705, SubBytesIns_Inst_Sbox_2_M36}), .c ({new_AGEMA_signal_7892, new_AGEMA_signal_7891, SubBytesIns_Inst_Sbox_2_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M41_U1 ( .a ({new_AGEMA_signal_7888, new_AGEMA_signal_7887, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_7892, new_AGEMA_signal_7891, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_8142, new_AGEMA_signal_8141, SubBytesIns_Inst_Sbox_2_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M42_U1 ( .a ({new_AGEMA_signal_7886, new_AGEMA_signal_7885, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_7890, new_AGEMA_signal_7889, SubBytesIns_Inst_Sbox_2_M39}), .c ({new_AGEMA_signal_8144, new_AGEMA_signal_8143, SubBytesIns_Inst_Sbox_2_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M43_U1 ( .a ({new_AGEMA_signal_7886, new_AGEMA_signal_7885, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_7888, new_AGEMA_signal_7887, SubBytesIns_Inst_Sbox_2_M38}), .c ({new_AGEMA_signal_8146, new_AGEMA_signal_8145, SubBytesIns_Inst_Sbox_2_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M44_U1 ( .a ({new_AGEMA_signal_7890, new_AGEMA_signal_7889, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_7892, new_AGEMA_signal_7891, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_8148, new_AGEMA_signal_8147, SubBytesIns_Inst_Sbox_2_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M45_U1 ( .a ({new_AGEMA_signal_8144, new_AGEMA_signal_8143, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_8142, new_AGEMA_signal_8141, SubBytesIns_Inst_Sbox_2_M41}), .c ({new_AGEMA_signal_8622, new_AGEMA_signal_8621, SubBytesIns_Inst_Sbox_2_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M29_U1 ( .a ({new_AGEMA_signal_7512, new_AGEMA_signal_7511, SubBytesIns_Inst_Sbox_3_M28}), .b ({new_AGEMA_signal_7338, new_AGEMA_signal_7337, SubBytesIns_Inst_Sbox_3_M27}), .clk (clk), .r ({Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_7708, new_AGEMA_signal_7707, SubBytesIns_Inst_Sbox_3_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M30_U1 ( .a ({new_AGEMA_signal_7510, new_AGEMA_signal_7509, SubBytesIns_Inst_Sbox_3_M26}), .b ({new_AGEMA_signal_7508, new_AGEMA_signal_7507, SubBytesIns_Inst_Sbox_3_M24}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759]}), .c ({new_AGEMA_signal_7710, new_AGEMA_signal_7709, SubBytesIns_Inst_Sbox_3_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M32_U1 ( .a ({new_AGEMA_signal_7338, new_AGEMA_signal_7337, SubBytesIns_Inst_Sbox_3_M27}), .b ({new_AGEMA_signal_7514, new_AGEMA_signal_7513, SubBytesIns_Inst_Sbox_3_M31}), .clk (clk), .r ({Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_7712, new_AGEMA_signal_7711, SubBytesIns_Inst_Sbox_3_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M35_U1 ( .a ({new_AGEMA_signal_7508, new_AGEMA_signal_7507, SubBytesIns_Inst_Sbox_3_M24}), .b ({new_AGEMA_signal_7340, new_AGEMA_signal_7339, SubBytesIns_Inst_Sbox_3_M34}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765]}), .c ({new_AGEMA_signal_7714, new_AGEMA_signal_7713, SubBytesIns_Inst_Sbox_3_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M37_U1 ( .a ({new_AGEMA_signal_7178, new_AGEMA_signal_7177, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_7708, new_AGEMA_signal_7707, SubBytesIns_Inst_Sbox_3_M29}), .c ({new_AGEMA_signal_7894, new_AGEMA_signal_7893, SubBytesIns_Inst_Sbox_3_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M38_U1 ( .a ({new_AGEMA_signal_7712, new_AGEMA_signal_7711, SubBytesIns_Inst_Sbox_3_M32}), .b ({new_AGEMA_signal_7516, new_AGEMA_signal_7515, SubBytesIns_Inst_Sbox_3_M33}), .c ({new_AGEMA_signal_7896, new_AGEMA_signal_7895, SubBytesIns_Inst_Sbox_3_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M39_U1 ( .a ({new_AGEMA_signal_7334, new_AGEMA_signal_7333, SubBytesIns_Inst_Sbox_3_M23}), .b ({new_AGEMA_signal_7710, new_AGEMA_signal_7709, SubBytesIns_Inst_Sbox_3_M30}), .c ({new_AGEMA_signal_7898, new_AGEMA_signal_7897, SubBytesIns_Inst_Sbox_3_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M40_U1 ( .a ({new_AGEMA_signal_7714, new_AGEMA_signal_7713, SubBytesIns_Inst_Sbox_3_M35}), .b ({new_AGEMA_signal_7716, new_AGEMA_signal_7715, SubBytesIns_Inst_Sbox_3_M36}), .c ({new_AGEMA_signal_7900, new_AGEMA_signal_7899, SubBytesIns_Inst_Sbox_3_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M41_U1 ( .a ({new_AGEMA_signal_7896, new_AGEMA_signal_7895, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_7900, new_AGEMA_signal_7899, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_8166, new_AGEMA_signal_8165, SubBytesIns_Inst_Sbox_3_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M42_U1 ( .a ({new_AGEMA_signal_7894, new_AGEMA_signal_7893, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_7898, new_AGEMA_signal_7897, SubBytesIns_Inst_Sbox_3_M39}), .c ({new_AGEMA_signal_8168, new_AGEMA_signal_8167, SubBytesIns_Inst_Sbox_3_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M43_U1 ( .a ({new_AGEMA_signal_7894, new_AGEMA_signal_7893, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_7896, new_AGEMA_signal_7895, SubBytesIns_Inst_Sbox_3_M38}), .c ({new_AGEMA_signal_8170, new_AGEMA_signal_8169, SubBytesIns_Inst_Sbox_3_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M44_U1 ( .a ({new_AGEMA_signal_7898, new_AGEMA_signal_7897, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_7900, new_AGEMA_signal_7899, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_8172, new_AGEMA_signal_8171, SubBytesIns_Inst_Sbox_3_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M45_U1 ( .a ({new_AGEMA_signal_8168, new_AGEMA_signal_8167, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_8166, new_AGEMA_signal_8165, SubBytesIns_Inst_Sbox_3_M41}), .c ({new_AGEMA_signal_8646, new_AGEMA_signal_8645, SubBytesIns_Inst_Sbox_3_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M29_U1 ( .a ({new_AGEMA_signal_7522, new_AGEMA_signal_7521, SubBytesIns_Inst_Sbox_4_M28}), .b ({new_AGEMA_signal_7346, new_AGEMA_signal_7345, SubBytesIns_Inst_Sbox_4_M27}), .clk (clk), .r ({Fresh[770], Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_7718, new_AGEMA_signal_7717, SubBytesIns_Inst_Sbox_4_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M30_U1 ( .a ({new_AGEMA_signal_7520, new_AGEMA_signal_7519, SubBytesIns_Inst_Sbox_4_M26}), .b ({new_AGEMA_signal_7518, new_AGEMA_signal_7517, SubBytesIns_Inst_Sbox_4_M24}), .clk (clk), .r ({Fresh[773], Fresh[772], Fresh[771]}), .c ({new_AGEMA_signal_7720, new_AGEMA_signal_7719, SubBytesIns_Inst_Sbox_4_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M32_U1 ( .a ({new_AGEMA_signal_7346, new_AGEMA_signal_7345, SubBytesIns_Inst_Sbox_4_M27}), .b ({new_AGEMA_signal_7524, new_AGEMA_signal_7523, SubBytesIns_Inst_Sbox_4_M31}), .clk (clk), .r ({Fresh[776], Fresh[775], Fresh[774]}), .c ({new_AGEMA_signal_7722, new_AGEMA_signal_7721, SubBytesIns_Inst_Sbox_4_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M35_U1 ( .a ({new_AGEMA_signal_7518, new_AGEMA_signal_7517, SubBytesIns_Inst_Sbox_4_M24}), .b ({new_AGEMA_signal_7348, new_AGEMA_signal_7347, SubBytesIns_Inst_Sbox_4_M34}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777]}), .c ({new_AGEMA_signal_7724, new_AGEMA_signal_7723, SubBytesIns_Inst_Sbox_4_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M37_U1 ( .a ({new_AGEMA_signal_7186, new_AGEMA_signal_7185, SubBytesIns_Inst_Sbox_4_M21}), .b ({new_AGEMA_signal_7718, new_AGEMA_signal_7717, SubBytesIns_Inst_Sbox_4_M29}), .c ({new_AGEMA_signal_7902, new_AGEMA_signal_7901, SubBytesIns_Inst_Sbox_4_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M38_U1 ( .a ({new_AGEMA_signal_7722, new_AGEMA_signal_7721, SubBytesIns_Inst_Sbox_4_M32}), .b ({new_AGEMA_signal_7526, new_AGEMA_signal_7525, SubBytesIns_Inst_Sbox_4_M33}), .c ({new_AGEMA_signal_7904, new_AGEMA_signal_7903, SubBytesIns_Inst_Sbox_4_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M39_U1 ( .a ({new_AGEMA_signal_7342, new_AGEMA_signal_7341, SubBytesIns_Inst_Sbox_4_M23}), .b ({new_AGEMA_signal_7720, new_AGEMA_signal_7719, SubBytesIns_Inst_Sbox_4_M30}), .c ({new_AGEMA_signal_7906, new_AGEMA_signal_7905, SubBytesIns_Inst_Sbox_4_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M40_U1 ( .a ({new_AGEMA_signal_7724, new_AGEMA_signal_7723, SubBytesIns_Inst_Sbox_4_M35}), .b ({new_AGEMA_signal_7726, new_AGEMA_signal_7725, SubBytesIns_Inst_Sbox_4_M36}), .c ({new_AGEMA_signal_7908, new_AGEMA_signal_7907, SubBytesIns_Inst_Sbox_4_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M41_U1 ( .a ({new_AGEMA_signal_7904, new_AGEMA_signal_7903, SubBytesIns_Inst_Sbox_4_M38}), .b ({new_AGEMA_signal_7908, new_AGEMA_signal_7907, SubBytesIns_Inst_Sbox_4_M40}), .c ({new_AGEMA_signal_8190, new_AGEMA_signal_8189, SubBytesIns_Inst_Sbox_4_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M42_U1 ( .a ({new_AGEMA_signal_7902, new_AGEMA_signal_7901, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_7906, new_AGEMA_signal_7905, SubBytesIns_Inst_Sbox_4_M39}), .c ({new_AGEMA_signal_8192, new_AGEMA_signal_8191, SubBytesIns_Inst_Sbox_4_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M43_U1 ( .a ({new_AGEMA_signal_7902, new_AGEMA_signal_7901, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_7904, new_AGEMA_signal_7903, SubBytesIns_Inst_Sbox_4_M38}), .c ({new_AGEMA_signal_8194, new_AGEMA_signal_8193, SubBytesIns_Inst_Sbox_4_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M44_U1 ( .a ({new_AGEMA_signal_7906, new_AGEMA_signal_7905, SubBytesIns_Inst_Sbox_4_M39}), .b ({new_AGEMA_signal_7908, new_AGEMA_signal_7907, SubBytesIns_Inst_Sbox_4_M40}), .c ({new_AGEMA_signal_8196, new_AGEMA_signal_8195, SubBytesIns_Inst_Sbox_4_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M45_U1 ( .a ({new_AGEMA_signal_8192, new_AGEMA_signal_8191, SubBytesIns_Inst_Sbox_4_M42}), .b ({new_AGEMA_signal_8190, new_AGEMA_signal_8189, SubBytesIns_Inst_Sbox_4_M41}), .c ({new_AGEMA_signal_8670, new_AGEMA_signal_8669, SubBytesIns_Inst_Sbox_4_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M29_U1 ( .a ({new_AGEMA_signal_7532, new_AGEMA_signal_7531, SubBytesIns_Inst_Sbox_5_M28}), .b ({new_AGEMA_signal_7354, new_AGEMA_signal_7353, SubBytesIns_Inst_Sbox_5_M27}), .clk (clk), .r ({Fresh[782], Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_7728, new_AGEMA_signal_7727, SubBytesIns_Inst_Sbox_5_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M30_U1 ( .a ({new_AGEMA_signal_7530, new_AGEMA_signal_7529, SubBytesIns_Inst_Sbox_5_M26}), .b ({new_AGEMA_signal_7528, new_AGEMA_signal_7527, SubBytesIns_Inst_Sbox_5_M24}), .clk (clk), .r ({Fresh[785], Fresh[784], Fresh[783]}), .c ({new_AGEMA_signal_7730, new_AGEMA_signal_7729, SubBytesIns_Inst_Sbox_5_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M32_U1 ( .a ({new_AGEMA_signal_7354, new_AGEMA_signal_7353, SubBytesIns_Inst_Sbox_5_M27}), .b ({new_AGEMA_signal_7534, new_AGEMA_signal_7533, SubBytesIns_Inst_Sbox_5_M31}), .clk (clk), .r ({Fresh[788], Fresh[787], Fresh[786]}), .c ({new_AGEMA_signal_7732, new_AGEMA_signal_7731, SubBytesIns_Inst_Sbox_5_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M35_U1 ( .a ({new_AGEMA_signal_7528, new_AGEMA_signal_7527, SubBytesIns_Inst_Sbox_5_M24}), .b ({new_AGEMA_signal_7356, new_AGEMA_signal_7355, SubBytesIns_Inst_Sbox_5_M34}), .clk (clk), .r ({Fresh[791], Fresh[790], Fresh[789]}), .c ({new_AGEMA_signal_7734, new_AGEMA_signal_7733, SubBytesIns_Inst_Sbox_5_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M37_U1 ( .a ({new_AGEMA_signal_7194, new_AGEMA_signal_7193, SubBytesIns_Inst_Sbox_5_M21}), .b ({new_AGEMA_signal_7728, new_AGEMA_signal_7727, SubBytesIns_Inst_Sbox_5_M29}), .c ({new_AGEMA_signal_7910, new_AGEMA_signal_7909, SubBytesIns_Inst_Sbox_5_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M38_U1 ( .a ({new_AGEMA_signal_7732, new_AGEMA_signal_7731, SubBytesIns_Inst_Sbox_5_M32}), .b ({new_AGEMA_signal_7536, new_AGEMA_signal_7535, SubBytesIns_Inst_Sbox_5_M33}), .c ({new_AGEMA_signal_7912, new_AGEMA_signal_7911, SubBytesIns_Inst_Sbox_5_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M39_U1 ( .a ({new_AGEMA_signal_7350, new_AGEMA_signal_7349, SubBytesIns_Inst_Sbox_5_M23}), .b ({new_AGEMA_signal_7730, new_AGEMA_signal_7729, SubBytesIns_Inst_Sbox_5_M30}), .c ({new_AGEMA_signal_7914, new_AGEMA_signal_7913, SubBytesIns_Inst_Sbox_5_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M40_U1 ( .a ({new_AGEMA_signal_7734, new_AGEMA_signal_7733, SubBytesIns_Inst_Sbox_5_M35}), .b ({new_AGEMA_signal_7736, new_AGEMA_signal_7735, SubBytesIns_Inst_Sbox_5_M36}), .c ({new_AGEMA_signal_7916, new_AGEMA_signal_7915, SubBytesIns_Inst_Sbox_5_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M41_U1 ( .a ({new_AGEMA_signal_7912, new_AGEMA_signal_7911, SubBytesIns_Inst_Sbox_5_M38}), .b ({new_AGEMA_signal_7916, new_AGEMA_signal_7915, SubBytesIns_Inst_Sbox_5_M40}), .c ({new_AGEMA_signal_8214, new_AGEMA_signal_8213, SubBytesIns_Inst_Sbox_5_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M42_U1 ( .a ({new_AGEMA_signal_7910, new_AGEMA_signal_7909, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_7914, new_AGEMA_signal_7913, SubBytesIns_Inst_Sbox_5_M39}), .c ({new_AGEMA_signal_8216, new_AGEMA_signal_8215, SubBytesIns_Inst_Sbox_5_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M43_U1 ( .a ({new_AGEMA_signal_7910, new_AGEMA_signal_7909, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_7912, new_AGEMA_signal_7911, SubBytesIns_Inst_Sbox_5_M38}), .c ({new_AGEMA_signal_8218, new_AGEMA_signal_8217, SubBytesIns_Inst_Sbox_5_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M44_U1 ( .a ({new_AGEMA_signal_7914, new_AGEMA_signal_7913, SubBytesIns_Inst_Sbox_5_M39}), .b ({new_AGEMA_signal_7916, new_AGEMA_signal_7915, SubBytesIns_Inst_Sbox_5_M40}), .c ({new_AGEMA_signal_8220, new_AGEMA_signal_8219, SubBytesIns_Inst_Sbox_5_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M45_U1 ( .a ({new_AGEMA_signal_8216, new_AGEMA_signal_8215, SubBytesIns_Inst_Sbox_5_M42}), .b ({new_AGEMA_signal_8214, new_AGEMA_signal_8213, SubBytesIns_Inst_Sbox_5_M41}), .c ({new_AGEMA_signal_8694, new_AGEMA_signal_8693, SubBytesIns_Inst_Sbox_5_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M29_U1 ( .a ({new_AGEMA_signal_7542, new_AGEMA_signal_7541, SubBytesIns_Inst_Sbox_6_M28}), .b ({new_AGEMA_signal_7362, new_AGEMA_signal_7361, SubBytesIns_Inst_Sbox_6_M27}), .clk (clk), .r ({Fresh[794], Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_7738, new_AGEMA_signal_7737, SubBytesIns_Inst_Sbox_6_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M30_U1 ( .a ({new_AGEMA_signal_7540, new_AGEMA_signal_7539, SubBytesIns_Inst_Sbox_6_M26}), .b ({new_AGEMA_signal_7538, new_AGEMA_signal_7537, SubBytesIns_Inst_Sbox_6_M24}), .clk (clk), .r ({Fresh[797], Fresh[796], Fresh[795]}), .c ({new_AGEMA_signal_7740, new_AGEMA_signal_7739, SubBytesIns_Inst_Sbox_6_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M32_U1 ( .a ({new_AGEMA_signal_7362, new_AGEMA_signal_7361, SubBytesIns_Inst_Sbox_6_M27}), .b ({new_AGEMA_signal_7544, new_AGEMA_signal_7543, SubBytesIns_Inst_Sbox_6_M31}), .clk (clk), .r ({Fresh[800], Fresh[799], Fresh[798]}), .c ({new_AGEMA_signal_7742, new_AGEMA_signal_7741, SubBytesIns_Inst_Sbox_6_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M35_U1 ( .a ({new_AGEMA_signal_7538, new_AGEMA_signal_7537, SubBytesIns_Inst_Sbox_6_M24}), .b ({new_AGEMA_signal_7364, new_AGEMA_signal_7363, SubBytesIns_Inst_Sbox_6_M34}), .clk (clk), .r ({Fresh[803], Fresh[802], Fresh[801]}), .c ({new_AGEMA_signal_7744, new_AGEMA_signal_7743, SubBytesIns_Inst_Sbox_6_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M37_U1 ( .a ({new_AGEMA_signal_7202, new_AGEMA_signal_7201, SubBytesIns_Inst_Sbox_6_M21}), .b ({new_AGEMA_signal_7738, new_AGEMA_signal_7737, SubBytesIns_Inst_Sbox_6_M29}), .c ({new_AGEMA_signal_7918, new_AGEMA_signal_7917, SubBytesIns_Inst_Sbox_6_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M38_U1 ( .a ({new_AGEMA_signal_7742, new_AGEMA_signal_7741, SubBytesIns_Inst_Sbox_6_M32}), .b ({new_AGEMA_signal_7546, new_AGEMA_signal_7545, SubBytesIns_Inst_Sbox_6_M33}), .c ({new_AGEMA_signal_7920, new_AGEMA_signal_7919, SubBytesIns_Inst_Sbox_6_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M39_U1 ( .a ({new_AGEMA_signal_7358, new_AGEMA_signal_7357, SubBytesIns_Inst_Sbox_6_M23}), .b ({new_AGEMA_signal_7740, new_AGEMA_signal_7739, SubBytesIns_Inst_Sbox_6_M30}), .c ({new_AGEMA_signal_7922, new_AGEMA_signal_7921, SubBytesIns_Inst_Sbox_6_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M40_U1 ( .a ({new_AGEMA_signal_7744, new_AGEMA_signal_7743, SubBytesIns_Inst_Sbox_6_M35}), .b ({new_AGEMA_signal_7746, new_AGEMA_signal_7745, SubBytesIns_Inst_Sbox_6_M36}), .c ({new_AGEMA_signal_7924, new_AGEMA_signal_7923, SubBytesIns_Inst_Sbox_6_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M41_U1 ( .a ({new_AGEMA_signal_7920, new_AGEMA_signal_7919, SubBytesIns_Inst_Sbox_6_M38}), .b ({new_AGEMA_signal_7924, new_AGEMA_signal_7923, SubBytesIns_Inst_Sbox_6_M40}), .c ({new_AGEMA_signal_8238, new_AGEMA_signal_8237, SubBytesIns_Inst_Sbox_6_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M42_U1 ( .a ({new_AGEMA_signal_7918, new_AGEMA_signal_7917, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_7922, new_AGEMA_signal_7921, SubBytesIns_Inst_Sbox_6_M39}), .c ({new_AGEMA_signal_8240, new_AGEMA_signal_8239, SubBytesIns_Inst_Sbox_6_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M43_U1 ( .a ({new_AGEMA_signal_7918, new_AGEMA_signal_7917, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_7920, new_AGEMA_signal_7919, SubBytesIns_Inst_Sbox_6_M38}), .c ({new_AGEMA_signal_8242, new_AGEMA_signal_8241, SubBytesIns_Inst_Sbox_6_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M44_U1 ( .a ({new_AGEMA_signal_7922, new_AGEMA_signal_7921, SubBytesIns_Inst_Sbox_6_M39}), .b ({new_AGEMA_signal_7924, new_AGEMA_signal_7923, SubBytesIns_Inst_Sbox_6_M40}), .c ({new_AGEMA_signal_8244, new_AGEMA_signal_8243, SubBytesIns_Inst_Sbox_6_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M45_U1 ( .a ({new_AGEMA_signal_8240, new_AGEMA_signal_8239, SubBytesIns_Inst_Sbox_6_M42}), .b ({new_AGEMA_signal_8238, new_AGEMA_signal_8237, SubBytesIns_Inst_Sbox_6_M41}), .c ({new_AGEMA_signal_8718, new_AGEMA_signal_8717, SubBytesIns_Inst_Sbox_6_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M29_U1 ( .a ({new_AGEMA_signal_7552, new_AGEMA_signal_7551, SubBytesIns_Inst_Sbox_7_M28}), .b ({new_AGEMA_signal_7370, new_AGEMA_signal_7369, SubBytesIns_Inst_Sbox_7_M27}), .clk (clk), .r ({Fresh[806], Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_7748, new_AGEMA_signal_7747, SubBytesIns_Inst_Sbox_7_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M30_U1 ( .a ({new_AGEMA_signal_7550, new_AGEMA_signal_7549, SubBytesIns_Inst_Sbox_7_M26}), .b ({new_AGEMA_signal_7548, new_AGEMA_signal_7547, SubBytesIns_Inst_Sbox_7_M24}), .clk (clk), .r ({Fresh[809], Fresh[808], Fresh[807]}), .c ({new_AGEMA_signal_7750, new_AGEMA_signal_7749, SubBytesIns_Inst_Sbox_7_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M32_U1 ( .a ({new_AGEMA_signal_7370, new_AGEMA_signal_7369, SubBytesIns_Inst_Sbox_7_M27}), .b ({new_AGEMA_signal_7554, new_AGEMA_signal_7553, SubBytesIns_Inst_Sbox_7_M31}), .clk (clk), .r ({Fresh[812], Fresh[811], Fresh[810]}), .c ({new_AGEMA_signal_7752, new_AGEMA_signal_7751, SubBytesIns_Inst_Sbox_7_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M35_U1 ( .a ({new_AGEMA_signal_7548, new_AGEMA_signal_7547, SubBytesIns_Inst_Sbox_7_M24}), .b ({new_AGEMA_signal_7372, new_AGEMA_signal_7371, SubBytesIns_Inst_Sbox_7_M34}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813]}), .c ({new_AGEMA_signal_7754, new_AGEMA_signal_7753, SubBytesIns_Inst_Sbox_7_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M37_U1 ( .a ({new_AGEMA_signal_7210, new_AGEMA_signal_7209, SubBytesIns_Inst_Sbox_7_M21}), .b ({new_AGEMA_signal_7748, new_AGEMA_signal_7747, SubBytesIns_Inst_Sbox_7_M29}), .c ({new_AGEMA_signal_7926, new_AGEMA_signal_7925, SubBytesIns_Inst_Sbox_7_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M38_U1 ( .a ({new_AGEMA_signal_7752, new_AGEMA_signal_7751, SubBytesIns_Inst_Sbox_7_M32}), .b ({new_AGEMA_signal_7556, new_AGEMA_signal_7555, SubBytesIns_Inst_Sbox_7_M33}), .c ({new_AGEMA_signal_7928, new_AGEMA_signal_7927, SubBytesIns_Inst_Sbox_7_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M39_U1 ( .a ({new_AGEMA_signal_7366, new_AGEMA_signal_7365, SubBytesIns_Inst_Sbox_7_M23}), .b ({new_AGEMA_signal_7750, new_AGEMA_signal_7749, SubBytesIns_Inst_Sbox_7_M30}), .c ({new_AGEMA_signal_7930, new_AGEMA_signal_7929, SubBytesIns_Inst_Sbox_7_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M40_U1 ( .a ({new_AGEMA_signal_7754, new_AGEMA_signal_7753, SubBytesIns_Inst_Sbox_7_M35}), .b ({new_AGEMA_signal_7756, new_AGEMA_signal_7755, SubBytesIns_Inst_Sbox_7_M36}), .c ({new_AGEMA_signal_7932, new_AGEMA_signal_7931, SubBytesIns_Inst_Sbox_7_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M41_U1 ( .a ({new_AGEMA_signal_7928, new_AGEMA_signal_7927, SubBytesIns_Inst_Sbox_7_M38}), .b ({new_AGEMA_signal_7932, new_AGEMA_signal_7931, SubBytesIns_Inst_Sbox_7_M40}), .c ({new_AGEMA_signal_8262, new_AGEMA_signal_8261, SubBytesIns_Inst_Sbox_7_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M42_U1 ( .a ({new_AGEMA_signal_7926, new_AGEMA_signal_7925, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_7930, new_AGEMA_signal_7929, SubBytesIns_Inst_Sbox_7_M39}), .c ({new_AGEMA_signal_8264, new_AGEMA_signal_8263, SubBytesIns_Inst_Sbox_7_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M43_U1 ( .a ({new_AGEMA_signal_7926, new_AGEMA_signal_7925, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_7928, new_AGEMA_signal_7927, SubBytesIns_Inst_Sbox_7_M38}), .c ({new_AGEMA_signal_8266, new_AGEMA_signal_8265, SubBytesIns_Inst_Sbox_7_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M44_U1 ( .a ({new_AGEMA_signal_7930, new_AGEMA_signal_7929, SubBytesIns_Inst_Sbox_7_M39}), .b ({new_AGEMA_signal_7932, new_AGEMA_signal_7931, SubBytesIns_Inst_Sbox_7_M40}), .c ({new_AGEMA_signal_8268, new_AGEMA_signal_8267, SubBytesIns_Inst_Sbox_7_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M45_U1 ( .a ({new_AGEMA_signal_8264, new_AGEMA_signal_8263, SubBytesIns_Inst_Sbox_7_M42}), .b ({new_AGEMA_signal_8262, new_AGEMA_signal_8261, SubBytesIns_Inst_Sbox_7_M41}), .c ({new_AGEMA_signal_8742, new_AGEMA_signal_8741, SubBytesIns_Inst_Sbox_7_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M29_U1 ( .a ({new_AGEMA_signal_7562, new_AGEMA_signal_7561, SubBytesIns_Inst_Sbox_8_M28}), .b ({new_AGEMA_signal_7378, new_AGEMA_signal_7377, SubBytesIns_Inst_Sbox_8_M27}), .clk (clk), .r ({Fresh[818], Fresh[817], Fresh[816]}), .c ({new_AGEMA_signal_7758, new_AGEMA_signal_7757, SubBytesIns_Inst_Sbox_8_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M30_U1 ( .a ({new_AGEMA_signal_7560, new_AGEMA_signal_7559, SubBytesIns_Inst_Sbox_8_M26}), .b ({new_AGEMA_signal_7558, new_AGEMA_signal_7557, SubBytesIns_Inst_Sbox_8_M24}), .clk (clk), .r ({Fresh[821], Fresh[820], Fresh[819]}), .c ({new_AGEMA_signal_7760, new_AGEMA_signal_7759, SubBytesIns_Inst_Sbox_8_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M32_U1 ( .a ({new_AGEMA_signal_7378, new_AGEMA_signal_7377, SubBytesIns_Inst_Sbox_8_M27}), .b ({new_AGEMA_signal_7564, new_AGEMA_signal_7563, SubBytesIns_Inst_Sbox_8_M31}), .clk (clk), .r ({Fresh[824], Fresh[823], Fresh[822]}), .c ({new_AGEMA_signal_7762, new_AGEMA_signal_7761, SubBytesIns_Inst_Sbox_8_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M35_U1 ( .a ({new_AGEMA_signal_7558, new_AGEMA_signal_7557, SubBytesIns_Inst_Sbox_8_M24}), .b ({new_AGEMA_signal_7380, new_AGEMA_signal_7379, SubBytesIns_Inst_Sbox_8_M34}), .clk (clk), .r ({Fresh[827], Fresh[826], Fresh[825]}), .c ({new_AGEMA_signal_7764, new_AGEMA_signal_7763, SubBytesIns_Inst_Sbox_8_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M37_U1 ( .a ({new_AGEMA_signal_7218, new_AGEMA_signal_7217, SubBytesIns_Inst_Sbox_8_M21}), .b ({new_AGEMA_signal_7758, new_AGEMA_signal_7757, SubBytesIns_Inst_Sbox_8_M29}), .c ({new_AGEMA_signal_7934, new_AGEMA_signal_7933, SubBytesIns_Inst_Sbox_8_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M38_U1 ( .a ({new_AGEMA_signal_7762, new_AGEMA_signal_7761, SubBytesIns_Inst_Sbox_8_M32}), .b ({new_AGEMA_signal_7566, new_AGEMA_signal_7565, SubBytesIns_Inst_Sbox_8_M33}), .c ({new_AGEMA_signal_7936, new_AGEMA_signal_7935, SubBytesIns_Inst_Sbox_8_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M39_U1 ( .a ({new_AGEMA_signal_7374, new_AGEMA_signal_7373, SubBytesIns_Inst_Sbox_8_M23}), .b ({new_AGEMA_signal_7760, new_AGEMA_signal_7759, SubBytesIns_Inst_Sbox_8_M30}), .c ({new_AGEMA_signal_7938, new_AGEMA_signal_7937, SubBytesIns_Inst_Sbox_8_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M40_U1 ( .a ({new_AGEMA_signal_7764, new_AGEMA_signal_7763, SubBytesIns_Inst_Sbox_8_M35}), .b ({new_AGEMA_signal_7766, new_AGEMA_signal_7765, SubBytesIns_Inst_Sbox_8_M36}), .c ({new_AGEMA_signal_7940, new_AGEMA_signal_7939, SubBytesIns_Inst_Sbox_8_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M41_U1 ( .a ({new_AGEMA_signal_7936, new_AGEMA_signal_7935, SubBytesIns_Inst_Sbox_8_M38}), .b ({new_AGEMA_signal_7940, new_AGEMA_signal_7939, SubBytesIns_Inst_Sbox_8_M40}), .c ({new_AGEMA_signal_8286, new_AGEMA_signal_8285, SubBytesIns_Inst_Sbox_8_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M42_U1 ( .a ({new_AGEMA_signal_7934, new_AGEMA_signal_7933, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_7938, new_AGEMA_signal_7937, SubBytesIns_Inst_Sbox_8_M39}), .c ({new_AGEMA_signal_8288, new_AGEMA_signal_8287, SubBytesIns_Inst_Sbox_8_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M43_U1 ( .a ({new_AGEMA_signal_7934, new_AGEMA_signal_7933, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_7936, new_AGEMA_signal_7935, SubBytesIns_Inst_Sbox_8_M38}), .c ({new_AGEMA_signal_8290, new_AGEMA_signal_8289, SubBytesIns_Inst_Sbox_8_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M44_U1 ( .a ({new_AGEMA_signal_7938, new_AGEMA_signal_7937, SubBytesIns_Inst_Sbox_8_M39}), .b ({new_AGEMA_signal_7940, new_AGEMA_signal_7939, SubBytesIns_Inst_Sbox_8_M40}), .c ({new_AGEMA_signal_8292, new_AGEMA_signal_8291, SubBytesIns_Inst_Sbox_8_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M45_U1 ( .a ({new_AGEMA_signal_8288, new_AGEMA_signal_8287, SubBytesIns_Inst_Sbox_8_M42}), .b ({new_AGEMA_signal_8286, new_AGEMA_signal_8285, SubBytesIns_Inst_Sbox_8_M41}), .c ({new_AGEMA_signal_8766, new_AGEMA_signal_8765, SubBytesIns_Inst_Sbox_8_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M29_U1 ( .a ({new_AGEMA_signal_7572, new_AGEMA_signal_7571, SubBytesIns_Inst_Sbox_9_M28}), .b ({new_AGEMA_signal_7386, new_AGEMA_signal_7385, SubBytesIns_Inst_Sbox_9_M27}), .clk (clk), .r ({Fresh[830], Fresh[829], Fresh[828]}), .c ({new_AGEMA_signal_7768, new_AGEMA_signal_7767, SubBytesIns_Inst_Sbox_9_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M30_U1 ( .a ({new_AGEMA_signal_7570, new_AGEMA_signal_7569, SubBytesIns_Inst_Sbox_9_M26}), .b ({new_AGEMA_signal_7568, new_AGEMA_signal_7567, SubBytesIns_Inst_Sbox_9_M24}), .clk (clk), .r ({Fresh[833], Fresh[832], Fresh[831]}), .c ({new_AGEMA_signal_7770, new_AGEMA_signal_7769, SubBytesIns_Inst_Sbox_9_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M32_U1 ( .a ({new_AGEMA_signal_7386, new_AGEMA_signal_7385, SubBytesIns_Inst_Sbox_9_M27}), .b ({new_AGEMA_signal_7574, new_AGEMA_signal_7573, SubBytesIns_Inst_Sbox_9_M31}), .clk (clk), .r ({Fresh[836], Fresh[835], Fresh[834]}), .c ({new_AGEMA_signal_7772, new_AGEMA_signal_7771, SubBytesIns_Inst_Sbox_9_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M35_U1 ( .a ({new_AGEMA_signal_7568, new_AGEMA_signal_7567, SubBytesIns_Inst_Sbox_9_M24}), .b ({new_AGEMA_signal_7388, new_AGEMA_signal_7387, SubBytesIns_Inst_Sbox_9_M34}), .clk (clk), .r ({Fresh[839], Fresh[838], Fresh[837]}), .c ({new_AGEMA_signal_7774, new_AGEMA_signal_7773, SubBytesIns_Inst_Sbox_9_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M37_U1 ( .a ({new_AGEMA_signal_7226, new_AGEMA_signal_7225, SubBytesIns_Inst_Sbox_9_M21}), .b ({new_AGEMA_signal_7768, new_AGEMA_signal_7767, SubBytesIns_Inst_Sbox_9_M29}), .c ({new_AGEMA_signal_7942, new_AGEMA_signal_7941, SubBytesIns_Inst_Sbox_9_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M38_U1 ( .a ({new_AGEMA_signal_7772, new_AGEMA_signal_7771, SubBytesIns_Inst_Sbox_9_M32}), .b ({new_AGEMA_signal_7576, new_AGEMA_signal_7575, SubBytesIns_Inst_Sbox_9_M33}), .c ({new_AGEMA_signal_7944, new_AGEMA_signal_7943, SubBytesIns_Inst_Sbox_9_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M39_U1 ( .a ({new_AGEMA_signal_7382, new_AGEMA_signal_7381, SubBytesIns_Inst_Sbox_9_M23}), .b ({new_AGEMA_signal_7770, new_AGEMA_signal_7769, SubBytesIns_Inst_Sbox_9_M30}), .c ({new_AGEMA_signal_7946, new_AGEMA_signal_7945, SubBytesIns_Inst_Sbox_9_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M40_U1 ( .a ({new_AGEMA_signal_7774, new_AGEMA_signal_7773, SubBytesIns_Inst_Sbox_9_M35}), .b ({new_AGEMA_signal_7776, new_AGEMA_signal_7775, SubBytesIns_Inst_Sbox_9_M36}), .c ({new_AGEMA_signal_7948, new_AGEMA_signal_7947, SubBytesIns_Inst_Sbox_9_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M41_U1 ( .a ({new_AGEMA_signal_7944, new_AGEMA_signal_7943, SubBytesIns_Inst_Sbox_9_M38}), .b ({new_AGEMA_signal_7948, new_AGEMA_signal_7947, SubBytesIns_Inst_Sbox_9_M40}), .c ({new_AGEMA_signal_8310, new_AGEMA_signal_8309, SubBytesIns_Inst_Sbox_9_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M42_U1 ( .a ({new_AGEMA_signal_7942, new_AGEMA_signal_7941, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_7946, new_AGEMA_signal_7945, SubBytesIns_Inst_Sbox_9_M39}), .c ({new_AGEMA_signal_8312, new_AGEMA_signal_8311, SubBytesIns_Inst_Sbox_9_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M43_U1 ( .a ({new_AGEMA_signal_7942, new_AGEMA_signal_7941, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_7944, new_AGEMA_signal_7943, SubBytesIns_Inst_Sbox_9_M38}), .c ({new_AGEMA_signal_8314, new_AGEMA_signal_8313, SubBytesIns_Inst_Sbox_9_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M44_U1 ( .a ({new_AGEMA_signal_7946, new_AGEMA_signal_7945, SubBytesIns_Inst_Sbox_9_M39}), .b ({new_AGEMA_signal_7948, new_AGEMA_signal_7947, SubBytesIns_Inst_Sbox_9_M40}), .c ({new_AGEMA_signal_8316, new_AGEMA_signal_8315, SubBytesIns_Inst_Sbox_9_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M45_U1 ( .a ({new_AGEMA_signal_8312, new_AGEMA_signal_8311, SubBytesIns_Inst_Sbox_9_M42}), .b ({new_AGEMA_signal_8310, new_AGEMA_signal_8309, SubBytesIns_Inst_Sbox_9_M41}), .c ({new_AGEMA_signal_8790, new_AGEMA_signal_8789, SubBytesIns_Inst_Sbox_9_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M29_U1 ( .a ({new_AGEMA_signal_7582, new_AGEMA_signal_7581, SubBytesIns_Inst_Sbox_10_M28}), .b ({new_AGEMA_signal_7394, new_AGEMA_signal_7393, SubBytesIns_Inst_Sbox_10_M27}), .clk (clk), .r ({Fresh[842], Fresh[841], Fresh[840]}), .c ({new_AGEMA_signal_7778, new_AGEMA_signal_7777, SubBytesIns_Inst_Sbox_10_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M30_U1 ( .a ({new_AGEMA_signal_7580, new_AGEMA_signal_7579, SubBytesIns_Inst_Sbox_10_M26}), .b ({new_AGEMA_signal_7578, new_AGEMA_signal_7577, SubBytesIns_Inst_Sbox_10_M24}), .clk (clk), .r ({Fresh[845], Fresh[844], Fresh[843]}), .c ({new_AGEMA_signal_7780, new_AGEMA_signal_7779, SubBytesIns_Inst_Sbox_10_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M32_U1 ( .a ({new_AGEMA_signal_7394, new_AGEMA_signal_7393, SubBytesIns_Inst_Sbox_10_M27}), .b ({new_AGEMA_signal_7584, new_AGEMA_signal_7583, SubBytesIns_Inst_Sbox_10_M31}), .clk (clk), .r ({Fresh[848], Fresh[847], Fresh[846]}), .c ({new_AGEMA_signal_7782, new_AGEMA_signal_7781, SubBytesIns_Inst_Sbox_10_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M35_U1 ( .a ({new_AGEMA_signal_7578, new_AGEMA_signal_7577, SubBytesIns_Inst_Sbox_10_M24}), .b ({new_AGEMA_signal_7396, new_AGEMA_signal_7395, SubBytesIns_Inst_Sbox_10_M34}), .clk (clk), .r ({Fresh[851], Fresh[850], Fresh[849]}), .c ({new_AGEMA_signal_7784, new_AGEMA_signal_7783, SubBytesIns_Inst_Sbox_10_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M37_U1 ( .a ({new_AGEMA_signal_7234, new_AGEMA_signal_7233, SubBytesIns_Inst_Sbox_10_M21}), .b ({new_AGEMA_signal_7778, new_AGEMA_signal_7777, SubBytesIns_Inst_Sbox_10_M29}), .c ({new_AGEMA_signal_7950, new_AGEMA_signal_7949, SubBytesIns_Inst_Sbox_10_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M38_U1 ( .a ({new_AGEMA_signal_7782, new_AGEMA_signal_7781, SubBytesIns_Inst_Sbox_10_M32}), .b ({new_AGEMA_signal_7586, new_AGEMA_signal_7585, SubBytesIns_Inst_Sbox_10_M33}), .c ({new_AGEMA_signal_7952, new_AGEMA_signal_7951, SubBytesIns_Inst_Sbox_10_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M39_U1 ( .a ({new_AGEMA_signal_7390, new_AGEMA_signal_7389, SubBytesIns_Inst_Sbox_10_M23}), .b ({new_AGEMA_signal_7780, new_AGEMA_signal_7779, SubBytesIns_Inst_Sbox_10_M30}), .c ({new_AGEMA_signal_7954, new_AGEMA_signal_7953, SubBytesIns_Inst_Sbox_10_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M40_U1 ( .a ({new_AGEMA_signal_7784, new_AGEMA_signal_7783, SubBytesIns_Inst_Sbox_10_M35}), .b ({new_AGEMA_signal_7786, new_AGEMA_signal_7785, SubBytesIns_Inst_Sbox_10_M36}), .c ({new_AGEMA_signal_7956, new_AGEMA_signal_7955, SubBytesIns_Inst_Sbox_10_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M41_U1 ( .a ({new_AGEMA_signal_7952, new_AGEMA_signal_7951, SubBytesIns_Inst_Sbox_10_M38}), .b ({new_AGEMA_signal_7956, new_AGEMA_signal_7955, SubBytesIns_Inst_Sbox_10_M40}), .c ({new_AGEMA_signal_8334, new_AGEMA_signal_8333, SubBytesIns_Inst_Sbox_10_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M42_U1 ( .a ({new_AGEMA_signal_7950, new_AGEMA_signal_7949, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_7954, new_AGEMA_signal_7953, SubBytesIns_Inst_Sbox_10_M39}), .c ({new_AGEMA_signal_8336, new_AGEMA_signal_8335, SubBytesIns_Inst_Sbox_10_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M43_U1 ( .a ({new_AGEMA_signal_7950, new_AGEMA_signal_7949, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_7952, new_AGEMA_signal_7951, SubBytesIns_Inst_Sbox_10_M38}), .c ({new_AGEMA_signal_8338, new_AGEMA_signal_8337, SubBytesIns_Inst_Sbox_10_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M44_U1 ( .a ({new_AGEMA_signal_7954, new_AGEMA_signal_7953, SubBytesIns_Inst_Sbox_10_M39}), .b ({new_AGEMA_signal_7956, new_AGEMA_signal_7955, SubBytesIns_Inst_Sbox_10_M40}), .c ({new_AGEMA_signal_8340, new_AGEMA_signal_8339, SubBytesIns_Inst_Sbox_10_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M45_U1 ( .a ({new_AGEMA_signal_8336, new_AGEMA_signal_8335, SubBytesIns_Inst_Sbox_10_M42}), .b ({new_AGEMA_signal_8334, new_AGEMA_signal_8333, SubBytesIns_Inst_Sbox_10_M41}), .c ({new_AGEMA_signal_8814, new_AGEMA_signal_8813, SubBytesIns_Inst_Sbox_10_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M29_U1 ( .a ({new_AGEMA_signal_7592, new_AGEMA_signal_7591, SubBytesIns_Inst_Sbox_11_M28}), .b ({new_AGEMA_signal_7402, new_AGEMA_signal_7401, SubBytesIns_Inst_Sbox_11_M27}), .clk (clk), .r ({Fresh[854], Fresh[853], Fresh[852]}), .c ({new_AGEMA_signal_7788, new_AGEMA_signal_7787, SubBytesIns_Inst_Sbox_11_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M30_U1 ( .a ({new_AGEMA_signal_7590, new_AGEMA_signal_7589, SubBytesIns_Inst_Sbox_11_M26}), .b ({new_AGEMA_signal_7588, new_AGEMA_signal_7587, SubBytesIns_Inst_Sbox_11_M24}), .clk (clk), .r ({Fresh[857], Fresh[856], Fresh[855]}), .c ({new_AGEMA_signal_7790, new_AGEMA_signal_7789, SubBytesIns_Inst_Sbox_11_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M32_U1 ( .a ({new_AGEMA_signal_7402, new_AGEMA_signal_7401, SubBytesIns_Inst_Sbox_11_M27}), .b ({new_AGEMA_signal_7594, new_AGEMA_signal_7593, SubBytesIns_Inst_Sbox_11_M31}), .clk (clk), .r ({Fresh[860], Fresh[859], Fresh[858]}), .c ({new_AGEMA_signal_7792, new_AGEMA_signal_7791, SubBytesIns_Inst_Sbox_11_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M35_U1 ( .a ({new_AGEMA_signal_7588, new_AGEMA_signal_7587, SubBytesIns_Inst_Sbox_11_M24}), .b ({new_AGEMA_signal_7404, new_AGEMA_signal_7403, SubBytesIns_Inst_Sbox_11_M34}), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861]}), .c ({new_AGEMA_signal_7794, new_AGEMA_signal_7793, SubBytesIns_Inst_Sbox_11_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M37_U1 ( .a ({new_AGEMA_signal_7242, new_AGEMA_signal_7241, SubBytesIns_Inst_Sbox_11_M21}), .b ({new_AGEMA_signal_7788, new_AGEMA_signal_7787, SubBytesIns_Inst_Sbox_11_M29}), .c ({new_AGEMA_signal_7958, new_AGEMA_signal_7957, SubBytesIns_Inst_Sbox_11_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M38_U1 ( .a ({new_AGEMA_signal_7792, new_AGEMA_signal_7791, SubBytesIns_Inst_Sbox_11_M32}), .b ({new_AGEMA_signal_7596, new_AGEMA_signal_7595, SubBytesIns_Inst_Sbox_11_M33}), .c ({new_AGEMA_signal_7960, new_AGEMA_signal_7959, SubBytesIns_Inst_Sbox_11_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M39_U1 ( .a ({new_AGEMA_signal_7398, new_AGEMA_signal_7397, SubBytesIns_Inst_Sbox_11_M23}), .b ({new_AGEMA_signal_7790, new_AGEMA_signal_7789, SubBytesIns_Inst_Sbox_11_M30}), .c ({new_AGEMA_signal_7962, new_AGEMA_signal_7961, SubBytesIns_Inst_Sbox_11_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M40_U1 ( .a ({new_AGEMA_signal_7794, new_AGEMA_signal_7793, SubBytesIns_Inst_Sbox_11_M35}), .b ({new_AGEMA_signal_7796, new_AGEMA_signal_7795, SubBytesIns_Inst_Sbox_11_M36}), .c ({new_AGEMA_signal_7964, new_AGEMA_signal_7963, SubBytesIns_Inst_Sbox_11_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M41_U1 ( .a ({new_AGEMA_signal_7960, new_AGEMA_signal_7959, SubBytesIns_Inst_Sbox_11_M38}), .b ({new_AGEMA_signal_7964, new_AGEMA_signal_7963, SubBytesIns_Inst_Sbox_11_M40}), .c ({new_AGEMA_signal_8358, new_AGEMA_signal_8357, SubBytesIns_Inst_Sbox_11_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M42_U1 ( .a ({new_AGEMA_signal_7958, new_AGEMA_signal_7957, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_7962, new_AGEMA_signal_7961, SubBytesIns_Inst_Sbox_11_M39}), .c ({new_AGEMA_signal_8360, new_AGEMA_signal_8359, SubBytesIns_Inst_Sbox_11_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M43_U1 ( .a ({new_AGEMA_signal_7958, new_AGEMA_signal_7957, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_7960, new_AGEMA_signal_7959, SubBytesIns_Inst_Sbox_11_M38}), .c ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, SubBytesIns_Inst_Sbox_11_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M44_U1 ( .a ({new_AGEMA_signal_7962, new_AGEMA_signal_7961, SubBytesIns_Inst_Sbox_11_M39}), .b ({new_AGEMA_signal_7964, new_AGEMA_signal_7963, SubBytesIns_Inst_Sbox_11_M40}), .c ({new_AGEMA_signal_8364, new_AGEMA_signal_8363, SubBytesIns_Inst_Sbox_11_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M45_U1 ( .a ({new_AGEMA_signal_8360, new_AGEMA_signal_8359, SubBytesIns_Inst_Sbox_11_M42}), .b ({new_AGEMA_signal_8358, new_AGEMA_signal_8357, SubBytesIns_Inst_Sbox_11_M41}), .c ({new_AGEMA_signal_8838, new_AGEMA_signal_8837, SubBytesIns_Inst_Sbox_11_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M29_U1 ( .a ({new_AGEMA_signal_7602, new_AGEMA_signal_7601, SubBytesIns_Inst_Sbox_12_M28}), .b ({new_AGEMA_signal_7410, new_AGEMA_signal_7409, SubBytesIns_Inst_Sbox_12_M27}), .clk (clk), .r ({Fresh[866], Fresh[865], Fresh[864]}), .c ({new_AGEMA_signal_7798, new_AGEMA_signal_7797, SubBytesIns_Inst_Sbox_12_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M30_U1 ( .a ({new_AGEMA_signal_7600, new_AGEMA_signal_7599, SubBytesIns_Inst_Sbox_12_M26}), .b ({new_AGEMA_signal_7598, new_AGEMA_signal_7597, SubBytesIns_Inst_Sbox_12_M24}), .clk (clk), .r ({Fresh[869], Fresh[868], Fresh[867]}), .c ({new_AGEMA_signal_7800, new_AGEMA_signal_7799, SubBytesIns_Inst_Sbox_12_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M32_U1 ( .a ({new_AGEMA_signal_7410, new_AGEMA_signal_7409, SubBytesIns_Inst_Sbox_12_M27}), .b ({new_AGEMA_signal_7604, new_AGEMA_signal_7603, SubBytesIns_Inst_Sbox_12_M31}), .clk (clk), .r ({Fresh[872], Fresh[871], Fresh[870]}), .c ({new_AGEMA_signal_7802, new_AGEMA_signal_7801, SubBytesIns_Inst_Sbox_12_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M35_U1 ( .a ({new_AGEMA_signal_7598, new_AGEMA_signal_7597, SubBytesIns_Inst_Sbox_12_M24}), .b ({new_AGEMA_signal_7412, new_AGEMA_signal_7411, SubBytesIns_Inst_Sbox_12_M34}), .clk (clk), .r ({Fresh[875], Fresh[874], Fresh[873]}), .c ({new_AGEMA_signal_7804, new_AGEMA_signal_7803, SubBytesIns_Inst_Sbox_12_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M37_U1 ( .a ({new_AGEMA_signal_7250, new_AGEMA_signal_7249, SubBytesIns_Inst_Sbox_12_M21}), .b ({new_AGEMA_signal_7798, new_AGEMA_signal_7797, SubBytesIns_Inst_Sbox_12_M29}), .c ({new_AGEMA_signal_7966, new_AGEMA_signal_7965, SubBytesIns_Inst_Sbox_12_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M38_U1 ( .a ({new_AGEMA_signal_7802, new_AGEMA_signal_7801, SubBytesIns_Inst_Sbox_12_M32}), .b ({new_AGEMA_signal_7606, new_AGEMA_signal_7605, SubBytesIns_Inst_Sbox_12_M33}), .c ({new_AGEMA_signal_7968, new_AGEMA_signal_7967, SubBytesIns_Inst_Sbox_12_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M39_U1 ( .a ({new_AGEMA_signal_7406, new_AGEMA_signal_7405, SubBytesIns_Inst_Sbox_12_M23}), .b ({new_AGEMA_signal_7800, new_AGEMA_signal_7799, SubBytesIns_Inst_Sbox_12_M30}), .c ({new_AGEMA_signal_7970, new_AGEMA_signal_7969, SubBytesIns_Inst_Sbox_12_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M40_U1 ( .a ({new_AGEMA_signal_7804, new_AGEMA_signal_7803, SubBytesIns_Inst_Sbox_12_M35}), .b ({new_AGEMA_signal_7806, new_AGEMA_signal_7805, SubBytesIns_Inst_Sbox_12_M36}), .c ({new_AGEMA_signal_7972, new_AGEMA_signal_7971, SubBytesIns_Inst_Sbox_12_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M41_U1 ( .a ({new_AGEMA_signal_7968, new_AGEMA_signal_7967, SubBytesIns_Inst_Sbox_12_M38}), .b ({new_AGEMA_signal_7972, new_AGEMA_signal_7971, SubBytesIns_Inst_Sbox_12_M40}), .c ({new_AGEMA_signal_8382, new_AGEMA_signal_8381, SubBytesIns_Inst_Sbox_12_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M42_U1 ( .a ({new_AGEMA_signal_7966, new_AGEMA_signal_7965, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_7970, new_AGEMA_signal_7969, SubBytesIns_Inst_Sbox_12_M39}), .c ({new_AGEMA_signal_8384, new_AGEMA_signal_8383, SubBytesIns_Inst_Sbox_12_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M43_U1 ( .a ({new_AGEMA_signal_7966, new_AGEMA_signal_7965, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_7968, new_AGEMA_signal_7967, SubBytesIns_Inst_Sbox_12_M38}), .c ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, SubBytesIns_Inst_Sbox_12_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M44_U1 ( .a ({new_AGEMA_signal_7970, new_AGEMA_signal_7969, SubBytesIns_Inst_Sbox_12_M39}), .b ({new_AGEMA_signal_7972, new_AGEMA_signal_7971, SubBytesIns_Inst_Sbox_12_M40}), .c ({new_AGEMA_signal_8388, new_AGEMA_signal_8387, SubBytesIns_Inst_Sbox_12_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M45_U1 ( .a ({new_AGEMA_signal_8384, new_AGEMA_signal_8383, SubBytesIns_Inst_Sbox_12_M42}), .b ({new_AGEMA_signal_8382, new_AGEMA_signal_8381, SubBytesIns_Inst_Sbox_12_M41}), .c ({new_AGEMA_signal_8862, new_AGEMA_signal_8861, SubBytesIns_Inst_Sbox_12_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M29_U1 ( .a ({new_AGEMA_signal_7612, new_AGEMA_signal_7611, SubBytesIns_Inst_Sbox_13_M28}), .b ({new_AGEMA_signal_7418, new_AGEMA_signal_7417, SubBytesIns_Inst_Sbox_13_M27}), .clk (clk), .r ({Fresh[878], Fresh[877], Fresh[876]}), .c ({new_AGEMA_signal_7808, new_AGEMA_signal_7807, SubBytesIns_Inst_Sbox_13_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M30_U1 ( .a ({new_AGEMA_signal_7610, new_AGEMA_signal_7609, SubBytesIns_Inst_Sbox_13_M26}), .b ({new_AGEMA_signal_7608, new_AGEMA_signal_7607, SubBytesIns_Inst_Sbox_13_M24}), .clk (clk), .r ({Fresh[881], Fresh[880], Fresh[879]}), .c ({new_AGEMA_signal_7810, new_AGEMA_signal_7809, SubBytesIns_Inst_Sbox_13_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M32_U1 ( .a ({new_AGEMA_signal_7418, new_AGEMA_signal_7417, SubBytesIns_Inst_Sbox_13_M27}), .b ({new_AGEMA_signal_7614, new_AGEMA_signal_7613, SubBytesIns_Inst_Sbox_13_M31}), .clk (clk), .r ({Fresh[884], Fresh[883], Fresh[882]}), .c ({new_AGEMA_signal_7812, new_AGEMA_signal_7811, SubBytesIns_Inst_Sbox_13_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M35_U1 ( .a ({new_AGEMA_signal_7608, new_AGEMA_signal_7607, SubBytesIns_Inst_Sbox_13_M24}), .b ({new_AGEMA_signal_7420, new_AGEMA_signal_7419, SubBytesIns_Inst_Sbox_13_M34}), .clk (clk), .r ({Fresh[887], Fresh[886], Fresh[885]}), .c ({new_AGEMA_signal_7814, new_AGEMA_signal_7813, SubBytesIns_Inst_Sbox_13_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M37_U1 ( .a ({new_AGEMA_signal_7258, new_AGEMA_signal_7257, SubBytesIns_Inst_Sbox_13_M21}), .b ({new_AGEMA_signal_7808, new_AGEMA_signal_7807, SubBytesIns_Inst_Sbox_13_M29}), .c ({new_AGEMA_signal_7974, new_AGEMA_signal_7973, SubBytesIns_Inst_Sbox_13_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M38_U1 ( .a ({new_AGEMA_signal_7812, new_AGEMA_signal_7811, SubBytesIns_Inst_Sbox_13_M32}), .b ({new_AGEMA_signal_7616, new_AGEMA_signal_7615, SubBytesIns_Inst_Sbox_13_M33}), .c ({new_AGEMA_signal_7976, new_AGEMA_signal_7975, SubBytesIns_Inst_Sbox_13_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M39_U1 ( .a ({new_AGEMA_signal_7414, new_AGEMA_signal_7413, SubBytesIns_Inst_Sbox_13_M23}), .b ({new_AGEMA_signal_7810, new_AGEMA_signal_7809, SubBytesIns_Inst_Sbox_13_M30}), .c ({new_AGEMA_signal_7978, new_AGEMA_signal_7977, SubBytesIns_Inst_Sbox_13_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M40_U1 ( .a ({new_AGEMA_signal_7814, new_AGEMA_signal_7813, SubBytesIns_Inst_Sbox_13_M35}), .b ({new_AGEMA_signal_7816, new_AGEMA_signal_7815, SubBytesIns_Inst_Sbox_13_M36}), .c ({new_AGEMA_signal_7980, new_AGEMA_signal_7979, SubBytesIns_Inst_Sbox_13_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M41_U1 ( .a ({new_AGEMA_signal_7976, new_AGEMA_signal_7975, SubBytesIns_Inst_Sbox_13_M38}), .b ({new_AGEMA_signal_7980, new_AGEMA_signal_7979, SubBytesIns_Inst_Sbox_13_M40}), .c ({new_AGEMA_signal_8406, new_AGEMA_signal_8405, SubBytesIns_Inst_Sbox_13_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M42_U1 ( .a ({new_AGEMA_signal_7974, new_AGEMA_signal_7973, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_7978, new_AGEMA_signal_7977, SubBytesIns_Inst_Sbox_13_M39}), .c ({new_AGEMA_signal_8408, new_AGEMA_signal_8407, SubBytesIns_Inst_Sbox_13_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M43_U1 ( .a ({new_AGEMA_signal_7974, new_AGEMA_signal_7973, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_7976, new_AGEMA_signal_7975, SubBytesIns_Inst_Sbox_13_M38}), .c ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, SubBytesIns_Inst_Sbox_13_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M44_U1 ( .a ({new_AGEMA_signal_7978, new_AGEMA_signal_7977, SubBytesIns_Inst_Sbox_13_M39}), .b ({new_AGEMA_signal_7980, new_AGEMA_signal_7979, SubBytesIns_Inst_Sbox_13_M40}), .c ({new_AGEMA_signal_8412, new_AGEMA_signal_8411, SubBytesIns_Inst_Sbox_13_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M45_U1 ( .a ({new_AGEMA_signal_8408, new_AGEMA_signal_8407, SubBytesIns_Inst_Sbox_13_M42}), .b ({new_AGEMA_signal_8406, new_AGEMA_signal_8405, SubBytesIns_Inst_Sbox_13_M41}), .c ({new_AGEMA_signal_8886, new_AGEMA_signal_8885, SubBytesIns_Inst_Sbox_13_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M29_U1 ( .a ({new_AGEMA_signal_7622, new_AGEMA_signal_7621, SubBytesIns_Inst_Sbox_14_M28}), .b ({new_AGEMA_signal_7426, new_AGEMA_signal_7425, SubBytesIns_Inst_Sbox_14_M27}), .clk (clk), .r ({Fresh[890], Fresh[889], Fresh[888]}), .c ({new_AGEMA_signal_7818, new_AGEMA_signal_7817, SubBytesIns_Inst_Sbox_14_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M30_U1 ( .a ({new_AGEMA_signal_7620, new_AGEMA_signal_7619, SubBytesIns_Inst_Sbox_14_M26}), .b ({new_AGEMA_signal_7618, new_AGEMA_signal_7617, SubBytesIns_Inst_Sbox_14_M24}), .clk (clk), .r ({Fresh[893], Fresh[892], Fresh[891]}), .c ({new_AGEMA_signal_7820, new_AGEMA_signal_7819, SubBytesIns_Inst_Sbox_14_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M32_U1 ( .a ({new_AGEMA_signal_7426, new_AGEMA_signal_7425, SubBytesIns_Inst_Sbox_14_M27}), .b ({new_AGEMA_signal_7624, new_AGEMA_signal_7623, SubBytesIns_Inst_Sbox_14_M31}), .clk (clk), .r ({Fresh[896], Fresh[895], Fresh[894]}), .c ({new_AGEMA_signal_7822, new_AGEMA_signal_7821, SubBytesIns_Inst_Sbox_14_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M35_U1 ( .a ({new_AGEMA_signal_7618, new_AGEMA_signal_7617, SubBytesIns_Inst_Sbox_14_M24}), .b ({new_AGEMA_signal_7428, new_AGEMA_signal_7427, SubBytesIns_Inst_Sbox_14_M34}), .clk (clk), .r ({Fresh[899], Fresh[898], Fresh[897]}), .c ({new_AGEMA_signal_7824, new_AGEMA_signal_7823, SubBytesIns_Inst_Sbox_14_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M37_U1 ( .a ({new_AGEMA_signal_7266, new_AGEMA_signal_7265, SubBytesIns_Inst_Sbox_14_M21}), .b ({new_AGEMA_signal_7818, new_AGEMA_signal_7817, SubBytesIns_Inst_Sbox_14_M29}), .c ({new_AGEMA_signal_7982, new_AGEMA_signal_7981, SubBytesIns_Inst_Sbox_14_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M38_U1 ( .a ({new_AGEMA_signal_7822, new_AGEMA_signal_7821, SubBytesIns_Inst_Sbox_14_M32}), .b ({new_AGEMA_signal_7626, new_AGEMA_signal_7625, SubBytesIns_Inst_Sbox_14_M33}), .c ({new_AGEMA_signal_7984, new_AGEMA_signal_7983, SubBytesIns_Inst_Sbox_14_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M39_U1 ( .a ({new_AGEMA_signal_7422, new_AGEMA_signal_7421, SubBytesIns_Inst_Sbox_14_M23}), .b ({new_AGEMA_signal_7820, new_AGEMA_signal_7819, SubBytesIns_Inst_Sbox_14_M30}), .c ({new_AGEMA_signal_7986, new_AGEMA_signal_7985, SubBytesIns_Inst_Sbox_14_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M40_U1 ( .a ({new_AGEMA_signal_7824, new_AGEMA_signal_7823, SubBytesIns_Inst_Sbox_14_M35}), .b ({new_AGEMA_signal_7826, new_AGEMA_signal_7825, SubBytesIns_Inst_Sbox_14_M36}), .c ({new_AGEMA_signal_7988, new_AGEMA_signal_7987, SubBytesIns_Inst_Sbox_14_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M41_U1 ( .a ({new_AGEMA_signal_7984, new_AGEMA_signal_7983, SubBytesIns_Inst_Sbox_14_M38}), .b ({new_AGEMA_signal_7988, new_AGEMA_signal_7987, SubBytesIns_Inst_Sbox_14_M40}), .c ({new_AGEMA_signal_8430, new_AGEMA_signal_8429, SubBytesIns_Inst_Sbox_14_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M42_U1 ( .a ({new_AGEMA_signal_7982, new_AGEMA_signal_7981, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_7986, new_AGEMA_signal_7985, SubBytesIns_Inst_Sbox_14_M39}), .c ({new_AGEMA_signal_8432, new_AGEMA_signal_8431, SubBytesIns_Inst_Sbox_14_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M43_U1 ( .a ({new_AGEMA_signal_7982, new_AGEMA_signal_7981, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_7984, new_AGEMA_signal_7983, SubBytesIns_Inst_Sbox_14_M38}), .c ({new_AGEMA_signal_8434, new_AGEMA_signal_8433, SubBytesIns_Inst_Sbox_14_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M44_U1 ( .a ({new_AGEMA_signal_7986, new_AGEMA_signal_7985, SubBytesIns_Inst_Sbox_14_M39}), .b ({new_AGEMA_signal_7988, new_AGEMA_signal_7987, SubBytesIns_Inst_Sbox_14_M40}), .c ({new_AGEMA_signal_8436, new_AGEMA_signal_8435, SubBytesIns_Inst_Sbox_14_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M45_U1 ( .a ({new_AGEMA_signal_8432, new_AGEMA_signal_8431, SubBytesIns_Inst_Sbox_14_M42}), .b ({new_AGEMA_signal_8430, new_AGEMA_signal_8429, SubBytesIns_Inst_Sbox_14_M41}), .c ({new_AGEMA_signal_8910, new_AGEMA_signal_8909, SubBytesIns_Inst_Sbox_14_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M29_U1 ( .a ({new_AGEMA_signal_7632, new_AGEMA_signal_7631, SubBytesIns_Inst_Sbox_15_M28}), .b ({new_AGEMA_signal_7434, new_AGEMA_signal_7433, SubBytesIns_Inst_Sbox_15_M27}), .clk (clk), .r ({Fresh[902], Fresh[901], Fresh[900]}), .c ({new_AGEMA_signal_7828, new_AGEMA_signal_7827, SubBytesIns_Inst_Sbox_15_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M30_U1 ( .a ({new_AGEMA_signal_7630, new_AGEMA_signal_7629, SubBytesIns_Inst_Sbox_15_M26}), .b ({new_AGEMA_signal_7628, new_AGEMA_signal_7627, SubBytesIns_Inst_Sbox_15_M24}), .clk (clk), .r ({Fresh[905], Fresh[904], Fresh[903]}), .c ({new_AGEMA_signal_7830, new_AGEMA_signal_7829, SubBytesIns_Inst_Sbox_15_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M32_U1 ( .a ({new_AGEMA_signal_7434, new_AGEMA_signal_7433, SubBytesIns_Inst_Sbox_15_M27}), .b ({new_AGEMA_signal_7634, new_AGEMA_signal_7633, SubBytesIns_Inst_Sbox_15_M31}), .clk (clk), .r ({Fresh[908], Fresh[907], Fresh[906]}), .c ({new_AGEMA_signal_7832, new_AGEMA_signal_7831, SubBytesIns_Inst_Sbox_15_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M35_U1 ( .a ({new_AGEMA_signal_7628, new_AGEMA_signal_7627, SubBytesIns_Inst_Sbox_15_M24}), .b ({new_AGEMA_signal_7436, new_AGEMA_signal_7435, SubBytesIns_Inst_Sbox_15_M34}), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909]}), .c ({new_AGEMA_signal_7834, new_AGEMA_signal_7833, SubBytesIns_Inst_Sbox_15_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M37_U1 ( .a ({new_AGEMA_signal_7274, new_AGEMA_signal_7273, SubBytesIns_Inst_Sbox_15_M21}), .b ({new_AGEMA_signal_7828, new_AGEMA_signal_7827, SubBytesIns_Inst_Sbox_15_M29}), .c ({new_AGEMA_signal_7990, new_AGEMA_signal_7989, SubBytesIns_Inst_Sbox_15_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M38_U1 ( .a ({new_AGEMA_signal_7832, new_AGEMA_signal_7831, SubBytesIns_Inst_Sbox_15_M32}), .b ({new_AGEMA_signal_7636, new_AGEMA_signal_7635, SubBytesIns_Inst_Sbox_15_M33}), .c ({new_AGEMA_signal_7992, new_AGEMA_signal_7991, SubBytesIns_Inst_Sbox_15_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M39_U1 ( .a ({new_AGEMA_signal_7430, new_AGEMA_signal_7429, SubBytesIns_Inst_Sbox_15_M23}), .b ({new_AGEMA_signal_7830, new_AGEMA_signal_7829, SubBytesIns_Inst_Sbox_15_M30}), .c ({new_AGEMA_signal_7994, new_AGEMA_signal_7993, SubBytesIns_Inst_Sbox_15_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M40_U1 ( .a ({new_AGEMA_signal_7834, new_AGEMA_signal_7833, SubBytesIns_Inst_Sbox_15_M35}), .b ({new_AGEMA_signal_7836, new_AGEMA_signal_7835, SubBytesIns_Inst_Sbox_15_M36}), .c ({new_AGEMA_signal_7996, new_AGEMA_signal_7995, SubBytesIns_Inst_Sbox_15_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M41_U1 ( .a ({new_AGEMA_signal_7992, new_AGEMA_signal_7991, SubBytesIns_Inst_Sbox_15_M38}), .b ({new_AGEMA_signal_7996, new_AGEMA_signal_7995, SubBytesIns_Inst_Sbox_15_M40}), .c ({new_AGEMA_signal_8454, new_AGEMA_signal_8453, SubBytesIns_Inst_Sbox_15_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M42_U1 ( .a ({new_AGEMA_signal_7990, new_AGEMA_signal_7989, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_7994, new_AGEMA_signal_7993, SubBytesIns_Inst_Sbox_15_M39}), .c ({new_AGEMA_signal_8456, new_AGEMA_signal_8455, SubBytesIns_Inst_Sbox_15_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M43_U1 ( .a ({new_AGEMA_signal_7990, new_AGEMA_signal_7989, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_7992, new_AGEMA_signal_7991, SubBytesIns_Inst_Sbox_15_M38}), .c ({new_AGEMA_signal_8458, new_AGEMA_signal_8457, SubBytesIns_Inst_Sbox_15_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M44_U1 ( .a ({new_AGEMA_signal_7994, new_AGEMA_signal_7993, SubBytesIns_Inst_Sbox_15_M39}), .b ({new_AGEMA_signal_7996, new_AGEMA_signal_7995, SubBytesIns_Inst_Sbox_15_M40}), .c ({new_AGEMA_signal_8460, new_AGEMA_signal_8459, SubBytesIns_Inst_Sbox_15_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M45_U1 ( .a ({new_AGEMA_signal_8456, new_AGEMA_signal_8455, SubBytesIns_Inst_Sbox_15_M42}), .b ({new_AGEMA_signal_8454, new_AGEMA_signal_8453, SubBytesIns_Inst_Sbox_15_M41}), .c ({new_AGEMA_signal_8934, new_AGEMA_signal_8933, SubBytesIns_Inst_Sbox_15_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M29_U1 ( .a ({new_AGEMA_signal_7442, new_AGEMA_signal_7441, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28}), .b ({new_AGEMA_signal_7282, new_AGEMA_signal_7281, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27}), .clk (clk), .r ({Fresh[914], Fresh[913], Fresh[912]}), .c ({new_AGEMA_signal_7638, new_AGEMA_signal_7637, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M30_U1 ( .a ({new_AGEMA_signal_7440, new_AGEMA_signal_7439, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26}), .b ({new_AGEMA_signal_7438, new_AGEMA_signal_7437, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24}), .clk (clk), .r ({Fresh[917], Fresh[916], Fresh[915]}), .c ({new_AGEMA_signal_7640, new_AGEMA_signal_7639, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M32_U1 ( .a ({new_AGEMA_signal_7282, new_AGEMA_signal_7281, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27}), .b ({new_AGEMA_signal_7444, new_AGEMA_signal_7443, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31}), .clk (clk), .r ({Fresh[920], Fresh[919], Fresh[918]}), .c ({new_AGEMA_signal_7642, new_AGEMA_signal_7641, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M35_U1 ( .a ({new_AGEMA_signal_7438, new_AGEMA_signal_7437, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24}), .b ({new_AGEMA_signal_7284, new_AGEMA_signal_7283, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34}), .clk (clk), .r ({Fresh[923], Fresh[922], Fresh[921]}), .c ({new_AGEMA_signal_7644, new_AGEMA_signal_7643, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M37_U1 ( .a ({new_AGEMA_signal_7122, new_AGEMA_signal_7121, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_7638, new_AGEMA_signal_7637, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29}), .c ({new_AGEMA_signal_7838, new_AGEMA_signal_7837, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M38_U1 ( .a ({new_AGEMA_signal_7642, new_AGEMA_signal_7641, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32}), .b ({new_AGEMA_signal_7446, new_AGEMA_signal_7445, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33}), .c ({new_AGEMA_signal_7840, new_AGEMA_signal_7839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M39_U1 ( .a ({new_AGEMA_signal_7278, new_AGEMA_signal_7277, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}), .b ({new_AGEMA_signal_7640, new_AGEMA_signal_7639, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30}), .c ({new_AGEMA_signal_7842, new_AGEMA_signal_7841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M40_U1 ( .a ({new_AGEMA_signal_7644, new_AGEMA_signal_7643, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35}), .b ({new_AGEMA_signal_7646, new_AGEMA_signal_7645, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36}), .c ({new_AGEMA_signal_7844, new_AGEMA_signal_7843, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M41_U1 ( .a ({new_AGEMA_signal_7840, new_AGEMA_signal_7839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_7844, new_AGEMA_signal_7843, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_7998, new_AGEMA_signal_7997, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M42_U1 ( .a ({new_AGEMA_signal_7838, new_AGEMA_signal_7837, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_7842, new_AGEMA_signal_7841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .c ({new_AGEMA_signal_8000, new_AGEMA_signal_7999, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M43_U1 ( .a ({new_AGEMA_signal_7838, new_AGEMA_signal_7837, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_7840, new_AGEMA_signal_7839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .c ({new_AGEMA_signal_8002, new_AGEMA_signal_8001, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M44_U1 ( .a ({new_AGEMA_signal_7842, new_AGEMA_signal_7841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_7844, new_AGEMA_signal_7843, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_8004, new_AGEMA_signal_8003, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M45_U1 ( .a ({new_AGEMA_signal_8000, new_AGEMA_signal_7999, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_7998, new_AGEMA_signal_7997, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}), .c ({new_AGEMA_signal_8478, new_AGEMA_signal_8477, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M29_U1 ( .a ({new_AGEMA_signal_7452, new_AGEMA_signal_7451, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28}), .b ({new_AGEMA_signal_7290, new_AGEMA_signal_7289, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27}), .clk (clk), .r ({Fresh[926], Fresh[925], Fresh[924]}), .c ({new_AGEMA_signal_7648, new_AGEMA_signal_7647, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M30_U1 ( .a ({new_AGEMA_signal_7450, new_AGEMA_signal_7449, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26}), .b ({new_AGEMA_signal_7448, new_AGEMA_signal_7447, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24}), .clk (clk), .r ({Fresh[929], Fresh[928], Fresh[927]}), .c ({new_AGEMA_signal_7650, new_AGEMA_signal_7649, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M32_U1 ( .a ({new_AGEMA_signal_7290, new_AGEMA_signal_7289, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27}), .b ({new_AGEMA_signal_7454, new_AGEMA_signal_7453, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31}), .clk (clk), .r ({Fresh[932], Fresh[931], Fresh[930]}), .c ({new_AGEMA_signal_7652, new_AGEMA_signal_7651, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M35_U1 ( .a ({new_AGEMA_signal_7448, new_AGEMA_signal_7447, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24}), .b ({new_AGEMA_signal_7292, new_AGEMA_signal_7291, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34}), .clk (clk), .r ({Fresh[935], Fresh[934], Fresh[933]}), .c ({new_AGEMA_signal_7654, new_AGEMA_signal_7653, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M37_U1 ( .a ({new_AGEMA_signal_7130, new_AGEMA_signal_7129, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_7648, new_AGEMA_signal_7647, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29}), .c ({new_AGEMA_signal_7846, new_AGEMA_signal_7845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M38_U1 ( .a ({new_AGEMA_signal_7652, new_AGEMA_signal_7651, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32}), .b ({new_AGEMA_signal_7456, new_AGEMA_signal_7455, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33}), .c ({new_AGEMA_signal_7848, new_AGEMA_signal_7847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M39_U1 ( .a ({new_AGEMA_signal_7286, new_AGEMA_signal_7285, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}), .b ({new_AGEMA_signal_7650, new_AGEMA_signal_7649, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30}), .c ({new_AGEMA_signal_7850, new_AGEMA_signal_7849, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M40_U1 ( .a ({new_AGEMA_signal_7654, new_AGEMA_signal_7653, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35}), .b ({new_AGEMA_signal_7656, new_AGEMA_signal_7655, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36}), .c ({new_AGEMA_signal_7852, new_AGEMA_signal_7851, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M41_U1 ( .a ({new_AGEMA_signal_7848, new_AGEMA_signal_7847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_7852, new_AGEMA_signal_7851, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_8022, new_AGEMA_signal_8021, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M42_U1 ( .a ({new_AGEMA_signal_7846, new_AGEMA_signal_7845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_7850, new_AGEMA_signal_7849, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .c ({new_AGEMA_signal_8024, new_AGEMA_signal_8023, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M43_U1 ( .a ({new_AGEMA_signal_7846, new_AGEMA_signal_7845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_7848, new_AGEMA_signal_7847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .c ({new_AGEMA_signal_8026, new_AGEMA_signal_8025, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M44_U1 ( .a ({new_AGEMA_signal_7850, new_AGEMA_signal_7849, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_7852, new_AGEMA_signal_7851, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_8028, new_AGEMA_signal_8027, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M45_U1 ( .a ({new_AGEMA_signal_8024, new_AGEMA_signal_8023, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_8022, new_AGEMA_signal_8021, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}), .c ({new_AGEMA_signal_8502, new_AGEMA_signal_8501, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M29_U1 ( .a ({new_AGEMA_signal_7462, new_AGEMA_signal_7461, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28}), .b ({new_AGEMA_signal_7298, new_AGEMA_signal_7297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27}), .clk (clk), .r ({Fresh[938], Fresh[937], Fresh[936]}), .c ({new_AGEMA_signal_7658, new_AGEMA_signal_7657, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M30_U1 ( .a ({new_AGEMA_signal_7460, new_AGEMA_signal_7459, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26}), .b ({new_AGEMA_signal_7458, new_AGEMA_signal_7457, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24}), .clk (clk), .r ({Fresh[941], Fresh[940], Fresh[939]}), .c ({new_AGEMA_signal_7660, new_AGEMA_signal_7659, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M32_U1 ( .a ({new_AGEMA_signal_7298, new_AGEMA_signal_7297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27}), .b ({new_AGEMA_signal_7464, new_AGEMA_signal_7463, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31}), .clk (clk), .r ({Fresh[944], Fresh[943], Fresh[942]}), .c ({new_AGEMA_signal_7662, new_AGEMA_signal_7661, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M35_U1 ( .a ({new_AGEMA_signal_7458, new_AGEMA_signal_7457, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24}), .b ({new_AGEMA_signal_7300, new_AGEMA_signal_7299, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34}), .clk (clk), .r ({Fresh[947], Fresh[946], Fresh[945]}), .c ({new_AGEMA_signal_7664, new_AGEMA_signal_7663, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M37_U1 ( .a ({new_AGEMA_signal_7138, new_AGEMA_signal_7137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_7658, new_AGEMA_signal_7657, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29}), .c ({new_AGEMA_signal_7854, new_AGEMA_signal_7853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M38_U1 ( .a ({new_AGEMA_signal_7662, new_AGEMA_signal_7661, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32}), .b ({new_AGEMA_signal_7466, new_AGEMA_signal_7465, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33}), .c ({new_AGEMA_signal_7856, new_AGEMA_signal_7855, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M39_U1 ( .a ({new_AGEMA_signal_7294, new_AGEMA_signal_7293, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}), .b ({new_AGEMA_signal_7660, new_AGEMA_signal_7659, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30}), .c ({new_AGEMA_signal_7858, new_AGEMA_signal_7857, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M40_U1 ( .a ({new_AGEMA_signal_7664, new_AGEMA_signal_7663, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35}), .b ({new_AGEMA_signal_7666, new_AGEMA_signal_7665, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36}), .c ({new_AGEMA_signal_7860, new_AGEMA_signal_7859, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M41_U1 ( .a ({new_AGEMA_signal_7856, new_AGEMA_signal_7855, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_7860, new_AGEMA_signal_7859, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_8046, new_AGEMA_signal_8045, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M42_U1 ( .a ({new_AGEMA_signal_7854, new_AGEMA_signal_7853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_7858, new_AGEMA_signal_7857, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .c ({new_AGEMA_signal_8048, new_AGEMA_signal_8047, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M43_U1 ( .a ({new_AGEMA_signal_7854, new_AGEMA_signal_7853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_7856, new_AGEMA_signal_7855, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .c ({new_AGEMA_signal_8050, new_AGEMA_signal_8049, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M44_U1 ( .a ({new_AGEMA_signal_7858, new_AGEMA_signal_7857, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_7860, new_AGEMA_signal_7859, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_8052, new_AGEMA_signal_8051, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M45_U1 ( .a ({new_AGEMA_signal_8048, new_AGEMA_signal_8047, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_8046, new_AGEMA_signal_8045, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}), .c ({new_AGEMA_signal_8526, new_AGEMA_signal_8525, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M29_U1 ( .a ({new_AGEMA_signal_7472, new_AGEMA_signal_7471, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28}), .b ({new_AGEMA_signal_7306, new_AGEMA_signal_7305, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27}), .clk (clk), .r ({Fresh[950], Fresh[949], Fresh[948]}), .c ({new_AGEMA_signal_7668, new_AGEMA_signal_7667, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M30_U1 ( .a ({new_AGEMA_signal_7470, new_AGEMA_signal_7469, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26}), .b ({new_AGEMA_signal_7468, new_AGEMA_signal_7467, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24}), .clk (clk), .r ({Fresh[953], Fresh[952], Fresh[951]}), .c ({new_AGEMA_signal_7670, new_AGEMA_signal_7669, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M32_U1 ( .a ({new_AGEMA_signal_7306, new_AGEMA_signal_7305, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27}), .b ({new_AGEMA_signal_7474, new_AGEMA_signal_7473, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31}), .clk (clk), .r ({Fresh[956], Fresh[955], Fresh[954]}), .c ({new_AGEMA_signal_7672, new_AGEMA_signal_7671, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M35_U1 ( .a ({new_AGEMA_signal_7468, new_AGEMA_signal_7467, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24}), .b ({new_AGEMA_signal_7308, new_AGEMA_signal_7307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957]}), .c ({new_AGEMA_signal_7674, new_AGEMA_signal_7673, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M37_U1 ( .a ({new_AGEMA_signal_7146, new_AGEMA_signal_7145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_7668, new_AGEMA_signal_7667, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29}), .c ({new_AGEMA_signal_7862, new_AGEMA_signal_7861, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M38_U1 ( .a ({new_AGEMA_signal_7672, new_AGEMA_signal_7671, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32}), .b ({new_AGEMA_signal_7476, new_AGEMA_signal_7475, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33}), .c ({new_AGEMA_signal_7864, new_AGEMA_signal_7863, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M39_U1 ( .a ({new_AGEMA_signal_7302, new_AGEMA_signal_7301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}), .b ({new_AGEMA_signal_7670, new_AGEMA_signal_7669, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30}), .c ({new_AGEMA_signal_7866, new_AGEMA_signal_7865, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M40_U1 ( .a ({new_AGEMA_signal_7674, new_AGEMA_signal_7673, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35}), .b ({new_AGEMA_signal_7676, new_AGEMA_signal_7675, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36}), .c ({new_AGEMA_signal_7868, new_AGEMA_signal_7867, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M41_U1 ( .a ({new_AGEMA_signal_7864, new_AGEMA_signal_7863, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_7868, new_AGEMA_signal_7867, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_8070, new_AGEMA_signal_8069, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M42_U1 ( .a ({new_AGEMA_signal_7862, new_AGEMA_signal_7861, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_7866, new_AGEMA_signal_7865, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .c ({new_AGEMA_signal_8072, new_AGEMA_signal_8071, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M43_U1 ( .a ({new_AGEMA_signal_7862, new_AGEMA_signal_7861, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_7864, new_AGEMA_signal_7863, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .c ({new_AGEMA_signal_8074, new_AGEMA_signal_8073, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M44_U1 ( .a ({new_AGEMA_signal_7866, new_AGEMA_signal_7865, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_7868, new_AGEMA_signal_7867, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_8076, new_AGEMA_signal_8075, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M45_U1 ( .a ({new_AGEMA_signal_8072, new_AGEMA_signal_8071, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_8070, new_AGEMA_signal_8069, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}), .c ({new_AGEMA_signal_8550, new_AGEMA_signal_8549, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_masked #(.security_order(2), .pipeline(0)) U858 ( .s (n321), .b ({new_AGEMA_signal_9914, new_AGEMA_signal_9913, MixColumnsInput[0]}), .a ({new_AGEMA_signal_11644, new_AGEMA_signal_11643, MixColumnsOutput[0]}), .c ({new_AGEMA_signal_11832, new_AGEMA_signal_11831, RoundOutput[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U859 ( .s (n321), .b ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .a ({new_AGEMA_signal_11994, new_AGEMA_signal_11993, MixColumnsOutput[100]}), .c ({new_AGEMA_signal_12218, new_AGEMA_signal_12217, RoundOutput[100]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U860 ( .s (n321), .b ({new_AGEMA_signal_10226, new_AGEMA_signal_10225, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, MixColumnsOutput[101]}), .c ({new_AGEMA_signal_11834, new_AGEMA_signal_11833, RoundOutput[101]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U861 ( .s (n321), .b ({new_AGEMA_signal_10224, new_AGEMA_signal_10223, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .a ({new_AGEMA_signal_11396, new_AGEMA_signal_11395, MixColumnsOutput[102]}), .c ({new_AGEMA_signal_11836, new_AGEMA_signal_11835, RoundOutput[102]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U862 ( .s (n321), .b ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .a ({new_AGEMA_signal_11394, new_AGEMA_signal_11393, MixColumnsOutput[103]}), .c ({new_AGEMA_signal_11838, new_AGEMA_signal_11837, RoundOutput[103]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U863 ( .s (n321), .b ({new_AGEMA_signal_9936, new_AGEMA_signal_9935, MixColumnsInput[104]}), .a ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, MixColumnsOutput[104]}), .c ({new_AGEMA_signal_11840, new_AGEMA_signal_11839, RoundOutput[104]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U864 ( .s (n321), .b ({new_AGEMA_signal_10304, new_AGEMA_signal_10303, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .a ({new_AGEMA_signal_11992, new_AGEMA_signal_11991, MixColumnsOutput[105]}), .c ({new_AGEMA_signal_12220, new_AGEMA_signal_12219, RoundOutput[105]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U865 ( .s (n321), .b ({new_AGEMA_signal_10302, new_AGEMA_signal_10301, MixColumnsInput[106]}), .a ({new_AGEMA_signal_11450, new_AGEMA_signal_11449, MixColumnsOutput[106]}), .c ({new_AGEMA_signal_11842, new_AGEMA_signal_11841, RoundOutput[106]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U866 ( .s (n315), .b ({new_AGEMA_signal_10300, new_AGEMA_signal_10299, MixColumnsInput[107]}), .a ({new_AGEMA_signal_12014, new_AGEMA_signal_12013, MixColumnsOutput[107]}), .c ({new_AGEMA_signal_12222, new_AGEMA_signal_12221, RoundOutput[107]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U867 ( .s (n316), .b ({new_AGEMA_signal_10298, new_AGEMA_signal_10297, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .a ({new_AGEMA_signal_12012, new_AGEMA_signal_12011, MixColumnsOutput[108]}), .c ({new_AGEMA_signal_12224, new_AGEMA_signal_12223, RoundOutput[108]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U868 ( .s (n317), .b ({new_AGEMA_signal_10296, new_AGEMA_signal_10295, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .a ({new_AGEMA_signal_11444, new_AGEMA_signal_11443, MixColumnsOutput[109]}), .c ({new_AGEMA_signal_11844, new_AGEMA_signal_11843, RoundOutput[109]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U869 ( .s (n318), .b ({new_AGEMA_signal_10358, new_AGEMA_signal_10357, MixColumnsInput[10]}), .a ({new_AGEMA_signal_11642, new_AGEMA_signal_11641, MixColumnsOutput[10]}), .c ({new_AGEMA_signal_11846, new_AGEMA_signal_11845, RoundOutput[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U870 ( .s (n319), .b ({new_AGEMA_signal_10294, new_AGEMA_signal_10293, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .a ({new_AGEMA_signal_11442, new_AGEMA_signal_11441, MixColumnsOutput[110]}), .c ({new_AGEMA_signal_11848, new_AGEMA_signal_11847, RoundOutput[110]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U871 ( .s (n320), .b ({new_AGEMA_signal_10292, new_AGEMA_signal_10291, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .a ({new_AGEMA_signal_11440, new_AGEMA_signal_11439, MixColumnsOutput[111]}), .c ({new_AGEMA_signal_11850, new_AGEMA_signal_11849, RoundOutput[111]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U872 ( .s (n319), .b ({new_AGEMA_signal_10046, new_AGEMA_signal_10045, MixColumnsInput[112]}), .a ({new_AGEMA_signal_11438, new_AGEMA_signal_11437, MixColumnsOutput[112]}), .c ({new_AGEMA_signal_11852, new_AGEMA_signal_11851, RoundOutput[112]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U873 ( .s (n318), .b ({new_AGEMA_signal_10374, new_AGEMA_signal_10373, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .a ({new_AGEMA_signal_12010, new_AGEMA_signal_12009, MixColumnsOutput[113]}), .c ({new_AGEMA_signal_12226, new_AGEMA_signal_12225, RoundOutput[113]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U874 ( .s (n318), .b ({new_AGEMA_signal_10372, new_AGEMA_signal_10371, MixColumnsInput[114]}), .a ({new_AGEMA_signal_11434, new_AGEMA_signal_11433, MixColumnsOutput[114]}), .c ({new_AGEMA_signal_11854, new_AGEMA_signal_11853, RoundOutput[114]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U875 ( .s (n315), .b ({new_AGEMA_signal_10370, new_AGEMA_signal_10369, MixColumnsInput[115]}), .a ({new_AGEMA_signal_12008, new_AGEMA_signal_12007, MixColumnsOutput[115]}), .c ({new_AGEMA_signal_12228, new_AGEMA_signal_12227, RoundOutput[115]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U876 ( .s (n316), .b ({new_AGEMA_signal_10368, new_AGEMA_signal_10367, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .a ({new_AGEMA_signal_12004, new_AGEMA_signal_12003, MixColumnsOutput[116]}), .c ({new_AGEMA_signal_12230, new_AGEMA_signal_12229, RoundOutput[116]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U877 ( .s (n317), .b ({new_AGEMA_signal_10366, new_AGEMA_signal_10365, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .a ({new_AGEMA_signal_11426, new_AGEMA_signal_11425, MixColumnsOutput[117]}), .c ({new_AGEMA_signal_11856, new_AGEMA_signal_11855, RoundOutput[117]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U878 ( .s (n319), .b ({new_AGEMA_signal_10364, new_AGEMA_signal_10363, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .a ({new_AGEMA_signal_11424, new_AGEMA_signal_11423, MixColumnsOutput[118]}), .c ({new_AGEMA_signal_11858, new_AGEMA_signal_11857, RoundOutput[118]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U879 ( .s (n320), .b ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .a ({new_AGEMA_signal_11422, new_AGEMA_signal_11421, MixColumnsOutput[119]}), .c ({new_AGEMA_signal_11860, new_AGEMA_signal_11859, RoundOutput[119]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U880 ( .s (n320), .b ({new_AGEMA_signal_10356, new_AGEMA_signal_10355, MixColumnsInput[11]}), .a ({new_AGEMA_signal_12086, new_AGEMA_signal_12085, MixColumnsOutput[11]}), .c ({new_AGEMA_signal_12232, new_AGEMA_signal_12231, RoundOutput[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U881 ( .s (n319), .b ({new_AGEMA_signal_10156, new_AGEMA_signal_10155, MixColumnsInput[120]}), .a ({new_AGEMA_signal_11420, new_AGEMA_signal_11419, MixColumnsOutput[120]}), .c ({new_AGEMA_signal_11862, new_AGEMA_signal_11861, RoundOutput[120]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U882 ( .s (n318), .b ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .a ({new_AGEMA_signal_12002, new_AGEMA_signal_12001, MixColumnsOutput[121]}), .c ({new_AGEMA_signal_12234, new_AGEMA_signal_12233, RoundOutput[121]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U883 ( .s (n319), .b ({new_AGEMA_signal_10442, new_AGEMA_signal_10441, MixColumnsInput[122]}), .a ({new_AGEMA_signal_11416, new_AGEMA_signal_11415, MixColumnsOutput[122]}), .c ({new_AGEMA_signal_11864, new_AGEMA_signal_11863, RoundOutput[122]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U884 ( .s (n320), .b ({new_AGEMA_signal_10440, new_AGEMA_signal_10439, MixColumnsInput[123]}), .a ({new_AGEMA_signal_12000, new_AGEMA_signal_11999, MixColumnsOutput[123]}), .c ({new_AGEMA_signal_12236, new_AGEMA_signal_12235, RoundOutput[123]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U885 ( .s (n316), .b ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .a ({new_AGEMA_signal_11998, new_AGEMA_signal_11997, MixColumnsOutput[124]}), .c ({new_AGEMA_signal_12238, new_AGEMA_signal_12237, RoundOutput[124]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U886 ( .s (n320), .b ({new_AGEMA_signal_10436, new_AGEMA_signal_10435, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .a ({new_AGEMA_signal_11410, new_AGEMA_signal_11409, MixColumnsOutput[125]}), .c ({new_AGEMA_signal_11866, new_AGEMA_signal_11865, RoundOutput[125]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U887 ( .s (n316), .b ({new_AGEMA_signal_10434, new_AGEMA_signal_10433, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .a ({new_AGEMA_signal_11406, new_AGEMA_signal_11405, MixColumnsOutput[126]}), .c ({new_AGEMA_signal_11868, new_AGEMA_signal_11867, RoundOutput[126]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U888 ( .s (n317), .b ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .a ({new_AGEMA_signal_11404, new_AGEMA_signal_11403, MixColumnsOutput[127]}), .c ({new_AGEMA_signal_11870, new_AGEMA_signal_11869, RoundOutput[127]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U889 ( .s (n315), .b ({new_AGEMA_signal_10354, new_AGEMA_signal_10353, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .a ({new_AGEMA_signal_12084, new_AGEMA_signal_12083, MixColumnsOutput[12]}), .c ({new_AGEMA_signal_12240, new_AGEMA_signal_12239, RoundOutput[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U890 ( .s (n317), .b ({new_AGEMA_signal_10352, new_AGEMA_signal_10351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .a ({new_AGEMA_signal_11636, new_AGEMA_signal_11635, MixColumnsOutput[13]}), .c ({new_AGEMA_signal_11872, new_AGEMA_signal_11871, RoundOutput[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U891 ( .s (n316), .b ({new_AGEMA_signal_10350, new_AGEMA_signal_10349, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .a ({new_AGEMA_signal_11634, new_AGEMA_signal_11633, MixColumnsOutput[14]}), .c ({new_AGEMA_signal_11874, new_AGEMA_signal_11873, RoundOutput[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U892 ( .s (n317), .b ({new_AGEMA_signal_10348, new_AGEMA_signal_10347, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .a ({new_AGEMA_signal_11632, new_AGEMA_signal_11631, MixColumnsOutput[15]}), .c ({new_AGEMA_signal_11876, new_AGEMA_signal_11875, RoundOutput[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U893 ( .s (n315), .b ({new_AGEMA_signal_10134, new_AGEMA_signal_10133, MixColumnsInput[16]}), .a ({new_AGEMA_signal_11630, new_AGEMA_signal_11629, MixColumnsOutput[16]}), .c ({new_AGEMA_signal_11878, new_AGEMA_signal_11877, RoundOutput[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U894 ( .s (n318), .b ({new_AGEMA_signal_10430, new_AGEMA_signal_10429, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .a ({new_AGEMA_signal_12082, new_AGEMA_signal_12081, MixColumnsOutput[17]}), .c ({new_AGEMA_signal_12242, new_AGEMA_signal_12241, RoundOutput[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U895 ( .s (n319), .b ({new_AGEMA_signal_10428, new_AGEMA_signal_10427, MixColumnsInput[18]}), .a ({new_AGEMA_signal_11626, new_AGEMA_signal_11625, MixColumnsOutput[18]}), .c ({new_AGEMA_signal_11880, new_AGEMA_signal_11879, RoundOutput[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U896 ( .s (n320), .b ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, MixColumnsInput[19]}), .a ({new_AGEMA_signal_12080, new_AGEMA_signal_12079, MixColumnsOutput[19]}), .c ({new_AGEMA_signal_12244, new_AGEMA_signal_12243, RoundOutput[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U897 ( .s (n318), .b ({new_AGEMA_signal_10290, new_AGEMA_signal_10289, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .a ({new_AGEMA_signal_12078, new_AGEMA_signal_12077, MixColumnsOutput[1]}), .c ({new_AGEMA_signal_12246, new_AGEMA_signal_12245, RoundOutput[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U898 ( .s (n319), .b ({new_AGEMA_signal_10424, new_AGEMA_signal_10423, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .a ({new_AGEMA_signal_12076, new_AGEMA_signal_12075, MixColumnsOutput[20]}), .c ({new_AGEMA_signal_12248, new_AGEMA_signal_12247, RoundOutput[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U899 ( .s (n316), .b ({new_AGEMA_signal_10422, new_AGEMA_signal_10421, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .a ({new_AGEMA_signal_11618, new_AGEMA_signal_11617, MixColumnsOutput[21]}), .c ({new_AGEMA_signal_11882, new_AGEMA_signal_11881, RoundOutput[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U900 ( .s (n317), .b ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .a ({new_AGEMA_signal_11616, new_AGEMA_signal_11615, MixColumnsOutput[22]}), .c ({new_AGEMA_signal_11884, new_AGEMA_signal_11883, RoundOutput[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U901 ( .s (n315), .b ({new_AGEMA_signal_10418, new_AGEMA_signal_10417, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .a ({new_AGEMA_signal_11614, new_AGEMA_signal_11613, MixColumnsOutput[23]}), .c ({new_AGEMA_signal_11886, new_AGEMA_signal_11885, RoundOutput[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U902 ( .s (n320), .b ({new_AGEMA_signal_9892, new_AGEMA_signal_9891, MixColumnsInput[24]}), .a ({new_AGEMA_signal_11612, new_AGEMA_signal_11611, MixColumnsOutput[24]}), .c ({new_AGEMA_signal_11888, new_AGEMA_signal_11887, RoundOutput[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U903 ( .s (n318), .b ({new_AGEMA_signal_10276, new_AGEMA_signal_10275, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .a ({new_AGEMA_signal_12074, new_AGEMA_signal_12073, MixColumnsOutput[25]}), .c ({new_AGEMA_signal_12250, new_AGEMA_signal_12249, RoundOutput[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U904 ( .s (n316), .b ({new_AGEMA_signal_10274, new_AGEMA_signal_10273, MixColumnsInput[26]}), .a ({new_AGEMA_signal_11608, new_AGEMA_signal_11607, MixColumnsOutput[26]}), .c ({new_AGEMA_signal_11890, new_AGEMA_signal_11889, RoundOutput[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U905 ( .s (n317), .b ({new_AGEMA_signal_10272, new_AGEMA_signal_10271, MixColumnsInput[27]}), .a ({new_AGEMA_signal_12072, new_AGEMA_signal_12071, MixColumnsOutput[27]}), .c ({new_AGEMA_signal_12252, new_AGEMA_signal_12251, RoundOutput[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U906 ( .s (n315), .b ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .a ({new_AGEMA_signal_12070, new_AGEMA_signal_12069, MixColumnsOutput[28]}), .c ({new_AGEMA_signal_12254, new_AGEMA_signal_12253, RoundOutput[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U907 ( .s (n319), .b ({new_AGEMA_signal_10268, new_AGEMA_signal_10267, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .a ({new_AGEMA_signal_11602, new_AGEMA_signal_11601, MixColumnsOutput[29]}), .c ({new_AGEMA_signal_11892, new_AGEMA_signal_11891, RoundOutput[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U908 ( .s (n315), .b ({new_AGEMA_signal_10288, new_AGEMA_signal_10287, MixColumnsInput[2]}), .a ({new_AGEMA_signal_11600, new_AGEMA_signal_11599, MixColumnsOutput[2]}), .c ({new_AGEMA_signal_11894, new_AGEMA_signal_11893, RoundOutput[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U909 ( .s (n320), .b ({new_AGEMA_signal_10266, new_AGEMA_signal_10265, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .a ({new_AGEMA_signal_11598, new_AGEMA_signal_11597, MixColumnsOutput[30]}), .c ({new_AGEMA_signal_11896, new_AGEMA_signal_11895, RoundOutput[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U910 ( .s (n318), .b ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .a ({new_AGEMA_signal_11596, new_AGEMA_signal_11595, MixColumnsOutput[31]}), .c ({new_AGEMA_signal_11898, new_AGEMA_signal_11897, RoundOutput[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U911 ( .s (n316), .b ({new_AGEMA_signal_10002, new_AGEMA_signal_10001, MixColumnsInput[32]}), .a ({new_AGEMA_signal_11580, new_AGEMA_signal_11579, MixColumnsOutput[32]}), .c ({new_AGEMA_signal_11900, new_AGEMA_signal_11899, RoundOutput[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U912 ( .s (n317), .b ({new_AGEMA_signal_10346, new_AGEMA_signal_10345, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .a ({new_AGEMA_signal_12054, new_AGEMA_signal_12053, MixColumnsOutput[33]}), .c ({new_AGEMA_signal_12256, new_AGEMA_signal_12255, RoundOutput[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U913 ( .s (n315), .b ({new_AGEMA_signal_10344, new_AGEMA_signal_10343, MixColumnsInput[34]}), .a ({new_AGEMA_signal_11536, new_AGEMA_signal_11535, MixColumnsOutput[34]}), .c ({new_AGEMA_signal_11902, new_AGEMA_signal_11901, RoundOutput[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U914 ( .s (n320), .b ({new_AGEMA_signal_10342, new_AGEMA_signal_10341, MixColumnsInput[35]}), .a ({new_AGEMA_signal_12044, new_AGEMA_signal_12043, MixColumnsOutput[35]}), .c ({new_AGEMA_signal_12258, new_AGEMA_signal_12257, RoundOutput[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U915 ( .s (n320), .b ({new_AGEMA_signal_10340, new_AGEMA_signal_10339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .a ({new_AGEMA_signal_12042, new_AGEMA_signal_12041, MixColumnsOutput[36]}), .c ({new_AGEMA_signal_12260, new_AGEMA_signal_12259, RoundOutput[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U916 ( .s (n320), .b ({new_AGEMA_signal_10338, new_AGEMA_signal_10337, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .a ({new_AGEMA_signal_11526, new_AGEMA_signal_11525, MixColumnsOutput[37]}), .c ({new_AGEMA_signal_11904, new_AGEMA_signal_11903, RoundOutput[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U917 ( .s (n320), .b ({new_AGEMA_signal_10336, new_AGEMA_signal_10335, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .a ({new_AGEMA_signal_11524, new_AGEMA_signal_11523, MixColumnsOutput[38]}), .c ({new_AGEMA_signal_11906, new_AGEMA_signal_11905, RoundOutput[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U918 ( .s (n320), .b ({new_AGEMA_signal_10334, new_AGEMA_signal_10333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .a ({new_AGEMA_signal_11522, new_AGEMA_signal_11521, MixColumnsOutput[39]}), .c ({new_AGEMA_signal_11908, new_AGEMA_signal_11907, RoundOutput[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U919 ( .s (n320), .b ({new_AGEMA_signal_10286, new_AGEMA_signal_10285, MixColumnsInput[3]}), .a ({new_AGEMA_signal_12068, new_AGEMA_signal_12067, MixColumnsOutput[3]}), .c ({new_AGEMA_signal_12262, new_AGEMA_signal_12261, RoundOutput[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U920 ( .s (n320), .b ({new_AGEMA_signal_10112, new_AGEMA_signal_10111, MixColumnsInput[40]}), .a ({new_AGEMA_signal_11520, new_AGEMA_signal_11519, MixColumnsOutput[40]}), .c ({new_AGEMA_signal_11910, new_AGEMA_signal_11909, RoundOutput[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U921 ( .s (n320), .b ({new_AGEMA_signal_10416, new_AGEMA_signal_10415, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .a ({new_AGEMA_signal_12040, new_AGEMA_signal_12039, MixColumnsOutput[41]}), .c ({new_AGEMA_signal_12264, new_AGEMA_signal_12263, RoundOutput[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U922 ( .s (n320), .b ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, MixColumnsInput[42]}), .a ({new_AGEMA_signal_11578, new_AGEMA_signal_11577, MixColumnsOutput[42]}), .c ({new_AGEMA_signal_11912, new_AGEMA_signal_11911, RoundOutput[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U923 ( .s (n320), .b ({new_AGEMA_signal_10412, new_AGEMA_signal_10411, MixColumnsInput[43]}), .a ({new_AGEMA_signal_12062, new_AGEMA_signal_12061, MixColumnsOutput[43]}), .c ({new_AGEMA_signal_12266, new_AGEMA_signal_12265, RoundOutput[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U924 ( .s (n320), .b ({new_AGEMA_signal_10410, new_AGEMA_signal_10409, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .a ({new_AGEMA_signal_12060, new_AGEMA_signal_12059, MixColumnsOutput[44]}), .c ({new_AGEMA_signal_12268, new_AGEMA_signal_12267, RoundOutput[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U925 ( .s (n320), .b ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .a ({new_AGEMA_signal_11572, new_AGEMA_signal_11571, MixColumnsOutput[45]}), .c ({new_AGEMA_signal_11914, new_AGEMA_signal_11913, RoundOutput[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U926 ( .s (n319), .b ({new_AGEMA_signal_10406, new_AGEMA_signal_10405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .a ({new_AGEMA_signal_11570, new_AGEMA_signal_11569, MixColumnsOutput[46]}), .c ({new_AGEMA_signal_11916, new_AGEMA_signal_11915, RoundOutput[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U927 ( .s (n319), .b ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .a ({new_AGEMA_signal_11568, new_AGEMA_signal_11567, MixColumnsOutput[47]}), .c ({new_AGEMA_signal_11918, new_AGEMA_signal_11917, RoundOutput[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U928 ( .s (n319), .b ({new_AGEMA_signal_9870, new_AGEMA_signal_9869, MixColumnsInput[48]}), .a ({new_AGEMA_signal_11566, new_AGEMA_signal_11565, MixColumnsOutput[48]}), .c ({new_AGEMA_signal_11920, new_AGEMA_signal_11919, RoundOutput[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U929 ( .s (n319), .b ({new_AGEMA_signal_10262, new_AGEMA_signal_10261, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .a ({new_AGEMA_signal_12058, new_AGEMA_signal_12057, MixColumnsOutput[49]}), .c ({new_AGEMA_signal_12270, new_AGEMA_signal_12269, RoundOutput[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U930 ( .s (n319), .b ({new_AGEMA_signal_10284, new_AGEMA_signal_10283, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .a ({new_AGEMA_signal_12066, new_AGEMA_signal_12065, MixColumnsOutput[4]}), .c ({new_AGEMA_signal_12272, new_AGEMA_signal_12271, RoundOutput[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U931 ( .s (n319), .b ({new_AGEMA_signal_10260, new_AGEMA_signal_10259, MixColumnsInput[50]}), .a ({new_AGEMA_signal_11562, new_AGEMA_signal_11561, MixColumnsOutput[50]}), .c ({new_AGEMA_signal_11922, new_AGEMA_signal_11921, RoundOutput[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U932 ( .s (n319), .b ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, MixColumnsInput[51]}), .a ({new_AGEMA_signal_12056, new_AGEMA_signal_12055, MixColumnsOutput[51]}), .c ({new_AGEMA_signal_12274, new_AGEMA_signal_12273, RoundOutput[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U933 ( .s (n319), .b ({new_AGEMA_signal_10256, new_AGEMA_signal_10255, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .a ({new_AGEMA_signal_12052, new_AGEMA_signal_12051, MixColumnsOutput[52]}), .c ({new_AGEMA_signal_12276, new_AGEMA_signal_12275, RoundOutput[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U934 ( .s (n319), .b ({new_AGEMA_signal_10254, new_AGEMA_signal_10253, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .a ({new_AGEMA_signal_11554, new_AGEMA_signal_11553, MixColumnsOutput[53]}), .c ({new_AGEMA_signal_11924, new_AGEMA_signal_11923, RoundOutput[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U935 ( .s (n319), .b ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .a ({new_AGEMA_signal_11552, new_AGEMA_signal_11551, MixColumnsOutput[54]}), .c ({new_AGEMA_signal_11926, new_AGEMA_signal_11925, RoundOutput[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U936 ( .s (n319), .b ({new_AGEMA_signal_10250, new_AGEMA_signal_10249, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .a ({new_AGEMA_signal_11550, new_AGEMA_signal_11549, MixColumnsOutput[55]}), .c ({new_AGEMA_signal_11928, new_AGEMA_signal_11927, RoundOutput[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U937 ( .s (n319), .b ({new_AGEMA_signal_9980, new_AGEMA_signal_9979, MixColumnsInput[56]}), .a ({new_AGEMA_signal_11548, new_AGEMA_signal_11547, MixColumnsOutput[56]}), .c ({new_AGEMA_signal_11930, new_AGEMA_signal_11929, RoundOutput[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U938 ( .s (n318), .b ({new_AGEMA_signal_10332, new_AGEMA_signal_10331, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .a ({new_AGEMA_signal_12050, new_AGEMA_signal_12049, MixColumnsOutput[57]}), .c ({new_AGEMA_signal_12278, new_AGEMA_signal_12277, RoundOutput[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U939 ( .s (n318), .b ({new_AGEMA_signal_10330, new_AGEMA_signal_10329, MixColumnsInput[58]}), .a ({new_AGEMA_signal_11544, new_AGEMA_signal_11543, MixColumnsOutput[58]}), .c ({new_AGEMA_signal_11932, new_AGEMA_signal_11931, RoundOutput[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U940 ( .s (n318), .b ({new_AGEMA_signal_10328, new_AGEMA_signal_10327, MixColumnsInput[59]}), .a ({new_AGEMA_signal_12048, new_AGEMA_signal_12047, MixColumnsOutput[59]}), .c ({new_AGEMA_signal_12280, new_AGEMA_signal_12279, RoundOutput[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U941 ( .s (n318), .b ({new_AGEMA_signal_10282, new_AGEMA_signal_10281, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .a ({new_AGEMA_signal_11590, new_AGEMA_signal_11589, MixColumnsOutput[5]}), .c ({new_AGEMA_signal_11934, new_AGEMA_signal_11933, RoundOutput[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U942 ( .s (n318), .b ({new_AGEMA_signal_10326, new_AGEMA_signal_10325, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .a ({new_AGEMA_signal_12046, new_AGEMA_signal_12045, MixColumnsOutput[60]}), .c ({new_AGEMA_signal_12282, new_AGEMA_signal_12281, RoundOutput[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U943 ( .s (n318), .b ({new_AGEMA_signal_10324, new_AGEMA_signal_10323, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .a ({new_AGEMA_signal_11538, new_AGEMA_signal_11537, MixColumnsOutput[61]}), .c ({new_AGEMA_signal_11936, new_AGEMA_signal_11935, RoundOutput[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U944 ( .s (n318), .b ({new_AGEMA_signal_10322, new_AGEMA_signal_10321, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .a ({new_AGEMA_signal_11534, new_AGEMA_signal_11533, MixColumnsOutput[62]}), .c ({new_AGEMA_signal_11938, new_AGEMA_signal_11937, RoundOutput[62]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U945 ( .s (n318), .b ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .a ({new_AGEMA_signal_11532, new_AGEMA_signal_11531, MixColumnsOutput[63]}), .c ({new_AGEMA_signal_11940, new_AGEMA_signal_11939, RoundOutput[63]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U946 ( .s (n318), .b ({new_AGEMA_signal_10090, new_AGEMA_signal_10089, MixColumnsInput[64]}), .a ({new_AGEMA_signal_11516, new_AGEMA_signal_11515, MixColumnsOutput[64]}), .c ({new_AGEMA_signal_11942, new_AGEMA_signal_11941, RoundOutput[64]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U947 ( .s (n318), .b ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .a ({new_AGEMA_signal_12030, new_AGEMA_signal_12029, MixColumnsOutput[65]}), .c ({new_AGEMA_signal_12284, new_AGEMA_signal_12283, RoundOutput[65]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U948 ( .s (n318), .b ({new_AGEMA_signal_10400, new_AGEMA_signal_10399, MixColumnsInput[66]}), .a ({new_AGEMA_signal_11472, new_AGEMA_signal_11471, MixColumnsOutput[66]}), .c ({new_AGEMA_signal_11944, new_AGEMA_signal_11943, RoundOutput[66]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U949 ( .s (n318), .b ({new_AGEMA_signal_10398, new_AGEMA_signal_10397, MixColumnsInput[67]}), .a ({new_AGEMA_signal_12020, new_AGEMA_signal_12019, MixColumnsOutput[67]}), .c ({new_AGEMA_signal_12286, new_AGEMA_signal_12285, RoundOutput[67]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U950 ( .s (n317), .b ({new_AGEMA_signal_10396, new_AGEMA_signal_10395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .a ({new_AGEMA_signal_12018, new_AGEMA_signal_12017, MixColumnsOutput[68]}), .c ({new_AGEMA_signal_12288, new_AGEMA_signal_12287, RoundOutput[68]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U951 ( .s (n317), .b ({new_AGEMA_signal_10394, new_AGEMA_signal_10393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .a ({new_AGEMA_signal_11462, new_AGEMA_signal_11461, MixColumnsOutput[69]}), .c ({new_AGEMA_signal_11946, new_AGEMA_signal_11945, RoundOutput[69]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U952 ( .s (n317), .b ({new_AGEMA_signal_10280, new_AGEMA_signal_10279, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .a ({new_AGEMA_signal_11588, new_AGEMA_signal_11587, MixColumnsOutput[6]}), .c ({new_AGEMA_signal_11948, new_AGEMA_signal_11947, RoundOutput[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U953 ( .s (n317), .b ({new_AGEMA_signal_10392, new_AGEMA_signal_10391, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .a ({new_AGEMA_signal_11460, new_AGEMA_signal_11459, MixColumnsOutput[70]}), .c ({new_AGEMA_signal_11950, new_AGEMA_signal_11949, RoundOutput[70]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U954 ( .s (n317), .b ({new_AGEMA_signal_10390, new_AGEMA_signal_10389, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .a ({new_AGEMA_signal_11458, new_AGEMA_signal_11457, MixColumnsOutput[71]}), .c ({new_AGEMA_signal_11952, new_AGEMA_signal_11951, RoundOutput[71]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U955 ( .s (n317), .b ({new_AGEMA_signal_9848, new_AGEMA_signal_9847, MixColumnsInput[72]}), .a ({new_AGEMA_signal_11456, new_AGEMA_signal_11455, MixColumnsOutput[72]}), .c ({new_AGEMA_signal_11954, new_AGEMA_signal_11953, RoundOutput[72]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U956 ( .s (n317), .b ({new_AGEMA_signal_10248, new_AGEMA_signal_10247, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .a ({new_AGEMA_signal_12016, new_AGEMA_signal_12015, MixColumnsOutput[73]}), .c ({new_AGEMA_signal_12290, new_AGEMA_signal_12289, RoundOutput[73]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U957 ( .s (n317), .b ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, MixColumnsInput[74]}), .a ({new_AGEMA_signal_11514, new_AGEMA_signal_11513, MixColumnsOutput[74]}), .c ({new_AGEMA_signal_11956, new_AGEMA_signal_11955, RoundOutput[74]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U958 ( .s (n317), .b ({new_AGEMA_signal_10244, new_AGEMA_signal_10243, MixColumnsInput[75]}), .a ({new_AGEMA_signal_12038, new_AGEMA_signal_12037, MixColumnsOutput[75]}), .c ({new_AGEMA_signal_12292, new_AGEMA_signal_12291, RoundOutput[75]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U959 ( .s (n317), .b ({new_AGEMA_signal_10242, new_AGEMA_signal_10241, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .a ({new_AGEMA_signal_12036, new_AGEMA_signal_12035, MixColumnsOutput[76]}), .c ({new_AGEMA_signal_12294, new_AGEMA_signal_12293, RoundOutput[76]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U960 ( .s (n317), .b ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .a ({new_AGEMA_signal_11508, new_AGEMA_signal_11507, MixColumnsOutput[77]}), .c ({new_AGEMA_signal_11958, new_AGEMA_signal_11957, RoundOutput[77]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U961 ( .s (n317), .b ({new_AGEMA_signal_10238, new_AGEMA_signal_10237, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .a ({new_AGEMA_signal_11506, new_AGEMA_signal_11505, MixColumnsOutput[78]}), .c ({new_AGEMA_signal_11960, new_AGEMA_signal_11959, RoundOutput[78]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U962 ( .s (n316), .b ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .a ({new_AGEMA_signal_11504, new_AGEMA_signal_11503, MixColumnsOutput[79]}), .c ({new_AGEMA_signal_11962, new_AGEMA_signal_11961, RoundOutput[79]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U963 ( .s (n316), .b ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .a ({new_AGEMA_signal_11586, new_AGEMA_signal_11585, MixColumnsOutput[7]}), .c ({new_AGEMA_signal_11964, new_AGEMA_signal_11963, RoundOutput[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U964 ( .s (n316), .b ({new_AGEMA_signal_9958, new_AGEMA_signal_9957, MixColumnsInput[80]}), .a ({new_AGEMA_signal_11502, new_AGEMA_signal_11501, MixColumnsOutput[80]}), .c ({new_AGEMA_signal_11966, new_AGEMA_signal_11965, RoundOutput[80]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U965 ( .s (n316), .b ({new_AGEMA_signal_10318, new_AGEMA_signal_10317, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .a ({new_AGEMA_signal_12034, new_AGEMA_signal_12033, MixColumnsOutput[81]}), .c ({new_AGEMA_signal_12296, new_AGEMA_signal_12295, RoundOutput[81]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U966 ( .s (n316), .b ({new_AGEMA_signal_10316, new_AGEMA_signal_10315, MixColumnsInput[82]}), .a ({new_AGEMA_signal_11498, new_AGEMA_signal_11497, MixColumnsOutput[82]}), .c ({new_AGEMA_signal_11968, new_AGEMA_signal_11967, RoundOutput[82]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U967 ( .s (n316), .b ({new_AGEMA_signal_10314, new_AGEMA_signal_10313, MixColumnsInput[83]}), .a ({new_AGEMA_signal_12032, new_AGEMA_signal_12031, MixColumnsOutput[83]}), .c ({new_AGEMA_signal_12298, new_AGEMA_signal_12297, RoundOutput[83]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U968 ( .s (n316), .b ({new_AGEMA_signal_10312, new_AGEMA_signal_10311, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .a ({new_AGEMA_signal_12028, new_AGEMA_signal_12027, MixColumnsOutput[84]}), .c ({new_AGEMA_signal_12300, new_AGEMA_signal_12299, RoundOutput[84]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U969 ( .s (n316), .b ({new_AGEMA_signal_10310, new_AGEMA_signal_10309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .a ({new_AGEMA_signal_11490, new_AGEMA_signal_11489, MixColumnsOutput[85]}), .c ({new_AGEMA_signal_11970, new_AGEMA_signal_11969, RoundOutput[85]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U970 ( .s (n316), .b ({new_AGEMA_signal_10308, new_AGEMA_signal_10307, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .a ({new_AGEMA_signal_11488, new_AGEMA_signal_11487, MixColumnsOutput[86]}), .c ({new_AGEMA_signal_11972, new_AGEMA_signal_11971, RoundOutput[86]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U971 ( .s (n316), .b ({new_AGEMA_signal_10306, new_AGEMA_signal_10305, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .a ({new_AGEMA_signal_11486, new_AGEMA_signal_11485, MixColumnsOutput[87]}), .c ({new_AGEMA_signal_11974, new_AGEMA_signal_11973, RoundOutput[87]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U972 ( .s (n316), .b ({new_AGEMA_signal_10068, new_AGEMA_signal_10067, MixColumnsInput[88]}), .a ({new_AGEMA_signal_11484, new_AGEMA_signal_11483, MixColumnsOutput[88]}), .c ({new_AGEMA_signal_11976, new_AGEMA_signal_11975, RoundOutput[88]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U973 ( .s (n316), .b ({new_AGEMA_signal_10388, new_AGEMA_signal_10387, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .a ({new_AGEMA_signal_12026, new_AGEMA_signal_12025, MixColumnsOutput[89]}), .c ({new_AGEMA_signal_12302, new_AGEMA_signal_12301, RoundOutput[89]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U974 ( .s (n315), .b ({new_AGEMA_signal_10024, new_AGEMA_signal_10023, MixColumnsInput[8]}), .a ({new_AGEMA_signal_11584, new_AGEMA_signal_11583, MixColumnsOutput[8]}), .c ({new_AGEMA_signal_11978, new_AGEMA_signal_11977, RoundOutput[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U975 ( .s (n315), .b ({new_AGEMA_signal_10386, new_AGEMA_signal_10385, MixColumnsInput[90]}), .a ({new_AGEMA_signal_11480, new_AGEMA_signal_11479, MixColumnsOutput[90]}), .c ({new_AGEMA_signal_11980, new_AGEMA_signal_11979, RoundOutput[90]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U976 ( .s (n315), .b ({new_AGEMA_signal_10384, new_AGEMA_signal_10383, MixColumnsInput[91]}), .a ({new_AGEMA_signal_12024, new_AGEMA_signal_12023, MixColumnsOutput[91]}), .c ({new_AGEMA_signal_12304, new_AGEMA_signal_12303, RoundOutput[91]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U977 ( .s (n315), .b ({new_AGEMA_signal_10382, new_AGEMA_signal_10381, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .a ({new_AGEMA_signal_12022, new_AGEMA_signal_12021, MixColumnsOutput[92]}), .c ({new_AGEMA_signal_12306, new_AGEMA_signal_12305, RoundOutput[92]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U978 ( .s (n315), .b ({new_AGEMA_signal_10380, new_AGEMA_signal_10379, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .a ({new_AGEMA_signal_11474, new_AGEMA_signal_11473, MixColumnsOutput[93]}), .c ({new_AGEMA_signal_11982, new_AGEMA_signal_11981, RoundOutput[93]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U979 ( .s (n315), .b ({new_AGEMA_signal_10378, new_AGEMA_signal_10377, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .a ({new_AGEMA_signal_11470, new_AGEMA_signal_11469, MixColumnsOutput[94]}), .c ({new_AGEMA_signal_11984, new_AGEMA_signal_11983, RoundOutput[94]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U980 ( .s (n315), .b ({new_AGEMA_signal_10376, new_AGEMA_signal_10375, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .a ({new_AGEMA_signal_11468, new_AGEMA_signal_11467, MixColumnsOutput[95]}), .c ({new_AGEMA_signal_11986, new_AGEMA_signal_11985, RoundOutput[95]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U981 ( .s (n315), .b ({new_AGEMA_signal_9826, new_AGEMA_signal_9825, MixColumnsInput[96]}), .a ({new_AGEMA_signal_11452, new_AGEMA_signal_11451, MixColumnsOutput[96]}), .c ({new_AGEMA_signal_11988, new_AGEMA_signal_11987, RoundOutput[96]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U982 ( .s (n315), .b ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .a ({new_AGEMA_signal_12006, new_AGEMA_signal_12005, MixColumnsOutput[97]}), .c ({new_AGEMA_signal_12308, new_AGEMA_signal_12307, RoundOutput[97]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U983 ( .s (n315), .b ({new_AGEMA_signal_10232, new_AGEMA_signal_10231, MixColumnsInput[98]}), .a ({new_AGEMA_signal_11408, new_AGEMA_signal_11407, MixColumnsOutput[98]}), .c ({new_AGEMA_signal_11990, new_AGEMA_signal_11989, RoundOutput[98]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U984 ( .s (n315), .b ({new_AGEMA_signal_10230, new_AGEMA_signal_10229, MixColumnsInput[99]}), .a ({new_AGEMA_signal_11996, new_AGEMA_signal_11995, MixColumnsOutput[99]}), .c ({new_AGEMA_signal_12310, new_AGEMA_signal_12309, RoundOutput[99]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) U985 ( .s (n315), .b ({new_AGEMA_signal_10360, new_AGEMA_signal_10359, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .a ({new_AGEMA_signal_12064, new_AGEMA_signal_12063, MixColumnsOutput[9]}), .c ({new_AGEMA_signal_12312, new_AGEMA_signal_12311, RoundOutput[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11832, new_AGEMA_signal_11831, RoundOutput[0]}), .a ({plaintext_s2[0], plaintext_s1[0], plaintext_s0[0]}), .c ({new_AGEMA_signal_12316, new_AGEMA_signal_12315, RoundReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12246, new_AGEMA_signal_12245, RoundOutput[1]}), .a ({plaintext_s2[1], plaintext_s1[1], plaintext_s0[1]}), .c ({new_AGEMA_signal_12664, new_AGEMA_signal_12663, RoundReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11894, new_AGEMA_signal_11893, RoundOutput[2]}), .a ({plaintext_s2[2], plaintext_s1[2], plaintext_s0[2]}), .c ({new_AGEMA_signal_12320, new_AGEMA_signal_12319, RoundReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12262, new_AGEMA_signal_12261, RoundOutput[3]}), .a ({plaintext_s2[3], plaintext_s1[3], plaintext_s0[3]}), .c ({new_AGEMA_signal_12668, new_AGEMA_signal_12667, RoundReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12272, new_AGEMA_signal_12271, RoundOutput[4]}), .a ({plaintext_s2[4], plaintext_s1[4], plaintext_s0[4]}), .c ({new_AGEMA_signal_12672, new_AGEMA_signal_12671, RoundReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11934, new_AGEMA_signal_11933, RoundOutput[5]}), .a ({plaintext_s2[5], plaintext_s1[5], plaintext_s0[5]}), .c ({new_AGEMA_signal_12324, new_AGEMA_signal_12323, RoundReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11948, new_AGEMA_signal_11947, RoundOutput[6]}), .a ({plaintext_s2[6], plaintext_s1[6], plaintext_s0[6]}), .c ({new_AGEMA_signal_12328, new_AGEMA_signal_12327, RoundReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11964, new_AGEMA_signal_11963, RoundOutput[7]}), .a ({plaintext_s2[7], plaintext_s1[7], plaintext_s0[7]}), .c ({new_AGEMA_signal_12332, new_AGEMA_signal_12331, RoundReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11978, new_AGEMA_signal_11977, RoundOutput[8]}), .a ({plaintext_s2[8], plaintext_s1[8], plaintext_s0[8]}), .c ({new_AGEMA_signal_12336, new_AGEMA_signal_12335, RoundReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12312, new_AGEMA_signal_12311, RoundOutput[9]}), .a ({plaintext_s2[9], plaintext_s1[9], plaintext_s0[9]}), .c ({new_AGEMA_signal_12676, new_AGEMA_signal_12675, RoundReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11846, new_AGEMA_signal_11845, RoundOutput[10]}), .a ({plaintext_s2[10], plaintext_s1[10], plaintext_s0[10]}), .c ({new_AGEMA_signal_12340, new_AGEMA_signal_12339, RoundReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12232, new_AGEMA_signal_12231, RoundOutput[11]}), .a ({plaintext_s2[11], plaintext_s1[11], plaintext_s0[11]}), .c ({new_AGEMA_signal_12680, new_AGEMA_signal_12679, RoundReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12240, new_AGEMA_signal_12239, RoundOutput[12]}), .a ({plaintext_s2[12], plaintext_s1[12], plaintext_s0[12]}), .c ({new_AGEMA_signal_12684, new_AGEMA_signal_12683, RoundReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11872, new_AGEMA_signal_11871, RoundOutput[13]}), .a ({plaintext_s2[13], plaintext_s1[13], plaintext_s0[13]}), .c ({new_AGEMA_signal_12344, new_AGEMA_signal_12343, RoundReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11874, new_AGEMA_signal_11873, RoundOutput[14]}), .a ({plaintext_s2[14], plaintext_s1[14], plaintext_s0[14]}), .c ({new_AGEMA_signal_12348, new_AGEMA_signal_12347, RoundReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11876, new_AGEMA_signal_11875, RoundOutput[15]}), .a ({plaintext_s2[15], plaintext_s1[15], plaintext_s0[15]}), .c ({new_AGEMA_signal_12352, new_AGEMA_signal_12351, RoundReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11878, new_AGEMA_signal_11877, RoundOutput[16]}), .a ({plaintext_s2[16], plaintext_s1[16], plaintext_s0[16]}), .c ({new_AGEMA_signal_12356, new_AGEMA_signal_12355, RoundReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12242, new_AGEMA_signal_12241, RoundOutput[17]}), .a ({plaintext_s2[17], plaintext_s1[17], plaintext_s0[17]}), .c ({new_AGEMA_signal_12688, new_AGEMA_signal_12687, RoundReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11880, new_AGEMA_signal_11879, RoundOutput[18]}), .a ({plaintext_s2[18], plaintext_s1[18], plaintext_s0[18]}), .c ({new_AGEMA_signal_12360, new_AGEMA_signal_12359, RoundReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12244, new_AGEMA_signal_12243, RoundOutput[19]}), .a ({plaintext_s2[19], plaintext_s1[19], plaintext_s0[19]}), .c ({new_AGEMA_signal_12692, new_AGEMA_signal_12691, RoundReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12248, new_AGEMA_signal_12247, RoundOutput[20]}), .a ({plaintext_s2[20], plaintext_s1[20], plaintext_s0[20]}), .c ({new_AGEMA_signal_12696, new_AGEMA_signal_12695, RoundReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11882, new_AGEMA_signal_11881, RoundOutput[21]}), .a ({plaintext_s2[21], plaintext_s1[21], plaintext_s0[21]}), .c ({new_AGEMA_signal_12364, new_AGEMA_signal_12363, RoundReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11884, new_AGEMA_signal_11883, RoundOutput[22]}), .a ({plaintext_s2[22], plaintext_s1[22], plaintext_s0[22]}), .c ({new_AGEMA_signal_12368, new_AGEMA_signal_12367, RoundReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11886, new_AGEMA_signal_11885, RoundOutput[23]}), .a ({plaintext_s2[23], plaintext_s1[23], plaintext_s0[23]}), .c ({new_AGEMA_signal_12372, new_AGEMA_signal_12371, RoundReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11888, new_AGEMA_signal_11887, RoundOutput[24]}), .a ({plaintext_s2[24], plaintext_s1[24], plaintext_s0[24]}), .c ({new_AGEMA_signal_12376, new_AGEMA_signal_12375, RoundReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12250, new_AGEMA_signal_12249, RoundOutput[25]}), .a ({plaintext_s2[25], plaintext_s1[25], plaintext_s0[25]}), .c ({new_AGEMA_signal_12700, new_AGEMA_signal_12699, RoundReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11890, new_AGEMA_signal_11889, RoundOutput[26]}), .a ({plaintext_s2[26], plaintext_s1[26], plaintext_s0[26]}), .c ({new_AGEMA_signal_12380, new_AGEMA_signal_12379, RoundReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12252, new_AGEMA_signal_12251, RoundOutput[27]}), .a ({plaintext_s2[27], plaintext_s1[27], plaintext_s0[27]}), .c ({new_AGEMA_signal_12704, new_AGEMA_signal_12703, RoundReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12254, new_AGEMA_signal_12253, RoundOutput[28]}), .a ({plaintext_s2[28], plaintext_s1[28], plaintext_s0[28]}), .c ({new_AGEMA_signal_12708, new_AGEMA_signal_12707, RoundReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11892, new_AGEMA_signal_11891, RoundOutput[29]}), .a ({plaintext_s2[29], plaintext_s1[29], plaintext_s0[29]}), .c ({new_AGEMA_signal_12384, new_AGEMA_signal_12383, RoundReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11896, new_AGEMA_signal_11895, RoundOutput[30]}), .a ({plaintext_s2[30], plaintext_s1[30], plaintext_s0[30]}), .c ({new_AGEMA_signal_12388, new_AGEMA_signal_12387, RoundReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11898, new_AGEMA_signal_11897, RoundOutput[31]}), .a ({plaintext_s2[31], plaintext_s1[31], plaintext_s0[31]}), .c ({new_AGEMA_signal_12392, new_AGEMA_signal_12391, RoundReg_Inst_ff_SDE_31_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11900, new_AGEMA_signal_11899, RoundOutput[32]}), .a ({plaintext_s2[32], plaintext_s1[32], plaintext_s0[32]}), .c ({new_AGEMA_signal_12396, new_AGEMA_signal_12395, RoundReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12256, new_AGEMA_signal_12255, RoundOutput[33]}), .a ({plaintext_s2[33], plaintext_s1[33], plaintext_s0[33]}), .c ({new_AGEMA_signal_12712, new_AGEMA_signal_12711, RoundReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11902, new_AGEMA_signal_11901, RoundOutput[34]}), .a ({plaintext_s2[34], plaintext_s1[34], plaintext_s0[34]}), .c ({new_AGEMA_signal_12400, new_AGEMA_signal_12399, RoundReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12258, new_AGEMA_signal_12257, RoundOutput[35]}), .a ({plaintext_s2[35], plaintext_s1[35], plaintext_s0[35]}), .c ({new_AGEMA_signal_12716, new_AGEMA_signal_12715, RoundReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12260, new_AGEMA_signal_12259, RoundOutput[36]}), .a ({plaintext_s2[36], plaintext_s1[36], plaintext_s0[36]}), .c ({new_AGEMA_signal_12720, new_AGEMA_signal_12719, RoundReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11904, new_AGEMA_signal_11903, RoundOutput[37]}), .a ({plaintext_s2[37], plaintext_s1[37], plaintext_s0[37]}), .c ({new_AGEMA_signal_12404, new_AGEMA_signal_12403, RoundReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11906, new_AGEMA_signal_11905, RoundOutput[38]}), .a ({plaintext_s2[38], plaintext_s1[38], plaintext_s0[38]}), .c ({new_AGEMA_signal_12408, new_AGEMA_signal_12407, RoundReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11908, new_AGEMA_signal_11907, RoundOutput[39]}), .a ({plaintext_s2[39], plaintext_s1[39], plaintext_s0[39]}), .c ({new_AGEMA_signal_12412, new_AGEMA_signal_12411, RoundReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11910, new_AGEMA_signal_11909, RoundOutput[40]}), .a ({plaintext_s2[40], plaintext_s1[40], plaintext_s0[40]}), .c ({new_AGEMA_signal_12416, new_AGEMA_signal_12415, RoundReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12264, new_AGEMA_signal_12263, RoundOutput[41]}), .a ({plaintext_s2[41], plaintext_s1[41], plaintext_s0[41]}), .c ({new_AGEMA_signal_12724, new_AGEMA_signal_12723, RoundReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11912, new_AGEMA_signal_11911, RoundOutput[42]}), .a ({plaintext_s2[42], plaintext_s1[42], plaintext_s0[42]}), .c ({new_AGEMA_signal_12420, new_AGEMA_signal_12419, RoundReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12266, new_AGEMA_signal_12265, RoundOutput[43]}), .a ({plaintext_s2[43], plaintext_s1[43], plaintext_s0[43]}), .c ({new_AGEMA_signal_12728, new_AGEMA_signal_12727, RoundReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12268, new_AGEMA_signal_12267, RoundOutput[44]}), .a ({plaintext_s2[44], plaintext_s1[44], plaintext_s0[44]}), .c ({new_AGEMA_signal_12732, new_AGEMA_signal_12731, RoundReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11914, new_AGEMA_signal_11913, RoundOutput[45]}), .a ({plaintext_s2[45], plaintext_s1[45], plaintext_s0[45]}), .c ({new_AGEMA_signal_12424, new_AGEMA_signal_12423, RoundReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11916, new_AGEMA_signal_11915, RoundOutput[46]}), .a ({plaintext_s2[46], plaintext_s1[46], plaintext_s0[46]}), .c ({new_AGEMA_signal_12428, new_AGEMA_signal_12427, RoundReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11918, new_AGEMA_signal_11917, RoundOutput[47]}), .a ({plaintext_s2[47], plaintext_s1[47], plaintext_s0[47]}), .c ({new_AGEMA_signal_12432, new_AGEMA_signal_12431, RoundReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11920, new_AGEMA_signal_11919, RoundOutput[48]}), .a ({plaintext_s2[48], plaintext_s1[48], plaintext_s0[48]}), .c ({new_AGEMA_signal_12436, new_AGEMA_signal_12435, RoundReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12270, new_AGEMA_signal_12269, RoundOutput[49]}), .a ({plaintext_s2[49], plaintext_s1[49], plaintext_s0[49]}), .c ({new_AGEMA_signal_12736, new_AGEMA_signal_12735, RoundReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11922, new_AGEMA_signal_11921, RoundOutput[50]}), .a ({plaintext_s2[50], plaintext_s1[50], plaintext_s0[50]}), .c ({new_AGEMA_signal_12440, new_AGEMA_signal_12439, RoundReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12274, new_AGEMA_signal_12273, RoundOutput[51]}), .a ({plaintext_s2[51], plaintext_s1[51], plaintext_s0[51]}), .c ({new_AGEMA_signal_12740, new_AGEMA_signal_12739, RoundReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12276, new_AGEMA_signal_12275, RoundOutput[52]}), .a ({plaintext_s2[52], plaintext_s1[52], plaintext_s0[52]}), .c ({new_AGEMA_signal_12744, new_AGEMA_signal_12743, RoundReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11924, new_AGEMA_signal_11923, RoundOutput[53]}), .a ({plaintext_s2[53], plaintext_s1[53], plaintext_s0[53]}), .c ({new_AGEMA_signal_12444, new_AGEMA_signal_12443, RoundReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11926, new_AGEMA_signal_11925, RoundOutput[54]}), .a ({plaintext_s2[54], plaintext_s1[54], plaintext_s0[54]}), .c ({new_AGEMA_signal_12448, new_AGEMA_signal_12447, RoundReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11928, new_AGEMA_signal_11927, RoundOutput[55]}), .a ({plaintext_s2[55], plaintext_s1[55], plaintext_s0[55]}), .c ({new_AGEMA_signal_12452, new_AGEMA_signal_12451, RoundReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11930, new_AGEMA_signal_11929, RoundOutput[56]}), .a ({plaintext_s2[56], plaintext_s1[56], plaintext_s0[56]}), .c ({new_AGEMA_signal_12456, new_AGEMA_signal_12455, RoundReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12278, new_AGEMA_signal_12277, RoundOutput[57]}), .a ({plaintext_s2[57], plaintext_s1[57], plaintext_s0[57]}), .c ({new_AGEMA_signal_12748, new_AGEMA_signal_12747, RoundReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11932, new_AGEMA_signal_11931, RoundOutput[58]}), .a ({plaintext_s2[58], plaintext_s1[58], plaintext_s0[58]}), .c ({new_AGEMA_signal_12460, new_AGEMA_signal_12459, RoundReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12280, new_AGEMA_signal_12279, RoundOutput[59]}), .a ({plaintext_s2[59], plaintext_s1[59], plaintext_s0[59]}), .c ({new_AGEMA_signal_12752, new_AGEMA_signal_12751, RoundReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12282, new_AGEMA_signal_12281, RoundOutput[60]}), .a ({plaintext_s2[60], plaintext_s1[60], plaintext_s0[60]}), .c ({new_AGEMA_signal_12756, new_AGEMA_signal_12755, RoundReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11936, new_AGEMA_signal_11935, RoundOutput[61]}), .a ({plaintext_s2[61], plaintext_s1[61], plaintext_s0[61]}), .c ({new_AGEMA_signal_12464, new_AGEMA_signal_12463, RoundReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11938, new_AGEMA_signal_11937, RoundOutput[62]}), .a ({plaintext_s2[62], plaintext_s1[62], plaintext_s0[62]}), .c ({new_AGEMA_signal_12468, new_AGEMA_signal_12467, RoundReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11940, new_AGEMA_signal_11939, RoundOutput[63]}), .a ({plaintext_s2[63], plaintext_s1[63], plaintext_s0[63]}), .c ({new_AGEMA_signal_12472, new_AGEMA_signal_12471, RoundReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11942, new_AGEMA_signal_11941, RoundOutput[64]}), .a ({plaintext_s2[64], plaintext_s1[64], plaintext_s0[64]}), .c ({new_AGEMA_signal_12476, new_AGEMA_signal_12475, RoundReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12284, new_AGEMA_signal_12283, RoundOutput[65]}), .a ({plaintext_s2[65], plaintext_s1[65], plaintext_s0[65]}), .c ({new_AGEMA_signal_12760, new_AGEMA_signal_12759, RoundReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11944, new_AGEMA_signal_11943, RoundOutput[66]}), .a ({plaintext_s2[66], plaintext_s1[66], plaintext_s0[66]}), .c ({new_AGEMA_signal_12480, new_AGEMA_signal_12479, RoundReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12286, new_AGEMA_signal_12285, RoundOutput[67]}), .a ({plaintext_s2[67], plaintext_s1[67], plaintext_s0[67]}), .c ({new_AGEMA_signal_12764, new_AGEMA_signal_12763, RoundReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12288, new_AGEMA_signal_12287, RoundOutput[68]}), .a ({plaintext_s2[68], plaintext_s1[68], plaintext_s0[68]}), .c ({new_AGEMA_signal_12768, new_AGEMA_signal_12767, RoundReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11946, new_AGEMA_signal_11945, RoundOutput[69]}), .a ({plaintext_s2[69], plaintext_s1[69], plaintext_s0[69]}), .c ({new_AGEMA_signal_12484, new_AGEMA_signal_12483, RoundReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11950, new_AGEMA_signal_11949, RoundOutput[70]}), .a ({plaintext_s2[70], plaintext_s1[70], plaintext_s0[70]}), .c ({new_AGEMA_signal_12488, new_AGEMA_signal_12487, RoundReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11952, new_AGEMA_signal_11951, RoundOutput[71]}), .a ({plaintext_s2[71], plaintext_s1[71], plaintext_s0[71]}), .c ({new_AGEMA_signal_12492, new_AGEMA_signal_12491, RoundReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11954, new_AGEMA_signal_11953, RoundOutput[72]}), .a ({plaintext_s2[72], plaintext_s1[72], plaintext_s0[72]}), .c ({new_AGEMA_signal_12496, new_AGEMA_signal_12495, RoundReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12290, new_AGEMA_signal_12289, RoundOutput[73]}), .a ({plaintext_s2[73], plaintext_s1[73], plaintext_s0[73]}), .c ({new_AGEMA_signal_12772, new_AGEMA_signal_12771, RoundReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11956, new_AGEMA_signal_11955, RoundOutput[74]}), .a ({plaintext_s2[74], plaintext_s1[74], plaintext_s0[74]}), .c ({new_AGEMA_signal_12500, new_AGEMA_signal_12499, RoundReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12292, new_AGEMA_signal_12291, RoundOutput[75]}), .a ({plaintext_s2[75], plaintext_s1[75], plaintext_s0[75]}), .c ({new_AGEMA_signal_12776, new_AGEMA_signal_12775, RoundReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12294, new_AGEMA_signal_12293, RoundOutput[76]}), .a ({plaintext_s2[76], plaintext_s1[76], plaintext_s0[76]}), .c ({new_AGEMA_signal_12780, new_AGEMA_signal_12779, RoundReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11958, new_AGEMA_signal_11957, RoundOutput[77]}), .a ({plaintext_s2[77], plaintext_s1[77], plaintext_s0[77]}), .c ({new_AGEMA_signal_12504, new_AGEMA_signal_12503, RoundReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11960, new_AGEMA_signal_11959, RoundOutput[78]}), .a ({plaintext_s2[78], plaintext_s1[78], plaintext_s0[78]}), .c ({new_AGEMA_signal_12508, new_AGEMA_signal_12507, RoundReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11962, new_AGEMA_signal_11961, RoundOutput[79]}), .a ({plaintext_s2[79], plaintext_s1[79], plaintext_s0[79]}), .c ({new_AGEMA_signal_12512, new_AGEMA_signal_12511, RoundReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11966, new_AGEMA_signal_11965, RoundOutput[80]}), .a ({plaintext_s2[80], plaintext_s1[80], plaintext_s0[80]}), .c ({new_AGEMA_signal_12516, new_AGEMA_signal_12515, RoundReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12296, new_AGEMA_signal_12295, RoundOutput[81]}), .a ({plaintext_s2[81], plaintext_s1[81], plaintext_s0[81]}), .c ({new_AGEMA_signal_12784, new_AGEMA_signal_12783, RoundReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11968, new_AGEMA_signal_11967, RoundOutput[82]}), .a ({plaintext_s2[82], plaintext_s1[82], plaintext_s0[82]}), .c ({new_AGEMA_signal_12520, new_AGEMA_signal_12519, RoundReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12298, new_AGEMA_signal_12297, RoundOutput[83]}), .a ({plaintext_s2[83], plaintext_s1[83], plaintext_s0[83]}), .c ({new_AGEMA_signal_12788, new_AGEMA_signal_12787, RoundReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12300, new_AGEMA_signal_12299, RoundOutput[84]}), .a ({plaintext_s2[84], plaintext_s1[84], plaintext_s0[84]}), .c ({new_AGEMA_signal_12792, new_AGEMA_signal_12791, RoundReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11970, new_AGEMA_signal_11969, RoundOutput[85]}), .a ({plaintext_s2[85], plaintext_s1[85], plaintext_s0[85]}), .c ({new_AGEMA_signal_12524, new_AGEMA_signal_12523, RoundReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11972, new_AGEMA_signal_11971, RoundOutput[86]}), .a ({plaintext_s2[86], plaintext_s1[86], plaintext_s0[86]}), .c ({new_AGEMA_signal_12528, new_AGEMA_signal_12527, RoundReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11974, new_AGEMA_signal_11973, RoundOutput[87]}), .a ({plaintext_s2[87], plaintext_s1[87], plaintext_s0[87]}), .c ({new_AGEMA_signal_12532, new_AGEMA_signal_12531, RoundReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11976, new_AGEMA_signal_11975, RoundOutput[88]}), .a ({plaintext_s2[88], plaintext_s1[88], plaintext_s0[88]}), .c ({new_AGEMA_signal_12536, new_AGEMA_signal_12535, RoundReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12302, new_AGEMA_signal_12301, RoundOutput[89]}), .a ({plaintext_s2[89], plaintext_s1[89], plaintext_s0[89]}), .c ({new_AGEMA_signal_12796, new_AGEMA_signal_12795, RoundReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11980, new_AGEMA_signal_11979, RoundOutput[90]}), .a ({plaintext_s2[90], plaintext_s1[90], plaintext_s0[90]}), .c ({new_AGEMA_signal_12540, new_AGEMA_signal_12539, RoundReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12304, new_AGEMA_signal_12303, RoundOutput[91]}), .a ({plaintext_s2[91], plaintext_s1[91], plaintext_s0[91]}), .c ({new_AGEMA_signal_12800, new_AGEMA_signal_12799, RoundReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12306, new_AGEMA_signal_12305, RoundOutput[92]}), .a ({plaintext_s2[92], plaintext_s1[92], plaintext_s0[92]}), .c ({new_AGEMA_signal_12804, new_AGEMA_signal_12803, RoundReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11982, new_AGEMA_signal_11981, RoundOutput[93]}), .a ({plaintext_s2[93], plaintext_s1[93], plaintext_s0[93]}), .c ({new_AGEMA_signal_12544, new_AGEMA_signal_12543, RoundReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11984, new_AGEMA_signal_11983, RoundOutput[94]}), .a ({plaintext_s2[94], plaintext_s1[94], plaintext_s0[94]}), .c ({new_AGEMA_signal_12548, new_AGEMA_signal_12547, RoundReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11986, new_AGEMA_signal_11985, RoundOutput[95]}), .a ({plaintext_s2[95], plaintext_s1[95], plaintext_s0[95]}), .c ({new_AGEMA_signal_12552, new_AGEMA_signal_12551, RoundReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11988, new_AGEMA_signal_11987, RoundOutput[96]}), .a ({plaintext_s2[96], plaintext_s1[96], plaintext_s0[96]}), .c ({new_AGEMA_signal_12556, new_AGEMA_signal_12555, RoundReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12308, new_AGEMA_signal_12307, RoundOutput[97]}), .a ({plaintext_s2[97], plaintext_s1[97], plaintext_s0[97]}), .c ({new_AGEMA_signal_12808, new_AGEMA_signal_12807, RoundReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11990, new_AGEMA_signal_11989, RoundOutput[98]}), .a ({plaintext_s2[98], plaintext_s1[98], plaintext_s0[98]}), .c ({new_AGEMA_signal_12560, new_AGEMA_signal_12559, RoundReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12310, new_AGEMA_signal_12309, RoundOutput[99]}), .a ({plaintext_s2[99], plaintext_s1[99], plaintext_s0[99]}), .c ({new_AGEMA_signal_12812, new_AGEMA_signal_12811, RoundReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12218, new_AGEMA_signal_12217, RoundOutput[100]}), .a ({plaintext_s2[100], plaintext_s1[100], plaintext_s0[100]}), .c ({new_AGEMA_signal_12816, new_AGEMA_signal_12815, RoundReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11834, new_AGEMA_signal_11833, RoundOutput[101]}), .a ({plaintext_s2[101], plaintext_s1[101], plaintext_s0[101]}), .c ({new_AGEMA_signal_12564, new_AGEMA_signal_12563, RoundReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11836, new_AGEMA_signal_11835, RoundOutput[102]}), .a ({plaintext_s2[102], plaintext_s1[102], plaintext_s0[102]}), .c ({new_AGEMA_signal_12568, new_AGEMA_signal_12567, RoundReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11838, new_AGEMA_signal_11837, RoundOutput[103]}), .a ({plaintext_s2[103], plaintext_s1[103], plaintext_s0[103]}), .c ({new_AGEMA_signal_12572, new_AGEMA_signal_12571, RoundReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11840, new_AGEMA_signal_11839, RoundOutput[104]}), .a ({plaintext_s2[104], plaintext_s1[104], plaintext_s0[104]}), .c ({new_AGEMA_signal_12576, new_AGEMA_signal_12575, RoundReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12220, new_AGEMA_signal_12219, RoundOutput[105]}), .a ({plaintext_s2[105], plaintext_s1[105], plaintext_s0[105]}), .c ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, RoundReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11842, new_AGEMA_signal_11841, RoundOutput[106]}), .a ({plaintext_s2[106], plaintext_s1[106], plaintext_s0[106]}), .c ({new_AGEMA_signal_12580, new_AGEMA_signal_12579, RoundReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12222, new_AGEMA_signal_12221, RoundOutput[107]}), .a ({plaintext_s2[107], plaintext_s1[107], plaintext_s0[107]}), .c ({new_AGEMA_signal_12824, new_AGEMA_signal_12823, RoundReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12224, new_AGEMA_signal_12223, RoundOutput[108]}), .a ({plaintext_s2[108], plaintext_s1[108], plaintext_s0[108]}), .c ({new_AGEMA_signal_12828, new_AGEMA_signal_12827, RoundReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11844, new_AGEMA_signal_11843, RoundOutput[109]}), .a ({plaintext_s2[109], plaintext_s1[109], plaintext_s0[109]}), .c ({new_AGEMA_signal_12584, new_AGEMA_signal_12583, RoundReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11848, new_AGEMA_signal_11847, RoundOutput[110]}), .a ({plaintext_s2[110], plaintext_s1[110], plaintext_s0[110]}), .c ({new_AGEMA_signal_12588, new_AGEMA_signal_12587, RoundReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11850, new_AGEMA_signal_11849, RoundOutput[111]}), .a ({plaintext_s2[111], plaintext_s1[111], plaintext_s0[111]}), .c ({new_AGEMA_signal_12592, new_AGEMA_signal_12591, RoundReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11852, new_AGEMA_signal_11851, RoundOutput[112]}), .a ({plaintext_s2[112], plaintext_s1[112], plaintext_s0[112]}), .c ({new_AGEMA_signal_12596, new_AGEMA_signal_12595, RoundReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12226, new_AGEMA_signal_12225, RoundOutput[113]}), .a ({plaintext_s2[113], plaintext_s1[113], plaintext_s0[113]}), .c ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, RoundReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11854, new_AGEMA_signal_11853, RoundOutput[114]}), .a ({plaintext_s2[114], plaintext_s1[114], plaintext_s0[114]}), .c ({new_AGEMA_signal_12600, new_AGEMA_signal_12599, RoundReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12228, new_AGEMA_signal_12227, RoundOutput[115]}), .a ({plaintext_s2[115], plaintext_s1[115], plaintext_s0[115]}), .c ({new_AGEMA_signal_12836, new_AGEMA_signal_12835, RoundReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12230, new_AGEMA_signal_12229, RoundOutput[116]}), .a ({plaintext_s2[116], plaintext_s1[116], plaintext_s0[116]}), .c ({new_AGEMA_signal_12840, new_AGEMA_signal_12839, RoundReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11856, new_AGEMA_signal_11855, RoundOutput[117]}), .a ({plaintext_s2[117], plaintext_s1[117], plaintext_s0[117]}), .c ({new_AGEMA_signal_12604, new_AGEMA_signal_12603, RoundReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11858, new_AGEMA_signal_11857, RoundOutput[118]}), .a ({plaintext_s2[118], plaintext_s1[118], plaintext_s0[118]}), .c ({new_AGEMA_signal_12608, new_AGEMA_signal_12607, RoundReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11860, new_AGEMA_signal_11859, RoundOutput[119]}), .a ({plaintext_s2[119], plaintext_s1[119], plaintext_s0[119]}), .c ({new_AGEMA_signal_12612, new_AGEMA_signal_12611, RoundReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11862, new_AGEMA_signal_11861, RoundOutput[120]}), .a ({plaintext_s2[120], plaintext_s1[120], plaintext_s0[120]}), .c ({new_AGEMA_signal_12616, new_AGEMA_signal_12615, RoundReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12234, new_AGEMA_signal_12233, RoundOutput[121]}), .a ({plaintext_s2[121], plaintext_s1[121], plaintext_s0[121]}), .c ({new_AGEMA_signal_12844, new_AGEMA_signal_12843, RoundReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11864, new_AGEMA_signal_11863, RoundOutput[122]}), .a ({plaintext_s2[122], plaintext_s1[122], plaintext_s0[122]}), .c ({new_AGEMA_signal_12620, new_AGEMA_signal_12619, RoundReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12236, new_AGEMA_signal_12235, RoundOutput[123]}), .a ({plaintext_s2[123], plaintext_s1[123], plaintext_s0[123]}), .c ({new_AGEMA_signal_12848, new_AGEMA_signal_12847, RoundReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12238, new_AGEMA_signal_12237, RoundOutput[124]}), .a ({plaintext_s2[124], plaintext_s1[124], plaintext_s0[124]}), .c ({new_AGEMA_signal_12852, new_AGEMA_signal_12851, RoundReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11866, new_AGEMA_signal_11865, RoundOutput[125]}), .a ({plaintext_s2[125], plaintext_s1[125], plaintext_s0[125]}), .c ({new_AGEMA_signal_12624, new_AGEMA_signal_12623, RoundReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11868, new_AGEMA_signal_11867, RoundOutput[126]}), .a ({plaintext_s2[126], plaintext_s1[126], plaintext_s0[126]}), .c ({new_AGEMA_signal_12628, new_AGEMA_signal_12627, RoundReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11870, new_AGEMA_signal_11869, RoundOutput[127]}), .a ({plaintext_s2[127], plaintext_s1[127], plaintext_s0[127]}), .c ({new_AGEMA_signal_12632, new_AGEMA_signal_12631, RoundReg_Inst_ff_SDE_127_next_state}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M46_U1 ( .a ({new_AGEMA_signal_8100, new_AGEMA_signal_8099, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_5782, new_AGEMA_signal_5781, SubBytesIns_Inst_Sbox_0_T6}), .clk (clk), .r ({Fresh[962], Fresh[961], Fresh[960]}), .c ({new_AGEMA_signal_8576, new_AGEMA_signal_8575, SubBytesIns_Inst_Sbox_0_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M47_U1 ( .a ({new_AGEMA_signal_7876, new_AGEMA_signal_7875, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_6142, new_AGEMA_signal_6141, SubBytesIns_Inst_Sbox_0_T8}), .clk (clk), .r ({Fresh[965], Fresh[964], Fresh[963]}), .c ({new_AGEMA_signal_8102, new_AGEMA_signal_8101, SubBytesIns_Inst_Sbox_0_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M48_U1 ( .a ({new_AGEMA_signal_7874, new_AGEMA_signal_7873, SubBytesIns_Inst_Sbox_0_M39}), .b ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .clk (clk), .r ({Fresh[968], Fresh[967], Fresh[966]}), .c ({new_AGEMA_signal_8104, new_AGEMA_signal_8103, SubBytesIns_Inst_Sbox_0_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M49_U1 ( .a ({new_AGEMA_signal_8098, new_AGEMA_signal_8097, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_5790, new_AGEMA_signal_5789, SubBytesIns_Inst_Sbox_0_T16}), .clk (clk), .r ({Fresh[971], Fresh[970], Fresh[969]}), .c ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, SubBytesIns_Inst_Sbox_0_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M50_U1 ( .a ({new_AGEMA_signal_7872, new_AGEMA_signal_7871, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_5784, new_AGEMA_signal_5783, SubBytesIns_Inst_Sbox_0_T9}), .clk (clk), .r ({Fresh[974], Fresh[973], Fresh[972]}), .c ({new_AGEMA_signal_8106, new_AGEMA_signal_8105, SubBytesIns_Inst_Sbox_0_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M51_U1 ( .a ({new_AGEMA_signal_7870, new_AGEMA_signal_7869, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_6148, new_AGEMA_signal_6147, SubBytesIns_Inst_Sbox_0_T17}), .clk (clk), .r ({Fresh[977], Fresh[976], Fresh[975]}), .c ({new_AGEMA_signal_8108, new_AGEMA_signal_8107, SubBytesIns_Inst_Sbox_0_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M52_U1 ( .a ({new_AGEMA_signal_8096, new_AGEMA_signal_8095, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_5788, new_AGEMA_signal_5787, SubBytesIns_Inst_Sbox_0_T15}), .clk (clk), .r ({Fresh[980], Fresh[979], Fresh[978]}), .c ({new_AGEMA_signal_8580, new_AGEMA_signal_8579, SubBytesIns_Inst_Sbox_0_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M53_U1 ( .a ({new_AGEMA_signal_8574, new_AGEMA_signal_8573, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_5796, new_AGEMA_signal_5795, SubBytesIns_Inst_Sbox_0_T27}), .clk (clk), .r ({Fresh[983], Fresh[982], Fresh[981]}), .c ({new_AGEMA_signal_9038, new_AGEMA_signal_9037, SubBytesIns_Inst_Sbox_0_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M54_U1 ( .a ({new_AGEMA_signal_8094, new_AGEMA_signal_8093, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_6144, new_AGEMA_signal_6143, SubBytesIns_Inst_Sbox_0_T10}), .clk (clk), .r ({Fresh[986], Fresh[985], Fresh[984]}), .c ({new_AGEMA_signal_8582, new_AGEMA_signal_8581, SubBytesIns_Inst_Sbox_0_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M55_U1 ( .a ({new_AGEMA_signal_8100, new_AGEMA_signal_8099, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_5786, new_AGEMA_signal_5785, SubBytesIns_Inst_Sbox_0_T13}), .clk (clk), .r ({Fresh[989], Fresh[988], Fresh[987]}), .c ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, SubBytesIns_Inst_Sbox_0_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M56_U1 ( .a ({new_AGEMA_signal_7876, new_AGEMA_signal_7875, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_6152, new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_0_T23}), .clk (clk), .r ({Fresh[992], Fresh[991], Fresh[990]}), .c ({new_AGEMA_signal_8110, new_AGEMA_signal_8109, SubBytesIns_Inst_Sbox_0_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M57_U1 ( .a ({new_AGEMA_signal_7874, new_AGEMA_signal_7873, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_5792, new_AGEMA_signal_5791, SubBytesIns_Inst_Sbox_0_T19}), .clk (clk), .r ({Fresh[995], Fresh[994], Fresh[993]}), .c ({new_AGEMA_signal_8112, new_AGEMA_signal_8111, SubBytesIns_Inst_Sbox_0_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M58_U1 ( .a ({new_AGEMA_signal_8098, new_AGEMA_signal_8097, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_5402, new_AGEMA_signal_5401, SubBytesIns_Inst_Sbox_0_T3}), .clk (clk), .r ({Fresh[998], Fresh[997], Fresh[996]}), .c ({new_AGEMA_signal_8586, new_AGEMA_signal_8585, SubBytesIns_Inst_Sbox_0_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M59_U1 ( .a ({new_AGEMA_signal_7872, new_AGEMA_signal_7871, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_5794, new_AGEMA_signal_5793, SubBytesIns_Inst_Sbox_0_T22}), .clk (clk), .r ({Fresh[1001], Fresh[1000], Fresh[999]}), .c ({new_AGEMA_signal_8114, new_AGEMA_signal_8113, SubBytesIns_Inst_Sbox_0_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M60_U1 ( .a ({new_AGEMA_signal_7870, new_AGEMA_signal_7869, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_6150, new_AGEMA_signal_6149, SubBytesIns_Inst_Sbox_0_T20}), .clk (clk), .r ({Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({new_AGEMA_signal_8116, new_AGEMA_signal_8115, SubBytesIns_Inst_Sbox_0_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M61_U1 ( .a ({new_AGEMA_signal_8096, new_AGEMA_signal_8095, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_5398, new_AGEMA_signal_5397, SubBytesIns_Inst_Sbox_0_T1}), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005]}), .c ({new_AGEMA_signal_8588, new_AGEMA_signal_8587, SubBytesIns_Inst_Sbox_0_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M62_U1 ( .a ({new_AGEMA_signal_8574, new_AGEMA_signal_8573, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_5404, new_AGEMA_signal_5403, SubBytesIns_Inst_Sbox_0_T4}), .clk (clk), .r ({Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({new_AGEMA_signal_9040, new_AGEMA_signal_9039, SubBytesIns_Inst_Sbox_0_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M63_U1 ( .a ({new_AGEMA_signal_8094, new_AGEMA_signal_8093, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, SubBytesIns_Inst_Sbox_0_T2}), .clk (clk), .r ({Fresh[1013], Fresh[1012], Fresh[1011]}), .c ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, SubBytesIns_Inst_Sbox_0_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L0_U1 ( .a ({new_AGEMA_signal_8588, new_AGEMA_signal_8587, SubBytesIns_Inst_Sbox_0_M61}), .b ({new_AGEMA_signal_9040, new_AGEMA_signal_9039, SubBytesIns_Inst_Sbox_0_M62}), .c ({new_AGEMA_signal_9430, new_AGEMA_signal_9429, SubBytesIns_Inst_Sbox_0_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L1_U1 ( .a ({new_AGEMA_signal_8106, new_AGEMA_signal_8105, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_8110, new_AGEMA_signal_8109, SubBytesIns_Inst_Sbox_0_M56}), .c ({new_AGEMA_signal_8592, new_AGEMA_signal_8591, SubBytesIns_Inst_Sbox_0_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L2_U1 ( .a ({new_AGEMA_signal_8576, new_AGEMA_signal_8575, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_8104, new_AGEMA_signal_8103, SubBytesIns_Inst_Sbox_0_M48}), .c ({new_AGEMA_signal_9042, new_AGEMA_signal_9041, SubBytesIns_Inst_Sbox_0_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L3_U1 ( .a ({new_AGEMA_signal_8102, new_AGEMA_signal_8101, SubBytesIns_Inst_Sbox_0_M47}), .b ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, SubBytesIns_Inst_Sbox_0_M55}), .c ({new_AGEMA_signal_9044, new_AGEMA_signal_9043, SubBytesIns_Inst_Sbox_0_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L4_U1 ( .a ({new_AGEMA_signal_8582, new_AGEMA_signal_8581, SubBytesIns_Inst_Sbox_0_M54}), .b ({new_AGEMA_signal_8586, new_AGEMA_signal_8585, SubBytesIns_Inst_Sbox_0_M58}), .c ({new_AGEMA_signal_9046, new_AGEMA_signal_9045, SubBytesIns_Inst_Sbox_0_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L5_U1 ( .a ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, SubBytesIns_Inst_Sbox_0_M49}), .b ({new_AGEMA_signal_8588, new_AGEMA_signal_8587, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_9048, new_AGEMA_signal_9047, SubBytesIns_Inst_Sbox_0_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L6_U1 ( .a ({new_AGEMA_signal_9040, new_AGEMA_signal_9039, SubBytesIns_Inst_Sbox_0_M62}), .b ({new_AGEMA_signal_9048, new_AGEMA_signal_9047, SubBytesIns_Inst_Sbox_0_L5}), .c ({new_AGEMA_signal_9432, new_AGEMA_signal_9431, SubBytesIns_Inst_Sbox_0_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L7_U1 ( .a ({new_AGEMA_signal_8576, new_AGEMA_signal_8575, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_9044, new_AGEMA_signal_9043, SubBytesIns_Inst_Sbox_0_L3}), .c ({new_AGEMA_signal_9434, new_AGEMA_signal_9433, SubBytesIns_Inst_Sbox_0_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L8_U1 ( .a ({new_AGEMA_signal_8108, new_AGEMA_signal_8107, SubBytesIns_Inst_Sbox_0_M51}), .b ({new_AGEMA_signal_8114, new_AGEMA_signal_8113, SubBytesIns_Inst_Sbox_0_M59}), .c ({new_AGEMA_signal_8594, new_AGEMA_signal_8593, SubBytesIns_Inst_Sbox_0_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L9_U1 ( .a ({new_AGEMA_signal_8580, new_AGEMA_signal_8579, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_9038, new_AGEMA_signal_9037, SubBytesIns_Inst_Sbox_0_M53}), .c ({new_AGEMA_signal_9436, new_AGEMA_signal_9435, SubBytesIns_Inst_Sbox_0_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L10_U1 ( .a ({new_AGEMA_signal_9038, new_AGEMA_signal_9037, SubBytesIns_Inst_Sbox_0_M53}), .b ({new_AGEMA_signal_9046, new_AGEMA_signal_9045, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_9438, new_AGEMA_signal_9437, SubBytesIns_Inst_Sbox_0_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L11_U1 ( .a ({new_AGEMA_signal_8116, new_AGEMA_signal_8115, SubBytesIns_Inst_Sbox_0_M60}), .b ({new_AGEMA_signal_9042, new_AGEMA_signal_9041, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_9440, new_AGEMA_signal_9439, SubBytesIns_Inst_Sbox_0_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L12_U1 ( .a ({new_AGEMA_signal_8104, new_AGEMA_signal_8103, SubBytesIns_Inst_Sbox_0_M48}), .b ({new_AGEMA_signal_8108, new_AGEMA_signal_8107, SubBytesIns_Inst_Sbox_0_M51}), .c ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, SubBytesIns_Inst_Sbox_0_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L13_U1 ( .a ({new_AGEMA_signal_8106, new_AGEMA_signal_8105, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_9430, new_AGEMA_signal_9429, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_9806, new_AGEMA_signal_9805, SubBytesIns_Inst_Sbox_0_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L14_U1 ( .a ({new_AGEMA_signal_8580, new_AGEMA_signal_8579, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_8588, new_AGEMA_signal_8587, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_9050, new_AGEMA_signal_9049, SubBytesIns_Inst_Sbox_0_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L15_U1 ( .a ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, SubBytesIns_Inst_Sbox_0_M55}), .b ({new_AGEMA_signal_8592, new_AGEMA_signal_8591, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_9052, new_AGEMA_signal_9051, SubBytesIns_Inst_Sbox_0_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L16_U1 ( .a ({new_AGEMA_signal_8110, new_AGEMA_signal_8109, SubBytesIns_Inst_Sbox_0_M56}), .b ({new_AGEMA_signal_9430, new_AGEMA_signal_9429, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_9808, new_AGEMA_signal_9807, SubBytesIns_Inst_Sbox_0_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L17_U1 ( .a ({new_AGEMA_signal_8112, new_AGEMA_signal_8111, SubBytesIns_Inst_Sbox_0_M57}), .b ({new_AGEMA_signal_8592, new_AGEMA_signal_8591, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_9054, new_AGEMA_signal_9053, SubBytesIns_Inst_Sbox_0_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L18_U1 ( .a ({new_AGEMA_signal_8586, new_AGEMA_signal_8585, SubBytesIns_Inst_Sbox_0_M58}), .b ({new_AGEMA_signal_8594, new_AGEMA_signal_8593, SubBytesIns_Inst_Sbox_0_L8}), .c ({new_AGEMA_signal_9056, new_AGEMA_signal_9055, SubBytesIns_Inst_Sbox_0_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L19_U1 ( .a ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, SubBytesIns_Inst_Sbox_0_M63}), .b ({new_AGEMA_signal_9046, new_AGEMA_signal_9045, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_9442, new_AGEMA_signal_9441, SubBytesIns_Inst_Sbox_0_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L20_U1 ( .a ({new_AGEMA_signal_9430, new_AGEMA_signal_9429, SubBytesIns_Inst_Sbox_0_L0}), .b ({new_AGEMA_signal_8592, new_AGEMA_signal_8591, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_9810, new_AGEMA_signal_9809, SubBytesIns_Inst_Sbox_0_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L21_U1 ( .a ({new_AGEMA_signal_8592, new_AGEMA_signal_8591, SubBytesIns_Inst_Sbox_0_L1}), .b ({new_AGEMA_signal_9434, new_AGEMA_signal_9433, SubBytesIns_Inst_Sbox_0_L7}), .c ({new_AGEMA_signal_9812, new_AGEMA_signal_9811, SubBytesIns_Inst_Sbox_0_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L22_U1 ( .a ({new_AGEMA_signal_9044, new_AGEMA_signal_9043, SubBytesIns_Inst_Sbox_0_L3}), .b ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, SubBytesIns_Inst_Sbox_0_L12}), .c ({new_AGEMA_signal_9444, new_AGEMA_signal_9443, SubBytesIns_Inst_Sbox_0_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L23_U1 ( .a ({new_AGEMA_signal_9056, new_AGEMA_signal_9055, SubBytesIns_Inst_Sbox_0_L18}), .b ({new_AGEMA_signal_9042, new_AGEMA_signal_9041, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_9446, new_AGEMA_signal_9445, SubBytesIns_Inst_Sbox_0_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L24_U1 ( .a ({new_AGEMA_signal_9052, new_AGEMA_signal_9051, SubBytesIns_Inst_Sbox_0_L15}), .b ({new_AGEMA_signal_9436, new_AGEMA_signal_9435, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_9814, new_AGEMA_signal_9813, SubBytesIns_Inst_Sbox_0_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L25_U1 ( .a ({new_AGEMA_signal_9432, new_AGEMA_signal_9431, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_9438, new_AGEMA_signal_9437, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_9816, new_AGEMA_signal_9815, SubBytesIns_Inst_Sbox_0_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L26_U1 ( .a ({new_AGEMA_signal_9434, new_AGEMA_signal_9433, SubBytesIns_Inst_Sbox_0_L7}), .b ({new_AGEMA_signal_9436, new_AGEMA_signal_9435, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_9818, new_AGEMA_signal_9817, SubBytesIns_Inst_Sbox_0_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L27_U1 ( .a ({new_AGEMA_signal_8594, new_AGEMA_signal_8593, SubBytesIns_Inst_Sbox_0_L8}), .b ({new_AGEMA_signal_9438, new_AGEMA_signal_9437, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_9820, new_AGEMA_signal_9819, SubBytesIns_Inst_Sbox_0_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L28_U1 ( .a ({new_AGEMA_signal_9440, new_AGEMA_signal_9439, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_9050, new_AGEMA_signal_9049, SubBytesIns_Inst_Sbox_0_L14}), .c ({new_AGEMA_signal_9822, new_AGEMA_signal_9821, SubBytesIns_Inst_Sbox_0_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L29_U1 ( .a ({new_AGEMA_signal_9440, new_AGEMA_signal_9439, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_9054, new_AGEMA_signal_9053, SubBytesIns_Inst_Sbox_0_L17}), .c ({new_AGEMA_signal_9824, new_AGEMA_signal_9823, SubBytesIns_Inst_Sbox_0_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S0_U1 ( .a ({new_AGEMA_signal_9432, new_AGEMA_signal_9431, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_9814, new_AGEMA_signal_9813, SubBytesIns_Inst_Sbox_0_L24}), .c ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S1_U1 ( .a ({new_AGEMA_signal_9808, new_AGEMA_signal_9807, SubBytesIns_Inst_Sbox_0_L16}), .b ({new_AGEMA_signal_9818, new_AGEMA_signal_9817, SubBytesIns_Inst_Sbox_0_L26}), .c ({new_AGEMA_signal_10224, new_AGEMA_signal_10223, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S2_U1 ( .a ({new_AGEMA_signal_9442, new_AGEMA_signal_9441, SubBytesIns_Inst_Sbox_0_L19}), .b ({new_AGEMA_signal_9822, new_AGEMA_signal_9821, SubBytesIns_Inst_Sbox_0_L28}), .c ({new_AGEMA_signal_10226, new_AGEMA_signal_10225, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S3_U1 ( .a ({new_AGEMA_signal_9432, new_AGEMA_signal_9431, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_9812, new_AGEMA_signal_9811, SubBytesIns_Inst_Sbox_0_L21}), .c ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S4_U1 ( .a ({new_AGEMA_signal_9810, new_AGEMA_signal_9809, SubBytesIns_Inst_Sbox_0_L20}), .b ({new_AGEMA_signal_9444, new_AGEMA_signal_9443, SubBytesIns_Inst_Sbox_0_L22}), .c ({new_AGEMA_signal_10230, new_AGEMA_signal_10229, MixColumnsInput[99]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S5_U1 ( .a ({new_AGEMA_signal_9816, new_AGEMA_signal_9815, SubBytesIns_Inst_Sbox_0_L25}), .b ({new_AGEMA_signal_9824, new_AGEMA_signal_9823, SubBytesIns_Inst_Sbox_0_L29}), .c ({new_AGEMA_signal_10232, new_AGEMA_signal_10231, MixColumnsInput[98]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S6_U1 ( .a ({new_AGEMA_signal_9806, new_AGEMA_signal_9805, SubBytesIns_Inst_Sbox_0_L13}), .b ({new_AGEMA_signal_9820, new_AGEMA_signal_9819, SubBytesIns_Inst_Sbox_0_L27}), .c ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S7_U1 ( .a ({new_AGEMA_signal_9432, new_AGEMA_signal_9431, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_9446, new_AGEMA_signal_9445, SubBytesIns_Inst_Sbox_0_L23}), .c ({new_AGEMA_signal_9826, new_AGEMA_signal_9825, MixColumnsInput[96]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M46_U1 ( .a ({new_AGEMA_signal_8124, new_AGEMA_signal_8123, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_5798, new_AGEMA_signal_5797, SubBytesIns_Inst_Sbox_1_T6}), .clk (clk), .r ({Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({new_AGEMA_signal_8600, new_AGEMA_signal_8599, SubBytesIns_Inst_Sbox_1_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M47_U1 ( .a ({new_AGEMA_signal_7884, new_AGEMA_signal_7883, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_6168, new_AGEMA_signal_6167, SubBytesIns_Inst_Sbox_1_T8}), .clk (clk), .r ({Fresh[1019], Fresh[1018], Fresh[1017]}), .c ({new_AGEMA_signal_8126, new_AGEMA_signal_8125, SubBytesIns_Inst_Sbox_1_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M48_U1 ( .a ({new_AGEMA_signal_7882, new_AGEMA_signal_7881, SubBytesIns_Inst_Sbox_1_M39}), .b ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .clk (clk), .r ({Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({new_AGEMA_signal_8128, new_AGEMA_signal_8127, SubBytesIns_Inst_Sbox_1_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M49_U1 ( .a ({new_AGEMA_signal_8122, new_AGEMA_signal_8121, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_5806, new_AGEMA_signal_5805, SubBytesIns_Inst_Sbox_1_T16}), .clk (clk), .r ({Fresh[1025], Fresh[1024], Fresh[1023]}), .c ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, SubBytesIns_Inst_Sbox_1_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M50_U1 ( .a ({new_AGEMA_signal_7880, new_AGEMA_signal_7879, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_5800, new_AGEMA_signal_5799, SubBytesIns_Inst_Sbox_1_T9}), .clk (clk), .r ({Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({new_AGEMA_signal_8130, new_AGEMA_signal_8129, SubBytesIns_Inst_Sbox_1_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M51_U1 ( .a ({new_AGEMA_signal_7878, new_AGEMA_signal_7877, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_6174, new_AGEMA_signal_6173, SubBytesIns_Inst_Sbox_1_T17}), .clk (clk), .r ({Fresh[1031], Fresh[1030], Fresh[1029]}), .c ({new_AGEMA_signal_8132, new_AGEMA_signal_8131, SubBytesIns_Inst_Sbox_1_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M52_U1 ( .a ({new_AGEMA_signal_8120, new_AGEMA_signal_8119, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_5804, new_AGEMA_signal_5803, SubBytesIns_Inst_Sbox_1_T15}), .clk (clk), .r ({Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({new_AGEMA_signal_8604, new_AGEMA_signal_8603, SubBytesIns_Inst_Sbox_1_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M53_U1 ( .a ({new_AGEMA_signal_8598, new_AGEMA_signal_8597, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_5812, new_AGEMA_signal_5811, SubBytesIns_Inst_Sbox_1_T27}), .clk (clk), .r ({Fresh[1037], Fresh[1036], Fresh[1035]}), .c ({new_AGEMA_signal_9058, new_AGEMA_signal_9057, SubBytesIns_Inst_Sbox_1_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M54_U1 ( .a ({new_AGEMA_signal_8118, new_AGEMA_signal_8117, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_6170, new_AGEMA_signal_6169, SubBytesIns_Inst_Sbox_1_T10}), .clk (clk), .r ({Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({new_AGEMA_signal_8606, new_AGEMA_signal_8605, SubBytesIns_Inst_Sbox_1_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M55_U1 ( .a ({new_AGEMA_signal_8124, new_AGEMA_signal_8123, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_5802, new_AGEMA_signal_5801, SubBytesIns_Inst_Sbox_1_T13}), .clk (clk), .r ({Fresh[1043], Fresh[1042], Fresh[1041]}), .c ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, SubBytesIns_Inst_Sbox_1_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M56_U1 ( .a ({new_AGEMA_signal_7884, new_AGEMA_signal_7883, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_6178, new_AGEMA_signal_6177, SubBytesIns_Inst_Sbox_1_T23}), .clk (clk), .r ({Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({new_AGEMA_signal_8134, new_AGEMA_signal_8133, SubBytesIns_Inst_Sbox_1_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M57_U1 ( .a ({new_AGEMA_signal_7882, new_AGEMA_signal_7881, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_5808, new_AGEMA_signal_5807, SubBytesIns_Inst_Sbox_1_T19}), .clk (clk), .r ({Fresh[1049], Fresh[1048], Fresh[1047]}), .c ({new_AGEMA_signal_8136, new_AGEMA_signal_8135, SubBytesIns_Inst_Sbox_1_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M58_U1 ( .a ({new_AGEMA_signal_8122, new_AGEMA_signal_8121, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_5422, new_AGEMA_signal_5421, SubBytesIns_Inst_Sbox_1_T3}), .clk (clk), .r ({Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({new_AGEMA_signal_8610, new_AGEMA_signal_8609, SubBytesIns_Inst_Sbox_1_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M59_U1 ( .a ({new_AGEMA_signal_7880, new_AGEMA_signal_7879, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_5810, new_AGEMA_signal_5809, SubBytesIns_Inst_Sbox_1_T22}), .clk (clk), .r ({Fresh[1055], Fresh[1054], Fresh[1053]}), .c ({new_AGEMA_signal_8138, new_AGEMA_signal_8137, SubBytesIns_Inst_Sbox_1_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M60_U1 ( .a ({new_AGEMA_signal_7878, new_AGEMA_signal_7877, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_6176, new_AGEMA_signal_6175, SubBytesIns_Inst_Sbox_1_T20}), .clk (clk), .r ({Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({new_AGEMA_signal_8140, new_AGEMA_signal_8139, SubBytesIns_Inst_Sbox_1_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M61_U1 ( .a ({new_AGEMA_signal_8120, new_AGEMA_signal_8119, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_5418, new_AGEMA_signal_5417, SubBytesIns_Inst_Sbox_1_T1}), .clk (clk), .r ({Fresh[1061], Fresh[1060], Fresh[1059]}), .c ({new_AGEMA_signal_8612, new_AGEMA_signal_8611, SubBytesIns_Inst_Sbox_1_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M62_U1 ( .a ({new_AGEMA_signal_8598, new_AGEMA_signal_8597, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_5424, new_AGEMA_signal_5423, SubBytesIns_Inst_Sbox_1_T4}), .clk (clk), .r ({Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({new_AGEMA_signal_9060, new_AGEMA_signal_9059, SubBytesIns_Inst_Sbox_1_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M63_U1 ( .a ({new_AGEMA_signal_8118, new_AGEMA_signal_8117, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_5420, new_AGEMA_signal_5419, SubBytesIns_Inst_Sbox_1_T2}), .clk (clk), .r ({Fresh[1067], Fresh[1066], Fresh[1065]}), .c ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, SubBytesIns_Inst_Sbox_1_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L0_U1 ( .a ({new_AGEMA_signal_8612, new_AGEMA_signal_8611, SubBytesIns_Inst_Sbox_1_M61}), .b ({new_AGEMA_signal_9060, new_AGEMA_signal_9059, SubBytesIns_Inst_Sbox_1_M62}), .c ({new_AGEMA_signal_9448, new_AGEMA_signal_9447, SubBytesIns_Inst_Sbox_1_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L1_U1 ( .a ({new_AGEMA_signal_8130, new_AGEMA_signal_8129, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_8134, new_AGEMA_signal_8133, SubBytesIns_Inst_Sbox_1_M56}), .c ({new_AGEMA_signal_8616, new_AGEMA_signal_8615, SubBytesIns_Inst_Sbox_1_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L2_U1 ( .a ({new_AGEMA_signal_8600, new_AGEMA_signal_8599, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_8128, new_AGEMA_signal_8127, SubBytesIns_Inst_Sbox_1_M48}), .c ({new_AGEMA_signal_9062, new_AGEMA_signal_9061, SubBytesIns_Inst_Sbox_1_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L3_U1 ( .a ({new_AGEMA_signal_8126, new_AGEMA_signal_8125, SubBytesIns_Inst_Sbox_1_M47}), .b ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, SubBytesIns_Inst_Sbox_1_M55}), .c ({new_AGEMA_signal_9064, new_AGEMA_signal_9063, SubBytesIns_Inst_Sbox_1_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L4_U1 ( .a ({new_AGEMA_signal_8606, new_AGEMA_signal_8605, SubBytesIns_Inst_Sbox_1_M54}), .b ({new_AGEMA_signal_8610, new_AGEMA_signal_8609, SubBytesIns_Inst_Sbox_1_M58}), .c ({new_AGEMA_signal_9066, new_AGEMA_signal_9065, SubBytesIns_Inst_Sbox_1_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L5_U1 ( .a ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, SubBytesIns_Inst_Sbox_1_M49}), .b ({new_AGEMA_signal_8612, new_AGEMA_signal_8611, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_9068, new_AGEMA_signal_9067, SubBytesIns_Inst_Sbox_1_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L6_U1 ( .a ({new_AGEMA_signal_9060, new_AGEMA_signal_9059, SubBytesIns_Inst_Sbox_1_M62}), .b ({new_AGEMA_signal_9068, new_AGEMA_signal_9067, SubBytesIns_Inst_Sbox_1_L5}), .c ({new_AGEMA_signal_9450, new_AGEMA_signal_9449, SubBytesIns_Inst_Sbox_1_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L7_U1 ( .a ({new_AGEMA_signal_8600, new_AGEMA_signal_8599, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_9064, new_AGEMA_signal_9063, SubBytesIns_Inst_Sbox_1_L3}), .c ({new_AGEMA_signal_9452, new_AGEMA_signal_9451, SubBytesIns_Inst_Sbox_1_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L8_U1 ( .a ({new_AGEMA_signal_8132, new_AGEMA_signal_8131, SubBytesIns_Inst_Sbox_1_M51}), .b ({new_AGEMA_signal_8138, new_AGEMA_signal_8137, SubBytesIns_Inst_Sbox_1_M59}), .c ({new_AGEMA_signal_8618, new_AGEMA_signal_8617, SubBytesIns_Inst_Sbox_1_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L9_U1 ( .a ({new_AGEMA_signal_8604, new_AGEMA_signal_8603, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_9058, new_AGEMA_signal_9057, SubBytesIns_Inst_Sbox_1_M53}), .c ({new_AGEMA_signal_9454, new_AGEMA_signal_9453, SubBytesIns_Inst_Sbox_1_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L10_U1 ( .a ({new_AGEMA_signal_9058, new_AGEMA_signal_9057, SubBytesIns_Inst_Sbox_1_M53}), .b ({new_AGEMA_signal_9066, new_AGEMA_signal_9065, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_9456, new_AGEMA_signal_9455, SubBytesIns_Inst_Sbox_1_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L11_U1 ( .a ({new_AGEMA_signal_8140, new_AGEMA_signal_8139, SubBytesIns_Inst_Sbox_1_M60}), .b ({new_AGEMA_signal_9062, new_AGEMA_signal_9061, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_9458, new_AGEMA_signal_9457, SubBytesIns_Inst_Sbox_1_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L12_U1 ( .a ({new_AGEMA_signal_8128, new_AGEMA_signal_8127, SubBytesIns_Inst_Sbox_1_M48}), .b ({new_AGEMA_signal_8132, new_AGEMA_signal_8131, SubBytesIns_Inst_Sbox_1_M51}), .c ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, SubBytesIns_Inst_Sbox_1_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L13_U1 ( .a ({new_AGEMA_signal_8130, new_AGEMA_signal_8129, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_9448, new_AGEMA_signal_9447, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_9828, new_AGEMA_signal_9827, SubBytesIns_Inst_Sbox_1_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L14_U1 ( .a ({new_AGEMA_signal_8604, new_AGEMA_signal_8603, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_8612, new_AGEMA_signal_8611, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_9070, new_AGEMA_signal_9069, SubBytesIns_Inst_Sbox_1_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L15_U1 ( .a ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, SubBytesIns_Inst_Sbox_1_M55}), .b ({new_AGEMA_signal_8616, new_AGEMA_signal_8615, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_9072, new_AGEMA_signal_9071, SubBytesIns_Inst_Sbox_1_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L16_U1 ( .a ({new_AGEMA_signal_8134, new_AGEMA_signal_8133, SubBytesIns_Inst_Sbox_1_M56}), .b ({new_AGEMA_signal_9448, new_AGEMA_signal_9447, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_9830, new_AGEMA_signal_9829, SubBytesIns_Inst_Sbox_1_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L17_U1 ( .a ({new_AGEMA_signal_8136, new_AGEMA_signal_8135, SubBytesIns_Inst_Sbox_1_M57}), .b ({new_AGEMA_signal_8616, new_AGEMA_signal_8615, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_9074, new_AGEMA_signal_9073, SubBytesIns_Inst_Sbox_1_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L18_U1 ( .a ({new_AGEMA_signal_8610, new_AGEMA_signal_8609, SubBytesIns_Inst_Sbox_1_M58}), .b ({new_AGEMA_signal_8618, new_AGEMA_signal_8617, SubBytesIns_Inst_Sbox_1_L8}), .c ({new_AGEMA_signal_9076, new_AGEMA_signal_9075, SubBytesIns_Inst_Sbox_1_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L19_U1 ( .a ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, SubBytesIns_Inst_Sbox_1_M63}), .b ({new_AGEMA_signal_9066, new_AGEMA_signal_9065, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_9460, new_AGEMA_signal_9459, SubBytesIns_Inst_Sbox_1_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L20_U1 ( .a ({new_AGEMA_signal_9448, new_AGEMA_signal_9447, SubBytesIns_Inst_Sbox_1_L0}), .b ({new_AGEMA_signal_8616, new_AGEMA_signal_8615, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_9832, new_AGEMA_signal_9831, SubBytesIns_Inst_Sbox_1_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L21_U1 ( .a ({new_AGEMA_signal_8616, new_AGEMA_signal_8615, SubBytesIns_Inst_Sbox_1_L1}), .b ({new_AGEMA_signal_9452, new_AGEMA_signal_9451, SubBytesIns_Inst_Sbox_1_L7}), .c ({new_AGEMA_signal_9834, new_AGEMA_signal_9833, SubBytesIns_Inst_Sbox_1_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L22_U1 ( .a ({new_AGEMA_signal_9064, new_AGEMA_signal_9063, SubBytesIns_Inst_Sbox_1_L3}), .b ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, SubBytesIns_Inst_Sbox_1_L12}), .c ({new_AGEMA_signal_9462, new_AGEMA_signal_9461, SubBytesIns_Inst_Sbox_1_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L23_U1 ( .a ({new_AGEMA_signal_9076, new_AGEMA_signal_9075, SubBytesIns_Inst_Sbox_1_L18}), .b ({new_AGEMA_signal_9062, new_AGEMA_signal_9061, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_9464, new_AGEMA_signal_9463, SubBytesIns_Inst_Sbox_1_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L24_U1 ( .a ({new_AGEMA_signal_9072, new_AGEMA_signal_9071, SubBytesIns_Inst_Sbox_1_L15}), .b ({new_AGEMA_signal_9454, new_AGEMA_signal_9453, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_9836, new_AGEMA_signal_9835, SubBytesIns_Inst_Sbox_1_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L25_U1 ( .a ({new_AGEMA_signal_9450, new_AGEMA_signal_9449, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_9456, new_AGEMA_signal_9455, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_9838, new_AGEMA_signal_9837, SubBytesIns_Inst_Sbox_1_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L26_U1 ( .a ({new_AGEMA_signal_9452, new_AGEMA_signal_9451, SubBytesIns_Inst_Sbox_1_L7}), .b ({new_AGEMA_signal_9454, new_AGEMA_signal_9453, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_9840, new_AGEMA_signal_9839, SubBytesIns_Inst_Sbox_1_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L27_U1 ( .a ({new_AGEMA_signal_8618, new_AGEMA_signal_8617, SubBytesIns_Inst_Sbox_1_L8}), .b ({new_AGEMA_signal_9456, new_AGEMA_signal_9455, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_9842, new_AGEMA_signal_9841, SubBytesIns_Inst_Sbox_1_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L28_U1 ( .a ({new_AGEMA_signal_9458, new_AGEMA_signal_9457, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_9070, new_AGEMA_signal_9069, SubBytesIns_Inst_Sbox_1_L14}), .c ({new_AGEMA_signal_9844, new_AGEMA_signal_9843, SubBytesIns_Inst_Sbox_1_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L29_U1 ( .a ({new_AGEMA_signal_9458, new_AGEMA_signal_9457, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_9074, new_AGEMA_signal_9073, SubBytesIns_Inst_Sbox_1_L17}), .c ({new_AGEMA_signal_9846, new_AGEMA_signal_9845, SubBytesIns_Inst_Sbox_1_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S0_U1 ( .a ({new_AGEMA_signal_9450, new_AGEMA_signal_9449, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_9836, new_AGEMA_signal_9835, SubBytesIns_Inst_Sbox_1_L24}), .c ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S1_U1 ( .a ({new_AGEMA_signal_9830, new_AGEMA_signal_9829, SubBytesIns_Inst_Sbox_1_L16}), .b ({new_AGEMA_signal_9840, new_AGEMA_signal_9839, SubBytesIns_Inst_Sbox_1_L26}), .c ({new_AGEMA_signal_10238, new_AGEMA_signal_10237, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S2_U1 ( .a ({new_AGEMA_signal_9460, new_AGEMA_signal_9459, SubBytesIns_Inst_Sbox_1_L19}), .b ({new_AGEMA_signal_9844, new_AGEMA_signal_9843, SubBytesIns_Inst_Sbox_1_L28}), .c ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S3_U1 ( .a ({new_AGEMA_signal_9450, new_AGEMA_signal_9449, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_9834, new_AGEMA_signal_9833, SubBytesIns_Inst_Sbox_1_L21}), .c ({new_AGEMA_signal_10242, new_AGEMA_signal_10241, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S4_U1 ( .a ({new_AGEMA_signal_9832, new_AGEMA_signal_9831, SubBytesIns_Inst_Sbox_1_L20}), .b ({new_AGEMA_signal_9462, new_AGEMA_signal_9461, SubBytesIns_Inst_Sbox_1_L22}), .c ({new_AGEMA_signal_10244, new_AGEMA_signal_10243, MixColumnsInput[75]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S5_U1 ( .a ({new_AGEMA_signal_9838, new_AGEMA_signal_9837, SubBytesIns_Inst_Sbox_1_L25}), .b ({new_AGEMA_signal_9846, new_AGEMA_signal_9845, SubBytesIns_Inst_Sbox_1_L29}), .c ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, MixColumnsInput[74]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S6_U1 ( .a ({new_AGEMA_signal_9828, new_AGEMA_signal_9827, SubBytesIns_Inst_Sbox_1_L13}), .b ({new_AGEMA_signal_9842, new_AGEMA_signal_9841, SubBytesIns_Inst_Sbox_1_L27}), .c ({new_AGEMA_signal_10248, new_AGEMA_signal_10247, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S7_U1 ( .a ({new_AGEMA_signal_9450, new_AGEMA_signal_9449, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_9464, new_AGEMA_signal_9463, SubBytesIns_Inst_Sbox_1_L23}), .c ({new_AGEMA_signal_9848, new_AGEMA_signal_9847, MixColumnsInput[72]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M46_U1 ( .a ({new_AGEMA_signal_8148, new_AGEMA_signal_8147, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_5814, new_AGEMA_signal_5813, SubBytesIns_Inst_Sbox_2_T6}), .clk (clk), .r ({Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({new_AGEMA_signal_8624, new_AGEMA_signal_8623, SubBytesIns_Inst_Sbox_2_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M47_U1 ( .a ({new_AGEMA_signal_7892, new_AGEMA_signal_7891, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_6194, new_AGEMA_signal_6193, SubBytesIns_Inst_Sbox_2_T8}), .clk (clk), .r ({Fresh[1073], Fresh[1072], Fresh[1071]}), .c ({new_AGEMA_signal_8150, new_AGEMA_signal_8149, SubBytesIns_Inst_Sbox_2_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M48_U1 ( .a ({new_AGEMA_signal_7890, new_AGEMA_signal_7889, SubBytesIns_Inst_Sbox_2_M39}), .b ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .clk (clk), .r ({Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({new_AGEMA_signal_8152, new_AGEMA_signal_8151, SubBytesIns_Inst_Sbox_2_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M49_U1 ( .a ({new_AGEMA_signal_8146, new_AGEMA_signal_8145, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_2_T16}), .clk (clk), .r ({Fresh[1079], Fresh[1078], Fresh[1077]}), .c ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, SubBytesIns_Inst_Sbox_2_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M50_U1 ( .a ({new_AGEMA_signal_7888, new_AGEMA_signal_7887, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_5816, new_AGEMA_signal_5815, SubBytesIns_Inst_Sbox_2_T9}), .clk (clk), .r ({Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({new_AGEMA_signal_8154, new_AGEMA_signal_8153, SubBytesIns_Inst_Sbox_2_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M51_U1 ( .a ({new_AGEMA_signal_7886, new_AGEMA_signal_7885, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_6200, new_AGEMA_signal_6199, SubBytesIns_Inst_Sbox_2_T17}), .clk (clk), .r ({Fresh[1085], Fresh[1084], Fresh[1083]}), .c ({new_AGEMA_signal_8156, new_AGEMA_signal_8155, SubBytesIns_Inst_Sbox_2_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M52_U1 ( .a ({new_AGEMA_signal_8144, new_AGEMA_signal_8143, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_5820, new_AGEMA_signal_5819, SubBytesIns_Inst_Sbox_2_T15}), .clk (clk), .r ({Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({new_AGEMA_signal_8628, new_AGEMA_signal_8627, SubBytesIns_Inst_Sbox_2_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M53_U1 ( .a ({new_AGEMA_signal_8622, new_AGEMA_signal_8621, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_5828, new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_2_T27}), .clk (clk), .r ({Fresh[1091], Fresh[1090], Fresh[1089]}), .c ({new_AGEMA_signal_9078, new_AGEMA_signal_9077, SubBytesIns_Inst_Sbox_2_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M54_U1 ( .a ({new_AGEMA_signal_8142, new_AGEMA_signal_8141, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_6196, new_AGEMA_signal_6195, SubBytesIns_Inst_Sbox_2_T10}), .clk (clk), .r ({Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({new_AGEMA_signal_8630, new_AGEMA_signal_8629, SubBytesIns_Inst_Sbox_2_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M55_U1 ( .a ({new_AGEMA_signal_8148, new_AGEMA_signal_8147, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_5818, new_AGEMA_signal_5817, SubBytesIns_Inst_Sbox_2_T13}), .clk (clk), .r ({Fresh[1097], Fresh[1096], Fresh[1095]}), .c ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, SubBytesIns_Inst_Sbox_2_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M56_U1 ( .a ({new_AGEMA_signal_7892, new_AGEMA_signal_7891, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_6204, new_AGEMA_signal_6203, SubBytesIns_Inst_Sbox_2_T23}), .clk (clk), .r ({Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({new_AGEMA_signal_8158, new_AGEMA_signal_8157, SubBytesIns_Inst_Sbox_2_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M57_U1 ( .a ({new_AGEMA_signal_7890, new_AGEMA_signal_7889, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_5824, new_AGEMA_signal_5823, SubBytesIns_Inst_Sbox_2_T19}), .clk (clk), .r ({Fresh[1103], Fresh[1102], Fresh[1101]}), .c ({new_AGEMA_signal_8160, new_AGEMA_signal_8159, SubBytesIns_Inst_Sbox_2_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M58_U1 ( .a ({new_AGEMA_signal_8146, new_AGEMA_signal_8145, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_5442, new_AGEMA_signal_5441, SubBytesIns_Inst_Sbox_2_T3}), .clk (clk), .r ({Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({new_AGEMA_signal_8634, new_AGEMA_signal_8633, SubBytesIns_Inst_Sbox_2_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M59_U1 ( .a ({new_AGEMA_signal_7888, new_AGEMA_signal_7887, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_5826, new_AGEMA_signal_5825, SubBytesIns_Inst_Sbox_2_T22}), .clk (clk), .r ({Fresh[1109], Fresh[1108], Fresh[1107]}), .c ({new_AGEMA_signal_8162, new_AGEMA_signal_8161, SubBytesIns_Inst_Sbox_2_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M60_U1 ( .a ({new_AGEMA_signal_7886, new_AGEMA_signal_7885, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_6202, new_AGEMA_signal_6201, SubBytesIns_Inst_Sbox_2_T20}), .clk (clk), .r ({Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({new_AGEMA_signal_8164, new_AGEMA_signal_8163, SubBytesIns_Inst_Sbox_2_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M61_U1 ( .a ({new_AGEMA_signal_8144, new_AGEMA_signal_8143, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_5438, new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_2_T1}), .clk (clk), .r ({Fresh[1115], Fresh[1114], Fresh[1113]}), .c ({new_AGEMA_signal_8636, new_AGEMA_signal_8635, SubBytesIns_Inst_Sbox_2_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M62_U1 ( .a ({new_AGEMA_signal_8622, new_AGEMA_signal_8621, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_5444, new_AGEMA_signal_5443, SubBytesIns_Inst_Sbox_2_T4}), .clk (clk), .r ({Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({new_AGEMA_signal_9080, new_AGEMA_signal_9079, SubBytesIns_Inst_Sbox_2_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M63_U1 ( .a ({new_AGEMA_signal_8142, new_AGEMA_signal_8141, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_5440, new_AGEMA_signal_5439, SubBytesIns_Inst_Sbox_2_T2}), .clk (clk), .r ({Fresh[1121], Fresh[1120], Fresh[1119]}), .c ({new_AGEMA_signal_8638, new_AGEMA_signal_8637, SubBytesIns_Inst_Sbox_2_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L0_U1 ( .a ({new_AGEMA_signal_8636, new_AGEMA_signal_8635, SubBytesIns_Inst_Sbox_2_M61}), .b ({new_AGEMA_signal_9080, new_AGEMA_signal_9079, SubBytesIns_Inst_Sbox_2_M62}), .c ({new_AGEMA_signal_9466, new_AGEMA_signal_9465, SubBytesIns_Inst_Sbox_2_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L1_U1 ( .a ({new_AGEMA_signal_8154, new_AGEMA_signal_8153, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_8158, new_AGEMA_signal_8157, SubBytesIns_Inst_Sbox_2_M56}), .c ({new_AGEMA_signal_8640, new_AGEMA_signal_8639, SubBytesIns_Inst_Sbox_2_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L2_U1 ( .a ({new_AGEMA_signal_8624, new_AGEMA_signal_8623, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_8152, new_AGEMA_signal_8151, SubBytesIns_Inst_Sbox_2_M48}), .c ({new_AGEMA_signal_9082, new_AGEMA_signal_9081, SubBytesIns_Inst_Sbox_2_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L3_U1 ( .a ({new_AGEMA_signal_8150, new_AGEMA_signal_8149, SubBytesIns_Inst_Sbox_2_M47}), .b ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, SubBytesIns_Inst_Sbox_2_M55}), .c ({new_AGEMA_signal_9084, new_AGEMA_signal_9083, SubBytesIns_Inst_Sbox_2_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L4_U1 ( .a ({new_AGEMA_signal_8630, new_AGEMA_signal_8629, SubBytesIns_Inst_Sbox_2_M54}), .b ({new_AGEMA_signal_8634, new_AGEMA_signal_8633, SubBytesIns_Inst_Sbox_2_M58}), .c ({new_AGEMA_signal_9086, new_AGEMA_signal_9085, SubBytesIns_Inst_Sbox_2_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L5_U1 ( .a ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, SubBytesIns_Inst_Sbox_2_M49}), .b ({new_AGEMA_signal_8636, new_AGEMA_signal_8635, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_9088, new_AGEMA_signal_9087, SubBytesIns_Inst_Sbox_2_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L6_U1 ( .a ({new_AGEMA_signal_9080, new_AGEMA_signal_9079, SubBytesIns_Inst_Sbox_2_M62}), .b ({new_AGEMA_signal_9088, new_AGEMA_signal_9087, SubBytesIns_Inst_Sbox_2_L5}), .c ({new_AGEMA_signal_9468, new_AGEMA_signal_9467, SubBytesIns_Inst_Sbox_2_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L7_U1 ( .a ({new_AGEMA_signal_8624, new_AGEMA_signal_8623, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_9084, new_AGEMA_signal_9083, SubBytesIns_Inst_Sbox_2_L3}), .c ({new_AGEMA_signal_9470, new_AGEMA_signal_9469, SubBytesIns_Inst_Sbox_2_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L8_U1 ( .a ({new_AGEMA_signal_8156, new_AGEMA_signal_8155, SubBytesIns_Inst_Sbox_2_M51}), .b ({new_AGEMA_signal_8162, new_AGEMA_signal_8161, SubBytesIns_Inst_Sbox_2_M59}), .c ({new_AGEMA_signal_8642, new_AGEMA_signal_8641, SubBytesIns_Inst_Sbox_2_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L9_U1 ( .a ({new_AGEMA_signal_8628, new_AGEMA_signal_8627, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_9078, new_AGEMA_signal_9077, SubBytesIns_Inst_Sbox_2_M53}), .c ({new_AGEMA_signal_9472, new_AGEMA_signal_9471, SubBytesIns_Inst_Sbox_2_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L10_U1 ( .a ({new_AGEMA_signal_9078, new_AGEMA_signal_9077, SubBytesIns_Inst_Sbox_2_M53}), .b ({new_AGEMA_signal_9086, new_AGEMA_signal_9085, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_9474, new_AGEMA_signal_9473, SubBytesIns_Inst_Sbox_2_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L11_U1 ( .a ({new_AGEMA_signal_8164, new_AGEMA_signal_8163, SubBytesIns_Inst_Sbox_2_M60}), .b ({new_AGEMA_signal_9082, new_AGEMA_signal_9081, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_9476, new_AGEMA_signal_9475, SubBytesIns_Inst_Sbox_2_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L12_U1 ( .a ({new_AGEMA_signal_8152, new_AGEMA_signal_8151, SubBytesIns_Inst_Sbox_2_M48}), .b ({new_AGEMA_signal_8156, new_AGEMA_signal_8155, SubBytesIns_Inst_Sbox_2_M51}), .c ({new_AGEMA_signal_8644, new_AGEMA_signal_8643, SubBytesIns_Inst_Sbox_2_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L13_U1 ( .a ({new_AGEMA_signal_8154, new_AGEMA_signal_8153, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_9466, new_AGEMA_signal_9465, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_9850, new_AGEMA_signal_9849, SubBytesIns_Inst_Sbox_2_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L14_U1 ( .a ({new_AGEMA_signal_8628, new_AGEMA_signal_8627, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_8636, new_AGEMA_signal_8635, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_9090, new_AGEMA_signal_9089, SubBytesIns_Inst_Sbox_2_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L15_U1 ( .a ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, SubBytesIns_Inst_Sbox_2_M55}), .b ({new_AGEMA_signal_8640, new_AGEMA_signal_8639, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_9092, new_AGEMA_signal_9091, SubBytesIns_Inst_Sbox_2_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L16_U1 ( .a ({new_AGEMA_signal_8158, new_AGEMA_signal_8157, SubBytesIns_Inst_Sbox_2_M56}), .b ({new_AGEMA_signal_9466, new_AGEMA_signal_9465, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_9852, new_AGEMA_signal_9851, SubBytesIns_Inst_Sbox_2_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L17_U1 ( .a ({new_AGEMA_signal_8160, new_AGEMA_signal_8159, SubBytesIns_Inst_Sbox_2_M57}), .b ({new_AGEMA_signal_8640, new_AGEMA_signal_8639, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_9094, new_AGEMA_signal_9093, SubBytesIns_Inst_Sbox_2_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L18_U1 ( .a ({new_AGEMA_signal_8634, new_AGEMA_signal_8633, SubBytesIns_Inst_Sbox_2_M58}), .b ({new_AGEMA_signal_8642, new_AGEMA_signal_8641, SubBytesIns_Inst_Sbox_2_L8}), .c ({new_AGEMA_signal_9096, new_AGEMA_signal_9095, SubBytesIns_Inst_Sbox_2_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L19_U1 ( .a ({new_AGEMA_signal_8638, new_AGEMA_signal_8637, SubBytesIns_Inst_Sbox_2_M63}), .b ({new_AGEMA_signal_9086, new_AGEMA_signal_9085, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_9478, new_AGEMA_signal_9477, SubBytesIns_Inst_Sbox_2_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L20_U1 ( .a ({new_AGEMA_signal_9466, new_AGEMA_signal_9465, SubBytesIns_Inst_Sbox_2_L0}), .b ({new_AGEMA_signal_8640, new_AGEMA_signal_8639, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_9854, new_AGEMA_signal_9853, SubBytesIns_Inst_Sbox_2_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L21_U1 ( .a ({new_AGEMA_signal_8640, new_AGEMA_signal_8639, SubBytesIns_Inst_Sbox_2_L1}), .b ({new_AGEMA_signal_9470, new_AGEMA_signal_9469, SubBytesIns_Inst_Sbox_2_L7}), .c ({new_AGEMA_signal_9856, new_AGEMA_signal_9855, SubBytesIns_Inst_Sbox_2_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L22_U1 ( .a ({new_AGEMA_signal_9084, new_AGEMA_signal_9083, SubBytesIns_Inst_Sbox_2_L3}), .b ({new_AGEMA_signal_8644, new_AGEMA_signal_8643, SubBytesIns_Inst_Sbox_2_L12}), .c ({new_AGEMA_signal_9480, new_AGEMA_signal_9479, SubBytesIns_Inst_Sbox_2_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L23_U1 ( .a ({new_AGEMA_signal_9096, new_AGEMA_signal_9095, SubBytesIns_Inst_Sbox_2_L18}), .b ({new_AGEMA_signal_9082, new_AGEMA_signal_9081, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_9482, new_AGEMA_signal_9481, SubBytesIns_Inst_Sbox_2_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L24_U1 ( .a ({new_AGEMA_signal_9092, new_AGEMA_signal_9091, SubBytesIns_Inst_Sbox_2_L15}), .b ({new_AGEMA_signal_9472, new_AGEMA_signal_9471, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_9858, new_AGEMA_signal_9857, SubBytesIns_Inst_Sbox_2_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L25_U1 ( .a ({new_AGEMA_signal_9468, new_AGEMA_signal_9467, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_9474, new_AGEMA_signal_9473, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_9860, new_AGEMA_signal_9859, SubBytesIns_Inst_Sbox_2_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L26_U1 ( .a ({new_AGEMA_signal_9470, new_AGEMA_signal_9469, SubBytesIns_Inst_Sbox_2_L7}), .b ({new_AGEMA_signal_9472, new_AGEMA_signal_9471, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_9862, new_AGEMA_signal_9861, SubBytesIns_Inst_Sbox_2_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L27_U1 ( .a ({new_AGEMA_signal_8642, new_AGEMA_signal_8641, SubBytesIns_Inst_Sbox_2_L8}), .b ({new_AGEMA_signal_9474, new_AGEMA_signal_9473, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_9864, new_AGEMA_signal_9863, SubBytesIns_Inst_Sbox_2_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L28_U1 ( .a ({new_AGEMA_signal_9476, new_AGEMA_signal_9475, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_9090, new_AGEMA_signal_9089, SubBytesIns_Inst_Sbox_2_L14}), .c ({new_AGEMA_signal_9866, new_AGEMA_signal_9865, SubBytesIns_Inst_Sbox_2_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L29_U1 ( .a ({new_AGEMA_signal_9476, new_AGEMA_signal_9475, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_9094, new_AGEMA_signal_9093, SubBytesIns_Inst_Sbox_2_L17}), .c ({new_AGEMA_signal_9868, new_AGEMA_signal_9867, SubBytesIns_Inst_Sbox_2_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S0_U1 ( .a ({new_AGEMA_signal_9468, new_AGEMA_signal_9467, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_9858, new_AGEMA_signal_9857, SubBytesIns_Inst_Sbox_2_L24}), .c ({new_AGEMA_signal_10250, new_AGEMA_signal_10249, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S1_U1 ( .a ({new_AGEMA_signal_9852, new_AGEMA_signal_9851, SubBytesIns_Inst_Sbox_2_L16}), .b ({new_AGEMA_signal_9862, new_AGEMA_signal_9861, SubBytesIns_Inst_Sbox_2_L26}), .c ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S2_U1 ( .a ({new_AGEMA_signal_9478, new_AGEMA_signal_9477, SubBytesIns_Inst_Sbox_2_L19}), .b ({new_AGEMA_signal_9866, new_AGEMA_signal_9865, SubBytesIns_Inst_Sbox_2_L28}), .c ({new_AGEMA_signal_10254, new_AGEMA_signal_10253, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S3_U1 ( .a ({new_AGEMA_signal_9468, new_AGEMA_signal_9467, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_9856, new_AGEMA_signal_9855, SubBytesIns_Inst_Sbox_2_L21}), .c ({new_AGEMA_signal_10256, new_AGEMA_signal_10255, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S4_U1 ( .a ({new_AGEMA_signal_9854, new_AGEMA_signal_9853, SubBytesIns_Inst_Sbox_2_L20}), .b ({new_AGEMA_signal_9480, new_AGEMA_signal_9479, SubBytesIns_Inst_Sbox_2_L22}), .c ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, MixColumnsInput[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S5_U1 ( .a ({new_AGEMA_signal_9860, new_AGEMA_signal_9859, SubBytesIns_Inst_Sbox_2_L25}), .b ({new_AGEMA_signal_9868, new_AGEMA_signal_9867, SubBytesIns_Inst_Sbox_2_L29}), .c ({new_AGEMA_signal_10260, new_AGEMA_signal_10259, MixColumnsInput[50]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S6_U1 ( .a ({new_AGEMA_signal_9850, new_AGEMA_signal_9849, SubBytesIns_Inst_Sbox_2_L13}), .b ({new_AGEMA_signal_9864, new_AGEMA_signal_9863, SubBytesIns_Inst_Sbox_2_L27}), .c ({new_AGEMA_signal_10262, new_AGEMA_signal_10261, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S7_U1 ( .a ({new_AGEMA_signal_9468, new_AGEMA_signal_9467, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_9482, new_AGEMA_signal_9481, SubBytesIns_Inst_Sbox_2_L23}), .c ({new_AGEMA_signal_9870, new_AGEMA_signal_9869, MixColumnsInput[48]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M46_U1 ( .a ({new_AGEMA_signal_8172, new_AGEMA_signal_8171, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, SubBytesIns_Inst_Sbox_3_T6}), .clk (clk), .r ({Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({new_AGEMA_signal_8648, new_AGEMA_signal_8647, SubBytesIns_Inst_Sbox_3_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M47_U1 ( .a ({new_AGEMA_signal_7900, new_AGEMA_signal_7899, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_6220, new_AGEMA_signal_6219, SubBytesIns_Inst_Sbox_3_T8}), .clk (clk), .r ({Fresh[1127], Fresh[1126], Fresh[1125]}), .c ({new_AGEMA_signal_8174, new_AGEMA_signal_8173, SubBytesIns_Inst_Sbox_3_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M48_U1 ( .a ({new_AGEMA_signal_7898, new_AGEMA_signal_7897, SubBytesIns_Inst_Sbox_3_M39}), .b ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .clk (clk), .r ({Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({new_AGEMA_signal_8176, new_AGEMA_signal_8175, SubBytesIns_Inst_Sbox_3_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M49_U1 ( .a ({new_AGEMA_signal_8170, new_AGEMA_signal_8169, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, SubBytesIns_Inst_Sbox_3_T16}), .clk (clk), .r ({Fresh[1133], Fresh[1132], Fresh[1131]}), .c ({new_AGEMA_signal_8650, new_AGEMA_signal_8649, SubBytesIns_Inst_Sbox_3_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M50_U1 ( .a ({new_AGEMA_signal_7896, new_AGEMA_signal_7895, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_5832, new_AGEMA_signal_5831, SubBytesIns_Inst_Sbox_3_T9}), .clk (clk), .r ({Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({new_AGEMA_signal_8178, new_AGEMA_signal_8177, SubBytesIns_Inst_Sbox_3_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M51_U1 ( .a ({new_AGEMA_signal_7894, new_AGEMA_signal_7893, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_6226, new_AGEMA_signal_6225, SubBytesIns_Inst_Sbox_3_T17}), .clk (clk), .r ({Fresh[1139], Fresh[1138], Fresh[1137]}), .c ({new_AGEMA_signal_8180, new_AGEMA_signal_8179, SubBytesIns_Inst_Sbox_3_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M52_U1 ( .a ({new_AGEMA_signal_8168, new_AGEMA_signal_8167, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_5836, new_AGEMA_signal_5835, SubBytesIns_Inst_Sbox_3_T15}), .clk (clk), .r ({Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({new_AGEMA_signal_8652, new_AGEMA_signal_8651, SubBytesIns_Inst_Sbox_3_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M53_U1 ( .a ({new_AGEMA_signal_8646, new_AGEMA_signal_8645, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_5844, new_AGEMA_signal_5843, SubBytesIns_Inst_Sbox_3_T27}), .clk (clk), .r ({Fresh[1145], Fresh[1144], Fresh[1143]}), .c ({new_AGEMA_signal_9098, new_AGEMA_signal_9097, SubBytesIns_Inst_Sbox_3_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M54_U1 ( .a ({new_AGEMA_signal_8166, new_AGEMA_signal_8165, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_6222, new_AGEMA_signal_6221, SubBytesIns_Inst_Sbox_3_T10}), .clk (clk), .r ({Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({new_AGEMA_signal_8654, new_AGEMA_signal_8653, SubBytesIns_Inst_Sbox_3_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M55_U1 ( .a ({new_AGEMA_signal_8172, new_AGEMA_signal_8171, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_5834, new_AGEMA_signal_5833, SubBytesIns_Inst_Sbox_3_T13}), .clk (clk), .r ({Fresh[1151], Fresh[1150], Fresh[1149]}), .c ({new_AGEMA_signal_8656, new_AGEMA_signal_8655, SubBytesIns_Inst_Sbox_3_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M56_U1 ( .a ({new_AGEMA_signal_7900, new_AGEMA_signal_7899, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_6230, new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_3_T23}), .clk (clk), .r ({Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({new_AGEMA_signal_8182, new_AGEMA_signal_8181, SubBytesIns_Inst_Sbox_3_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M57_U1 ( .a ({new_AGEMA_signal_7898, new_AGEMA_signal_7897, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_5840, new_AGEMA_signal_5839, SubBytesIns_Inst_Sbox_3_T19}), .clk (clk), .r ({Fresh[1157], Fresh[1156], Fresh[1155]}), .c ({new_AGEMA_signal_8184, new_AGEMA_signal_8183, SubBytesIns_Inst_Sbox_3_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M58_U1 ( .a ({new_AGEMA_signal_8170, new_AGEMA_signal_8169, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_5462, new_AGEMA_signal_5461, SubBytesIns_Inst_Sbox_3_T3}), .clk (clk), .r ({Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({new_AGEMA_signal_8658, new_AGEMA_signal_8657, SubBytesIns_Inst_Sbox_3_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M59_U1 ( .a ({new_AGEMA_signal_7896, new_AGEMA_signal_7895, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_5842, new_AGEMA_signal_5841, SubBytesIns_Inst_Sbox_3_T22}), .clk (clk), .r ({Fresh[1163], Fresh[1162], Fresh[1161]}), .c ({new_AGEMA_signal_8186, new_AGEMA_signal_8185, SubBytesIns_Inst_Sbox_3_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M60_U1 ( .a ({new_AGEMA_signal_7894, new_AGEMA_signal_7893, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, SubBytesIns_Inst_Sbox_3_T20}), .clk (clk), .r ({Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({new_AGEMA_signal_8188, new_AGEMA_signal_8187, SubBytesIns_Inst_Sbox_3_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M61_U1 ( .a ({new_AGEMA_signal_8168, new_AGEMA_signal_8167, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_5458, new_AGEMA_signal_5457, SubBytesIns_Inst_Sbox_3_T1}), .clk (clk), .r ({Fresh[1169], Fresh[1168], Fresh[1167]}), .c ({new_AGEMA_signal_8660, new_AGEMA_signal_8659, SubBytesIns_Inst_Sbox_3_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M62_U1 ( .a ({new_AGEMA_signal_8646, new_AGEMA_signal_8645, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_5464, new_AGEMA_signal_5463, SubBytesIns_Inst_Sbox_3_T4}), .clk (clk), .r ({Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({new_AGEMA_signal_9100, new_AGEMA_signal_9099, SubBytesIns_Inst_Sbox_3_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M63_U1 ( .a ({new_AGEMA_signal_8166, new_AGEMA_signal_8165, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_5460, new_AGEMA_signal_5459, SubBytesIns_Inst_Sbox_3_T2}), .clk (clk), .r ({Fresh[1175], Fresh[1174], Fresh[1173]}), .c ({new_AGEMA_signal_8662, new_AGEMA_signal_8661, SubBytesIns_Inst_Sbox_3_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L0_U1 ( .a ({new_AGEMA_signal_8660, new_AGEMA_signal_8659, SubBytesIns_Inst_Sbox_3_M61}), .b ({new_AGEMA_signal_9100, new_AGEMA_signal_9099, SubBytesIns_Inst_Sbox_3_M62}), .c ({new_AGEMA_signal_9484, new_AGEMA_signal_9483, SubBytesIns_Inst_Sbox_3_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L1_U1 ( .a ({new_AGEMA_signal_8178, new_AGEMA_signal_8177, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_8182, new_AGEMA_signal_8181, SubBytesIns_Inst_Sbox_3_M56}), .c ({new_AGEMA_signal_8664, new_AGEMA_signal_8663, SubBytesIns_Inst_Sbox_3_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L2_U1 ( .a ({new_AGEMA_signal_8648, new_AGEMA_signal_8647, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_8176, new_AGEMA_signal_8175, SubBytesIns_Inst_Sbox_3_M48}), .c ({new_AGEMA_signal_9102, new_AGEMA_signal_9101, SubBytesIns_Inst_Sbox_3_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L3_U1 ( .a ({new_AGEMA_signal_8174, new_AGEMA_signal_8173, SubBytesIns_Inst_Sbox_3_M47}), .b ({new_AGEMA_signal_8656, new_AGEMA_signal_8655, SubBytesIns_Inst_Sbox_3_M55}), .c ({new_AGEMA_signal_9104, new_AGEMA_signal_9103, SubBytesIns_Inst_Sbox_3_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L4_U1 ( .a ({new_AGEMA_signal_8654, new_AGEMA_signal_8653, SubBytesIns_Inst_Sbox_3_M54}), .b ({new_AGEMA_signal_8658, new_AGEMA_signal_8657, SubBytesIns_Inst_Sbox_3_M58}), .c ({new_AGEMA_signal_9106, new_AGEMA_signal_9105, SubBytesIns_Inst_Sbox_3_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L5_U1 ( .a ({new_AGEMA_signal_8650, new_AGEMA_signal_8649, SubBytesIns_Inst_Sbox_3_M49}), .b ({new_AGEMA_signal_8660, new_AGEMA_signal_8659, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_9108, new_AGEMA_signal_9107, SubBytesIns_Inst_Sbox_3_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L6_U1 ( .a ({new_AGEMA_signal_9100, new_AGEMA_signal_9099, SubBytesIns_Inst_Sbox_3_M62}), .b ({new_AGEMA_signal_9108, new_AGEMA_signal_9107, SubBytesIns_Inst_Sbox_3_L5}), .c ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, SubBytesIns_Inst_Sbox_3_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L7_U1 ( .a ({new_AGEMA_signal_8648, new_AGEMA_signal_8647, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_9104, new_AGEMA_signal_9103, SubBytesIns_Inst_Sbox_3_L3}), .c ({new_AGEMA_signal_9488, new_AGEMA_signal_9487, SubBytesIns_Inst_Sbox_3_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L8_U1 ( .a ({new_AGEMA_signal_8180, new_AGEMA_signal_8179, SubBytesIns_Inst_Sbox_3_M51}), .b ({new_AGEMA_signal_8186, new_AGEMA_signal_8185, SubBytesIns_Inst_Sbox_3_M59}), .c ({new_AGEMA_signal_8666, new_AGEMA_signal_8665, SubBytesIns_Inst_Sbox_3_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L9_U1 ( .a ({new_AGEMA_signal_8652, new_AGEMA_signal_8651, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_9098, new_AGEMA_signal_9097, SubBytesIns_Inst_Sbox_3_M53}), .c ({new_AGEMA_signal_9490, new_AGEMA_signal_9489, SubBytesIns_Inst_Sbox_3_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L10_U1 ( .a ({new_AGEMA_signal_9098, new_AGEMA_signal_9097, SubBytesIns_Inst_Sbox_3_M53}), .b ({new_AGEMA_signal_9106, new_AGEMA_signal_9105, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_9492, new_AGEMA_signal_9491, SubBytesIns_Inst_Sbox_3_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L11_U1 ( .a ({new_AGEMA_signal_8188, new_AGEMA_signal_8187, SubBytesIns_Inst_Sbox_3_M60}), .b ({new_AGEMA_signal_9102, new_AGEMA_signal_9101, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_9494, new_AGEMA_signal_9493, SubBytesIns_Inst_Sbox_3_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L12_U1 ( .a ({new_AGEMA_signal_8176, new_AGEMA_signal_8175, SubBytesIns_Inst_Sbox_3_M48}), .b ({new_AGEMA_signal_8180, new_AGEMA_signal_8179, SubBytesIns_Inst_Sbox_3_M51}), .c ({new_AGEMA_signal_8668, new_AGEMA_signal_8667, SubBytesIns_Inst_Sbox_3_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L13_U1 ( .a ({new_AGEMA_signal_8178, new_AGEMA_signal_8177, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_9484, new_AGEMA_signal_9483, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_9872, new_AGEMA_signal_9871, SubBytesIns_Inst_Sbox_3_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L14_U1 ( .a ({new_AGEMA_signal_8652, new_AGEMA_signal_8651, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_8660, new_AGEMA_signal_8659, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_9110, new_AGEMA_signal_9109, SubBytesIns_Inst_Sbox_3_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L15_U1 ( .a ({new_AGEMA_signal_8656, new_AGEMA_signal_8655, SubBytesIns_Inst_Sbox_3_M55}), .b ({new_AGEMA_signal_8664, new_AGEMA_signal_8663, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_9112, new_AGEMA_signal_9111, SubBytesIns_Inst_Sbox_3_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L16_U1 ( .a ({new_AGEMA_signal_8182, new_AGEMA_signal_8181, SubBytesIns_Inst_Sbox_3_M56}), .b ({new_AGEMA_signal_9484, new_AGEMA_signal_9483, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_9874, new_AGEMA_signal_9873, SubBytesIns_Inst_Sbox_3_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L17_U1 ( .a ({new_AGEMA_signal_8184, new_AGEMA_signal_8183, SubBytesIns_Inst_Sbox_3_M57}), .b ({new_AGEMA_signal_8664, new_AGEMA_signal_8663, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_9114, new_AGEMA_signal_9113, SubBytesIns_Inst_Sbox_3_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L18_U1 ( .a ({new_AGEMA_signal_8658, new_AGEMA_signal_8657, SubBytesIns_Inst_Sbox_3_M58}), .b ({new_AGEMA_signal_8666, new_AGEMA_signal_8665, SubBytesIns_Inst_Sbox_3_L8}), .c ({new_AGEMA_signal_9116, new_AGEMA_signal_9115, SubBytesIns_Inst_Sbox_3_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L19_U1 ( .a ({new_AGEMA_signal_8662, new_AGEMA_signal_8661, SubBytesIns_Inst_Sbox_3_M63}), .b ({new_AGEMA_signal_9106, new_AGEMA_signal_9105, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_9496, new_AGEMA_signal_9495, SubBytesIns_Inst_Sbox_3_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L20_U1 ( .a ({new_AGEMA_signal_9484, new_AGEMA_signal_9483, SubBytesIns_Inst_Sbox_3_L0}), .b ({new_AGEMA_signal_8664, new_AGEMA_signal_8663, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_9876, new_AGEMA_signal_9875, SubBytesIns_Inst_Sbox_3_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L21_U1 ( .a ({new_AGEMA_signal_8664, new_AGEMA_signal_8663, SubBytesIns_Inst_Sbox_3_L1}), .b ({new_AGEMA_signal_9488, new_AGEMA_signal_9487, SubBytesIns_Inst_Sbox_3_L7}), .c ({new_AGEMA_signal_9878, new_AGEMA_signal_9877, SubBytesIns_Inst_Sbox_3_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L22_U1 ( .a ({new_AGEMA_signal_9104, new_AGEMA_signal_9103, SubBytesIns_Inst_Sbox_3_L3}), .b ({new_AGEMA_signal_8668, new_AGEMA_signal_8667, SubBytesIns_Inst_Sbox_3_L12}), .c ({new_AGEMA_signal_9498, new_AGEMA_signal_9497, SubBytesIns_Inst_Sbox_3_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L23_U1 ( .a ({new_AGEMA_signal_9116, new_AGEMA_signal_9115, SubBytesIns_Inst_Sbox_3_L18}), .b ({new_AGEMA_signal_9102, new_AGEMA_signal_9101, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_9500, new_AGEMA_signal_9499, SubBytesIns_Inst_Sbox_3_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L24_U1 ( .a ({new_AGEMA_signal_9112, new_AGEMA_signal_9111, SubBytesIns_Inst_Sbox_3_L15}), .b ({new_AGEMA_signal_9490, new_AGEMA_signal_9489, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_9880, new_AGEMA_signal_9879, SubBytesIns_Inst_Sbox_3_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L25_U1 ( .a ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_9492, new_AGEMA_signal_9491, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_9882, new_AGEMA_signal_9881, SubBytesIns_Inst_Sbox_3_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L26_U1 ( .a ({new_AGEMA_signal_9488, new_AGEMA_signal_9487, SubBytesIns_Inst_Sbox_3_L7}), .b ({new_AGEMA_signal_9490, new_AGEMA_signal_9489, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_9884, new_AGEMA_signal_9883, SubBytesIns_Inst_Sbox_3_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L27_U1 ( .a ({new_AGEMA_signal_8666, new_AGEMA_signal_8665, SubBytesIns_Inst_Sbox_3_L8}), .b ({new_AGEMA_signal_9492, new_AGEMA_signal_9491, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_9886, new_AGEMA_signal_9885, SubBytesIns_Inst_Sbox_3_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L28_U1 ( .a ({new_AGEMA_signal_9494, new_AGEMA_signal_9493, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_9110, new_AGEMA_signal_9109, SubBytesIns_Inst_Sbox_3_L14}), .c ({new_AGEMA_signal_9888, new_AGEMA_signal_9887, SubBytesIns_Inst_Sbox_3_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L29_U1 ( .a ({new_AGEMA_signal_9494, new_AGEMA_signal_9493, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_9114, new_AGEMA_signal_9113, SubBytesIns_Inst_Sbox_3_L17}), .c ({new_AGEMA_signal_9890, new_AGEMA_signal_9889, SubBytesIns_Inst_Sbox_3_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S0_U1 ( .a ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_9880, new_AGEMA_signal_9879, SubBytesIns_Inst_Sbox_3_L24}), .c ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S1_U1 ( .a ({new_AGEMA_signal_9874, new_AGEMA_signal_9873, SubBytesIns_Inst_Sbox_3_L16}), .b ({new_AGEMA_signal_9884, new_AGEMA_signal_9883, SubBytesIns_Inst_Sbox_3_L26}), .c ({new_AGEMA_signal_10266, new_AGEMA_signal_10265, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S2_U1 ( .a ({new_AGEMA_signal_9496, new_AGEMA_signal_9495, SubBytesIns_Inst_Sbox_3_L19}), .b ({new_AGEMA_signal_9888, new_AGEMA_signal_9887, SubBytesIns_Inst_Sbox_3_L28}), .c ({new_AGEMA_signal_10268, new_AGEMA_signal_10267, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S3_U1 ( .a ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_9878, new_AGEMA_signal_9877, SubBytesIns_Inst_Sbox_3_L21}), .c ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S4_U1 ( .a ({new_AGEMA_signal_9876, new_AGEMA_signal_9875, SubBytesIns_Inst_Sbox_3_L20}), .b ({new_AGEMA_signal_9498, new_AGEMA_signal_9497, SubBytesIns_Inst_Sbox_3_L22}), .c ({new_AGEMA_signal_10272, new_AGEMA_signal_10271, MixColumnsInput[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S5_U1 ( .a ({new_AGEMA_signal_9882, new_AGEMA_signal_9881, SubBytesIns_Inst_Sbox_3_L25}), .b ({new_AGEMA_signal_9890, new_AGEMA_signal_9889, SubBytesIns_Inst_Sbox_3_L29}), .c ({new_AGEMA_signal_10274, new_AGEMA_signal_10273, MixColumnsInput[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S6_U1 ( .a ({new_AGEMA_signal_9872, new_AGEMA_signal_9871, SubBytesIns_Inst_Sbox_3_L13}), .b ({new_AGEMA_signal_9886, new_AGEMA_signal_9885, SubBytesIns_Inst_Sbox_3_L27}), .c ({new_AGEMA_signal_10276, new_AGEMA_signal_10275, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S7_U1 ( .a ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_9500, new_AGEMA_signal_9499, SubBytesIns_Inst_Sbox_3_L23}), .c ({new_AGEMA_signal_9892, new_AGEMA_signal_9891, MixColumnsInput[24]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M46_U1 ( .a ({new_AGEMA_signal_8196, new_AGEMA_signal_8195, SubBytesIns_Inst_Sbox_4_M44}), .b ({new_AGEMA_signal_5846, new_AGEMA_signal_5845, SubBytesIns_Inst_Sbox_4_T6}), .clk (clk), .r ({Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({new_AGEMA_signal_8672, new_AGEMA_signal_8671, SubBytesIns_Inst_Sbox_4_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M47_U1 ( .a ({new_AGEMA_signal_7908, new_AGEMA_signal_7907, SubBytesIns_Inst_Sbox_4_M40}), .b ({new_AGEMA_signal_6246, new_AGEMA_signal_6245, SubBytesIns_Inst_Sbox_4_T8}), .clk (clk), .r ({Fresh[1181], Fresh[1180], Fresh[1179]}), .c ({new_AGEMA_signal_8198, new_AGEMA_signal_8197, SubBytesIns_Inst_Sbox_4_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M48_U1 ( .a ({new_AGEMA_signal_7906, new_AGEMA_signal_7905, SubBytesIns_Inst_Sbox_4_M39}), .b ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .clk (clk), .r ({Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({new_AGEMA_signal_8200, new_AGEMA_signal_8199, SubBytesIns_Inst_Sbox_4_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M49_U1 ( .a ({new_AGEMA_signal_8194, new_AGEMA_signal_8193, SubBytesIns_Inst_Sbox_4_M43}), .b ({new_AGEMA_signal_5854, new_AGEMA_signal_5853, SubBytesIns_Inst_Sbox_4_T16}), .clk (clk), .r ({Fresh[1187], Fresh[1186], Fresh[1185]}), .c ({new_AGEMA_signal_8674, new_AGEMA_signal_8673, SubBytesIns_Inst_Sbox_4_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M50_U1 ( .a ({new_AGEMA_signal_7904, new_AGEMA_signal_7903, SubBytesIns_Inst_Sbox_4_M38}), .b ({new_AGEMA_signal_5848, new_AGEMA_signal_5847, SubBytesIns_Inst_Sbox_4_T9}), .clk (clk), .r ({Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({new_AGEMA_signal_8202, new_AGEMA_signal_8201, SubBytesIns_Inst_Sbox_4_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M51_U1 ( .a ({new_AGEMA_signal_7902, new_AGEMA_signal_7901, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_6252, new_AGEMA_signal_6251, SubBytesIns_Inst_Sbox_4_T17}), .clk (clk), .r ({Fresh[1193], Fresh[1192], Fresh[1191]}), .c ({new_AGEMA_signal_8204, new_AGEMA_signal_8203, SubBytesIns_Inst_Sbox_4_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M52_U1 ( .a ({new_AGEMA_signal_8192, new_AGEMA_signal_8191, SubBytesIns_Inst_Sbox_4_M42}), .b ({new_AGEMA_signal_5852, new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_4_T15}), .clk (clk), .r ({Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({new_AGEMA_signal_8676, new_AGEMA_signal_8675, SubBytesIns_Inst_Sbox_4_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M53_U1 ( .a ({new_AGEMA_signal_8670, new_AGEMA_signal_8669, SubBytesIns_Inst_Sbox_4_M45}), .b ({new_AGEMA_signal_5860, new_AGEMA_signal_5859, SubBytesIns_Inst_Sbox_4_T27}), .clk (clk), .r ({Fresh[1199], Fresh[1198], Fresh[1197]}), .c ({new_AGEMA_signal_9118, new_AGEMA_signal_9117, SubBytesIns_Inst_Sbox_4_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M54_U1 ( .a ({new_AGEMA_signal_8190, new_AGEMA_signal_8189, SubBytesIns_Inst_Sbox_4_M41}), .b ({new_AGEMA_signal_6248, new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_4_T10}), .clk (clk), .r ({Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({new_AGEMA_signal_8678, new_AGEMA_signal_8677, SubBytesIns_Inst_Sbox_4_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M55_U1 ( .a ({new_AGEMA_signal_8196, new_AGEMA_signal_8195, SubBytesIns_Inst_Sbox_4_M44}), .b ({new_AGEMA_signal_5850, new_AGEMA_signal_5849, SubBytesIns_Inst_Sbox_4_T13}), .clk (clk), .r ({Fresh[1205], Fresh[1204], Fresh[1203]}), .c ({new_AGEMA_signal_8680, new_AGEMA_signal_8679, SubBytesIns_Inst_Sbox_4_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M56_U1 ( .a ({new_AGEMA_signal_7908, new_AGEMA_signal_7907, SubBytesIns_Inst_Sbox_4_M40}), .b ({new_AGEMA_signal_6256, new_AGEMA_signal_6255, SubBytesIns_Inst_Sbox_4_T23}), .clk (clk), .r ({Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({new_AGEMA_signal_8206, new_AGEMA_signal_8205, SubBytesIns_Inst_Sbox_4_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M57_U1 ( .a ({new_AGEMA_signal_7906, new_AGEMA_signal_7905, SubBytesIns_Inst_Sbox_4_M39}), .b ({new_AGEMA_signal_5856, new_AGEMA_signal_5855, SubBytesIns_Inst_Sbox_4_T19}), .clk (clk), .r ({Fresh[1211], Fresh[1210], Fresh[1209]}), .c ({new_AGEMA_signal_8208, new_AGEMA_signal_8207, SubBytesIns_Inst_Sbox_4_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M58_U1 ( .a ({new_AGEMA_signal_8194, new_AGEMA_signal_8193, SubBytesIns_Inst_Sbox_4_M43}), .b ({new_AGEMA_signal_5482, new_AGEMA_signal_5481, SubBytesIns_Inst_Sbox_4_T3}), .clk (clk), .r ({Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({new_AGEMA_signal_8682, new_AGEMA_signal_8681, SubBytesIns_Inst_Sbox_4_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M59_U1 ( .a ({new_AGEMA_signal_7904, new_AGEMA_signal_7903, SubBytesIns_Inst_Sbox_4_M38}), .b ({new_AGEMA_signal_5858, new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_4_T22}), .clk (clk), .r ({Fresh[1217], Fresh[1216], Fresh[1215]}), .c ({new_AGEMA_signal_8210, new_AGEMA_signal_8209, SubBytesIns_Inst_Sbox_4_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M60_U1 ( .a ({new_AGEMA_signal_7902, new_AGEMA_signal_7901, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_6254, new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_4_T20}), .clk (clk), .r ({Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({new_AGEMA_signal_8212, new_AGEMA_signal_8211, SubBytesIns_Inst_Sbox_4_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M61_U1 ( .a ({new_AGEMA_signal_8192, new_AGEMA_signal_8191, SubBytesIns_Inst_Sbox_4_M42}), .b ({new_AGEMA_signal_5478, new_AGEMA_signal_5477, SubBytesIns_Inst_Sbox_4_T1}), .clk (clk), .r ({Fresh[1223], Fresh[1222], Fresh[1221]}), .c ({new_AGEMA_signal_8684, new_AGEMA_signal_8683, SubBytesIns_Inst_Sbox_4_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M62_U1 ( .a ({new_AGEMA_signal_8670, new_AGEMA_signal_8669, SubBytesIns_Inst_Sbox_4_M45}), .b ({new_AGEMA_signal_5484, new_AGEMA_signal_5483, SubBytesIns_Inst_Sbox_4_T4}), .clk (clk), .r ({Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({new_AGEMA_signal_9120, new_AGEMA_signal_9119, SubBytesIns_Inst_Sbox_4_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M63_U1 ( .a ({new_AGEMA_signal_8190, new_AGEMA_signal_8189, SubBytesIns_Inst_Sbox_4_M41}), .b ({new_AGEMA_signal_5480, new_AGEMA_signal_5479, SubBytesIns_Inst_Sbox_4_T2}), .clk (clk), .r ({Fresh[1229], Fresh[1228], Fresh[1227]}), .c ({new_AGEMA_signal_8686, new_AGEMA_signal_8685, SubBytesIns_Inst_Sbox_4_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L0_U1 ( .a ({new_AGEMA_signal_8684, new_AGEMA_signal_8683, SubBytesIns_Inst_Sbox_4_M61}), .b ({new_AGEMA_signal_9120, new_AGEMA_signal_9119, SubBytesIns_Inst_Sbox_4_M62}), .c ({new_AGEMA_signal_9502, new_AGEMA_signal_9501, SubBytesIns_Inst_Sbox_4_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L1_U1 ( .a ({new_AGEMA_signal_8202, new_AGEMA_signal_8201, SubBytesIns_Inst_Sbox_4_M50}), .b ({new_AGEMA_signal_8206, new_AGEMA_signal_8205, SubBytesIns_Inst_Sbox_4_M56}), .c ({new_AGEMA_signal_8688, new_AGEMA_signal_8687, SubBytesIns_Inst_Sbox_4_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L2_U1 ( .a ({new_AGEMA_signal_8672, new_AGEMA_signal_8671, SubBytesIns_Inst_Sbox_4_M46}), .b ({new_AGEMA_signal_8200, new_AGEMA_signal_8199, SubBytesIns_Inst_Sbox_4_M48}), .c ({new_AGEMA_signal_9122, new_AGEMA_signal_9121, SubBytesIns_Inst_Sbox_4_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L3_U1 ( .a ({new_AGEMA_signal_8198, new_AGEMA_signal_8197, SubBytesIns_Inst_Sbox_4_M47}), .b ({new_AGEMA_signal_8680, new_AGEMA_signal_8679, SubBytesIns_Inst_Sbox_4_M55}), .c ({new_AGEMA_signal_9124, new_AGEMA_signal_9123, SubBytesIns_Inst_Sbox_4_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L4_U1 ( .a ({new_AGEMA_signal_8678, new_AGEMA_signal_8677, SubBytesIns_Inst_Sbox_4_M54}), .b ({new_AGEMA_signal_8682, new_AGEMA_signal_8681, SubBytesIns_Inst_Sbox_4_M58}), .c ({new_AGEMA_signal_9126, new_AGEMA_signal_9125, SubBytesIns_Inst_Sbox_4_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L5_U1 ( .a ({new_AGEMA_signal_8674, new_AGEMA_signal_8673, SubBytesIns_Inst_Sbox_4_M49}), .b ({new_AGEMA_signal_8684, new_AGEMA_signal_8683, SubBytesIns_Inst_Sbox_4_M61}), .c ({new_AGEMA_signal_9128, new_AGEMA_signal_9127, SubBytesIns_Inst_Sbox_4_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L6_U1 ( .a ({new_AGEMA_signal_9120, new_AGEMA_signal_9119, SubBytesIns_Inst_Sbox_4_M62}), .b ({new_AGEMA_signal_9128, new_AGEMA_signal_9127, SubBytesIns_Inst_Sbox_4_L5}), .c ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, SubBytesIns_Inst_Sbox_4_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L7_U1 ( .a ({new_AGEMA_signal_8672, new_AGEMA_signal_8671, SubBytesIns_Inst_Sbox_4_M46}), .b ({new_AGEMA_signal_9124, new_AGEMA_signal_9123, SubBytesIns_Inst_Sbox_4_L3}), .c ({new_AGEMA_signal_9506, new_AGEMA_signal_9505, SubBytesIns_Inst_Sbox_4_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L8_U1 ( .a ({new_AGEMA_signal_8204, new_AGEMA_signal_8203, SubBytesIns_Inst_Sbox_4_M51}), .b ({new_AGEMA_signal_8210, new_AGEMA_signal_8209, SubBytesIns_Inst_Sbox_4_M59}), .c ({new_AGEMA_signal_8690, new_AGEMA_signal_8689, SubBytesIns_Inst_Sbox_4_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L9_U1 ( .a ({new_AGEMA_signal_8676, new_AGEMA_signal_8675, SubBytesIns_Inst_Sbox_4_M52}), .b ({new_AGEMA_signal_9118, new_AGEMA_signal_9117, SubBytesIns_Inst_Sbox_4_M53}), .c ({new_AGEMA_signal_9508, new_AGEMA_signal_9507, SubBytesIns_Inst_Sbox_4_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L10_U1 ( .a ({new_AGEMA_signal_9118, new_AGEMA_signal_9117, SubBytesIns_Inst_Sbox_4_M53}), .b ({new_AGEMA_signal_9126, new_AGEMA_signal_9125, SubBytesIns_Inst_Sbox_4_L4}), .c ({new_AGEMA_signal_9510, new_AGEMA_signal_9509, SubBytesIns_Inst_Sbox_4_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L11_U1 ( .a ({new_AGEMA_signal_8212, new_AGEMA_signal_8211, SubBytesIns_Inst_Sbox_4_M60}), .b ({new_AGEMA_signal_9122, new_AGEMA_signal_9121, SubBytesIns_Inst_Sbox_4_L2}), .c ({new_AGEMA_signal_9512, new_AGEMA_signal_9511, SubBytesIns_Inst_Sbox_4_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L12_U1 ( .a ({new_AGEMA_signal_8200, new_AGEMA_signal_8199, SubBytesIns_Inst_Sbox_4_M48}), .b ({new_AGEMA_signal_8204, new_AGEMA_signal_8203, SubBytesIns_Inst_Sbox_4_M51}), .c ({new_AGEMA_signal_8692, new_AGEMA_signal_8691, SubBytesIns_Inst_Sbox_4_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L13_U1 ( .a ({new_AGEMA_signal_8202, new_AGEMA_signal_8201, SubBytesIns_Inst_Sbox_4_M50}), .b ({new_AGEMA_signal_9502, new_AGEMA_signal_9501, SubBytesIns_Inst_Sbox_4_L0}), .c ({new_AGEMA_signal_9894, new_AGEMA_signal_9893, SubBytesIns_Inst_Sbox_4_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L14_U1 ( .a ({new_AGEMA_signal_8676, new_AGEMA_signal_8675, SubBytesIns_Inst_Sbox_4_M52}), .b ({new_AGEMA_signal_8684, new_AGEMA_signal_8683, SubBytesIns_Inst_Sbox_4_M61}), .c ({new_AGEMA_signal_9130, new_AGEMA_signal_9129, SubBytesIns_Inst_Sbox_4_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L15_U1 ( .a ({new_AGEMA_signal_8680, new_AGEMA_signal_8679, SubBytesIns_Inst_Sbox_4_M55}), .b ({new_AGEMA_signal_8688, new_AGEMA_signal_8687, SubBytesIns_Inst_Sbox_4_L1}), .c ({new_AGEMA_signal_9132, new_AGEMA_signal_9131, SubBytesIns_Inst_Sbox_4_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L16_U1 ( .a ({new_AGEMA_signal_8206, new_AGEMA_signal_8205, SubBytesIns_Inst_Sbox_4_M56}), .b ({new_AGEMA_signal_9502, new_AGEMA_signal_9501, SubBytesIns_Inst_Sbox_4_L0}), .c ({new_AGEMA_signal_9896, new_AGEMA_signal_9895, SubBytesIns_Inst_Sbox_4_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L17_U1 ( .a ({new_AGEMA_signal_8208, new_AGEMA_signal_8207, SubBytesIns_Inst_Sbox_4_M57}), .b ({new_AGEMA_signal_8688, new_AGEMA_signal_8687, SubBytesIns_Inst_Sbox_4_L1}), .c ({new_AGEMA_signal_9134, new_AGEMA_signal_9133, SubBytesIns_Inst_Sbox_4_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L18_U1 ( .a ({new_AGEMA_signal_8682, new_AGEMA_signal_8681, SubBytesIns_Inst_Sbox_4_M58}), .b ({new_AGEMA_signal_8690, new_AGEMA_signal_8689, SubBytesIns_Inst_Sbox_4_L8}), .c ({new_AGEMA_signal_9136, new_AGEMA_signal_9135, SubBytesIns_Inst_Sbox_4_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L19_U1 ( .a ({new_AGEMA_signal_8686, new_AGEMA_signal_8685, SubBytesIns_Inst_Sbox_4_M63}), .b ({new_AGEMA_signal_9126, new_AGEMA_signal_9125, SubBytesIns_Inst_Sbox_4_L4}), .c ({new_AGEMA_signal_9514, new_AGEMA_signal_9513, SubBytesIns_Inst_Sbox_4_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L20_U1 ( .a ({new_AGEMA_signal_9502, new_AGEMA_signal_9501, SubBytesIns_Inst_Sbox_4_L0}), .b ({new_AGEMA_signal_8688, new_AGEMA_signal_8687, SubBytesIns_Inst_Sbox_4_L1}), .c ({new_AGEMA_signal_9898, new_AGEMA_signal_9897, SubBytesIns_Inst_Sbox_4_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L21_U1 ( .a ({new_AGEMA_signal_8688, new_AGEMA_signal_8687, SubBytesIns_Inst_Sbox_4_L1}), .b ({new_AGEMA_signal_9506, new_AGEMA_signal_9505, SubBytesIns_Inst_Sbox_4_L7}), .c ({new_AGEMA_signal_9900, new_AGEMA_signal_9899, SubBytesIns_Inst_Sbox_4_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L22_U1 ( .a ({new_AGEMA_signal_9124, new_AGEMA_signal_9123, SubBytesIns_Inst_Sbox_4_L3}), .b ({new_AGEMA_signal_8692, new_AGEMA_signal_8691, SubBytesIns_Inst_Sbox_4_L12}), .c ({new_AGEMA_signal_9516, new_AGEMA_signal_9515, SubBytesIns_Inst_Sbox_4_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L23_U1 ( .a ({new_AGEMA_signal_9136, new_AGEMA_signal_9135, SubBytesIns_Inst_Sbox_4_L18}), .b ({new_AGEMA_signal_9122, new_AGEMA_signal_9121, SubBytesIns_Inst_Sbox_4_L2}), .c ({new_AGEMA_signal_9518, new_AGEMA_signal_9517, SubBytesIns_Inst_Sbox_4_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L24_U1 ( .a ({new_AGEMA_signal_9132, new_AGEMA_signal_9131, SubBytesIns_Inst_Sbox_4_L15}), .b ({new_AGEMA_signal_9508, new_AGEMA_signal_9507, SubBytesIns_Inst_Sbox_4_L9}), .c ({new_AGEMA_signal_9902, new_AGEMA_signal_9901, SubBytesIns_Inst_Sbox_4_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L25_U1 ( .a ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_9510, new_AGEMA_signal_9509, SubBytesIns_Inst_Sbox_4_L10}), .c ({new_AGEMA_signal_9904, new_AGEMA_signal_9903, SubBytesIns_Inst_Sbox_4_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L26_U1 ( .a ({new_AGEMA_signal_9506, new_AGEMA_signal_9505, SubBytesIns_Inst_Sbox_4_L7}), .b ({new_AGEMA_signal_9508, new_AGEMA_signal_9507, SubBytesIns_Inst_Sbox_4_L9}), .c ({new_AGEMA_signal_9906, new_AGEMA_signal_9905, SubBytesIns_Inst_Sbox_4_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L27_U1 ( .a ({new_AGEMA_signal_8690, new_AGEMA_signal_8689, SubBytesIns_Inst_Sbox_4_L8}), .b ({new_AGEMA_signal_9510, new_AGEMA_signal_9509, SubBytesIns_Inst_Sbox_4_L10}), .c ({new_AGEMA_signal_9908, new_AGEMA_signal_9907, SubBytesIns_Inst_Sbox_4_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L28_U1 ( .a ({new_AGEMA_signal_9512, new_AGEMA_signal_9511, SubBytesIns_Inst_Sbox_4_L11}), .b ({new_AGEMA_signal_9130, new_AGEMA_signal_9129, SubBytesIns_Inst_Sbox_4_L14}), .c ({new_AGEMA_signal_9910, new_AGEMA_signal_9909, SubBytesIns_Inst_Sbox_4_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L29_U1 ( .a ({new_AGEMA_signal_9512, new_AGEMA_signal_9511, SubBytesIns_Inst_Sbox_4_L11}), .b ({new_AGEMA_signal_9134, new_AGEMA_signal_9133, SubBytesIns_Inst_Sbox_4_L17}), .c ({new_AGEMA_signal_9912, new_AGEMA_signal_9911, SubBytesIns_Inst_Sbox_4_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S0_U1 ( .a ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_9902, new_AGEMA_signal_9901, SubBytesIns_Inst_Sbox_4_L24}), .c ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S1_U1 ( .a ({new_AGEMA_signal_9896, new_AGEMA_signal_9895, SubBytesIns_Inst_Sbox_4_L16}), .b ({new_AGEMA_signal_9906, new_AGEMA_signal_9905, SubBytesIns_Inst_Sbox_4_L26}), .c ({new_AGEMA_signal_10280, new_AGEMA_signal_10279, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S2_U1 ( .a ({new_AGEMA_signal_9514, new_AGEMA_signal_9513, SubBytesIns_Inst_Sbox_4_L19}), .b ({new_AGEMA_signal_9910, new_AGEMA_signal_9909, SubBytesIns_Inst_Sbox_4_L28}), .c ({new_AGEMA_signal_10282, new_AGEMA_signal_10281, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S3_U1 ( .a ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_9900, new_AGEMA_signal_9899, SubBytesIns_Inst_Sbox_4_L21}), .c ({new_AGEMA_signal_10284, new_AGEMA_signal_10283, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S4_U1 ( .a ({new_AGEMA_signal_9898, new_AGEMA_signal_9897, SubBytesIns_Inst_Sbox_4_L20}), .b ({new_AGEMA_signal_9516, new_AGEMA_signal_9515, SubBytesIns_Inst_Sbox_4_L22}), .c ({new_AGEMA_signal_10286, new_AGEMA_signal_10285, MixColumnsInput[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S5_U1 ( .a ({new_AGEMA_signal_9904, new_AGEMA_signal_9903, SubBytesIns_Inst_Sbox_4_L25}), .b ({new_AGEMA_signal_9912, new_AGEMA_signal_9911, SubBytesIns_Inst_Sbox_4_L29}), .c ({new_AGEMA_signal_10288, new_AGEMA_signal_10287, MixColumnsInput[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S6_U1 ( .a ({new_AGEMA_signal_9894, new_AGEMA_signal_9893, SubBytesIns_Inst_Sbox_4_L13}), .b ({new_AGEMA_signal_9908, new_AGEMA_signal_9907, SubBytesIns_Inst_Sbox_4_L27}), .c ({new_AGEMA_signal_10290, new_AGEMA_signal_10289, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S7_U1 ( .a ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_9518, new_AGEMA_signal_9517, SubBytesIns_Inst_Sbox_4_L23}), .c ({new_AGEMA_signal_9914, new_AGEMA_signal_9913, MixColumnsInput[0]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M46_U1 ( .a ({new_AGEMA_signal_8220, new_AGEMA_signal_8219, SubBytesIns_Inst_Sbox_5_M44}), .b ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, SubBytesIns_Inst_Sbox_5_T6}), .clk (clk), .r ({Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({new_AGEMA_signal_8696, new_AGEMA_signal_8695, SubBytesIns_Inst_Sbox_5_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M47_U1 ( .a ({new_AGEMA_signal_7916, new_AGEMA_signal_7915, SubBytesIns_Inst_Sbox_5_M40}), .b ({new_AGEMA_signal_6272, new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_5_T8}), .clk (clk), .r ({Fresh[1235], Fresh[1234], Fresh[1233]}), .c ({new_AGEMA_signal_8222, new_AGEMA_signal_8221, SubBytesIns_Inst_Sbox_5_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M48_U1 ( .a ({new_AGEMA_signal_7914, new_AGEMA_signal_7913, SubBytesIns_Inst_Sbox_5_M39}), .b ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .clk (clk), .r ({Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({new_AGEMA_signal_8224, new_AGEMA_signal_8223, SubBytesIns_Inst_Sbox_5_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M49_U1 ( .a ({new_AGEMA_signal_8218, new_AGEMA_signal_8217, SubBytesIns_Inst_Sbox_5_M43}), .b ({new_AGEMA_signal_5870, new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_5_T16}), .clk (clk), .r ({Fresh[1241], Fresh[1240], Fresh[1239]}), .c ({new_AGEMA_signal_8698, new_AGEMA_signal_8697, SubBytesIns_Inst_Sbox_5_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M50_U1 ( .a ({new_AGEMA_signal_7912, new_AGEMA_signal_7911, SubBytesIns_Inst_Sbox_5_M38}), .b ({new_AGEMA_signal_5864, new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_5_T9}), .clk (clk), .r ({Fresh[1244], Fresh[1243], Fresh[1242]}), .c ({new_AGEMA_signal_8226, new_AGEMA_signal_8225, SubBytesIns_Inst_Sbox_5_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M51_U1 ( .a ({new_AGEMA_signal_7910, new_AGEMA_signal_7909, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_6278, new_AGEMA_signal_6277, SubBytesIns_Inst_Sbox_5_T17}), .clk (clk), .r ({Fresh[1247], Fresh[1246], Fresh[1245]}), .c ({new_AGEMA_signal_8228, new_AGEMA_signal_8227, SubBytesIns_Inst_Sbox_5_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M52_U1 ( .a ({new_AGEMA_signal_8216, new_AGEMA_signal_8215, SubBytesIns_Inst_Sbox_5_M42}), .b ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, SubBytesIns_Inst_Sbox_5_T15}), .clk (clk), .r ({Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({new_AGEMA_signal_8700, new_AGEMA_signal_8699, SubBytesIns_Inst_Sbox_5_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M53_U1 ( .a ({new_AGEMA_signal_8694, new_AGEMA_signal_8693, SubBytesIns_Inst_Sbox_5_M45}), .b ({new_AGEMA_signal_5876, new_AGEMA_signal_5875, SubBytesIns_Inst_Sbox_5_T27}), .clk (clk), .r ({Fresh[1253], Fresh[1252], Fresh[1251]}), .c ({new_AGEMA_signal_9138, new_AGEMA_signal_9137, SubBytesIns_Inst_Sbox_5_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M54_U1 ( .a ({new_AGEMA_signal_8214, new_AGEMA_signal_8213, SubBytesIns_Inst_Sbox_5_M41}), .b ({new_AGEMA_signal_6274, new_AGEMA_signal_6273, SubBytesIns_Inst_Sbox_5_T10}), .clk (clk), .r ({Fresh[1256], Fresh[1255], Fresh[1254]}), .c ({new_AGEMA_signal_8702, new_AGEMA_signal_8701, SubBytesIns_Inst_Sbox_5_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M55_U1 ( .a ({new_AGEMA_signal_8220, new_AGEMA_signal_8219, SubBytesIns_Inst_Sbox_5_M44}), .b ({new_AGEMA_signal_5866, new_AGEMA_signal_5865, SubBytesIns_Inst_Sbox_5_T13}), .clk (clk), .r ({Fresh[1259], Fresh[1258], Fresh[1257]}), .c ({new_AGEMA_signal_8704, new_AGEMA_signal_8703, SubBytesIns_Inst_Sbox_5_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M56_U1 ( .a ({new_AGEMA_signal_7916, new_AGEMA_signal_7915, SubBytesIns_Inst_Sbox_5_M40}), .b ({new_AGEMA_signal_6282, new_AGEMA_signal_6281, SubBytesIns_Inst_Sbox_5_T23}), .clk (clk), .r ({Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({new_AGEMA_signal_8230, new_AGEMA_signal_8229, SubBytesIns_Inst_Sbox_5_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M57_U1 ( .a ({new_AGEMA_signal_7914, new_AGEMA_signal_7913, SubBytesIns_Inst_Sbox_5_M39}), .b ({new_AGEMA_signal_5872, new_AGEMA_signal_5871, SubBytesIns_Inst_Sbox_5_T19}), .clk (clk), .r ({Fresh[1265], Fresh[1264], Fresh[1263]}), .c ({new_AGEMA_signal_8232, new_AGEMA_signal_8231, SubBytesIns_Inst_Sbox_5_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M58_U1 ( .a ({new_AGEMA_signal_8218, new_AGEMA_signal_8217, SubBytesIns_Inst_Sbox_5_M43}), .b ({new_AGEMA_signal_5502, new_AGEMA_signal_5501, SubBytesIns_Inst_Sbox_5_T3}), .clk (clk), .r ({Fresh[1268], Fresh[1267], Fresh[1266]}), .c ({new_AGEMA_signal_8706, new_AGEMA_signal_8705, SubBytesIns_Inst_Sbox_5_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M59_U1 ( .a ({new_AGEMA_signal_7912, new_AGEMA_signal_7911, SubBytesIns_Inst_Sbox_5_M38}), .b ({new_AGEMA_signal_5874, new_AGEMA_signal_5873, SubBytesIns_Inst_Sbox_5_T22}), .clk (clk), .r ({Fresh[1271], Fresh[1270], Fresh[1269]}), .c ({new_AGEMA_signal_8234, new_AGEMA_signal_8233, SubBytesIns_Inst_Sbox_5_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M60_U1 ( .a ({new_AGEMA_signal_7910, new_AGEMA_signal_7909, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_6280, new_AGEMA_signal_6279, SubBytesIns_Inst_Sbox_5_T20}), .clk (clk), .r ({Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({new_AGEMA_signal_8236, new_AGEMA_signal_8235, SubBytesIns_Inst_Sbox_5_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M61_U1 ( .a ({new_AGEMA_signal_8216, new_AGEMA_signal_8215, SubBytesIns_Inst_Sbox_5_M42}), .b ({new_AGEMA_signal_5498, new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_5_T1}), .clk (clk), .r ({Fresh[1277], Fresh[1276], Fresh[1275]}), .c ({new_AGEMA_signal_8708, new_AGEMA_signal_8707, SubBytesIns_Inst_Sbox_5_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M62_U1 ( .a ({new_AGEMA_signal_8694, new_AGEMA_signal_8693, SubBytesIns_Inst_Sbox_5_M45}), .b ({new_AGEMA_signal_5504, new_AGEMA_signal_5503, SubBytesIns_Inst_Sbox_5_T4}), .clk (clk), .r ({Fresh[1280], Fresh[1279], Fresh[1278]}), .c ({new_AGEMA_signal_9140, new_AGEMA_signal_9139, SubBytesIns_Inst_Sbox_5_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M63_U1 ( .a ({new_AGEMA_signal_8214, new_AGEMA_signal_8213, SubBytesIns_Inst_Sbox_5_M41}), .b ({new_AGEMA_signal_5500, new_AGEMA_signal_5499, SubBytesIns_Inst_Sbox_5_T2}), .clk (clk), .r ({Fresh[1283], Fresh[1282], Fresh[1281]}), .c ({new_AGEMA_signal_8710, new_AGEMA_signal_8709, SubBytesIns_Inst_Sbox_5_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L0_U1 ( .a ({new_AGEMA_signal_8708, new_AGEMA_signal_8707, SubBytesIns_Inst_Sbox_5_M61}), .b ({new_AGEMA_signal_9140, new_AGEMA_signal_9139, SubBytesIns_Inst_Sbox_5_M62}), .c ({new_AGEMA_signal_9520, new_AGEMA_signal_9519, SubBytesIns_Inst_Sbox_5_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L1_U1 ( .a ({new_AGEMA_signal_8226, new_AGEMA_signal_8225, SubBytesIns_Inst_Sbox_5_M50}), .b ({new_AGEMA_signal_8230, new_AGEMA_signal_8229, SubBytesIns_Inst_Sbox_5_M56}), .c ({new_AGEMA_signal_8712, new_AGEMA_signal_8711, SubBytesIns_Inst_Sbox_5_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L2_U1 ( .a ({new_AGEMA_signal_8696, new_AGEMA_signal_8695, SubBytesIns_Inst_Sbox_5_M46}), .b ({new_AGEMA_signal_8224, new_AGEMA_signal_8223, SubBytesIns_Inst_Sbox_5_M48}), .c ({new_AGEMA_signal_9142, new_AGEMA_signal_9141, SubBytesIns_Inst_Sbox_5_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L3_U1 ( .a ({new_AGEMA_signal_8222, new_AGEMA_signal_8221, SubBytesIns_Inst_Sbox_5_M47}), .b ({new_AGEMA_signal_8704, new_AGEMA_signal_8703, SubBytesIns_Inst_Sbox_5_M55}), .c ({new_AGEMA_signal_9144, new_AGEMA_signal_9143, SubBytesIns_Inst_Sbox_5_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L4_U1 ( .a ({new_AGEMA_signal_8702, new_AGEMA_signal_8701, SubBytesIns_Inst_Sbox_5_M54}), .b ({new_AGEMA_signal_8706, new_AGEMA_signal_8705, SubBytesIns_Inst_Sbox_5_M58}), .c ({new_AGEMA_signal_9146, new_AGEMA_signal_9145, SubBytesIns_Inst_Sbox_5_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L5_U1 ( .a ({new_AGEMA_signal_8698, new_AGEMA_signal_8697, SubBytesIns_Inst_Sbox_5_M49}), .b ({new_AGEMA_signal_8708, new_AGEMA_signal_8707, SubBytesIns_Inst_Sbox_5_M61}), .c ({new_AGEMA_signal_9148, new_AGEMA_signal_9147, SubBytesIns_Inst_Sbox_5_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L6_U1 ( .a ({new_AGEMA_signal_9140, new_AGEMA_signal_9139, SubBytesIns_Inst_Sbox_5_M62}), .b ({new_AGEMA_signal_9148, new_AGEMA_signal_9147, SubBytesIns_Inst_Sbox_5_L5}), .c ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, SubBytesIns_Inst_Sbox_5_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L7_U1 ( .a ({new_AGEMA_signal_8696, new_AGEMA_signal_8695, SubBytesIns_Inst_Sbox_5_M46}), .b ({new_AGEMA_signal_9144, new_AGEMA_signal_9143, SubBytesIns_Inst_Sbox_5_L3}), .c ({new_AGEMA_signal_9524, new_AGEMA_signal_9523, SubBytesIns_Inst_Sbox_5_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L8_U1 ( .a ({new_AGEMA_signal_8228, new_AGEMA_signal_8227, SubBytesIns_Inst_Sbox_5_M51}), .b ({new_AGEMA_signal_8234, new_AGEMA_signal_8233, SubBytesIns_Inst_Sbox_5_M59}), .c ({new_AGEMA_signal_8714, new_AGEMA_signal_8713, SubBytesIns_Inst_Sbox_5_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L9_U1 ( .a ({new_AGEMA_signal_8700, new_AGEMA_signal_8699, SubBytesIns_Inst_Sbox_5_M52}), .b ({new_AGEMA_signal_9138, new_AGEMA_signal_9137, SubBytesIns_Inst_Sbox_5_M53}), .c ({new_AGEMA_signal_9526, new_AGEMA_signal_9525, SubBytesIns_Inst_Sbox_5_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L10_U1 ( .a ({new_AGEMA_signal_9138, new_AGEMA_signal_9137, SubBytesIns_Inst_Sbox_5_M53}), .b ({new_AGEMA_signal_9146, new_AGEMA_signal_9145, SubBytesIns_Inst_Sbox_5_L4}), .c ({new_AGEMA_signal_9528, new_AGEMA_signal_9527, SubBytesIns_Inst_Sbox_5_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L11_U1 ( .a ({new_AGEMA_signal_8236, new_AGEMA_signal_8235, SubBytesIns_Inst_Sbox_5_M60}), .b ({new_AGEMA_signal_9142, new_AGEMA_signal_9141, SubBytesIns_Inst_Sbox_5_L2}), .c ({new_AGEMA_signal_9530, new_AGEMA_signal_9529, SubBytesIns_Inst_Sbox_5_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L12_U1 ( .a ({new_AGEMA_signal_8224, new_AGEMA_signal_8223, SubBytesIns_Inst_Sbox_5_M48}), .b ({new_AGEMA_signal_8228, new_AGEMA_signal_8227, SubBytesIns_Inst_Sbox_5_M51}), .c ({new_AGEMA_signal_8716, new_AGEMA_signal_8715, SubBytesIns_Inst_Sbox_5_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L13_U1 ( .a ({new_AGEMA_signal_8226, new_AGEMA_signal_8225, SubBytesIns_Inst_Sbox_5_M50}), .b ({new_AGEMA_signal_9520, new_AGEMA_signal_9519, SubBytesIns_Inst_Sbox_5_L0}), .c ({new_AGEMA_signal_9916, new_AGEMA_signal_9915, SubBytesIns_Inst_Sbox_5_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L14_U1 ( .a ({new_AGEMA_signal_8700, new_AGEMA_signal_8699, SubBytesIns_Inst_Sbox_5_M52}), .b ({new_AGEMA_signal_8708, new_AGEMA_signal_8707, SubBytesIns_Inst_Sbox_5_M61}), .c ({new_AGEMA_signal_9150, new_AGEMA_signal_9149, SubBytesIns_Inst_Sbox_5_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L15_U1 ( .a ({new_AGEMA_signal_8704, new_AGEMA_signal_8703, SubBytesIns_Inst_Sbox_5_M55}), .b ({new_AGEMA_signal_8712, new_AGEMA_signal_8711, SubBytesIns_Inst_Sbox_5_L1}), .c ({new_AGEMA_signal_9152, new_AGEMA_signal_9151, SubBytesIns_Inst_Sbox_5_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L16_U1 ( .a ({new_AGEMA_signal_8230, new_AGEMA_signal_8229, SubBytesIns_Inst_Sbox_5_M56}), .b ({new_AGEMA_signal_9520, new_AGEMA_signal_9519, SubBytesIns_Inst_Sbox_5_L0}), .c ({new_AGEMA_signal_9918, new_AGEMA_signal_9917, SubBytesIns_Inst_Sbox_5_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L17_U1 ( .a ({new_AGEMA_signal_8232, new_AGEMA_signal_8231, SubBytesIns_Inst_Sbox_5_M57}), .b ({new_AGEMA_signal_8712, new_AGEMA_signal_8711, SubBytesIns_Inst_Sbox_5_L1}), .c ({new_AGEMA_signal_9154, new_AGEMA_signal_9153, SubBytesIns_Inst_Sbox_5_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L18_U1 ( .a ({new_AGEMA_signal_8706, new_AGEMA_signal_8705, SubBytesIns_Inst_Sbox_5_M58}), .b ({new_AGEMA_signal_8714, new_AGEMA_signal_8713, SubBytesIns_Inst_Sbox_5_L8}), .c ({new_AGEMA_signal_9156, new_AGEMA_signal_9155, SubBytesIns_Inst_Sbox_5_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L19_U1 ( .a ({new_AGEMA_signal_8710, new_AGEMA_signal_8709, SubBytesIns_Inst_Sbox_5_M63}), .b ({new_AGEMA_signal_9146, new_AGEMA_signal_9145, SubBytesIns_Inst_Sbox_5_L4}), .c ({new_AGEMA_signal_9532, new_AGEMA_signal_9531, SubBytesIns_Inst_Sbox_5_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L20_U1 ( .a ({new_AGEMA_signal_9520, new_AGEMA_signal_9519, SubBytesIns_Inst_Sbox_5_L0}), .b ({new_AGEMA_signal_8712, new_AGEMA_signal_8711, SubBytesIns_Inst_Sbox_5_L1}), .c ({new_AGEMA_signal_9920, new_AGEMA_signal_9919, SubBytesIns_Inst_Sbox_5_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L21_U1 ( .a ({new_AGEMA_signal_8712, new_AGEMA_signal_8711, SubBytesIns_Inst_Sbox_5_L1}), .b ({new_AGEMA_signal_9524, new_AGEMA_signal_9523, SubBytesIns_Inst_Sbox_5_L7}), .c ({new_AGEMA_signal_9922, new_AGEMA_signal_9921, SubBytesIns_Inst_Sbox_5_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L22_U1 ( .a ({new_AGEMA_signal_9144, new_AGEMA_signal_9143, SubBytesIns_Inst_Sbox_5_L3}), .b ({new_AGEMA_signal_8716, new_AGEMA_signal_8715, SubBytesIns_Inst_Sbox_5_L12}), .c ({new_AGEMA_signal_9534, new_AGEMA_signal_9533, SubBytesIns_Inst_Sbox_5_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L23_U1 ( .a ({new_AGEMA_signal_9156, new_AGEMA_signal_9155, SubBytesIns_Inst_Sbox_5_L18}), .b ({new_AGEMA_signal_9142, new_AGEMA_signal_9141, SubBytesIns_Inst_Sbox_5_L2}), .c ({new_AGEMA_signal_9536, new_AGEMA_signal_9535, SubBytesIns_Inst_Sbox_5_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L24_U1 ( .a ({new_AGEMA_signal_9152, new_AGEMA_signal_9151, SubBytesIns_Inst_Sbox_5_L15}), .b ({new_AGEMA_signal_9526, new_AGEMA_signal_9525, SubBytesIns_Inst_Sbox_5_L9}), .c ({new_AGEMA_signal_9924, new_AGEMA_signal_9923, SubBytesIns_Inst_Sbox_5_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L25_U1 ( .a ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_9528, new_AGEMA_signal_9527, SubBytesIns_Inst_Sbox_5_L10}), .c ({new_AGEMA_signal_9926, new_AGEMA_signal_9925, SubBytesIns_Inst_Sbox_5_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L26_U1 ( .a ({new_AGEMA_signal_9524, new_AGEMA_signal_9523, SubBytesIns_Inst_Sbox_5_L7}), .b ({new_AGEMA_signal_9526, new_AGEMA_signal_9525, SubBytesIns_Inst_Sbox_5_L9}), .c ({new_AGEMA_signal_9928, new_AGEMA_signal_9927, SubBytesIns_Inst_Sbox_5_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L27_U1 ( .a ({new_AGEMA_signal_8714, new_AGEMA_signal_8713, SubBytesIns_Inst_Sbox_5_L8}), .b ({new_AGEMA_signal_9528, new_AGEMA_signal_9527, SubBytesIns_Inst_Sbox_5_L10}), .c ({new_AGEMA_signal_9930, new_AGEMA_signal_9929, SubBytesIns_Inst_Sbox_5_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L28_U1 ( .a ({new_AGEMA_signal_9530, new_AGEMA_signal_9529, SubBytesIns_Inst_Sbox_5_L11}), .b ({new_AGEMA_signal_9150, new_AGEMA_signal_9149, SubBytesIns_Inst_Sbox_5_L14}), .c ({new_AGEMA_signal_9932, new_AGEMA_signal_9931, SubBytesIns_Inst_Sbox_5_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L29_U1 ( .a ({new_AGEMA_signal_9530, new_AGEMA_signal_9529, SubBytesIns_Inst_Sbox_5_L11}), .b ({new_AGEMA_signal_9154, new_AGEMA_signal_9153, SubBytesIns_Inst_Sbox_5_L17}), .c ({new_AGEMA_signal_9934, new_AGEMA_signal_9933, SubBytesIns_Inst_Sbox_5_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S0_U1 ( .a ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_9924, new_AGEMA_signal_9923, SubBytesIns_Inst_Sbox_5_L24}), .c ({new_AGEMA_signal_10292, new_AGEMA_signal_10291, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S1_U1 ( .a ({new_AGEMA_signal_9918, new_AGEMA_signal_9917, SubBytesIns_Inst_Sbox_5_L16}), .b ({new_AGEMA_signal_9928, new_AGEMA_signal_9927, SubBytesIns_Inst_Sbox_5_L26}), .c ({new_AGEMA_signal_10294, new_AGEMA_signal_10293, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S2_U1 ( .a ({new_AGEMA_signal_9532, new_AGEMA_signal_9531, SubBytesIns_Inst_Sbox_5_L19}), .b ({new_AGEMA_signal_9932, new_AGEMA_signal_9931, SubBytesIns_Inst_Sbox_5_L28}), .c ({new_AGEMA_signal_10296, new_AGEMA_signal_10295, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S3_U1 ( .a ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_9922, new_AGEMA_signal_9921, SubBytesIns_Inst_Sbox_5_L21}), .c ({new_AGEMA_signal_10298, new_AGEMA_signal_10297, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S4_U1 ( .a ({new_AGEMA_signal_9920, new_AGEMA_signal_9919, SubBytesIns_Inst_Sbox_5_L20}), .b ({new_AGEMA_signal_9534, new_AGEMA_signal_9533, SubBytesIns_Inst_Sbox_5_L22}), .c ({new_AGEMA_signal_10300, new_AGEMA_signal_10299, MixColumnsInput[107]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S5_U1 ( .a ({new_AGEMA_signal_9926, new_AGEMA_signal_9925, SubBytesIns_Inst_Sbox_5_L25}), .b ({new_AGEMA_signal_9934, new_AGEMA_signal_9933, SubBytesIns_Inst_Sbox_5_L29}), .c ({new_AGEMA_signal_10302, new_AGEMA_signal_10301, MixColumnsInput[106]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S6_U1 ( .a ({new_AGEMA_signal_9916, new_AGEMA_signal_9915, SubBytesIns_Inst_Sbox_5_L13}), .b ({new_AGEMA_signal_9930, new_AGEMA_signal_9929, SubBytesIns_Inst_Sbox_5_L27}), .c ({new_AGEMA_signal_10304, new_AGEMA_signal_10303, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S7_U1 ( .a ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_9536, new_AGEMA_signal_9535, SubBytesIns_Inst_Sbox_5_L23}), .c ({new_AGEMA_signal_9936, new_AGEMA_signal_9935, MixColumnsInput[104]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M46_U1 ( .a ({new_AGEMA_signal_8244, new_AGEMA_signal_8243, SubBytesIns_Inst_Sbox_6_M44}), .b ({new_AGEMA_signal_5878, new_AGEMA_signal_5877, SubBytesIns_Inst_Sbox_6_T6}), .clk (clk), .r ({Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({new_AGEMA_signal_8720, new_AGEMA_signal_8719, SubBytesIns_Inst_Sbox_6_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M47_U1 ( .a ({new_AGEMA_signal_7924, new_AGEMA_signal_7923, SubBytesIns_Inst_Sbox_6_M40}), .b ({new_AGEMA_signal_6298, new_AGEMA_signal_6297, SubBytesIns_Inst_Sbox_6_T8}), .clk (clk), .r ({Fresh[1289], Fresh[1288], Fresh[1287]}), .c ({new_AGEMA_signal_8246, new_AGEMA_signal_8245, SubBytesIns_Inst_Sbox_6_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M48_U1 ( .a ({new_AGEMA_signal_7922, new_AGEMA_signal_7921, SubBytesIns_Inst_Sbox_6_M39}), .b ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .clk (clk), .r ({Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({new_AGEMA_signal_8248, new_AGEMA_signal_8247, SubBytesIns_Inst_Sbox_6_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M49_U1 ( .a ({new_AGEMA_signal_8242, new_AGEMA_signal_8241, SubBytesIns_Inst_Sbox_6_M43}), .b ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, SubBytesIns_Inst_Sbox_6_T16}), .clk (clk), .r ({Fresh[1295], Fresh[1294], Fresh[1293]}), .c ({new_AGEMA_signal_8722, new_AGEMA_signal_8721, SubBytesIns_Inst_Sbox_6_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M50_U1 ( .a ({new_AGEMA_signal_7920, new_AGEMA_signal_7919, SubBytesIns_Inst_Sbox_6_M38}), .b ({new_AGEMA_signal_5880, new_AGEMA_signal_5879, SubBytesIns_Inst_Sbox_6_T9}), .clk (clk), .r ({Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({new_AGEMA_signal_8250, new_AGEMA_signal_8249, SubBytesIns_Inst_Sbox_6_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M51_U1 ( .a ({new_AGEMA_signal_7918, new_AGEMA_signal_7917, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_6304, new_AGEMA_signal_6303, SubBytesIns_Inst_Sbox_6_T17}), .clk (clk), .r ({Fresh[1301], Fresh[1300], Fresh[1299]}), .c ({new_AGEMA_signal_8252, new_AGEMA_signal_8251, SubBytesIns_Inst_Sbox_6_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M52_U1 ( .a ({new_AGEMA_signal_8240, new_AGEMA_signal_8239, SubBytesIns_Inst_Sbox_6_M42}), .b ({new_AGEMA_signal_5884, new_AGEMA_signal_5883, SubBytesIns_Inst_Sbox_6_T15}), .clk (clk), .r ({Fresh[1304], Fresh[1303], Fresh[1302]}), .c ({new_AGEMA_signal_8724, new_AGEMA_signal_8723, SubBytesIns_Inst_Sbox_6_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M53_U1 ( .a ({new_AGEMA_signal_8718, new_AGEMA_signal_8717, SubBytesIns_Inst_Sbox_6_M45}), .b ({new_AGEMA_signal_5892, new_AGEMA_signal_5891, SubBytesIns_Inst_Sbox_6_T27}), .clk (clk), .r ({Fresh[1307], Fresh[1306], Fresh[1305]}), .c ({new_AGEMA_signal_9158, new_AGEMA_signal_9157, SubBytesIns_Inst_Sbox_6_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M54_U1 ( .a ({new_AGEMA_signal_8238, new_AGEMA_signal_8237, SubBytesIns_Inst_Sbox_6_M41}), .b ({new_AGEMA_signal_6300, new_AGEMA_signal_6299, SubBytesIns_Inst_Sbox_6_T10}), .clk (clk), .r ({Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({new_AGEMA_signal_8726, new_AGEMA_signal_8725, SubBytesIns_Inst_Sbox_6_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M55_U1 ( .a ({new_AGEMA_signal_8244, new_AGEMA_signal_8243, SubBytesIns_Inst_Sbox_6_M44}), .b ({new_AGEMA_signal_5882, new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_6_T13}), .clk (clk), .r ({Fresh[1313], Fresh[1312], Fresh[1311]}), .c ({new_AGEMA_signal_8728, new_AGEMA_signal_8727, SubBytesIns_Inst_Sbox_6_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M56_U1 ( .a ({new_AGEMA_signal_7924, new_AGEMA_signal_7923, SubBytesIns_Inst_Sbox_6_M40}), .b ({new_AGEMA_signal_6308, new_AGEMA_signal_6307, SubBytesIns_Inst_Sbox_6_T23}), .clk (clk), .r ({Fresh[1316], Fresh[1315], Fresh[1314]}), .c ({new_AGEMA_signal_8254, new_AGEMA_signal_8253, SubBytesIns_Inst_Sbox_6_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M57_U1 ( .a ({new_AGEMA_signal_7922, new_AGEMA_signal_7921, SubBytesIns_Inst_Sbox_6_M39}), .b ({new_AGEMA_signal_5888, new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_6_T19}), .clk (clk), .r ({Fresh[1319], Fresh[1318], Fresh[1317]}), .c ({new_AGEMA_signal_8256, new_AGEMA_signal_8255, SubBytesIns_Inst_Sbox_6_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M58_U1 ( .a ({new_AGEMA_signal_8242, new_AGEMA_signal_8241, SubBytesIns_Inst_Sbox_6_M43}), .b ({new_AGEMA_signal_5522, new_AGEMA_signal_5521, SubBytesIns_Inst_Sbox_6_T3}), .clk (clk), .r ({Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({new_AGEMA_signal_8730, new_AGEMA_signal_8729, SubBytesIns_Inst_Sbox_6_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M59_U1 ( .a ({new_AGEMA_signal_7920, new_AGEMA_signal_7919, SubBytesIns_Inst_Sbox_6_M38}), .b ({new_AGEMA_signal_5890, new_AGEMA_signal_5889, SubBytesIns_Inst_Sbox_6_T22}), .clk (clk), .r ({Fresh[1325], Fresh[1324], Fresh[1323]}), .c ({new_AGEMA_signal_8258, new_AGEMA_signal_8257, SubBytesIns_Inst_Sbox_6_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M60_U1 ( .a ({new_AGEMA_signal_7918, new_AGEMA_signal_7917, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_6306, new_AGEMA_signal_6305, SubBytesIns_Inst_Sbox_6_T20}), .clk (clk), .r ({Fresh[1328], Fresh[1327], Fresh[1326]}), .c ({new_AGEMA_signal_8260, new_AGEMA_signal_8259, SubBytesIns_Inst_Sbox_6_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M61_U1 ( .a ({new_AGEMA_signal_8240, new_AGEMA_signal_8239, SubBytesIns_Inst_Sbox_6_M42}), .b ({new_AGEMA_signal_5518, new_AGEMA_signal_5517, SubBytesIns_Inst_Sbox_6_T1}), .clk (clk), .r ({Fresh[1331], Fresh[1330], Fresh[1329]}), .c ({new_AGEMA_signal_8732, new_AGEMA_signal_8731, SubBytesIns_Inst_Sbox_6_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M62_U1 ( .a ({new_AGEMA_signal_8718, new_AGEMA_signal_8717, SubBytesIns_Inst_Sbox_6_M45}), .b ({new_AGEMA_signal_5524, new_AGEMA_signal_5523, SubBytesIns_Inst_Sbox_6_T4}), .clk (clk), .r ({Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({new_AGEMA_signal_9160, new_AGEMA_signal_9159, SubBytesIns_Inst_Sbox_6_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M63_U1 ( .a ({new_AGEMA_signal_8238, new_AGEMA_signal_8237, SubBytesIns_Inst_Sbox_6_M41}), .b ({new_AGEMA_signal_5520, new_AGEMA_signal_5519, SubBytesIns_Inst_Sbox_6_T2}), .clk (clk), .r ({Fresh[1337], Fresh[1336], Fresh[1335]}), .c ({new_AGEMA_signal_8734, new_AGEMA_signal_8733, SubBytesIns_Inst_Sbox_6_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L0_U1 ( .a ({new_AGEMA_signal_8732, new_AGEMA_signal_8731, SubBytesIns_Inst_Sbox_6_M61}), .b ({new_AGEMA_signal_9160, new_AGEMA_signal_9159, SubBytesIns_Inst_Sbox_6_M62}), .c ({new_AGEMA_signal_9538, new_AGEMA_signal_9537, SubBytesIns_Inst_Sbox_6_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L1_U1 ( .a ({new_AGEMA_signal_8250, new_AGEMA_signal_8249, SubBytesIns_Inst_Sbox_6_M50}), .b ({new_AGEMA_signal_8254, new_AGEMA_signal_8253, SubBytesIns_Inst_Sbox_6_M56}), .c ({new_AGEMA_signal_8736, new_AGEMA_signal_8735, SubBytesIns_Inst_Sbox_6_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L2_U1 ( .a ({new_AGEMA_signal_8720, new_AGEMA_signal_8719, SubBytesIns_Inst_Sbox_6_M46}), .b ({new_AGEMA_signal_8248, new_AGEMA_signal_8247, SubBytesIns_Inst_Sbox_6_M48}), .c ({new_AGEMA_signal_9162, new_AGEMA_signal_9161, SubBytesIns_Inst_Sbox_6_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L3_U1 ( .a ({new_AGEMA_signal_8246, new_AGEMA_signal_8245, SubBytesIns_Inst_Sbox_6_M47}), .b ({new_AGEMA_signal_8728, new_AGEMA_signal_8727, SubBytesIns_Inst_Sbox_6_M55}), .c ({new_AGEMA_signal_9164, new_AGEMA_signal_9163, SubBytesIns_Inst_Sbox_6_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L4_U1 ( .a ({new_AGEMA_signal_8726, new_AGEMA_signal_8725, SubBytesIns_Inst_Sbox_6_M54}), .b ({new_AGEMA_signal_8730, new_AGEMA_signal_8729, SubBytesIns_Inst_Sbox_6_M58}), .c ({new_AGEMA_signal_9166, new_AGEMA_signal_9165, SubBytesIns_Inst_Sbox_6_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L5_U1 ( .a ({new_AGEMA_signal_8722, new_AGEMA_signal_8721, SubBytesIns_Inst_Sbox_6_M49}), .b ({new_AGEMA_signal_8732, new_AGEMA_signal_8731, SubBytesIns_Inst_Sbox_6_M61}), .c ({new_AGEMA_signal_9168, new_AGEMA_signal_9167, SubBytesIns_Inst_Sbox_6_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L6_U1 ( .a ({new_AGEMA_signal_9160, new_AGEMA_signal_9159, SubBytesIns_Inst_Sbox_6_M62}), .b ({new_AGEMA_signal_9168, new_AGEMA_signal_9167, SubBytesIns_Inst_Sbox_6_L5}), .c ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, SubBytesIns_Inst_Sbox_6_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L7_U1 ( .a ({new_AGEMA_signal_8720, new_AGEMA_signal_8719, SubBytesIns_Inst_Sbox_6_M46}), .b ({new_AGEMA_signal_9164, new_AGEMA_signal_9163, SubBytesIns_Inst_Sbox_6_L3}), .c ({new_AGEMA_signal_9542, new_AGEMA_signal_9541, SubBytesIns_Inst_Sbox_6_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L8_U1 ( .a ({new_AGEMA_signal_8252, new_AGEMA_signal_8251, SubBytesIns_Inst_Sbox_6_M51}), .b ({new_AGEMA_signal_8258, new_AGEMA_signal_8257, SubBytesIns_Inst_Sbox_6_M59}), .c ({new_AGEMA_signal_8738, new_AGEMA_signal_8737, SubBytesIns_Inst_Sbox_6_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L9_U1 ( .a ({new_AGEMA_signal_8724, new_AGEMA_signal_8723, SubBytesIns_Inst_Sbox_6_M52}), .b ({new_AGEMA_signal_9158, new_AGEMA_signal_9157, SubBytesIns_Inst_Sbox_6_M53}), .c ({new_AGEMA_signal_9544, new_AGEMA_signal_9543, SubBytesIns_Inst_Sbox_6_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L10_U1 ( .a ({new_AGEMA_signal_9158, new_AGEMA_signal_9157, SubBytesIns_Inst_Sbox_6_M53}), .b ({new_AGEMA_signal_9166, new_AGEMA_signal_9165, SubBytesIns_Inst_Sbox_6_L4}), .c ({new_AGEMA_signal_9546, new_AGEMA_signal_9545, SubBytesIns_Inst_Sbox_6_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L11_U1 ( .a ({new_AGEMA_signal_8260, new_AGEMA_signal_8259, SubBytesIns_Inst_Sbox_6_M60}), .b ({new_AGEMA_signal_9162, new_AGEMA_signal_9161, SubBytesIns_Inst_Sbox_6_L2}), .c ({new_AGEMA_signal_9548, new_AGEMA_signal_9547, SubBytesIns_Inst_Sbox_6_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L12_U1 ( .a ({new_AGEMA_signal_8248, new_AGEMA_signal_8247, SubBytesIns_Inst_Sbox_6_M48}), .b ({new_AGEMA_signal_8252, new_AGEMA_signal_8251, SubBytesIns_Inst_Sbox_6_M51}), .c ({new_AGEMA_signal_8740, new_AGEMA_signal_8739, SubBytesIns_Inst_Sbox_6_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L13_U1 ( .a ({new_AGEMA_signal_8250, new_AGEMA_signal_8249, SubBytesIns_Inst_Sbox_6_M50}), .b ({new_AGEMA_signal_9538, new_AGEMA_signal_9537, SubBytesIns_Inst_Sbox_6_L0}), .c ({new_AGEMA_signal_9938, new_AGEMA_signal_9937, SubBytesIns_Inst_Sbox_6_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L14_U1 ( .a ({new_AGEMA_signal_8724, new_AGEMA_signal_8723, SubBytesIns_Inst_Sbox_6_M52}), .b ({new_AGEMA_signal_8732, new_AGEMA_signal_8731, SubBytesIns_Inst_Sbox_6_M61}), .c ({new_AGEMA_signal_9170, new_AGEMA_signal_9169, SubBytesIns_Inst_Sbox_6_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L15_U1 ( .a ({new_AGEMA_signal_8728, new_AGEMA_signal_8727, SubBytesIns_Inst_Sbox_6_M55}), .b ({new_AGEMA_signal_8736, new_AGEMA_signal_8735, SubBytesIns_Inst_Sbox_6_L1}), .c ({new_AGEMA_signal_9172, new_AGEMA_signal_9171, SubBytesIns_Inst_Sbox_6_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L16_U1 ( .a ({new_AGEMA_signal_8254, new_AGEMA_signal_8253, SubBytesIns_Inst_Sbox_6_M56}), .b ({new_AGEMA_signal_9538, new_AGEMA_signal_9537, SubBytesIns_Inst_Sbox_6_L0}), .c ({new_AGEMA_signal_9940, new_AGEMA_signal_9939, SubBytesIns_Inst_Sbox_6_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L17_U1 ( .a ({new_AGEMA_signal_8256, new_AGEMA_signal_8255, SubBytesIns_Inst_Sbox_6_M57}), .b ({new_AGEMA_signal_8736, new_AGEMA_signal_8735, SubBytesIns_Inst_Sbox_6_L1}), .c ({new_AGEMA_signal_9174, new_AGEMA_signal_9173, SubBytesIns_Inst_Sbox_6_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L18_U1 ( .a ({new_AGEMA_signal_8730, new_AGEMA_signal_8729, SubBytesIns_Inst_Sbox_6_M58}), .b ({new_AGEMA_signal_8738, new_AGEMA_signal_8737, SubBytesIns_Inst_Sbox_6_L8}), .c ({new_AGEMA_signal_9176, new_AGEMA_signal_9175, SubBytesIns_Inst_Sbox_6_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L19_U1 ( .a ({new_AGEMA_signal_8734, new_AGEMA_signal_8733, SubBytesIns_Inst_Sbox_6_M63}), .b ({new_AGEMA_signal_9166, new_AGEMA_signal_9165, SubBytesIns_Inst_Sbox_6_L4}), .c ({new_AGEMA_signal_9550, new_AGEMA_signal_9549, SubBytesIns_Inst_Sbox_6_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L20_U1 ( .a ({new_AGEMA_signal_9538, new_AGEMA_signal_9537, SubBytesIns_Inst_Sbox_6_L0}), .b ({new_AGEMA_signal_8736, new_AGEMA_signal_8735, SubBytesIns_Inst_Sbox_6_L1}), .c ({new_AGEMA_signal_9942, new_AGEMA_signal_9941, SubBytesIns_Inst_Sbox_6_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L21_U1 ( .a ({new_AGEMA_signal_8736, new_AGEMA_signal_8735, SubBytesIns_Inst_Sbox_6_L1}), .b ({new_AGEMA_signal_9542, new_AGEMA_signal_9541, SubBytesIns_Inst_Sbox_6_L7}), .c ({new_AGEMA_signal_9944, new_AGEMA_signal_9943, SubBytesIns_Inst_Sbox_6_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L22_U1 ( .a ({new_AGEMA_signal_9164, new_AGEMA_signal_9163, SubBytesIns_Inst_Sbox_6_L3}), .b ({new_AGEMA_signal_8740, new_AGEMA_signal_8739, SubBytesIns_Inst_Sbox_6_L12}), .c ({new_AGEMA_signal_9552, new_AGEMA_signal_9551, SubBytesIns_Inst_Sbox_6_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L23_U1 ( .a ({new_AGEMA_signal_9176, new_AGEMA_signal_9175, SubBytesIns_Inst_Sbox_6_L18}), .b ({new_AGEMA_signal_9162, new_AGEMA_signal_9161, SubBytesIns_Inst_Sbox_6_L2}), .c ({new_AGEMA_signal_9554, new_AGEMA_signal_9553, SubBytesIns_Inst_Sbox_6_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L24_U1 ( .a ({new_AGEMA_signal_9172, new_AGEMA_signal_9171, SubBytesIns_Inst_Sbox_6_L15}), .b ({new_AGEMA_signal_9544, new_AGEMA_signal_9543, SubBytesIns_Inst_Sbox_6_L9}), .c ({new_AGEMA_signal_9946, new_AGEMA_signal_9945, SubBytesIns_Inst_Sbox_6_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L25_U1 ( .a ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_9546, new_AGEMA_signal_9545, SubBytesIns_Inst_Sbox_6_L10}), .c ({new_AGEMA_signal_9948, new_AGEMA_signal_9947, SubBytesIns_Inst_Sbox_6_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L26_U1 ( .a ({new_AGEMA_signal_9542, new_AGEMA_signal_9541, SubBytesIns_Inst_Sbox_6_L7}), .b ({new_AGEMA_signal_9544, new_AGEMA_signal_9543, SubBytesIns_Inst_Sbox_6_L9}), .c ({new_AGEMA_signal_9950, new_AGEMA_signal_9949, SubBytesIns_Inst_Sbox_6_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L27_U1 ( .a ({new_AGEMA_signal_8738, new_AGEMA_signal_8737, SubBytesIns_Inst_Sbox_6_L8}), .b ({new_AGEMA_signal_9546, new_AGEMA_signal_9545, SubBytesIns_Inst_Sbox_6_L10}), .c ({new_AGEMA_signal_9952, new_AGEMA_signal_9951, SubBytesIns_Inst_Sbox_6_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L28_U1 ( .a ({new_AGEMA_signal_9548, new_AGEMA_signal_9547, SubBytesIns_Inst_Sbox_6_L11}), .b ({new_AGEMA_signal_9170, new_AGEMA_signal_9169, SubBytesIns_Inst_Sbox_6_L14}), .c ({new_AGEMA_signal_9954, new_AGEMA_signal_9953, SubBytesIns_Inst_Sbox_6_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L29_U1 ( .a ({new_AGEMA_signal_9548, new_AGEMA_signal_9547, SubBytesIns_Inst_Sbox_6_L11}), .b ({new_AGEMA_signal_9174, new_AGEMA_signal_9173, SubBytesIns_Inst_Sbox_6_L17}), .c ({new_AGEMA_signal_9956, new_AGEMA_signal_9955, SubBytesIns_Inst_Sbox_6_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S0_U1 ( .a ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_9946, new_AGEMA_signal_9945, SubBytesIns_Inst_Sbox_6_L24}), .c ({new_AGEMA_signal_10306, new_AGEMA_signal_10305, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S1_U1 ( .a ({new_AGEMA_signal_9940, new_AGEMA_signal_9939, SubBytesIns_Inst_Sbox_6_L16}), .b ({new_AGEMA_signal_9950, new_AGEMA_signal_9949, SubBytesIns_Inst_Sbox_6_L26}), .c ({new_AGEMA_signal_10308, new_AGEMA_signal_10307, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S2_U1 ( .a ({new_AGEMA_signal_9550, new_AGEMA_signal_9549, SubBytesIns_Inst_Sbox_6_L19}), .b ({new_AGEMA_signal_9954, new_AGEMA_signal_9953, SubBytesIns_Inst_Sbox_6_L28}), .c ({new_AGEMA_signal_10310, new_AGEMA_signal_10309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S3_U1 ( .a ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_9944, new_AGEMA_signal_9943, SubBytesIns_Inst_Sbox_6_L21}), .c ({new_AGEMA_signal_10312, new_AGEMA_signal_10311, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S4_U1 ( .a ({new_AGEMA_signal_9942, new_AGEMA_signal_9941, SubBytesIns_Inst_Sbox_6_L20}), .b ({new_AGEMA_signal_9552, new_AGEMA_signal_9551, SubBytesIns_Inst_Sbox_6_L22}), .c ({new_AGEMA_signal_10314, new_AGEMA_signal_10313, MixColumnsInput[83]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S5_U1 ( .a ({new_AGEMA_signal_9948, new_AGEMA_signal_9947, SubBytesIns_Inst_Sbox_6_L25}), .b ({new_AGEMA_signal_9956, new_AGEMA_signal_9955, SubBytesIns_Inst_Sbox_6_L29}), .c ({new_AGEMA_signal_10316, new_AGEMA_signal_10315, MixColumnsInput[82]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S6_U1 ( .a ({new_AGEMA_signal_9938, new_AGEMA_signal_9937, SubBytesIns_Inst_Sbox_6_L13}), .b ({new_AGEMA_signal_9952, new_AGEMA_signal_9951, SubBytesIns_Inst_Sbox_6_L27}), .c ({new_AGEMA_signal_10318, new_AGEMA_signal_10317, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S7_U1 ( .a ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_9554, new_AGEMA_signal_9553, SubBytesIns_Inst_Sbox_6_L23}), .c ({new_AGEMA_signal_9958, new_AGEMA_signal_9957, MixColumnsInput[80]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M46_U1 ( .a ({new_AGEMA_signal_8268, new_AGEMA_signal_8267, SubBytesIns_Inst_Sbox_7_M44}), .b ({new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_7_T6}), .clk (clk), .r ({Fresh[1340], Fresh[1339], Fresh[1338]}), .c ({new_AGEMA_signal_8744, new_AGEMA_signal_8743, SubBytesIns_Inst_Sbox_7_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M47_U1 ( .a ({new_AGEMA_signal_7932, new_AGEMA_signal_7931, SubBytesIns_Inst_Sbox_7_M40}), .b ({new_AGEMA_signal_6324, new_AGEMA_signal_6323, SubBytesIns_Inst_Sbox_7_T8}), .clk (clk), .r ({Fresh[1343], Fresh[1342], Fresh[1341]}), .c ({new_AGEMA_signal_8270, new_AGEMA_signal_8269, SubBytesIns_Inst_Sbox_7_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M48_U1 ( .a ({new_AGEMA_signal_7930, new_AGEMA_signal_7929, SubBytesIns_Inst_Sbox_7_M39}), .b ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .clk (clk), .r ({Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({new_AGEMA_signal_8272, new_AGEMA_signal_8271, SubBytesIns_Inst_Sbox_7_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M49_U1 ( .a ({new_AGEMA_signal_8266, new_AGEMA_signal_8265, SubBytesIns_Inst_Sbox_7_M43}), .b ({new_AGEMA_signal_5902, new_AGEMA_signal_5901, SubBytesIns_Inst_Sbox_7_T16}), .clk (clk), .r ({Fresh[1349], Fresh[1348], Fresh[1347]}), .c ({new_AGEMA_signal_8746, new_AGEMA_signal_8745, SubBytesIns_Inst_Sbox_7_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M50_U1 ( .a ({new_AGEMA_signal_7928, new_AGEMA_signal_7927, SubBytesIns_Inst_Sbox_7_M38}), .b ({new_AGEMA_signal_5896, new_AGEMA_signal_5895, SubBytesIns_Inst_Sbox_7_T9}), .clk (clk), .r ({Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({new_AGEMA_signal_8274, new_AGEMA_signal_8273, SubBytesIns_Inst_Sbox_7_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M51_U1 ( .a ({new_AGEMA_signal_7926, new_AGEMA_signal_7925, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_6330, new_AGEMA_signal_6329, SubBytesIns_Inst_Sbox_7_T17}), .clk (clk), .r ({Fresh[1355], Fresh[1354], Fresh[1353]}), .c ({new_AGEMA_signal_8276, new_AGEMA_signal_8275, SubBytesIns_Inst_Sbox_7_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M52_U1 ( .a ({new_AGEMA_signal_8264, new_AGEMA_signal_8263, SubBytesIns_Inst_Sbox_7_M42}), .b ({new_AGEMA_signal_5900, new_AGEMA_signal_5899, SubBytesIns_Inst_Sbox_7_T15}), .clk (clk), .r ({Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({new_AGEMA_signal_8748, new_AGEMA_signal_8747, SubBytesIns_Inst_Sbox_7_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M53_U1 ( .a ({new_AGEMA_signal_8742, new_AGEMA_signal_8741, SubBytesIns_Inst_Sbox_7_M45}), .b ({new_AGEMA_signal_5908, new_AGEMA_signal_5907, SubBytesIns_Inst_Sbox_7_T27}), .clk (clk), .r ({Fresh[1361], Fresh[1360], Fresh[1359]}), .c ({new_AGEMA_signal_9178, new_AGEMA_signal_9177, SubBytesIns_Inst_Sbox_7_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M54_U1 ( .a ({new_AGEMA_signal_8262, new_AGEMA_signal_8261, SubBytesIns_Inst_Sbox_7_M41}), .b ({new_AGEMA_signal_6326, new_AGEMA_signal_6325, SubBytesIns_Inst_Sbox_7_T10}), .clk (clk), .r ({Fresh[1364], Fresh[1363], Fresh[1362]}), .c ({new_AGEMA_signal_8750, new_AGEMA_signal_8749, SubBytesIns_Inst_Sbox_7_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M55_U1 ( .a ({new_AGEMA_signal_8268, new_AGEMA_signal_8267, SubBytesIns_Inst_Sbox_7_M44}), .b ({new_AGEMA_signal_5898, new_AGEMA_signal_5897, SubBytesIns_Inst_Sbox_7_T13}), .clk (clk), .r ({Fresh[1367], Fresh[1366], Fresh[1365]}), .c ({new_AGEMA_signal_8752, new_AGEMA_signal_8751, SubBytesIns_Inst_Sbox_7_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M56_U1 ( .a ({new_AGEMA_signal_7932, new_AGEMA_signal_7931, SubBytesIns_Inst_Sbox_7_M40}), .b ({new_AGEMA_signal_6334, new_AGEMA_signal_6333, SubBytesIns_Inst_Sbox_7_T23}), .clk (clk), .r ({Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({new_AGEMA_signal_8278, new_AGEMA_signal_8277, SubBytesIns_Inst_Sbox_7_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M57_U1 ( .a ({new_AGEMA_signal_7930, new_AGEMA_signal_7929, SubBytesIns_Inst_Sbox_7_M39}), .b ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, SubBytesIns_Inst_Sbox_7_T19}), .clk (clk), .r ({Fresh[1373], Fresh[1372], Fresh[1371]}), .c ({new_AGEMA_signal_8280, new_AGEMA_signal_8279, SubBytesIns_Inst_Sbox_7_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M58_U1 ( .a ({new_AGEMA_signal_8266, new_AGEMA_signal_8265, SubBytesIns_Inst_Sbox_7_M43}), .b ({new_AGEMA_signal_5542, new_AGEMA_signal_5541, SubBytesIns_Inst_Sbox_7_T3}), .clk (clk), .r ({Fresh[1376], Fresh[1375], Fresh[1374]}), .c ({new_AGEMA_signal_8754, new_AGEMA_signal_8753, SubBytesIns_Inst_Sbox_7_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M59_U1 ( .a ({new_AGEMA_signal_7928, new_AGEMA_signal_7927, SubBytesIns_Inst_Sbox_7_M38}), .b ({new_AGEMA_signal_5906, new_AGEMA_signal_5905, SubBytesIns_Inst_Sbox_7_T22}), .clk (clk), .r ({Fresh[1379], Fresh[1378], Fresh[1377]}), .c ({new_AGEMA_signal_8282, new_AGEMA_signal_8281, SubBytesIns_Inst_Sbox_7_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M60_U1 ( .a ({new_AGEMA_signal_7926, new_AGEMA_signal_7925, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_6332, new_AGEMA_signal_6331, SubBytesIns_Inst_Sbox_7_T20}), .clk (clk), .r ({Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({new_AGEMA_signal_8284, new_AGEMA_signal_8283, SubBytesIns_Inst_Sbox_7_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M61_U1 ( .a ({new_AGEMA_signal_8264, new_AGEMA_signal_8263, SubBytesIns_Inst_Sbox_7_M42}), .b ({new_AGEMA_signal_5538, new_AGEMA_signal_5537, SubBytesIns_Inst_Sbox_7_T1}), .clk (clk), .r ({Fresh[1385], Fresh[1384], Fresh[1383]}), .c ({new_AGEMA_signal_8756, new_AGEMA_signal_8755, SubBytesIns_Inst_Sbox_7_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M62_U1 ( .a ({new_AGEMA_signal_8742, new_AGEMA_signal_8741, SubBytesIns_Inst_Sbox_7_M45}), .b ({new_AGEMA_signal_5544, new_AGEMA_signal_5543, SubBytesIns_Inst_Sbox_7_T4}), .clk (clk), .r ({Fresh[1388], Fresh[1387], Fresh[1386]}), .c ({new_AGEMA_signal_9180, new_AGEMA_signal_9179, SubBytesIns_Inst_Sbox_7_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M63_U1 ( .a ({new_AGEMA_signal_8262, new_AGEMA_signal_8261, SubBytesIns_Inst_Sbox_7_M41}), .b ({new_AGEMA_signal_5540, new_AGEMA_signal_5539, SubBytesIns_Inst_Sbox_7_T2}), .clk (clk), .r ({Fresh[1391], Fresh[1390], Fresh[1389]}), .c ({new_AGEMA_signal_8758, new_AGEMA_signal_8757, SubBytesIns_Inst_Sbox_7_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L0_U1 ( .a ({new_AGEMA_signal_8756, new_AGEMA_signal_8755, SubBytesIns_Inst_Sbox_7_M61}), .b ({new_AGEMA_signal_9180, new_AGEMA_signal_9179, SubBytesIns_Inst_Sbox_7_M62}), .c ({new_AGEMA_signal_9556, new_AGEMA_signal_9555, SubBytesIns_Inst_Sbox_7_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L1_U1 ( .a ({new_AGEMA_signal_8274, new_AGEMA_signal_8273, SubBytesIns_Inst_Sbox_7_M50}), .b ({new_AGEMA_signal_8278, new_AGEMA_signal_8277, SubBytesIns_Inst_Sbox_7_M56}), .c ({new_AGEMA_signal_8760, new_AGEMA_signal_8759, SubBytesIns_Inst_Sbox_7_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L2_U1 ( .a ({new_AGEMA_signal_8744, new_AGEMA_signal_8743, SubBytesIns_Inst_Sbox_7_M46}), .b ({new_AGEMA_signal_8272, new_AGEMA_signal_8271, SubBytesIns_Inst_Sbox_7_M48}), .c ({new_AGEMA_signal_9182, new_AGEMA_signal_9181, SubBytesIns_Inst_Sbox_7_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L3_U1 ( .a ({new_AGEMA_signal_8270, new_AGEMA_signal_8269, SubBytesIns_Inst_Sbox_7_M47}), .b ({new_AGEMA_signal_8752, new_AGEMA_signal_8751, SubBytesIns_Inst_Sbox_7_M55}), .c ({new_AGEMA_signal_9184, new_AGEMA_signal_9183, SubBytesIns_Inst_Sbox_7_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L4_U1 ( .a ({new_AGEMA_signal_8750, new_AGEMA_signal_8749, SubBytesIns_Inst_Sbox_7_M54}), .b ({new_AGEMA_signal_8754, new_AGEMA_signal_8753, SubBytesIns_Inst_Sbox_7_M58}), .c ({new_AGEMA_signal_9186, new_AGEMA_signal_9185, SubBytesIns_Inst_Sbox_7_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L5_U1 ( .a ({new_AGEMA_signal_8746, new_AGEMA_signal_8745, SubBytesIns_Inst_Sbox_7_M49}), .b ({new_AGEMA_signal_8756, new_AGEMA_signal_8755, SubBytesIns_Inst_Sbox_7_M61}), .c ({new_AGEMA_signal_9188, new_AGEMA_signal_9187, SubBytesIns_Inst_Sbox_7_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L6_U1 ( .a ({new_AGEMA_signal_9180, new_AGEMA_signal_9179, SubBytesIns_Inst_Sbox_7_M62}), .b ({new_AGEMA_signal_9188, new_AGEMA_signal_9187, SubBytesIns_Inst_Sbox_7_L5}), .c ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, SubBytesIns_Inst_Sbox_7_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L7_U1 ( .a ({new_AGEMA_signal_8744, new_AGEMA_signal_8743, SubBytesIns_Inst_Sbox_7_M46}), .b ({new_AGEMA_signal_9184, new_AGEMA_signal_9183, SubBytesIns_Inst_Sbox_7_L3}), .c ({new_AGEMA_signal_9560, new_AGEMA_signal_9559, SubBytesIns_Inst_Sbox_7_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L8_U1 ( .a ({new_AGEMA_signal_8276, new_AGEMA_signal_8275, SubBytesIns_Inst_Sbox_7_M51}), .b ({new_AGEMA_signal_8282, new_AGEMA_signal_8281, SubBytesIns_Inst_Sbox_7_M59}), .c ({new_AGEMA_signal_8762, new_AGEMA_signal_8761, SubBytesIns_Inst_Sbox_7_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L9_U1 ( .a ({new_AGEMA_signal_8748, new_AGEMA_signal_8747, SubBytesIns_Inst_Sbox_7_M52}), .b ({new_AGEMA_signal_9178, new_AGEMA_signal_9177, SubBytesIns_Inst_Sbox_7_M53}), .c ({new_AGEMA_signal_9562, new_AGEMA_signal_9561, SubBytesIns_Inst_Sbox_7_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L10_U1 ( .a ({new_AGEMA_signal_9178, new_AGEMA_signal_9177, SubBytesIns_Inst_Sbox_7_M53}), .b ({new_AGEMA_signal_9186, new_AGEMA_signal_9185, SubBytesIns_Inst_Sbox_7_L4}), .c ({new_AGEMA_signal_9564, new_AGEMA_signal_9563, SubBytesIns_Inst_Sbox_7_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L11_U1 ( .a ({new_AGEMA_signal_8284, new_AGEMA_signal_8283, SubBytesIns_Inst_Sbox_7_M60}), .b ({new_AGEMA_signal_9182, new_AGEMA_signal_9181, SubBytesIns_Inst_Sbox_7_L2}), .c ({new_AGEMA_signal_9566, new_AGEMA_signal_9565, SubBytesIns_Inst_Sbox_7_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L12_U1 ( .a ({new_AGEMA_signal_8272, new_AGEMA_signal_8271, SubBytesIns_Inst_Sbox_7_M48}), .b ({new_AGEMA_signal_8276, new_AGEMA_signal_8275, SubBytesIns_Inst_Sbox_7_M51}), .c ({new_AGEMA_signal_8764, new_AGEMA_signal_8763, SubBytesIns_Inst_Sbox_7_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L13_U1 ( .a ({new_AGEMA_signal_8274, new_AGEMA_signal_8273, SubBytesIns_Inst_Sbox_7_M50}), .b ({new_AGEMA_signal_9556, new_AGEMA_signal_9555, SubBytesIns_Inst_Sbox_7_L0}), .c ({new_AGEMA_signal_9960, new_AGEMA_signal_9959, SubBytesIns_Inst_Sbox_7_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L14_U1 ( .a ({new_AGEMA_signal_8748, new_AGEMA_signal_8747, SubBytesIns_Inst_Sbox_7_M52}), .b ({new_AGEMA_signal_8756, new_AGEMA_signal_8755, SubBytesIns_Inst_Sbox_7_M61}), .c ({new_AGEMA_signal_9190, new_AGEMA_signal_9189, SubBytesIns_Inst_Sbox_7_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L15_U1 ( .a ({new_AGEMA_signal_8752, new_AGEMA_signal_8751, SubBytesIns_Inst_Sbox_7_M55}), .b ({new_AGEMA_signal_8760, new_AGEMA_signal_8759, SubBytesIns_Inst_Sbox_7_L1}), .c ({new_AGEMA_signal_9192, new_AGEMA_signal_9191, SubBytesIns_Inst_Sbox_7_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L16_U1 ( .a ({new_AGEMA_signal_8278, new_AGEMA_signal_8277, SubBytesIns_Inst_Sbox_7_M56}), .b ({new_AGEMA_signal_9556, new_AGEMA_signal_9555, SubBytesIns_Inst_Sbox_7_L0}), .c ({new_AGEMA_signal_9962, new_AGEMA_signal_9961, SubBytesIns_Inst_Sbox_7_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L17_U1 ( .a ({new_AGEMA_signal_8280, new_AGEMA_signal_8279, SubBytesIns_Inst_Sbox_7_M57}), .b ({new_AGEMA_signal_8760, new_AGEMA_signal_8759, SubBytesIns_Inst_Sbox_7_L1}), .c ({new_AGEMA_signal_9194, new_AGEMA_signal_9193, SubBytesIns_Inst_Sbox_7_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L18_U1 ( .a ({new_AGEMA_signal_8754, new_AGEMA_signal_8753, SubBytesIns_Inst_Sbox_7_M58}), .b ({new_AGEMA_signal_8762, new_AGEMA_signal_8761, SubBytesIns_Inst_Sbox_7_L8}), .c ({new_AGEMA_signal_9196, new_AGEMA_signal_9195, SubBytesIns_Inst_Sbox_7_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L19_U1 ( .a ({new_AGEMA_signal_8758, new_AGEMA_signal_8757, SubBytesIns_Inst_Sbox_7_M63}), .b ({new_AGEMA_signal_9186, new_AGEMA_signal_9185, SubBytesIns_Inst_Sbox_7_L4}), .c ({new_AGEMA_signal_9568, new_AGEMA_signal_9567, SubBytesIns_Inst_Sbox_7_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L20_U1 ( .a ({new_AGEMA_signal_9556, new_AGEMA_signal_9555, SubBytesIns_Inst_Sbox_7_L0}), .b ({new_AGEMA_signal_8760, new_AGEMA_signal_8759, SubBytesIns_Inst_Sbox_7_L1}), .c ({new_AGEMA_signal_9964, new_AGEMA_signal_9963, SubBytesIns_Inst_Sbox_7_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L21_U1 ( .a ({new_AGEMA_signal_8760, new_AGEMA_signal_8759, SubBytesIns_Inst_Sbox_7_L1}), .b ({new_AGEMA_signal_9560, new_AGEMA_signal_9559, SubBytesIns_Inst_Sbox_7_L7}), .c ({new_AGEMA_signal_9966, new_AGEMA_signal_9965, SubBytesIns_Inst_Sbox_7_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L22_U1 ( .a ({new_AGEMA_signal_9184, new_AGEMA_signal_9183, SubBytesIns_Inst_Sbox_7_L3}), .b ({new_AGEMA_signal_8764, new_AGEMA_signal_8763, SubBytesIns_Inst_Sbox_7_L12}), .c ({new_AGEMA_signal_9570, new_AGEMA_signal_9569, SubBytesIns_Inst_Sbox_7_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L23_U1 ( .a ({new_AGEMA_signal_9196, new_AGEMA_signal_9195, SubBytesIns_Inst_Sbox_7_L18}), .b ({new_AGEMA_signal_9182, new_AGEMA_signal_9181, SubBytesIns_Inst_Sbox_7_L2}), .c ({new_AGEMA_signal_9572, new_AGEMA_signal_9571, SubBytesIns_Inst_Sbox_7_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L24_U1 ( .a ({new_AGEMA_signal_9192, new_AGEMA_signal_9191, SubBytesIns_Inst_Sbox_7_L15}), .b ({new_AGEMA_signal_9562, new_AGEMA_signal_9561, SubBytesIns_Inst_Sbox_7_L9}), .c ({new_AGEMA_signal_9968, new_AGEMA_signal_9967, SubBytesIns_Inst_Sbox_7_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L25_U1 ( .a ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_9564, new_AGEMA_signal_9563, SubBytesIns_Inst_Sbox_7_L10}), .c ({new_AGEMA_signal_9970, new_AGEMA_signal_9969, SubBytesIns_Inst_Sbox_7_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L26_U1 ( .a ({new_AGEMA_signal_9560, new_AGEMA_signal_9559, SubBytesIns_Inst_Sbox_7_L7}), .b ({new_AGEMA_signal_9562, new_AGEMA_signal_9561, SubBytesIns_Inst_Sbox_7_L9}), .c ({new_AGEMA_signal_9972, new_AGEMA_signal_9971, SubBytesIns_Inst_Sbox_7_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L27_U1 ( .a ({new_AGEMA_signal_8762, new_AGEMA_signal_8761, SubBytesIns_Inst_Sbox_7_L8}), .b ({new_AGEMA_signal_9564, new_AGEMA_signal_9563, SubBytesIns_Inst_Sbox_7_L10}), .c ({new_AGEMA_signal_9974, new_AGEMA_signal_9973, SubBytesIns_Inst_Sbox_7_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L28_U1 ( .a ({new_AGEMA_signal_9566, new_AGEMA_signal_9565, SubBytesIns_Inst_Sbox_7_L11}), .b ({new_AGEMA_signal_9190, new_AGEMA_signal_9189, SubBytesIns_Inst_Sbox_7_L14}), .c ({new_AGEMA_signal_9976, new_AGEMA_signal_9975, SubBytesIns_Inst_Sbox_7_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L29_U1 ( .a ({new_AGEMA_signal_9566, new_AGEMA_signal_9565, SubBytesIns_Inst_Sbox_7_L11}), .b ({new_AGEMA_signal_9194, new_AGEMA_signal_9193, SubBytesIns_Inst_Sbox_7_L17}), .c ({new_AGEMA_signal_9978, new_AGEMA_signal_9977, SubBytesIns_Inst_Sbox_7_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S0_U1 ( .a ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_9968, new_AGEMA_signal_9967, SubBytesIns_Inst_Sbox_7_L24}), .c ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S1_U1 ( .a ({new_AGEMA_signal_9962, new_AGEMA_signal_9961, SubBytesIns_Inst_Sbox_7_L16}), .b ({new_AGEMA_signal_9972, new_AGEMA_signal_9971, SubBytesIns_Inst_Sbox_7_L26}), .c ({new_AGEMA_signal_10322, new_AGEMA_signal_10321, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S2_U1 ( .a ({new_AGEMA_signal_9568, new_AGEMA_signal_9567, SubBytesIns_Inst_Sbox_7_L19}), .b ({new_AGEMA_signal_9976, new_AGEMA_signal_9975, SubBytesIns_Inst_Sbox_7_L28}), .c ({new_AGEMA_signal_10324, new_AGEMA_signal_10323, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S3_U1 ( .a ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_9966, new_AGEMA_signal_9965, SubBytesIns_Inst_Sbox_7_L21}), .c ({new_AGEMA_signal_10326, new_AGEMA_signal_10325, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S4_U1 ( .a ({new_AGEMA_signal_9964, new_AGEMA_signal_9963, SubBytesIns_Inst_Sbox_7_L20}), .b ({new_AGEMA_signal_9570, new_AGEMA_signal_9569, SubBytesIns_Inst_Sbox_7_L22}), .c ({new_AGEMA_signal_10328, new_AGEMA_signal_10327, MixColumnsInput[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S5_U1 ( .a ({new_AGEMA_signal_9970, new_AGEMA_signal_9969, SubBytesIns_Inst_Sbox_7_L25}), .b ({new_AGEMA_signal_9978, new_AGEMA_signal_9977, SubBytesIns_Inst_Sbox_7_L29}), .c ({new_AGEMA_signal_10330, new_AGEMA_signal_10329, MixColumnsInput[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S6_U1 ( .a ({new_AGEMA_signal_9960, new_AGEMA_signal_9959, SubBytesIns_Inst_Sbox_7_L13}), .b ({new_AGEMA_signal_9974, new_AGEMA_signal_9973, SubBytesIns_Inst_Sbox_7_L27}), .c ({new_AGEMA_signal_10332, new_AGEMA_signal_10331, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S7_U1 ( .a ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_9572, new_AGEMA_signal_9571, SubBytesIns_Inst_Sbox_7_L23}), .c ({new_AGEMA_signal_9980, new_AGEMA_signal_9979, MixColumnsInput[56]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M46_U1 ( .a ({new_AGEMA_signal_8292, new_AGEMA_signal_8291, SubBytesIns_Inst_Sbox_8_M44}), .b ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, SubBytesIns_Inst_Sbox_8_T6}), .clk (clk), .r ({Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({new_AGEMA_signal_8768, new_AGEMA_signal_8767, SubBytesIns_Inst_Sbox_8_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M47_U1 ( .a ({new_AGEMA_signal_7940, new_AGEMA_signal_7939, SubBytesIns_Inst_Sbox_8_M40}), .b ({new_AGEMA_signal_6350, new_AGEMA_signal_6349, SubBytesIns_Inst_Sbox_8_T8}), .clk (clk), .r ({Fresh[1397], Fresh[1396], Fresh[1395]}), .c ({new_AGEMA_signal_8294, new_AGEMA_signal_8293, SubBytesIns_Inst_Sbox_8_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M48_U1 ( .a ({new_AGEMA_signal_7938, new_AGEMA_signal_7937, SubBytesIns_Inst_Sbox_8_M39}), .b ({ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .clk (clk), .r ({Fresh[1400], Fresh[1399], Fresh[1398]}), .c ({new_AGEMA_signal_8296, new_AGEMA_signal_8295, SubBytesIns_Inst_Sbox_8_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M49_U1 ( .a ({new_AGEMA_signal_8290, new_AGEMA_signal_8289, SubBytesIns_Inst_Sbox_8_M43}), .b ({new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesIns_Inst_Sbox_8_T16}), .clk (clk), .r ({Fresh[1403], Fresh[1402], Fresh[1401]}), .c ({new_AGEMA_signal_8770, new_AGEMA_signal_8769, SubBytesIns_Inst_Sbox_8_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M50_U1 ( .a ({new_AGEMA_signal_7936, new_AGEMA_signal_7935, SubBytesIns_Inst_Sbox_8_M38}), .b ({new_AGEMA_signal_5912, new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_8_T9}), .clk (clk), .r ({Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({new_AGEMA_signal_8298, new_AGEMA_signal_8297, SubBytesIns_Inst_Sbox_8_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M51_U1 ( .a ({new_AGEMA_signal_7934, new_AGEMA_signal_7933, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_6356, new_AGEMA_signal_6355, SubBytesIns_Inst_Sbox_8_T17}), .clk (clk), .r ({Fresh[1409], Fresh[1408], Fresh[1407]}), .c ({new_AGEMA_signal_8300, new_AGEMA_signal_8299, SubBytesIns_Inst_Sbox_8_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M52_U1 ( .a ({new_AGEMA_signal_8288, new_AGEMA_signal_8287, SubBytesIns_Inst_Sbox_8_M42}), .b ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, SubBytesIns_Inst_Sbox_8_T15}), .clk (clk), .r ({Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({new_AGEMA_signal_8772, new_AGEMA_signal_8771, SubBytesIns_Inst_Sbox_8_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M53_U1 ( .a ({new_AGEMA_signal_8766, new_AGEMA_signal_8765, SubBytesIns_Inst_Sbox_8_M45}), .b ({new_AGEMA_signal_5924, new_AGEMA_signal_5923, SubBytesIns_Inst_Sbox_8_T27}), .clk (clk), .r ({Fresh[1415], Fresh[1414], Fresh[1413]}), .c ({new_AGEMA_signal_9198, new_AGEMA_signal_9197, SubBytesIns_Inst_Sbox_8_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M54_U1 ( .a ({new_AGEMA_signal_8286, new_AGEMA_signal_8285, SubBytesIns_Inst_Sbox_8_M41}), .b ({new_AGEMA_signal_6352, new_AGEMA_signal_6351, SubBytesIns_Inst_Sbox_8_T10}), .clk (clk), .r ({Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({new_AGEMA_signal_8774, new_AGEMA_signal_8773, SubBytesIns_Inst_Sbox_8_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M55_U1 ( .a ({new_AGEMA_signal_8292, new_AGEMA_signal_8291, SubBytesIns_Inst_Sbox_8_M44}), .b ({new_AGEMA_signal_5914, new_AGEMA_signal_5913, SubBytesIns_Inst_Sbox_8_T13}), .clk (clk), .r ({Fresh[1421], Fresh[1420], Fresh[1419]}), .c ({new_AGEMA_signal_8776, new_AGEMA_signal_8775, SubBytesIns_Inst_Sbox_8_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M56_U1 ( .a ({new_AGEMA_signal_7940, new_AGEMA_signal_7939, SubBytesIns_Inst_Sbox_8_M40}), .b ({new_AGEMA_signal_6360, new_AGEMA_signal_6359, SubBytesIns_Inst_Sbox_8_T23}), .clk (clk), .r ({Fresh[1424], Fresh[1423], Fresh[1422]}), .c ({new_AGEMA_signal_8302, new_AGEMA_signal_8301, SubBytesIns_Inst_Sbox_8_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M57_U1 ( .a ({new_AGEMA_signal_7938, new_AGEMA_signal_7937, SubBytesIns_Inst_Sbox_8_M39}), .b ({new_AGEMA_signal_5920, new_AGEMA_signal_5919, SubBytesIns_Inst_Sbox_8_T19}), .clk (clk), .r ({Fresh[1427], Fresh[1426], Fresh[1425]}), .c ({new_AGEMA_signal_8304, new_AGEMA_signal_8303, SubBytesIns_Inst_Sbox_8_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M58_U1 ( .a ({new_AGEMA_signal_8290, new_AGEMA_signal_8289, SubBytesIns_Inst_Sbox_8_M43}), .b ({new_AGEMA_signal_5562, new_AGEMA_signal_5561, SubBytesIns_Inst_Sbox_8_T3}), .clk (clk), .r ({Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({new_AGEMA_signal_8778, new_AGEMA_signal_8777, SubBytesIns_Inst_Sbox_8_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M59_U1 ( .a ({new_AGEMA_signal_7936, new_AGEMA_signal_7935, SubBytesIns_Inst_Sbox_8_M38}), .b ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, SubBytesIns_Inst_Sbox_8_T22}), .clk (clk), .r ({Fresh[1433], Fresh[1432], Fresh[1431]}), .c ({new_AGEMA_signal_8306, new_AGEMA_signal_8305, SubBytesIns_Inst_Sbox_8_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M60_U1 ( .a ({new_AGEMA_signal_7934, new_AGEMA_signal_7933, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_6358, new_AGEMA_signal_6357, SubBytesIns_Inst_Sbox_8_T20}), .clk (clk), .r ({Fresh[1436], Fresh[1435], Fresh[1434]}), .c ({new_AGEMA_signal_8308, new_AGEMA_signal_8307, SubBytesIns_Inst_Sbox_8_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M61_U1 ( .a ({new_AGEMA_signal_8288, new_AGEMA_signal_8287, SubBytesIns_Inst_Sbox_8_M42}), .b ({new_AGEMA_signal_5558, new_AGEMA_signal_5557, SubBytesIns_Inst_Sbox_8_T1}), .clk (clk), .r ({Fresh[1439], Fresh[1438], Fresh[1437]}), .c ({new_AGEMA_signal_8780, new_AGEMA_signal_8779, SubBytesIns_Inst_Sbox_8_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M62_U1 ( .a ({new_AGEMA_signal_8766, new_AGEMA_signal_8765, SubBytesIns_Inst_Sbox_8_M45}), .b ({new_AGEMA_signal_5564, new_AGEMA_signal_5563, SubBytesIns_Inst_Sbox_8_T4}), .clk (clk), .r ({Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({new_AGEMA_signal_9200, new_AGEMA_signal_9199, SubBytesIns_Inst_Sbox_8_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M63_U1 ( .a ({new_AGEMA_signal_8286, new_AGEMA_signal_8285, SubBytesIns_Inst_Sbox_8_M41}), .b ({new_AGEMA_signal_5560, new_AGEMA_signal_5559, SubBytesIns_Inst_Sbox_8_T2}), .clk (clk), .r ({Fresh[1445], Fresh[1444], Fresh[1443]}), .c ({new_AGEMA_signal_8782, new_AGEMA_signal_8781, SubBytesIns_Inst_Sbox_8_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L0_U1 ( .a ({new_AGEMA_signal_8780, new_AGEMA_signal_8779, SubBytesIns_Inst_Sbox_8_M61}), .b ({new_AGEMA_signal_9200, new_AGEMA_signal_9199, SubBytesIns_Inst_Sbox_8_M62}), .c ({new_AGEMA_signal_9574, new_AGEMA_signal_9573, SubBytesIns_Inst_Sbox_8_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L1_U1 ( .a ({new_AGEMA_signal_8298, new_AGEMA_signal_8297, SubBytesIns_Inst_Sbox_8_M50}), .b ({new_AGEMA_signal_8302, new_AGEMA_signal_8301, SubBytesIns_Inst_Sbox_8_M56}), .c ({new_AGEMA_signal_8784, new_AGEMA_signal_8783, SubBytesIns_Inst_Sbox_8_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L2_U1 ( .a ({new_AGEMA_signal_8768, new_AGEMA_signal_8767, SubBytesIns_Inst_Sbox_8_M46}), .b ({new_AGEMA_signal_8296, new_AGEMA_signal_8295, SubBytesIns_Inst_Sbox_8_M48}), .c ({new_AGEMA_signal_9202, new_AGEMA_signal_9201, SubBytesIns_Inst_Sbox_8_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L3_U1 ( .a ({new_AGEMA_signal_8294, new_AGEMA_signal_8293, SubBytesIns_Inst_Sbox_8_M47}), .b ({new_AGEMA_signal_8776, new_AGEMA_signal_8775, SubBytesIns_Inst_Sbox_8_M55}), .c ({new_AGEMA_signal_9204, new_AGEMA_signal_9203, SubBytesIns_Inst_Sbox_8_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L4_U1 ( .a ({new_AGEMA_signal_8774, new_AGEMA_signal_8773, SubBytesIns_Inst_Sbox_8_M54}), .b ({new_AGEMA_signal_8778, new_AGEMA_signal_8777, SubBytesIns_Inst_Sbox_8_M58}), .c ({new_AGEMA_signal_9206, new_AGEMA_signal_9205, SubBytesIns_Inst_Sbox_8_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L5_U1 ( .a ({new_AGEMA_signal_8770, new_AGEMA_signal_8769, SubBytesIns_Inst_Sbox_8_M49}), .b ({new_AGEMA_signal_8780, new_AGEMA_signal_8779, SubBytesIns_Inst_Sbox_8_M61}), .c ({new_AGEMA_signal_9208, new_AGEMA_signal_9207, SubBytesIns_Inst_Sbox_8_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L6_U1 ( .a ({new_AGEMA_signal_9200, new_AGEMA_signal_9199, SubBytesIns_Inst_Sbox_8_M62}), .b ({new_AGEMA_signal_9208, new_AGEMA_signal_9207, SubBytesIns_Inst_Sbox_8_L5}), .c ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, SubBytesIns_Inst_Sbox_8_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L7_U1 ( .a ({new_AGEMA_signal_8768, new_AGEMA_signal_8767, SubBytesIns_Inst_Sbox_8_M46}), .b ({new_AGEMA_signal_9204, new_AGEMA_signal_9203, SubBytesIns_Inst_Sbox_8_L3}), .c ({new_AGEMA_signal_9578, new_AGEMA_signal_9577, SubBytesIns_Inst_Sbox_8_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L8_U1 ( .a ({new_AGEMA_signal_8300, new_AGEMA_signal_8299, SubBytesIns_Inst_Sbox_8_M51}), .b ({new_AGEMA_signal_8306, new_AGEMA_signal_8305, SubBytesIns_Inst_Sbox_8_M59}), .c ({new_AGEMA_signal_8786, new_AGEMA_signal_8785, SubBytesIns_Inst_Sbox_8_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L9_U1 ( .a ({new_AGEMA_signal_8772, new_AGEMA_signal_8771, SubBytesIns_Inst_Sbox_8_M52}), .b ({new_AGEMA_signal_9198, new_AGEMA_signal_9197, SubBytesIns_Inst_Sbox_8_M53}), .c ({new_AGEMA_signal_9580, new_AGEMA_signal_9579, SubBytesIns_Inst_Sbox_8_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L10_U1 ( .a ({new_AGEMA_signal_9198, new_AGEMA_signal_9197, SubBytesIns_Inst_Sbox_8_M53}), .b ({new_AGEMA_signal_9206, new_AGEMA_signal_9205, SubBytesIns_Inst_Sbox_8_L4}), .c ({new_AGEMA_signal_9582, new_AGEMA_signal_9581, SubBytesIns_Inst_Sbox_8_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L11_U1 ( .a ({new_AGEMA_signal_8308, new_AGEMA_signal_8307, SubBytesIns_Inst_Sbox_8_M60}), .b ({new_AGEMA_signal_9202, new_AGEMA_signal_9201, SubBytesIns_Inst_Sbox_8_L2}), .c ({new_AGEMA_signal_9584, new_AGEMA_signal_9583, SubBytesIns_Inst_Sbox_8_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L12_U1 ( .a ({new_AGEMA_signal_8296, new_AGEMA_signal_8295, SubBytesIns_Inst_Sbox_8_M48}), .b ({new_AGEMA_signal_8300, new_AGEMA_signal_8299, SubBytesIns_Inst_Sbox_8_M51}), .c ({new_AGEMA_signal_8788, new_AGEMA_signal_8787, SubBytesIns_Inst_Sbox_8_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L13_U1 ( .a ({new_AGEMA_signal_8298, new_AGEMA_signal_8297, SubBytesIns_Inst_Sbox_8_M50}), .b ({new_AGEMA_signal_9574, new_AGEMA_signal_9573, SubBytesIns_Inst_Sbox_8_L0}), .c ({new_AGEMA_signal_9982, new_AGEMA_signal_9981, SubBytesIns_Inst_Sbox_8_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L14_U1 ( .a ({new_AGEMA_signal_8772, new_AGEMA_signal_8771, SubBytesIns_Inst_Sbox_8_M52}), .b ({new_AGEMA_signal_8780, new_AGEMA_signal_8779, SubBytesIns_Inst_Sbox_8_M61}), .c ({new_AGEMA_signal_9210, new_AGEMA_signal_9209, SubBytesIns_Inst_Sbox_8_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L15_U1 ( .a ({new_AGEMA_signal_8776, new_AGEMA_signal_8775, SubBytesIns_Inst_Sbox_8_M55}), .b ({new_AGEMA_signal_8784, new_AGEMA_signal_8783, SubBytesIns_Inst_Sbox_8_L1}), .c ({new_AGEMA_signal_9212, new_AGEMA_signal_9211, SubBytesIns_Inst_Sbox_8_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L16_U1 ( .a ({new_AGEMA_signal_8302, new_AGEMA_signal_8301, SubBytesIns_Inst_Sbox_8_M56}), .b ({new_AGEMA_signal_9574, new_AGEMA_signal_9573, SubBytesIns_Inst_Sbox_8_L0}), .c ({new_AGEMA_signal_9984, new_AGEMA_signal_9983, SubBytesIns_Inst_Sbox_8_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L17_U1 ( .a ({new_AGEMA_signal_8304, new_AGEMA_signal_8303, SubBytesIns_Inst_Sbox_8_M57}), .b ({new_AGEMA_signal_8784, new_AGEMA_signal_8783, SubBytesIns_Inst_Sbox_8_L1}), .c ({new_AGEMA_signal_9214, new_AGEMA_signal_9213, SubBytesIns_Inst_Sbox_8_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L18_U1 ( .a ({new_AGEMA_signal_8778, new_AGEMA_signal_8777, SubBytesIns_Inst_Sbox_8_M58}), .b ({new_AGEMA_signal_8786, new_AGEMA_signal_8785, SubBytesIns_Inst_Sbox_8_L8}), .c ({new_AGEMA_signal_9216, new_AGEMA_signal_9215, SubBytesIns_Inst_Sbox_8_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L19_U1 ( .a ({new_AGEMA_signal_8782, new_AGEMA_signal_8781, SubBytesIns_Inst_Sbox_8_M63}), .b ({new_AGEMA_signal_9206, new_AGEMA_signal_9205, SubBytesIns_Inst_Sbox_8_L4}), .c ({new_AGEMA_signal_9586, new_AGEMA_signal_9585, SubBytesIns_Inst_Sbox_8_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L20_U1 ( .a ({new_AGEMA_signal_9574, new_AGEMA_signal_9573, SubBytesIns_Inst_Sbox_8_L0}), .b ({new_AGEMA_signal_8784, new_AGEMA_signal_8783, SubBytesIns_Inst_Sbox_8_L1}), .c ({new_AGEMA_signal_9986, new_AGEMA_signal_9985, SubBytesIns_Inst_Sbox_8_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L21_U1 ( .a ({new_AGEMA_signal_8784, new_AGEMA_signal_8783, SubBytesIns_Inst_Sbox_8_L1}), .b ({new_AGEMA_signal_9578, new_AGEMA_signal_9577, SubBytesIns_Inst_Sbox_8_L7}), .c ({new_AGEMA_signal_9988, new_AGEMA_signal_9987, SubBytesIns_Inst_Sbox_8_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L22_U1 ( .a ({new_AGEMA_signal_9204, new_AGEMA_signal_9203, SubBytesIns_Inst_Sbox_8_L3}), .b ({new_AGEMA_signal_8788, new_AGEMA_signal_8787, SubBytesIns_Inst_Sbox_8_L12}), .c ({new_AGEMA_signal_9588, new_AGEMA_signal_9587, SubBytesIns_Inst_Sbox_8_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L23_U1 ( .a ({new_AGEMA_signal_9216, new_AGEMA_signal_9215, SubBytesIns_Inst_Sbox_8_L18}), .b ({new_AGEMA_signal_9202, new_AGEMA_signal_9201, SubBytesIns_Inst_Sbox_8_L2}), .c ({new_AGEMA_signal_9590, new_AGEMA_signal_9589, SubBytesIns_Inst_Sbox_8_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L24_U1 ( .a ({new_AGEMA_signal_9212, new_AGEMA_signal_9211, SubBytesIns_Inst_Sbox_8_L15}), .b ({new_AGEMA_signal_9580, new_AGEMA_signal_9579, SubBytesIns_Inst_Sbox_8_L9}), .c ({new_AGEMA_signal_9990, new_AGEMA_signal_9989, SubBytesIns_Inst_Sbox_8_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L25_U1 ( .a ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_9582, new_AGEMA_signal_9581, SubBytesIns_Inst_Sbox_8_L10}), .c ({new_AGEMA_signal_9992, new_AGEMA_signal_9991, SubBytesIns_Inst_Sbox_8_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L26_U1 ( .a ({new_AGEMA_signal_9578, new_AGEMA_signal_9577, SubBytesIns_Inst_Sbox_8_L7}), .b ({new_AGEMA_signal_9580, new_AGEMA_signal_9579, SubBytesIns_Inst_Sbox_8_L9}), .c ({new_AGEMA_signal_9994, new_AGEMA_signal_9993, SubBytesIns_Inst_Sbox_8_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L27_U1 ( .a ({new_AGEMA_signal_8786, new_AGEMA_signal_8785, SubBytesIns_Inst_Sbox_8_L8}), .b ({new_AGEMA_signal_9582, new_AGEMA_signal_9581, SubBytesIns_Inst_Sbox_8_L10}), .c ({new_AGEMA_signal_9996, new_AGEMA_signal_9995, SubBytesIns_Inst_Sbox_8_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L28_U1 ( .a ({new_AGEMA_signal_9584, new_AGEMA_signal_9583, SubBytesIns_Inst_Sbox_8_L11}), .b ({new_AGEMA_signal_9210, new_AGEMA_signal_9209, SubBytesIns_Inst_Sbox_8_L14}), .c ({new_AGEMA_signal_9998, new_AGEMA_signal_9997, SubBytesIns_Inst_Sbox_8_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L29_U1 ( .a ({new_AGEMA_signal_9584, new_AGEMA_signal_9583, SubBytesIns_Inst_Sbox_8_L11}), .b ({new_AGEMA_signal_9214, new_AGEMA_signal_9213, SubBytesIns_Inst_Sbox_8_L17}), .c ({new_AGEMA_signal_10000, new_AGEMA_signal_9999, SubBytesIns_Inst_Sbox_8_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S0_U1 ( .a ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_9990, new_AGEMA_signal_9989, SubBytesIns_Inst_Sbox_8_L24}), .c ({new_AGEMA_signal_10334, new_AGEMA_signal_10333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S1_U1 ( .a ({new_AGEMA_signal_9984, new_AGEMA_signal_9983, SubBytesIns_Inst_Sbox_8_L16}), .b ({new_AGEMA_signal_9994, new_AGEMA_signal_9993, SubBytesIns_Inst_Sbox_8_L26}), .c ({new_AGEMA_signal_10336, new_AGEMA_signal_10335, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S2_U1 ( .a ({new_AGEMA_signal_9586, new_AGEMA_signal_9585, SubBytesIns_Inst_Sbox_8_L19}), .b ({new_AGEMA_signal_9998, new_AGEMA_signal_9997, SubBytesIns_Inst_Sbox_8_L28}), .c ({new_AGEMA_signal_10338, new_AGEMA_signal_10337, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S3_U1 ( .a ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_9988, new_AGEMA_signal_9987, SubBytesIns_Inst_Sbox_8_L21}), .c ({new_AGEMA_signal_10340, new_AGEMA_signal_10339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S4_U1 ( .a ({new_AGEMA_signal_9986, new_AGEMA_signal_9985, SubBytesIns_Inst_Sbox_8_L20}), .b ({new_AGEMA_signal_9588, new_AGEMA_signal_9587, SubBytesIns_Inst_Sbox_8_L22}), .c ({new_AGEMA_signal_10342, new_AGEMA_signal_10341, MixColumnsInput[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S5_U1 ( .a ({new_AGEMA_signal_9992, new_AGEMA_signal_9991, SubBytesIns_Inst_Sbox_8_L25}), .b ({new_AGEMA_signal_10000, new_AGEMA_signal_9999, SubBytesIns_Inst_Sbox_8_L29}), .c ({new_AGEMA_signal_10344, new_AGEMA_signal_10343, MixColumnsInput[34]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S6_U1 ( .a ({new_AGEMA_signal_9982, new_AGEMA_signal_9981, SubBytesIns_Inst_Sbox_8_L13}), .b ({new_AGEMA_signal_9996, new_AGEMA_signal_9995, SubBytesIns_Inst_Sbox_8_L27}), .c ({new_AGEMA_signal_10346, new_AGEMA_signal_10345, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S7_U1 ( .a ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_9590, new_AGEMA_signal_9589, SubBytesIns_Inst_Sbox_8_L23}), .c ({new_AGEMA_signal_10002, new_AGEMA_signal_10001, MixColumnsInput[32]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M46_U1 ( .a ({new_AGEMA_signal_8316, new_AGEMA_signal_8315, SubBytesIns_Inst_Sbox_9_M44}), .b ({new_AGEMA_signal_5926, new_AGEMA_signal_5925, SubBytesIns_Inst_Sbox_9_T6}), .clk (clk), .r ({Fresh[1448], Fresh[1447], Fresh[1446]}), .c ({new_AGEMA_signal_8792, new_AGEMA_signal_8791, SubBytesIns_Inst_Sbox_9_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M47_U1 ( .a ({new_AGEMA_signal_7948, new_AGEMA_signal_7947, SubBytesIns_Inst_Sbox_9_M40}), .b ({new_AGEMA_signal_6376, new_AGEMA_signal_6375, SubBytesIns_Inst_Sbox_9_T8}), .clk (clk), .r ({Fresh[1451], Fresh[1450], Fresh[1449]}), .c ({new_AGEMA_signal_8318, new_AGEMA_signal_8317, SubBytesIns_Inst_Sbox_9_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M48_U1 ( .a ({new_AGEMA_signal_7946, new_AGEMA_signal_7945, SubBytesIns_Inst_Sbox_9_M39}), .b ({ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .clk (clk), .r ({Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({new_AGEMA_signal_8320, new_AGEMA_signal_8319, SubBytesIns_Inst_Sbox_9_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M49_U1 ( .a ({new_AGEMA_signal_8314, new_AGEMA_signal_8313, SubBytesIns_Inst_Sbox_9_M43}), .b ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, SubBytesIns_Inst_Sbox_9_T16}), .clk (clk), .r ({Fresh[1457], Fresh[1456], Fresh[1455]}), .c ({new_AGEMA_signal_8794, new_AGEMA_signal_8793, SubBytesIns_Inst_Sbox_9_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M50_U1 ( .a ({new_AGEMA_signal_7944, new_AGEMA_signal_7943, SubBytesIns_Inst_Sbox_9_M38}), .b ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, SubBytesIns_Inst_Sbox_9_T9}), .clk (clk), .r ({Fresh[1460], Fresh[1459], Fresh[1458]}), .c ({new_AGEMA_signal_8322, new_AGEMA_signal_8321, SubBytesIns_Inst_Sbox_9_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M51_U1 ( .a ({new_AGEMA_signal_7942, new_AGEMA_signal_7941, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_6382, new_AGEMA_signal_6381, SubBytesIns_Inst_Sbox_9_T17}), .clk (clk), .r ({Fresh[1463], Fresh[1462], Fresh[1461]}), .c ({new_AGEMA_signal_8324, new_AGEMA_signal_8323, SubBytesIns_Inst_Sbox_9_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M52_U1 ( .a ({new_AGEMA_signal_8312, new_AGEMA_signal_8311, SubBytesIns_Inst_Sbox_9_M42}), .b ({new_AGEMA_signal_5932, new_AGEMA_signal_5931, SubBytesIns_Inst_Sbox_9_T15}), .clk (clk), .r ({Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({new_AGEMA_signal_8796, new_AGEMA_signal_8795, SubBytesIns_Inst_Sbox_9_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M53_U1 ( .a ({new_AGEMA_signal_8790, new_AGEMA_signal_8789, SubBytesIns_Inst_Sbox_9_M45}), .b ({new_AGEMA_signal_5940, new_AGEMA_signal_5939, SubBytesIns_Inst_Sbox_9_T27}), .clk (clk), .r ({Fresh[1469], Fresh[1468], Fresh[1467]}), .c ({new_AGEMA_signal_9218, new_AGEMA_signal_9217, SubBytesIns_Inst_Sbox_9_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M54_U1 ( .a ({new_AGEMA_signal_8310, new_AGEMA_signal_8309, SubBytesIns_Inst_Sbox_9_M41}), .b ({new_AGEMA_signal_6378, new_AGEMA_signal_6377, SubBytesIns_Inst_Sbox_9_T10}), .clk (clk), .r ({Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({new_AGEMA_signal_8798, new_AGEMA_signal_8797, SubBytesIns_Inst_Sbox_9_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M55_U1 ( .a ({new_AGEMA_signal_8316, new_AGEMA_signal_8315, SubBytesIns_Inst_Sbox_9_M44}), .b ({new_AGEMA_signal_5930, new_AGEMA_signal_5929, SubBytesIns_Inst_Sbox_9_T13}), .clk (clk), .r ({Fresh[1475], Fresh[1474], Fresh[1473]}), .c ({new_AGEMA_signal_8800, new_AGEMA_signal_8799, SubBytesIns_Inst_Sbox_9_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M56_U1 ( .a ({new_AGEMA_signal_7948, new_AGEMA_signal_7947, SubBytesIns_Inst_Sbox_9_M40}), .b ({new_AGEMA_signal_6386, new_AGEMA_signal_6385, SubBytesIns_Inst_Sbox_9_T23}), .clk (clk), .r ({Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({new_AGEMA_signal_8326, new_AGEMA_signal_8325, SubBytesIns_Inst_Sbox_9_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M57_U1 ( .a ({new_AGEMA_signal_7946, new_AGEMA_signal_7945, SubBytesIns_Inst_Sbox_9_M39}), .b ({new_AGEMA_signal_5936, new_AGEMA_signal_5935, SubBytesIns_Inst_Sbox_9_T19}), .clk (clk), .r ({Fresh[1481], Fresh[1480], Fresh[1479]}), .c ({new_AGEMA_signal_8328, new_AGEMA_signal_8327, SubBytesIns_Inst_Sbox_9_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M58_U1 ( .a ({new_AGEMA_signal_8314, new_AGEMA_signal_8313, SubBytesIns_Inst_Sbox_9_M43}), .b ({new_AGEMA_signal_5582, new_AGEMA_signal_5581, SubBytesIns_Inst_Sbox_9_T3}), .clk (clk), .r ({Fresh[1484], Fresh[1483], Fresh[1482]}), .c ({new_AGEMA_signal_8802, new_AGEMA_signal_8801, SubBytesIns_Inst_Sbox_9_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M59_U1 ( .a ({new_AGEMA_signal_7944, new_AGEMA_signal_7943, SubBytesIns_Inst_Sbox_9_M38}), .b ({new_AGEMA_signal_5938, new_AGEMA_signal_5937, SubBytesIns_Inst_Sbox_9_T22}), .clk (clk), .r ({Fresh[1487], Fresh[1486], Fresh[1485]}), .c ({new_AGEMA_signal_8330, new_AGEMA_signal_8329, SubBytesIns_Inst_Sbox_9_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M60_U1 ( .a ({new_AGEMA_signal_7942, new_AGEMA_signal_7941, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_6384, new_AGEMA_signal_6383, SubBytesIns_Inst_Sbox_9_T20}), .clk (clk), .r ({Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({new_AGEMA_signal_8332, new_AGEMA_signal_8331, SubBytesIns_Inst_Sbox_9_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M61_U1 ( .a ({new_AGEMA_signal_8312, new_AGEMA_signal_8311, SubBytesIns_Inst_Sbox_9_M42}), .b ({new_AGEMA_signal_5578, new_AGEMA_signal_5577, SubBytesIns_Inst_Sbox_9_T1}), .clk (clk), .r ({Fresh[1493], Fresh[1492], Fresh[1491]}), .c ({new_AGEMA_signal_8804, new_AGEMA_signal_8803, SubBytesIns_Inst_Sbox_9_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M62_U1 ( .a ({new_AGEMA_signal_8790, new_AGEMA_signal_8789, SubBytesIns_Inst_Sbox_9_M45}), .b ({new_AGEMA_signal_5584, new_AGEMA_signal_5583, SubBytesIns_Inst_Sbox_9_T4}), .clk (clk), .r ({Fresh[1496], Fresh[1495], Fresh[1494]}), .c ({new_AGEMA_signal_9220, new_AGEMA_signal_9219, SubBytesIns_Inst_Sbox_9_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M63_U1 ( .a ({new_AGEMA_signal_8310, new_AGEMA_signal_8309, SubBytesIns_Inst_Sbox_9_M41}), .b ({new_AGEMA_signal_5580, new_AGEMA_signal_5579, SubBytesIns_Inst_Sbox_9_T2}), .clk (clk), .r ({Fresh[1499], Fresh[1498], Fresh[1497]}), .c ({new_AGEMA_signal_8806, new_AGEMA_signal_8805, SubBytesIns_Inst_Sbox_9_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L0_U1 ( .a ({new_AGEMA_signal_8804, new_AGEMA_signal_8803, SubBytesIns_Inst_Sbox_9_M61}), .b ({new_AGEMA_signal_9220, new_AGEMA_signal_9219, SubBytesIns_Inst_Sbox_9_M62}), .c ({new_AGEMA_signal_9592, new_AGEMA_signal_9591, SubBytesIns_Inst_Sbox_9_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L1_U1 ( .a ({new_AGEMA_signal_8322, new_AGEMA_signal_8321, SubBytesIns_Inst_Sbox_9_M50}), .b ({new_AGEMA_signal_8326, new_AGEMA_signal_8325, SubBytesIns_Inst_Sbox_9_M56}), .c ({new_AGEMA_signal_8808, new_AGEMA_signal_8807, SubBytesIns_Inst_Sbox_9_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L2_U1 ( .a ({new_AGEMA_signal_8792, new_AGEMA_signal_8791, SubBytesIns_Inst_Sbox_9_M46}), .b ({new_AGEMA_signal_8320, new_AGEMA_signal_8319, SubBytesIns_Inst_Sbox_9_M48}), .c ({new_AGEMA_signal_9222, new_AGEMA_signal_9221, SubBytesIns_Inst_Sbox_9_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L3_U1 ( .a ({new_AGEMA_signal_8318, new_AGEMA_signal_8317, SubBytesIns_Inst_Sbox_9_M47}), .b ({new_AGEMA_signal_8800, new_AGEMA_signal_8799, SubBytesIns_Inst_Sbox_9_M55}), .c ({new_AGEMA_signal_9224, new_AGEMA_signal_9223, SubBytesIns_Inst_Sbox_9_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L4_U1 ( .a ({new_AGEMA_signal_8798, new_AGEMA_signal_8797, SubBytesIns_Inst_Sbox_9_M54}), .b ({new_AGEMA_signal_8802, new_AGEMA_signal_8801, SubBytesIns_Inst_Sbox_9_M58}), .c ({new_AGEMA_signal_9226, new_AGEMA_signal_9225, SubBytesIns_Inst_Sbox_9_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L5_U1 ( .a ({new_AGEMA_signal_8794, new_AGEMA_signal_8793, SubBytesIns_Inst_Sbox_9_M49}), .b ({new_AGEMA_signal_8804, new_AGEMA_signal_8803, SubBytesIns_Inst_Sbox_9_M61}), .c ({new_AGEMA_signal_9228, new_AGEMA_signal_9227, SubBytesIns_Inst_Sbox_9_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L6_U1 ( .a ({new_AGEMA_signal_9220, new_AGEMA_signal_9219, SubBytesIns_Inst_Sbox_9_M62}), .b ({new_AGEMA_signal_9228, new_AGEMA_signal_9227, SubBytesIns_Inst_Sbox_9_L5}), .c ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, SubBytesIns_Inst_Sbox_9_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L7_U1 ( .a ({new_AGEMA_signal_8792, new_AGEMA_signal_8791, SubBytesIns_Inst_Sbox_9_M46}), .b ({new_AGEMA_signal_9224, new_AGEMA_signal_9223, SubBytesIns_Inst_Sbox_9_L3}), .c ({new_AGEMA_signal_9596, new_AGEMA_signal_9595, SubBytesIns_Inst_Sbox_9_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L8_U1 ( .a ({new_AGEMA_signal_8324, new_AGEMA_signal_8323, SubBytesIns_Inst_Sbox_9_M51}), .b ({new_AGEMA_signal_8330, new_AGEMA_signal_8329, SubBytesIns_Inst_Sbox_9_M59}), .c ({new_AGEMA_signal_8810, new_AGEMA_signal_8809, SubBytesIns_Inst_Sbox_9_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L9_U1 ( .a ({new_AGEMA_signal_8796, new_AGEMA_signal_8795, SubBytesIns_Inst_Sbox_9_M52}), .b ({new_AGEMA_signal_9218, new_AGEMA_signal_9217, SubBytesIns_Inst_Sbox_9_M53}), .c ({new_AGEMA_signal_9598, new_AGEMA_signal_9597, SubBytesIns_Inst_Sbox_9_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L10_U1 ( .a ({new_AGEMA_signal_9218, new_AGEMA_signal_9217, SubBytesIns_Inst_Sbox_9_M53}), .b ({new_AGEMA_signal_9226, new_AGEMA_signal_9225, SubBytesIns_Inst_Sbox_9_L4}), .c ({new_AGEMA_signal_9600, new_AGEMA_signal_9599, SubBytesIns_Inst_Sbox_9_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L11_U1 ( .a ({new_AGEMA_signal_8332, new_AGEMA_signal_8331, SubBytesIns_Inst_Sbox_9_M60}), .b ({new_AGEMA_signal_9222, new_AGEMA_signal_9221, SubBytesIns_Inst_Sbox_9_L2}), .c ({new_AGEMA_signal_9602, new_AGEMA_signal_9601, SubBytesIns_Inst_Sbox_9_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L12_U1 ( .a ({new_AGEMA_signal_8320, new_AGEMA_signal_8319, SubBytesIns_Inst_Sbox_9_M48}), .b ({new_AGEMA_signal_8324, new_AGEMA_signal_8323, SubBytesIns_Inst_Sbox_9_M51}), .c ({new_AGEMA_signal_8812, new_AGEMA_signal_8811, SubBytesIns_Inst_Sbox_9_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L13_U1 ( .a ({new_AGEMA_signal_8322, new_AGEMA_signal_8321, SubBytesIns_Inst_Sbox_9_M50}), .b ({new_AGEMA_signal_9592, new_AGEMA_signal_9591, SubBytesIns_Inst_Sbox_9_L0}), .c ({new_AGEMA_signal_10004, new_AGEMA_signal_10003, SubBytesIns_Inst_Sbox_9_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L14_U1 ( .a ({new_AGEMA_signal_8796, new_AGEMA_signal_8795, SubBytesIns_Inst_Sbox_9_M52}), .b ({new_AGEMA_signal_8804, new_AGEMA_signal_8803, SubBytesIns_Inst_Sbox_9_M61}), .c ({new_AGEMA_signal_9230, new_AGEMA_signal_9229, SubBytesIns_Inst_Sbox_9_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L15_U1 ( .a ({new_AGEMA_signal_8800, new_AGEMA_signal_8799, SubBytesIns_Inst_Sbox_9_M55}), .b ({new_AGEMA_signal_8808, new_AGEMA_signal_8807, SubBytesIns_Inst_Sbox_9_L1}), .c ({new_AGEMA_signal_9232, new_AGEMA_signal_9231, SubBytesIns_Inst_Sbox_9_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L16_U1 ( .a ({new_AGEMA_signal_8326, new_AGEMA_signal_8325, SubBytesIns_Inst_Sbox_9_M56}), .b ({new_AGEMA_signal_9592, new_AGEMA_signal_9591, SubBytesIns_Inst_Sbox_9_L0}), .c ({new_AGEMA_signal_10006, new_AGEMA_signal_10005, SubBytesIns_Inst_Sbox_9_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L17_U1 ( .a ({new_AGEMA_signal_8328, new_AGEMA_signal_8327, SubBytesIns_Inst_Sbox_9_M57}), .b ({new_AGEMA_signal_8808, new_AGEMA_signal_8807, SubBytesIns_Inst_Sbox_9_L1}), .c ({new_AGEMA_signal_9234, new_AGEMA_signal_9233, SubBytesIns_Inst_Sbox_9_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L18_U1 ( .a ({new_AGEMA_signal_8802, new_AGEMA_signal_8801, SubBytesIns_Inst_Sbox_9_M58}), .b ({new_AGEMA_signal_8810, new_AGEMA_signal_8809, SubBytesIns_Inst_Sbox_9_L8}), .c ({new_AGEMA_signal_9236, new_AGEMA_signal_9235, SubBytesIns_Inst_Sbox_9_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L19_U1 ( .a ({new_AGEMA_signal_8806, new_AGEMA_signal_8805, SubBytesIns_Inst_Sbox_9_M63}), .b ({new_AGEMA_signal_9226, new_AGEMA_signal_9225, SubBytesIns_Inst_Sbox_9_L4}), .c ({new_AGEMA_signal_9604, new_AGEMA_signal_9603, SubBytesIns_Inst_Sbox_9_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L20_U1 ( .a ({new_AGEMA_signal_9592, new_AGEMA_signal_9591, SubBytesIns_Inst_Sbox_9_L0}), .b ({new_AGEMA_signal_8808, new_AGEMA_signal_8807, SubBytesIns_Inst_Sbox_9_L1}), .c ({new_AGEMA_signal_10008, new_AGEMA_signal_10007, SubBytesIns_Inst_Sbox_9_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L21_U1 ( .a ({new_AGEMA_signal_8808, new_AGEMA_signal_8807, SubBytesIns_Inst_Sbox_9_L1}), .b ({new_AGEMA_signal_9596, new_AGEMA_signal_9595, SubBytesIns_Inst_Sbox_9_L7}), .c ({new_AGEMA_signal_10010, new_AGEMA_signal_10009, SubBytesIns_Inst_Sbox_9_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L22_U1 ( .a ({new_AGEMA_signal_9224, new_AGEMA_signal_9223, SubBytesIns_Inst_Sbox_9_L3}), .b ({new_AGEMA_signal_8812, new_AGEMA_signal_8811, SubBytesIns_Inst_Sbox_9_L12}), .c ({new_AGEMA_signal_9606, new_AGEMA_signal_9605, SubBytesIns_Inst_Sbox_9_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L23_U1 ( .a ({new_AGEMA_signal_9236, new_AGEMA_signal_9235, SubBytesIns_Inst_Sbox_9_L18}), .b ({new_AGEMA_signal_9222, new_AGEMA_signal_9221, SubBytesIns_Inst_Sbox_9_L2}), .c ({new_AGEMA_signal_9608, new_AGEMA_signal_9607, SubBytesIns_Inst_Sbox_9_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L24_U1 ( .a ({new_AGEMA_signal_9232, new_AGEMA_signal_9231, SubBytesIns_Inst_Sbox_9_L15}), .b ({new_AGEMA_signal_9598, new_AGEMA_signal_9597, SubBytesIns_Inst_Sbox_9_L9}), .c ({new_AGEMA_signal_10012, new_AGEMA_signal_10011, SubBytesIns_Inst_Sbox_9_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L25_U1 ( .a ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_9600, new_AGEMA_signal_9599, SubBytesIns_Inst_Sbox_9_L10}), .c ({new_AGEMA_signal_10014, new_AGEMA_signal_10013, SubBytesIns_Inst_Sbox_9_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L26_U1 ( .a ({new_AGEMA_signal_9596, new_AGEMA_signal_9595, SubBytesIns_Inst_Sbox_9_L7}), .b ({new_AGEMA_signal_9598, new_AGEMA_signal_9597, SubBytesIns_Inst_Sbox_9_L9}), .c ({new_AGEMA_signal_10016, new_AGEMA_signal_10015, SubBytesIns_Inst_Sbox_9_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L27_U1 ( .a ({new_AGEMA_signal_8810, new_AGEMA_signal_8809, SubBytesIns_Inst_Sbox_9_L8}), .b ({new_AGEMA_signal_9600, new_AGEMA_signal_9599, SubBytesIns_Inst_Sbox_9_L10}), .c ({new_AGEMA_signal_10018, new_AGEMA_signal_10017, SubBytesIns_Inst_Sbox_9_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L28_U1 ( .a ({new_AGEMA_signal_9602, new_AGEMA_signal_9601, SubBytesIns_Inst_Sbox_9_L11}), .b ({new_AGEMA_signal_9230, new_AGEMA_signal_9229, SubBytesIns_Inst_Sbox_9_L14}), .c ({new_AGEMA_signal_10020, new_AGEMA_signal_10019, SubBytesIns_Inst_Sbox_9_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L29_U1 ( .a ({new_AGEMA_signal_9602, new_AGEMA_signal_9601, SubBytesIns_Inst_Sbox_9_L11}), .b ({new_AGEMA_signal_9234, new_AGEMA_signal_9233, SubBytesIns_Inst_Sbox_9_L17}), .c ({new_AGEMA_signal_10022, new_AGEMA_signal_10021, SubBytesIns_Inst_Sbox_9_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S0_U1 ( .a ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_10012, new_AGEMA_signal_10011, SubBytesIns_Inst_Sbox_9_L24}), .c ({new_AGEMA_signal_10348, new_AGEMA_signal_10347, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S1_U1 ( .a ({new_AGEMA_signal_10006, new_AGEMA_signal_10005, SubBytesIns_Inst_Sbox_9_L16}), .b ({new_AGEMA_signal_10016, new_AGEMA_signal_10015, SubBytesIns_Inst_Sbox_9_L26}), .c ({new_AGEMA_signal_10350, new_AGEMA_signal_10349, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S2_U1 ( .a ({new_AGEMA_signal_9604, new_AGEMA_signal_9603, SubBytesIns_Inst_Sbox_9_L19}), .b ({new_AGEMA_signal_10020, new_AGEMA_signal_10019, SubBytesIns_Inst_Sbox_9_L28}), .c ({new_AGEMA_signal_10352, new_AGEMA_signal_10351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S3_U1 ( .a ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_10010, new_AGEMA_signal_10009, SubBytesIns_Inst_Sbox_9_L21}), .c ({new_AGEMA_signal_10354, new_AGEMA_signal_10353, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S4_U1 ( .a ({new_AGEMA_signal_10008, new_AGEMA_signal_10007, SubBytesIns_Inst_Sbox_9_L20}), .b ({new_AGEMA_signal_9606, new_AGEMA_signal_9605, SubBytesIns_Inst_Sbox_9_L22}), .c ({new_AGEMA_signal_10356, new_AGEMA_signal_10355, MixColumnsInput[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S5_U1 ( .a ({new_AGEMA_signal_10014, new_AGEMA_signal_10013, SubBytesIns_Inst_Sbox_9_L25}), .b ({new_AGEMA_signal_10022, new_AGEMA_signal_10021, SubBytesIns_Inst_Sbox_9_L29}), .c ({new_AGEMA_signal_10358, new_AGEMA_signal_10357, MixColumnsInput[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S6_U1 ( .a ({new_AGEMA_signal_10004, new_AGEMA_signal_10003, SubBytesIns_Inst_Sbox_9_L13}), .b ({new_AGEMA_signal_10018, new_AGEMA_signal_10017, SubBytesIns_Inst_Sbox_9_L27}), .c ({new_AGEMA_signal_10360, new_AGEMA_signal_10359, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S7_U1 ( .a ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_9608, new_AGEMA_signal_9607, SubBytesIns_Inst_Sbox_9_L23}), .c ({new_AGEMA_signal_10024, new_AGEMA_signal_10023, MixColumnsInput[8]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M46_U1 ( .a ({new_AGEMA_signal_8340, new_AGEMA_signal_8339, SubBytesIns_Inst_Sbox_10_M44}), .b ({new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_10_T6}), .clk (clk), .r ({Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({new_AGEMA_signal_8816, new_AGEMA_signal_8815, SubBytesIns_Inst_Sbox_10_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M47_U1 ( .a ({new_AGEMA_signal_7956, new_AGEMA_signal_7955, SubBytesIns_Inst_Sbox_10_M40}), .b ({new_AGEMA_signal_6402, new_AGEMA_signal_6401, SubBytesIns_Inst_Sbox_10_T8}), .clk (clk), .r ({Fresh[1505], Fresh[1504], Fresh[1503]}), .c ({new_AGEMA_signal_8342, new_AGEMA_signal_8341, SubBytesIns_Inst_Sbox_10_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M48_U1 ( .a ({new_AGEMA_signal_7954, new_AGEMA_signal_7953, SubBytesIns_Inst_Sbox_10_M39}), .b ({ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .clk (clk), .r ({Fresh[1508], Fresh[1507], Fresh[1506]}), .c ({new_AGEMA_signal_8344, new_AGEMA_signal_8343, SubBytesIns_Inst_Sbox_10_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M49_U1 ( .a ({new_AGEMA_signal_8338, new_AGEMA_signal_8337, SubBytesIns_Inst_Sbox_10_M43}), .b ({new_AGEMA_signal_5950, new_AGEMA_signal_5949, SubBytesIns_Inst_Sbox_10_T16}), .clk (clk), .r ({Fresh[1511], Fresh[1510], Fresh[1509]}), .c ({new_AGEMA_signal_8818, new_AGEMA_signal_8817, SubBytesIns_Inst_Sbox_10_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M50_U1 ( .a ({new_AGEMA_signal_7952, new_AGEMA_signal_7951, SubBytesIns_Inst_Sbox_10_M38}), .b ({new_AGEMA_signal_5944, new_AGEMA_signal_5943, SubBytesIns_Inst_Sbox_10_T9}), .clk (clk), .r ({Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({new_AGEMA_signal_8346, new_AGEMA_signal_8345, SubBytesIns_Inst_Sbox_10_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M51_U1 ( .a ({new_AGEMA_signal_7950, new_AGEMA_signal_7949, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_6408, new_AGEMA_signal_6407, SubBytesIns_Inst_Sbox_10_T17}), .clk (clk), .r ({Fresh[1517], Fresh[1516], Fresh[1515]}), .c ({new_AGEMA_signal_8348, new_AGEMA_signal_8347, SubBytesIns_Inst_Sbox_10_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M52_U1 ( .a ({new_AGEMA_signal_8336, new_AGEMA_signal_8335, SubBytesIns_Inst_Sbox_10_M42}), .b ({new_AGEMA_signal_5948, new_AGEMA_signal_5947, SubBytesIns_Inst_Sbox_10_T15}), .clk (clk), .r ({Fresh[1520], Fresh[1519], Fresh[1518]}), .c ({new_AGEMA_signal_8820, new_AGEMA_signal_8819, SubBytesIns_Inst_Sbox_10_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M53_U1 ( .a ({new_AGEMA_signal_8814, new_AGEMA_signal_8813, SubBytesIns_Inst_Sbox_10_M45}), .b ({new_AGEMA_signal_5956, new_AGEMA_signal_5955, SubBytesIns_Inst_Sbox_10_T27}), .clk (clk), .r ({Fresh[1523], Fresh[1522], Fresh[1521]}), .c ({new_AGEMA_signal_9238, new_AGEMA_signal_9237, SubBytesIns_Inst_Sbox_10_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M54_U1 ( .a ({new_AGEMA_signal_8334, new_AGEMA_signal_8333, SubBytesIns_Inst_Sbox_10_M41}), .b ({new_AGEMA_signal_6404, new_AGEMA_signal_6403, SubBytesIns_Inst_Sbox_10_T10}), .clk (clk), .r ({Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({new_AGEMA_signal_8822, new_AGEMA_signal_8821, SubBytesIns_Inst_Sbox_10_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M55_U1 ( .a ({new_AGEMA_signal_8340, new_AGEMA_signal_8339, SubBytesIns_Inst_Sbox_10_M44}), .b ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, SubBytesIns_Inst_Sbox_10_T13}), .clk (clk), .r ({Fresh[1529], Fresh[1528], Fresh[1527]}), .c ({new_AGEMA_signal_8824, new_AGEMA_signal_8823, SubBytesIns_Inst_Sbox_10_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M56_U1 ( .a ({new_AGEMA_signal_7956, new_AGEMA_signal_7955, SubBytesIns_Inst_Sbox_10_M40}), .b ({new_AGEMA_signal_6412, new_AGEMA_signal_6411, SubBytesIns_Inst_Sbox_10_T23}), .clk (clk), .r ({Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({new_AGEMA_signal_8350, new_AGEMA_signal_8349, SubBytesIns_Inst_Sbox_10_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M57_U1 ( .a ({new_AGEMA_signal_7954, new_AGEMA_signal_7953, SubBytesIns_Inst_Sbox_10_M39}), .b ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, SubBytesIns_Inst_Sbox_10_T19}), .clk (clk), .r ({Fresh[1535], Fresh[1534], Fresh[1533]}), .c ({new_AGEMA_signal_8352, new_AGEMA_signal_8351, SubBytesIns_Inst_Sbox_10_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M58_U1 ( .a ({new_AGEMA_signal_8338, new_AGEMA_signal_8337, SubBytesIns_Inst_Sbox_10_M43}), .b ({new_AGEMA_signal_5602, new_AGEMA_signal_5601, SubBytesIns_Inst_Sbox_10_T3}), .clk (clk), .r ({Fresh[1538], Fresh[1537], Fresh[1536]}), .c ({new_AGEMA_signal_8826, new_AGEMA_signal_8825, SubBytesIns_Inst_Sbox_10_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M59_U1 ( .a ({new_AGEMA_signal_7952, new_AGEMA_signal_7951, SubBytesIns_Inst_Sbox_10_M38}), .b ({new_AGEMA_signal_5954, new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_10_T22}), .clk (clk), .r ({Fresh[1541], Fresh[1540], Fresh[1539]}), .c ({new_AGEMA_signal_8354, new_AGEMA_signal_8353, SubBytesIns_Inst_Sbox_10_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M60_U1 ( .a ({new_AGEMA_signal_7950, new_AGEMA_signal_7949, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_6410, new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_10_T20}), .clk (clk), .r ({Fresh[1544], Fresh[1543], Fresh[1542]}), .c ({new_AGEMA_signal_8356, new_AGEMA_signal_8355, SubBytesIns_Inst_Sbox_10_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M61_U1 ( .a ({new_AGEMA_signal_8336, new_AGEMA_signal_8335, SubBytesIns_Inst_Sbox_10_M42}), .b ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, SubBytesIns_Inst_Sbox_10_T1}), .clk (clk), .r ({Fresh[1547], Fresh[1546], Fresh[1545]}), .c ({new_AGEMA_signal_8828, new_AGEMA_signal_8827, SubBytesIns_Inst_Sbox_10_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M62_U1 ( .a ({new_AGEMA_signal_8814, new_AGEMA_signal_8813, SubBytesIns_Inst_Sbox_10_M45}), .b ({new_AGEMA_signal_5604, new_AGEMA_signal_5603, SubBytesIns_Inst_Sbox_10_T4}), .clk (clk), .r ({Fresh[1550], Fresh[1549], Fresh[1548]}), .c ({new_AGEMA_signal_9240, new_AGEMA_signal_9239, SubBytesIns_Inst_Sbox_10_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M63_U1 ( .a ({new_AGEMA_signal_8334, new_AGEMA_signal_8333, SubBytesIns_Inst_Sbox_10_M41}), .b ({new_AGEMA_signal_5600, new_AGEMA_signal_5599, SubBytesIns_Inst_Sbox_10_T2}), .clk (clk), .r ({Fresh[1553], Fresh[1552], Fresh[1551]}), .c ({new_AGEMA_signal_8830, new_AGEMA_signal_8829, SubBytesIns_Inst_Sbox_10_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L0_U1 ( .a ({new_AGEMA_signal_8828, new_AGEMA_signal_8827, SubBytesIns_Inst_Sbox_10_M61}), .b ({new_AGEMA_signal_9240, new_AGEMA_signal_9239, SubBytesIns_Inst_Sbox_10_M62}), .c ({new_AGEMA_signal_9610, new_AGEMA_signal_9609, SubBytesIns_Inst_Sbox_10_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L1_U1 ( .a ({new_AGEMA_signal_8346, new_AGEMA_signal_8345, SubBytesIns_Inst_Sbox_10_M50}), .b ({new_AGEMA_signal_8350, new_AGEMA_signal_8349, SubBytesIns_Inst_Sbox_10_M56}), .c ({new_AGEMA_signal_8832, new_AGEMA_signal_8831, SubBytesIns_Inst_Sbox_10_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L2_U1 ( .a ({new_AGEMA_signal_8816, new_AGEMA_signal_8815, SubBytesIns_Inst_Sbox_10_M46}), .b ({new_AGEMA_signal_8344, new_AGEMA_signal_8343, SubBytesIns_Inst_Sbox_10_M48}), .c ({new_AGEMA_signal_9242, new_AGEMA_signal_9241, SubBytesIns_Inst_Sbox_10_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L3_U1 ( .a ({new_AGEMA_signal_8342, new_AGEMA_signal_8341, SubBytesIns_Inst_Sbox_10_M47}), .b ({new_AGEMA_signal_8824, new_AGEMA_signal_8823, SubBytesIns_Inst_Sbox_10_M55}), .c ({new_AGEMA_signal_9244, new_AGEMA_signal_9243, SubBytesIns_Inst_Sbox_10_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L4_U1 ( .a ({new_AGEMA_signal_8822, new_AGEMA_signal_8821, SubBytesIns_Inst_Sbox_10_M54}), .b ({new_AGEMA_signal_8826, new_AGEMA_signal_8825, SubBytesIns_Inst_Sbox_10_M58}), .c ({new_AGEMA_signal_9246, new_AGEMA_signal_9245, SubBytesIns_Inst_Sbox_10_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L5_U1 ( .a ({new_AGEMA_signal_8818, new_AGEMA_signal_8817, SubBytesIns_Inst_Sbox_10_M49}), .b ({new_AGEMA_signal_8828, new_AGEMA_signal_8827, SubBytesIns_Inst_Sbox_10_M61}), .c ({new_AGEMA_signal_9248, new_AGEMA_signal_9247, SubBytesIns_Inst_Sbox_10_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L6_U1 ( .a ({new_AGEMA_signal_9240, new_AGEMA_signal_9239, SubBytesIns_Inst_Sbox_10_M62}), .b ({new_AGEMA_signal_9248, new_AGEMA_signal_9247, SubBytesIns_Inst_Sbox_10_L5}), .c ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, SubBytesIns_Inst_Sbox_10_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L7_U1 ( .a ({new_AGEMA_signal_8816, new_AGEMA_signal_8815, SubBytesIns_Inst_Sbox_10_M46}), .b ({new_AGEMA_signal_9244, new_AGEMA_signal_9243, SubBytesIns_Inst_Sbox_10_L3}), .c ({new_AGEMA_signal_9614, new_AGEMA_signal_9613, SubBytesIns_Inst_Sbox_10_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L8_U1 ( .a ({new_AGEMA_signal_8348, new_AGEMA_signal_8347, SubBytesIns_Inst_Sbox_10_M51}), .b ({new_AGEMA_signal_8354, new_AGEMA_signal_8353, SubBytesIns_Inst_Sbox_10_M59}), .c ({new_AGEMA_signal_8834, new_AGEMA_signal_8833, SubBytesIns_Inst_Sbox_10_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L9_U1 ( .a ({new_AGEMA_signal_8820, new_AGEMA_signal_8819, SubBytesIns_Inst_Sbox_10_M52}), .b ({new_AGEMA_signal_9238, new_AGEMA_signal_9237, SubBytesIns_Inst_Sbox_10_M53}), .c ({new_AGEMA_signal_9616, new_AGEMA_signal_9615, SubBytesIns_Inst_Sbox_10_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L10_U1 ( .a ({new_AGEMA_signal_9238, new_AGEMA_signal_9237, SubBytesIns_Inst_Sbox_10_M53}), .b ({new_AGEMA_signal_9246, new_AGEMA_signal_9245, SubBytesIns_Inst_Sbox_10_L4}), .c ({new_AGEMA_signal_9618, new_AGEMA_signal_9617, SubBytesIns_Inst_Sbox_10_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L11_U1 ( .a ({new_AGEMA_signal_8356, new_AGEMA_signal_8355, SubBytesIns_Inst_Sbox_10_M60}), .b ({new_AGEMA_signal_9242, new_AGEMA_signal_9241, SubBytesIns_Inst_Sbox_10_L2}), .c ({new_AGEMA_signal_9620, new_AGEMA_signal_9619, SubBytesIns_Inst_Sbox_10_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L12_U1 ( .a ({new_AGEMA_signal_8344, new_AGEMA_signal_8343, SubBytesIns_Inst_Sbox_10_M48}), .b ({new_AGEMA_signal_8348, new_AGEMA_signal_8347, SubBytesIns_Inst_Sbox_10_M51}), .c ({new_AGEMA_signal_8836, new_AGEMA_signal_8835, SubBytesIns_Inst_Sbox_10_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L13_U1 ( .a ({new_AGEMA_signal_8346, new_AGEMA_signal_8345, SubBytesIns_Inst_Sbox_10_M50}), .b ({new_AGEMA_signal_9610, new_AGEMA_signal_9609, SubBytesIns_Inst_Sbox_10_L0}), .c ({new_AGEMA_signal_10026, new_AGEMA_signal_10025, SubBytesIns_Inst_Sbox_10_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L14_U1 ( .a ({new_AGEMA_signal_8820, new_AGEMA_signal_8819, SubBytesIns_Inst_Sbox_10_M52}), .b ({new_AGEMA_signal_8828, new_AGEMA_signal_8827, SubBytesIns_Inst_Sbox_10_M61}), .c ({new_AGEMA_signal_9250, new_AGEMA_signal_9249, SubBytesIns_Inst_Sbox_10_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L15_U1 ( .a ({new_AGEMA_signal_8824, new_AGEMA_signal_8823, SubBytesIns_Inst_Sbox_10_M55}), .b ({new_AGEMA_signal_8832, new_AGEMA_signal_8831, SubBytesIns_Inst_Sbox_10_L1}), .c ({new_AGEMA_signal_9252, new_AGEMA_signal_9251, SubBytesIns_Inst_Sbox_10_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L16_U1 ( .a ({new_AGEMA_signal_8350, new_AGEMA_signal_8349, SubBytesIns_Inst_Sbox_10_M56}), .b ({new_AGEMA_signal_9610, new_AGEMA_signal_9609, SubBytesIns_Inst_Sbox_10_L0}), .c ({new_AGEMA_signal_10028, new_AGEMA_signal_10027, SubBytesIns_Inst_Sbox_10_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L17_U1 ( .a ({new_AGEMA_signal_8352, new_AGEMA_signal_8351, SubBytesIns_Inst_Sbox_10_M57}), .b ({new_AGEMA_signal_8832, new_AGEMA_signal_8831, SubBytesIns_Inst_Sbox_10_L1}), .c ({new_AGEMA_signal_9254, new_AGEMA_signal_9253, SubBytesIns_Inst_Sbox_10_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L18_U1 ( .a ({new_AGEMA_signal_8826, new_AGEMA_signal_8825, SubBytesIns_Inst_Sbox_10_M58}), .b ({new_AGEMA_signal_8834, new_AGEMA_signal_8833, SubBytesIns_Inst_Sbox_10_L8}), .c ({new_AGEMA_signal_9256, new_AGEMA_signal_9255, SubBytesIns_Inst_Sbox_10_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L19_U1 ( .a ({new_AGEMA_signal_8830, new_AGEMA_signal_8829, SubBytesIns_Inst_Sbox_10_M63}), .b ({new_AGEMA_signal_9246, new_AGEMA_signal_9245, SubBytesIns_Inst_Sbox_10_L4}), .c ({new_AGEMA_signal_9622, new_AGEMA_signal_9621, SubBytesIns_Inst_Sbox_10_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L20_U1 ( .a ({new_AGEMA_signal_9610, new_AGEMA_signal_9609, SubBytesIns_Inst_Sbox_10_L0}), .b ({new_AGEMA_signal_8832, new_AGEMA_signal_8831, SubBytesIns_Inst_Sbox_10_L1}), .c ({new_AGEMA_signal_10030, new_AGEMA_signal_10029, SubBytesIns_Inst_Sbox_10_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L21_U1 ( .a ({new_AGEMA_signal_8832, new_AGEMA_signal_8831, SubBytesIns_Inst_Sbox_10_L1}), .b ({new_AGEMA_signal_9614, new_AGEMA_signal_9613, SubBytesIns_Inst_Sbox_10_L7}), .c ({new_AGEMA_signal_10032, new_AGEMA_signal_10031, SubBytesIns_Inst_Sbox_10_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L22_U1 ( .a ({new_AGEMA_signal_9244, new_AGEMA_signal_9243, SubBytesIns_Inst_Sbox_10_L3}), .b ({new_AGEMA_signal_8836, new_AGEMA_signal_8835, SubBytesIns_Inst_Sbox_10_L12}), .c ({new_AGEMA_signal_9624, new_AGEMA_signal_9623, SubBytesIns_Inst_Sbox_10_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L23_U1 ( .a ({new_AGEMA_signal_9256, new_AGEMA_signal_9255, SubBytesIns_Inst_Sbox_10_L18}), .b ({new_AGEMA_signal_9242, new_AGEMA_signal_9241, SubBytesIns_Inst_Sbox_10_L2}), .c ({new_AGEMA_signal_9626, new_AGEMA_signal_9625, SubBytesIns_Inst_Sbox_10_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L24_U1 ( .a ({new_AGEMA_signal_9252, new_AGEMA_signal_9251, SubBytesIns_Inst_Sbox_10_L15}), .b ({new_AGEMA_signal_9616, new_AGEMA_signal_9615, SubBytesIns_Inst_Sbox_10_L9}), .c ({new_AGEMA_signal_10034, new_AGEMA_signal_10033, SubBytesIns_Inst_Sbox_10_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L25_U1 ( .a ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_9618, new_AGEMA_signal_9617, SubBytesIns_Inst_Sbox_10_L10}), .c ({new_AGEMA_signal_10036, new_AGEMA_signal_10035, SubBytesIns_Inst_Sbox_10_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L26_U1 ( .a ({new_AGEMA_signal_9614, new_AGEMA_signal_9613, SubBytesIns_Inst_Sbox_10_L7}), .b ({new_AGEMA_signal_9616, new_AGEMA_signal_9615, SubBytesIns_Inst_Sbox_10_L9}), .c ({new_AGEMA_signal_10038, new_AGEMA_signal_10037, SubBytesIns_Inst_Sbox_10_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L27_U1 ( .a ({new_AGEMA_signal_8834, new_AGEMA_signal_8833, SubBytesIns_Inst_Sbox_10_L8}), .b ({new_AGEMA_signal_9618, new_AGEMA_signal_9617, SubBytesIns_Inst_Sbox_10_L10}), .c ({new_AGEMA_signal_10040, new_AGEMA_signal_10039, SubBytesIns_Inst_Sbox_10_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L28_U1 ( .a ({new_AGEMA_signal_9620, new_AGEMA_signal_9619, SubBytesIns_Inst_Sbox_10_L11}), .b ({new_AGEMA_signal_9250, new_AGEMA_signal_9249, SubBytesIns_Inst_Sbox_10_L14}), .c ({new_AGEMA_signal_10042, new_AGEMA_signal_10041, SubBytesIns_Inst_Sbox_10_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L29_U1 ( .a ({new_AGEMA_signal_9620, new_AGEMA_signal_9619, SubBytesIns_Inst_Sbox_10_L11}), .b ({new_AGEMA_signal_9254, new_AGEMA_signal_9253, SubBytesIns_Inst_Sbox_10_L17}), .c ({new_AGEMA_signal_10044, new_AGEMA_signal_10043, SubBytesIns_Inst_Sbox_10_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S0_U1 ( .a ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_10034, new_AGEMA_signal_10033, SubBytesIns_Inst_Sbox_10_L24}), .c ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S1_U1 ( .a ({new_AGEMA_signal_10028, new_AGEMA_signal_10027, SubBytesIns_Inst_Sbox_10_L16}), .b ({new_AGEMA_signal_10038, new_AGEMA_signal_10037, SubBytesIns_Inst_Sbox_10_L26}), .c ({new_AGEMA_signal_10364, new_AGEMA_signal_10363, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S2_U1 ( .a ({new_AGEMA_signal_9622, new_AGEMA_signal_9621, SubBytesIns_Inst_Sbox_10_L19}), .b ({new_AGEMA_signal_10042, new_AGEMA_signal_10041, SubBytesIns_Inst_Sbox_10_L28}), .c ({new_AGEMA_signal_10366, new_AGEMA_signal_10365, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S3_U1 ( .a ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_10032, new_AGEMA_signal_10031, SubBytesIns_Inst_Sbox_10_L21}), .c ({new_AGEMA_signal_10368, new_AGEMA_signal_10367, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S4_U1 ( .a ({new_AGEMA_signal_10030, new_AGEMA_signal_10029, SubBytesIns_Inst_Sbox_10_L20}), .b ({new_AGEMA_signal_9624, new_AGEMA_signal_9623, SubBytesIns_Inst_Sbox_10_L22}), .c ({new_AGEMA_signal_10370, new_AGEMA_signal_10369, MixColumnsInput[115]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S5_U1 ( .a ({new_AGEMA_signal_10036, new_AGEMA_signal_10035, SubBytesIns_Inst_Sbox_10_L25}), .b ({new_AGEMA_signal_10044, new_AGEMA_signal_10043, SubBytesIns_Inst_Sbox_10_L29}), .c ({new_AGEMA_signal_10372, new_AGEMA_signal_10371, MixColumnsInput[114]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S6_U1 ( .a ({new_AGEMA_signal_10026, new_AGEMA_signal_10025, SubBytesIns_Inst_Sbox_10_L13}), .b ({new_AGEMA_signal_10040, new_AGEMA_signal_10039, SubBytesIns_Inst_Sbox_10_L27}), .c ({new_AGEMA_signal_10374, new_AGEMA_signal_10373, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S7_U1 ( .a ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_9626, new_AGEMA_signal_9625, SubBytesIns_Inst_Sbox_10_L23}), .c ({new_AGEMA_signal_10046, new_AGEMA_signal_10045, MixColumnsInput[112]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M46_U1 ( .a ({new_AGEMA_signal_8364, new_AGEMA_signal_8363, SubBytesIns_Inst_Sbox_11_M44}), .b ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, SubBytesIns_Inst_Sbox_11_T6}), .clk (clk), .r ({Fresh[1556], Fresh[1555], Fresh[1554]}), .c ({new_AGEMA_signal_8840, new_AGEMA_signal_8839, SubBytesIns_Inst_Sbox_11_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M47_U1 ( .a ({new_AGEMA_signal_7964, new_AGEMA_signal_7963, SubBytesIns_Inst_Sbox_11_M40}), .b ({new_AGEMA_signal_6428, new_AGEMA_signal_6427, SubBytesIns_Inst_Sbox_11_T8}), .clk (clk), .r ({Fresh[1559], Fresh[1558], Fresh[1557]}), .c ({new_AGEMA_signal_8366, new_AGEMA_signal_8365, SubBytesIns_Inst_Sbox_11_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M48_U1 ( .a ({new_AGEMA_signal_7962, new_AGEMA_signal_7961, SubBytesIns_Inst_Sbox_11_M39}), .b ({ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .clk (clk), .r ({Fresh[1562], Fresh[1561], Fresh[1560]}), .c ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, SubBytesIns_Inst_Sbox_11_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M49_U1 ( .a ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, SubBytesIns_Inst_Sbox_11_M43}), .b ({new_AGEMA_signal_5966, new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_11_T16}), .clk (clk), .r ({Fresh[1565], Fresh[1564], Fresh[1563]}), .c ({new_AGEMA_signal_8842, new_AGEMA_signal_8841, SubBytesIns_Inst_Sbox_11_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M50_U1 ( .a ({new_AGEMA_signal_7960, new_AGEMA_signal_7959, SubBytesIns_Inst_Sbox_11_M38}), .b ({new_AGEMA_signal_5960, new_AGEMA_signal_5959, SubBytesIns_Inst_Sbox_11_T9}), .clk (clk), .r ({Fresh[1568], Fresh[1567], Fresh[1566]}), .c ({new_AGEMA_signal_8370, new_AGEMA_signal_8369, SubBytesIns_Inst_Sbox_11_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M51_U1 ( .a ({new_AGEMA_signal_7958, new_AGEMA_signal_7957, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_6434, new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_11_T17}), .clk (clk), .r ({Fresh[1571], Fresh[1570], Fresh[1569]}), .c ({new_AGEMA_signal_8372, new_AGEMA_signal_8371, SubBytesIns_Inst_Sbox_11_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M52_U1 ( .a ({new_AGEMA_signal_8360, new_AGEMA_signal_8359, SubBytesIns_Inst_Sbox_11_M42}), .b ({new_AGEMA_signal_5964, new_AGEMA_signal_5963, SubBytesIns_Inst_Sbox_11_T15}), .clk (clk), .r ({Fresh[1574], Fresh[1573], Fresh[1572]}), .c ({new_AGEMA_signal_8844, new_AGEMA_signal_8843, SubBytesIns_Inst_Sbox_11_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M53_U1 ( .a ({new_AGEMA_signal_8838, new_AGEMA_signal_8837, SubBytesIns_Inst_Sbox_11_M45}), .b ({new_AGEMA_signal_5972, new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_11_T27}), .clk (clk), .r ({Fresh[1577], Fresh[1576], Fresh[1575]}), .c ({new_AGEMA_signal_9258, new_AGEMA_signal_9257, SubBytesIns_Inst_Sbox_11_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M54_U1 ( .a ({new_AGEMA_signal_8358, new_AGEMA_signal_8357, SubBytesIns_Inst_Sbox_11_M41}), .b ({new_AGEMA_signal_6430, new_AGEMA_signal_6429, SubBytesIns_Inst_Sbox_11_T10}), .clk (clk), .r ({Fresh[1580], Fresh[1579], Fresh[1578]}), .c ({new_AGEMA_signal_8846, new_AGEMA_signal_8845, SubBytesIns_Inst_Sbox_11_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M55_U1 ( .a ({new_AGEMA_signal_8364, new_AGEMA_signal_8363, SubBytesIns_Inst_Sbox_11_M44}), .b ({new_AGEMA_signal_5962, new_AGEMA_signal_5961, SubBytesIns_Inst_Sbox_11_T13}), .clk (clk), .r ({Fresh[1583], Fresh[1582], Fresh[1581]}), .c ({new_AGEMA_signal_8848, new_AGEMA_signal_8847, SubBytesIns_Inst_Sbox_11_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M56_U1 ( .a ({new_AGEMA_signal_7964, new_AGEMA_signal_7963, SubBytesIns_Inst_Sbox_11_M40}), .b ({new_AGEMA_signal_6438, new_AGEMA_signal_6437, SubBytesIns_Inst_Sbox_11_T23}), .clk (clk), .r ({Fresh[1586], Fresh[1585], Fresh[1584]}), .c ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, SubBytesIns_Inst_Sbox_11_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M57_U1 ( .a ({new_AGEMA_signal_7962, new_AGEMA_signal_7961, SubBytesIns_Inst_Sbox_11_M39}), .b ({new_AGEMA_signal_5968, new_AGEMA_signal_5967, SubBytesIns_Inst_Sbox_11_T19}), .clk (clk), .r ({Fresh[1589], Fresh[1588], Fresh[1587]}), .c ({new_AGEMA_signal_8376, new_AGEMA_signal_8375, SubBytesIns_Inst_Sbox_11_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M58_U1 ( .a ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, SubBytesIns_Inst_Sbox_11_M43}), .b ({new_AGEMA_signal_5622, new_AGEMA_signal_5621, SubBytesIns_Inst_Sbox_11_T3}), .clk (clk), .r ({Fresh[1592], Fresh[1591], Fresh[1590]}), .c ({new_AGEMA_signal_8850, new_AGEMA_signal_8849, SubBytesIns_Inst_Sbox_11_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M59_U1 ( .a ({new_AGEMA_signal_7960, new_AGEMA_signal_7959, SubBytesIns_Inst_Sbox_11_M38}), .b ({new_AGEMA_signal_5970, new_AGEMA_signal_5969, SubBytesIns_Inst_Sbox_11_T22}), .clk (clk), .r ({Fresh[1595], Fresh[1594], Fresh[1593]}), .c ({new_AGEMA_signal_8378, new_AGEMA_signal_8377, SubBytesIns_Inst_Sbox_11_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M60_U1 ( .a ({new_AGEMA_signal_7958, new_AGEMA_signal_7957, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_6436, new_AGEMA_signal_6435, SubBytesIns_Inst_Sbox_11_T20}), .clk (clk), .r ({Fresh[1598], Fresh[1597], Fresh[1596]}), .c ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, SubBytesIns_Inst_Sbox_11_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M61_U1 ( .a ({new_AGEMA_signal_8360, new_AGEMA_signal_8359, SubBytesIns_Inst_Sbox_11_M42}), .b ({new_AGEMA_signal_5618, new_AGEMA_signal_5617, SubBytesIns_Inst_Sbox_11_T1}), .clk (clk), .r ({Fresh[1601], Fresh[1600], Fresh[1599]}), .c ({new_AGEMA_signal_8852, new_AGEMA_signal_8851, SubBytesIns_Inst_Sbox_11_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M62_U1 ( .a ({new_AGEMA_signal_8838, new_AGEMA_signal_8837, SubBytesIns_Inst_Sbox_11_M45}), .b ({new_AGEMA_signal_5624, new_AGEMA_signal_5623, SubBytesIns_Inst_Sbox_11_T4}), .clk (clk), .r ({Fresh[1604], Fresh[1603], Fresh[1602]}), .c ({new_AGEMA_signal_9260, new_AGEMA_signal_9259, SubBytesIns_Inst_Sbox_11_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M63_U1 ( .a ({new_AGEMA_signal_8358, new_AGEMA_signal_8357, SubBytesIns_Inst_Sbox_11_M41}), .b ({new_AGEMA_signal_5620, new_AGEMA_signal_5619, SubBytesIns_Inst_Sbox_11_T2}), .clk (clk), .r ({Fresh[1607], Fresh[1606], Fresh[1605]}), .c ({new_AGEMA_signal_8854, new_AGEMA_signal_8853, SubBytesIns_Inst_Sbox_11_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L0_U1 ( .a ({new_AGEMA_signal_8852, new_AGEMA_signal_8851, SubBytesIns_Inst_Sbox_11_M61}), .b ({new_AGEMA_signal_9260, new_AGEMA_signal_9259, SubBytesIns_Inst_Sbox_11_M62}), .c ({new_AGEMA_signal_9628, new_AGEMA_signal_9627, SubBytesIns_Inst_Sbox_11_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L1_U1 ( .a ({new_AGEMA_signal_8370, new_AGEMA_signal_8369, SubBytesIns_Inst_Sbox_11_M50}), .b ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, SubBytesIns_Inst_Sbox_11_M56}), .c ({new_AGEMA_signal_8856, new_AGEMA_signal_8855, SubBytesIns_Inst_Sbox_11_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L2_U1 ( .a ({new_AGEMA_signal_8840, new_AGEMA_signal_8839, SubBytesIns_Inst_Sbox_11_M46}), .b ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, SubBytesIns_Inst_Sbox_11_M48}), .c ({new_AGEMA_signal_9262, new_AGEMA_signal_9261, SubBytesIns_Inst_Sbox_11_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L3_U1 ( .a ({new_AGEMA_signal_8366, new_AGEMA_signal_8365, SubBytesIns_Inst_Sbox_11_M47}), .b ({new_AGEMA_signal_8848, new_AGEMA_signal_8847, SubBytesIns_Inst_Sbox_11_M55}), .c ({new_AGEMA_signal_9264, new_AGEMA_signal_9263, SubBytesIns_Inst_Sbox_11_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L4_U1 ( .a ({new_AGEMA_signal_8846, new_AGEMA_signal_8845, SubBytesIns_Inst_Sbox_11_M54}), .b ({new_AGEMA_signal_8850, new_AGEMA_signal_8849, SubBytesIns_Inst_Sbox_11_M58}), .c ({new_AGEMA_signal_9266, new_AGEMA_signal_9265, SubBytesIns_Inst_Sbox_11_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L5_U1 ( .a ({new_AGEMA_signal_8842, new_AGEMA_signal_8841, SubBytesIns_Inst_Sbox_11_M49}), .b ({new_AGEMA_signal_8852, new_AGEMA_signal_8851, SubBytesIns_Inst_Sbox_11_M61}), .c ({new_AGEMA_signal_9268, new_AGEMA_signal_9267, SubBytesIns_Inst_Sbox_11_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L6_U1 ( .a ({new_AGEMA_signal_9260, new_AGEMA_signal_9259, SubBytesIns_Inst_Sbox_11_M62}), .b ({new_AGEMA_signal_9268, new_AGEMA_signal_9267, SubBytesIns_Inst_Sbox_11_L5}), .c ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, SubBytesIns_Inst_Sbox_11_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L7_U1 ( .a ({new_AGEMA_signal_8840, new_AGEMA_signal_8839, SubBytesIns_Inst_Sbox_11_M46}), .b ({new_AGEMA_signal_9264, new_AGEMA_signal_9263, SubBytesIns_Inst_Sbox_11_L3}), .c ({new_AGEMA_signal_9632, new_AGEMA_signal_9631, SubBytesIns_Inst_Sbox_11_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L8_U1 ( .a ({new_AGEMA_signal_8372, new_AGEMA_signal_8371, SubBytesIns_Inst_Sbox_11_M51}), .b ({new_AGEMA_signal_8378, new_AGEMA_signal_8377, SubBytesIns_Inst_Sbox_11_M59}), .c ({new_AGEMA_signal_8858, new_AGEMA_signal_8857, SubBytesIns_Inst_Sbox_11_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L9_U1 ( .a ({new_AGEMA_signal_8844, new_AGEMA_signal_8843, SubBytesIns_Inst_Sbox_11_M52}), .b ({new_AGEMA_signal_9258, new_AGEMA_signal_9257, SubBytesIns_Inst_Sbox_11_M53}), .c ({new_AGEMA_signal_9634, new_AGEMA_signal_9633, SubBytesIns_Inst_Sbox_11_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L10_U1 ( .a ({new_AGEMA_signal_9258, new_AGEMA_signal_9257, SubBytesIns_Inst_Sbox_11_M53}), .b ({new_AGEMA_signal_9266, new_AGEMA_signal_9265, SubBytesIns_Inst_Sbox_11_L4}), .c ({new_AGEMA_signal_9636, new_AGEMA_signal_9635, SubBytesIns_Inst_Sbox_11_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L11_U1 ( .a ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, SubBytesIns_Inst_Sbox_11_M60}), .b ({new_AGEMA_signal_9262, new_AGEMA_signal_9261, SubBytesIns_Inst_Sbox_11_L2}), .c ({new_AGEMA_signal_9638, new_AGEMA_signal_9637, SubBytesIns_Inst_Sbox_11_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L12_U1 ( .a ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, SubBytesIns_Inst_Sbox_11_M48}), .b ({new_AGEMA_signal_8372, new_AGEMA_signal_8371, SubBytesIns_Inst_Sbox_11_M51}), .c ({new_AGEMA_signal_8860, new_AGEMA_signal_8859, SubBytesIns_Inst_Sbox_11_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L13_U1 ( .a ({new_AGEMA_signal_8370, new_AGEMA_signal_8369, SubBytesIns_Inst_Sbox_11_M50}), .b ({new_AGEMA_signal_9628, new_AGEMA_signal_9627, SubBytesIns_Inst_Sbox_11_L0}), .c ({new_AGEMA_signal_10048, new_AGEMA_signal_10047, SubBytesIns_Inst_Sbox_11_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L14_U1 ( .a ({new_AGEMA_signal_8844, new_AGEMA_signal_8843, SubBytesIns_Inst_Sbox_11_M52}), .b ({new_AGEMA_signal_8852, new_AGEMA_signal_8851, SubBytesIns_Inst_Sbox_11_M61}), .c ({new_AGEMA_signal_9270, new_AGEMA_signal_9269, SubBytesIns_Inst_Sbox_11_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L15_U1 ( .a ({new_AGEMA_signal_8848, new_AGEMA_signal_8847, SubBytesIns_Inst_Sbox_11_M55}), .b ({new_AGEMA_signal_8856, new_AGEMA_signal_8855, SubBytesIns_Inst_Sbox_11_L1}), .c ({new_AGEMA_signal_9272, new_AGEMA_signal_9271, SubBytesIns_Inst_Sbox_11_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L16_U1 ( .a ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, SubBytesIns_Inst_Sbox_11_M56}), .b ({new_AGEMA_signal_9628, new_AGEMA_signal_9627, SubBytesIns_Inst_Sbox_11_L0}), .c ({new_AGEMA_signal_10050, new_AGEMA_signal_10049, SubBytesIns_Inst_Sbox_11_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L17_U1 ( .a ({new_AGEMA_signal_8376, new_AGEMA_signal_8375, SubBytesIns_Inst_Sbox_11_M57}), .b ({new_AGEMA_signal_8856, new_AGEMA_signal_8855, SubBytesIns_Inst_Sbox_11_L1}), .c ({new_AGEMA_signal_9274, new_AGEMA_signal_9273, SubBytesIns_Inst_Sbox_11_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L18_U1 ( .a ({new_AGEMA_signal_8850, new_AGEMA_signal_8849, SubBytesIns_Inst_Sbox_11_M58}), .b ({new_AGEMA_signal_8858, new_AGEMA_signal_8857, SubBytesIns_Inst_Sbox_11_L8}), .c ({new_AGEMA_signal_9276, new_AGEMA_signal_9275, SubBytesIns_Inst_Sbox_11_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L19_U1 ( .a ({new_AGEMA_signal_8854, new_AGEMA_signal_8853, SubBytesIns_Inst_Sbox_11_M63}), .b ({new_AGEMA_signal_9266, new_AGEMA_signal_9265, SubBytesIns_Inst_Sbox_11_L4}), .c ({new_AGEMA_signal_9640, new_AGEMA_signal_9639, SubBytesIns_Inst_Sbox_11_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L20_U1 ( .a ({new_AGEMA_signal_9628, new_AGEMA_signal_9627, SubBytesIns_Inst_Sbox_11_L0}), .b ({new_AGEMA_signal_8856, new_AGEMA_signal_8855, SubBytesIns_Inst_Sbox_11_L1}), .c ({new_AGEMA_signal_10052, new_AGEMA_signal_10051, SubBytesIns_Inst_Sbox_11_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L21_U1 ( .a ({new_AGEMA_signal_8856, new_AGEMA_signal_8855, SubBytesIns_Inst_Sbox_11_L1}), .b ({new_AGEMA_signal_9632, new_AGEMA_signal_9631, SubBytesIns_Inst_Sbox_11_L7}), .c ({new_AGEMA_signal_10054, new_AGEMA_signal_10053, SubBytesIns_Inst_Sbox_11_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L22_U1 ( .a ({new_AGEMA_signal_9264, new_AGEMA_signal_9263, SubBytesIns_Inst_Sbox_11_L3}), .b ({new_AGEMA_signal_8860, new_AGEMA_signal_8859, SubBytesIns_Inst_Sbox_11_L12}), .c ({new_AGEMA_signal_9642, new_AGEMA_signal_9641, SubBytesIns_Inst_Sbox_11_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L23_U1 ( .a ({new_AGEMA_signal_9276, new_AGEMA_signal_9275, SubBytesIns_Inst_Sbox_11_L18}), .b ({new_AGEMA_signal_9262, new_AGEMA_signal_9261, SubBytesIns_Inst_Sbox_11_L2}), .c ({new_AGEMA_signal_9644, new_AGEMA_signal_9643, SubBytesIns_Inst_Sbox_11_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L24_U1 ( .a ({new_AGEMA_signal_9272, new_AGEMA_signal_9271, SubBytesIns_Inst_Sbox_11_L15}), .b ({new_AGEMA_signal_9634, new_AGEMA_signal_9633, SubBytesIns_Inst_Sbox_11_L9}), .c ({new_AGEMA_signal_10056, new_AGEMA_signal_10055, SubBytesIns_Inst_Sbox_11_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L25_U1 ( .a ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_9636, new_AGEMA_signal_9635, SubBytesIns_Inst_Sbox_11_L10}), .c ({new_AGEMA_signal_10058, new_AGEMA_signal_10057, SubBytesIns_Inst_Sbox_11_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L26_U1 ( .a ({new_AGEMA_signal_9632, new_AGEMA_signal_9631, SubBytesIns_Inst_Sbox_11_L7}), .b ({new_AGEMA_signal_9634, new_AGEMA_signal_9633, SubBytesIns_Inst_Sbox_11_L9}), .c ({new_AGEMA_signal_10060, new_AGEMA_signal_10059, SubBytesIns_Inst_Sbox_11_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L27_U1 ( .a ({new_AGEMA_signal_8858, new_AGEMA_signal_8857, SubBytesIns_Inst_Sbox_11_L8}), .b ({new_AGEMA_signal_9636, new_AGEMA_signal_9635, SubBytesIns_Inst_Sbox_11_L10}), .c ({new_AGEMA_signal_10062, new_AGEMA_signal_10061, SubBytesIns_Inst_Sbox_11_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L28_U1 ( .a ({new_AGEMA_signal_9638, new_AGEMA_signal_9637, SubBytesIns_Inst_Sbox_11_L11}), .b ({new_AGEMA_signal_9270, new_AGEMA_signal_9269, SubBytesIns_Inst_Sbox_11_L14}), .c ({new_AGEMA_signal_10064, new_AGEMA_signal_10063, SubBytesIns_Inst_Sbox_11_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L29_U1 ( .a ({new_AGEMA_signal_9638, new_AGEMA_signal_9637, SubBytesIns_Inst_Sbox_11_L11}), .b ({new_AGEMA_signal_9274, new_AGEMA_signal_9273, SubBytesIns_Inst_Sbox_11_L17}), .c ({new_AGEMA_signal_10066, new_AGEMA_signal_10065, SubBytesIns_Inst_Sbox_11_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S0_U1 ( .a ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_10056, new_AGEMA_signal_10055, SubBytesIns_Inst_Sbox_11_L24}), .c ({new_AGEMA_signal_10376, new_AGEMA_signal_10375, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S1_U1 ( .a ({new_AGEMA_signal_10050, new_AGEMA_signal_10049, SubBytesIns_Inst_Sbox_11_L16}), .b ({new_AGEMA_signal_10060, new_AGEMA_signal_10059, SubBytesIns_Inst_Sbox_11_L26}), .c ({new_AGEMA_signal_10378, new_AGEMA_signal_10377, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S2_U1 ( .a ({new_AGEMA_signal_9640, new_AGEMA_signal_9639, SubBytesIns_Inst_Sbox_11_L19}), .b ({new_AGEMA_signal_10064, new_AGEMA_signal_10063, SubBytesIns_Inst_Sbox_11_L28}), .c ({new_AGEMA_signal_10380, new_AGEMA_signal_10379, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S3_U1 ( .a ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_10054, new_AGEMA_signal_10053, SubBytesIns_Inst_Sbox_11_L21}), .c ({new_AGEMA_signal_10382, new_AGEMA_signal_10381, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S4_U1 ( .a ({new_AGEMA_signal_10052, new_AGEMA_signal_10051, SubBytesIns_Inst_Sbox_11_L20}), .b ({new_AGEMA_signal_9642, new_AGEMA_signal_9641, SubBytesIns_Inst_Sbox_11_L22}), .c ({new_AGEMA_signal_10384, new_AGEMA_signal_10383, MixColumnsInput[91]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S5_U1 ( .a ({new_AGEMA_signal_10058, new_AGEMA_signal_10057, SubBytesIns_Inst_Sbox_11_L25}), .b ({new_AGEMA_signal_10066, new_AGEMA_signal_10065, SubBytesIns_Inst_Sbox_11_L29}), .c ({new_AGEMA_signal_10386, new_AGEMA_signal_10385, MixColumnsInput[90]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S6_U1 ( .a ({new_AGEMA_signal_10048, new_AGEMA_signal_10047, SubBytesIns_Inst_Sbox_11_L13}), .b ({new_AGEMA_signal_10062, new_AGEMA_signal_10061, SubBytesIns_Inst_Sbox_11_L27}), .c ({new_AGEMA_signal_10388, new_AGEMA_signal_10387, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S7_U1 ( .a ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_9644, new_AGEMA_signal_9643, SubBytesIns_Inst_Sbox_11_L23}), .c ({new_AGEMA_signal_10068, new_AGEMA_signal_10067, MixColumnsInput[88]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M46_U1 ( .a ({new_AGEMA_signal_8388, new_AGEMA_signal_8387, SubBytesIns_Inst_Sbox_12_M44}), .b ({new_AGEMA_signal_5974, new_AGEMA_signal_5973, SubBytesIns_Inst_Sbox_12_T6}), .clk (clk), .r ({Fresh[1610], Fresh[1609], Fresh[1608]}), .c ({new_AGEMA_signal_8864, new_AGEMA_signal_8863, SubBytesIns_Inst_Sbox_12_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M47_U1 ( .a ({new_AGEMA_signal_7972, new_AGEMA_signal_7971, SubBytesIns_Inst_Sbox_12_M40}), .b ({new_AGEMA_signal_6454, new_AGEMA_signal_6453, SubBytesIns_Inst_Sbox_12_T8}), .clk (clk), .r ({Fresh[1613], Fresh[1612], Fresh[1611]}), .c ({new_AGEMA_signal_8390, new_AGEMA_signal_8389, SubBytesIns_Inst_Sbox_12_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M48_U1 ( .a ({new_AGEMA_signal_7970, new_AGEMA_signal_7969, SubBytesIns_Inst_Sbox_12_M39}), .b ({ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .clk (clk), .r ({Fresh[1616], Fresh[1615], Fresh[1614]}), .c ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, SubBytesIns_Inst_Sbox_12_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M49_U1 ( .a ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, SubBytesIns_Inst_Sbox_12_M43}), .b ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, SubBytesIns_Inst_Sbox_12_T16}), .clk (clk), .r ({Fresh[1619], Fresh[1618], Fresh[1617]}), .c ({new_AGEMA_signal_8866, new_AGEMA_signal_8865, SubBytesIns_Inst_Sbox_12_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M50_U1 ( .a ({new_AGEMA_signal_7968, new_AGEMA_signal_7967, SubBytesIns_Inst_Sbox_12_M38}), .b ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, SubBytesIns_Inst_Sbox_12_T9}), .clk (clk), .r ({Fresh[1622], Fresh[1621], Fresh[1620]}), .c ({new_AGEMA_signal_8394, new_AGEMA_signal_8393, SubBytesIns_Inst_Sbox_12_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M51_U1 ( .a ({new_AGEMA_signal_7966, new_AGEMA_signal_7965, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_6460, new_AGEMA_signal_6459, SubBytesIns_Inst_Sbox_12_T17}), .clk (clk), .r ({Fresh[1625], Fresh[1624], Fresh[1623]}), .c ({new_AGEMA_signal_8396, new_AGEMA_signal_8395, SubBytesIns_Inst_Sbox_12_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M52_U1 ( .a ({new_AGEMA_signal_8384, new_AGEMA_signal_8383, SubBytesIns_Inst_Sbox_12_M42}), .b ({new_AGEMA_signal_5980, new_AGEMA_signal_5979, SubBytesIns_Inst_Sbox_12_T15}), .clk (clk), .r ({Fresh[1628], Fresh[1627], Fresh[1626]}), .c ({new_AGEMA_signal_8868, new_AGEMA_signal_8867, SubBytesIns_Inst_Sbox_12_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M53_U1 ( .a ({new_AGEMA_signal_8862, new_AGEMA_signal_8861, SubBytesIns_Inst_Sbox_12_M45}), .b ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, SubBytesIns_Inst_Sbox_12_T27}), .clk (clk), .r ({Fresh[1631], Fresh[1630], Fresh[1629]}), .c ({new_AGEMA_signal_9278, new_AGEMA_signal_9277, SubBytesIns_Inst_Sbox_12_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M54_U1 ( .a ({new_AGEMA_signal_8382, new_AGEMA_signal_8381, SubBytesIns_Inst_Sbox_12_M41}), .b ({new_AGEMA_signal_6456, new_AGEMA_signal_6455, SubBytesIns_Inst_Sbox_12_T10}), .clk (clk), .r ({Fresh[1634], Fresh[1633], Fresh[1632]}), .c ({new_AGEMA_signal_8870, new_AGEMA_signal_8869, SubBytesIns_Inst_Sbox_12_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M55_U1 ( .a ({new_AGEMA_signal_8388, new_AGEMA_signal_8387, SubBytesIns_Inst_Sbox_12_M44}), .b ({new_AGEMA_signal_5978, new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_12_T13}), .clk (clk), .r ({Fresh[1637], Fresh[1636], Fresh[1635]}), .c ({new_AGEMA_signal_8872, new_AGEMA_signal_8871, SubBytesIns_Inst_Sbox_12_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M56_U1 ( .a ({new_AGEMA_signal_7972, new_AGEMA_signal_7971, SubBytesIns_Inst_Sbox_12_M40}), .b ({new_AGEMA_signal_6464, new_AGEMA_signal_6463, SubBytesIns_Inst_Sbox_12_T23}), .clk (clk), .r ({Fresh[1640], Fresh[1639], Fresh[1638]}), .c ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, SubBytesIns_Inst_Sbox_12_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M57_U1 ( .a ({new_AGEMA_signal_7970, new_AGEMA_signal_7969, SubBytesIns_Inst_Sbox_12_M39}), .b ({new_AGEMA_signal_5984, new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_12_T19}), .clk (clk), .r ({Fresh[1643], Fresh[1642], Fresh[1641]}), .c ({new_AGEMA_signal_8400, new_AGEMA_signal_8399, SubBytesIns_Inst_Sbox_12_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M58_U1 ( .a ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, SubBytesIns_Inst_Sbox_12_M43}), .b ({new_AGEMA_signal_5642, new_AGEMA_signal_5641, SubBytesIns_Inst_Sbox_12_T3}), .clk (clk), .r ({Fresh[1646], Fresh[1645], Fresh[1644]}), .c ({new_AGEMA_signal_8874, new_AGEMA_signal_8873, SubBytesIns_Inst_Sbox_12_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M59_U1 ( .a ({new_AGEMA_signal_7968, new_AGEMA_signal_7967, SubBytesIns_Inst_Sbox_12_M38}), .b ({new_AGEMA_signal_5986, new_AGEMA_signal_5985, SubBytesIns_Inst_Sbox_12_T22}), .clk (clk), .r ({Fresh[1649], Fresh[1648], Fresh[1647]}), .c ({new_AGEMA_signal_8402, new_AGEMA_signal_8401, SubBytesIns_Inst_Sbox_12_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M60_U1 ( .a ({new_AGEMA_signal_7966, new_AGEMA_signal_7965, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_6462, new_AGEMA_signal_6461, SubBytesIns_Inst_Sbox_12_T20}), .clk (clk), .r ({Fresh[1652], Fresh[1651], Fresh[1650]}), .c ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, SubBytesIns_Inst_Sbox_12_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M61_U1 ( .a ({new_AGEMA_signal_8384, new_AGEMA_signal_8383, SubBytesIns_Inst_Sbox_12_M42}), .b ({new_AGEMA_signal_5638, new_AGEMA_signal_5637, SubBytesIns_Inst_Sbox_12_T1}), .clk (clk), .r ({Fresh[1655], Fresh[1654], Fresh[1653]}), .c ({new_AGEMA_signal_8876, new_AGEMA_signal_8875, SubBytesIns_Inst_Sbox_12_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M62_U1 ( .a ({new_AGEMA_signal_8862, new_AGEMA_signal_8861, SubBytesIns_Inst_Sbox_12_M45}), .b ({new_AGEMA_signal_5644, new_AGEMA_signal_5643, SubBytesIns_Inst_Sbox_12_T4}), .clk (clk), .r ({Fresh[1658], Fresh[1657], Fresh[1656]}), .c ({new_AGEMA_signal_9280, new_AGEMA_signal_9279, SubBytesIns_Inst_Sbox_12_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M63_U1 ( .a ({new_AGEMA_signal_8382, new_AGEMA_signal_8381, SubBytesIns_Inst_Sbox_12_M41}), .b ({new_AGEMA_signal_5640, new_AGEMA_signal_5639, SubBytesIns_Inst_Sbox_12_T2}), .clk (clk), .r ({Fresh[1661], Fresh[1660], Fresh[1659]}), .c ({new_AGEMA_signal_8878, new_AGEMA_signal_8877, SubBytesIns_Inst_Sbox_12_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L0_U1 ( .a ({new_AGEMA_signal_8876, new_AGEMA_signal_8875, SubBytesIns_Inst_Sbox_12_M61}), .b ({new_AGEMA_signal_9280, new_AGEMA_signal_9279, SubBytesIns_Inst_Sbox_12_M62}), .c ({new_AGEMA_signal_9646, new_AGEMA_signal_9645, SubBytesIns_Inst_Sbox_12_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L1_U1 ( .a ({new_AGEMA_signal_8394, new_AGEMA_signal_8393, SubBytesIns_Inst_Sbox_12_M50}), .b ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, SubBytesIns_Inst_Sbox_12_M56}), .c ({new_AGEMA_signal_8880, new_AGEMA_signal_8879, SubBytesIns_Inst_Sbox_12_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L2_U1 ( .a ({new_AGEMA_signal_8864, new_AGEMA_signal_8863, SubBytesIns_Inst_Sbox_12_M46}), .b ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, SubBytesIns_Inst_Sbox_12_M48}), .c ({new_AGEMA_signal_9282, new_AGEMA_signal_9281, SubBytesIns_Inst_Sbox_12_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L3_U1 ( .a ({new_AGEMA_signal_8390, new_AGEMA_signal_8389, SubBytesIns_Inst_Sbox_12_M47}), .b ({new_AGEMA_signal_8872, new_AGEMA_signal_8871, SubBytesIns_Inst_Sbox_12_M55}), .c ({new_AGEMA_signal_9284, new_AGEMA_signal_9283, SubBytesIns_Inst_Sbox_12_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L4_U1 ( .a ({new_AGEMA_signal_8870, new_AGEMA_signal_8869, SubBytesIns_Inst_Sbox_12_M54}), .b ({new_AGEMA_signal_8874, new_AGEMA_signal_8873, SubBytesIns_Inst_Sbox_12_M58}), .c ({new_AGEMA_signal_9286, new_AGEMA_signal_9285, SubBytesIns_Inst_Sbox_12_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L5_U1 ( .a ({new_AGEMA_signal_8866, new_AGEMA_signal_8865, SubBytesIns_Inst_Sbox_12_M49}), .b ({new_AGEMA_signal_8876, new_AGEMA_signal_8875, SubBytesIns_Inst_Sbox_12_M61}), .c ({new_AGEMA_signal_9288, new_AGEMA_signal_9287, SubBytesIns_Inst_Sbox_12_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L6_U1 ( .a ({new_AGEMA_signal_9280, new_AGEMA_signal_9279, SubBytesIns_Inst_Sbox_12_M62}), .b ({new_AGEMA_signal_9288, new_AGEMA_signal_9287, SubBytesIns_Inst_Sbox_12_L5}), .c ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, SubBytesIns_Inst_Sbox_12_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L7_U1 ( .a ({new_AGEMA_signal_8864, new_AGEMA_signal_8863, SubBytesIns_Inst_Sbox_12_M46}), .b ({new_AGEMA_signal_9284, new_AGEMA_signal_9283, SubBytesIns_Inst_Sbox_12_L3}), .c ({new_AGEMA_signal_9650, new_AGEMA_signal_9649, SubBytesIns_Inst_Sbox_12_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L8_U1 ( .a ({new_AGEMA_signal_8396, new_AGEMA_signal_8395, SubBytesIns_Inst_Sbox_12_M51}), .b ({new_AGEMA_signal_8402, new_AGEMA_signal_8401, SubBytesIns_Inst_Sbox_12_M59}), .c ({new_AGEMA_signal_8882, new_AGEMA_signal_8881, SubBytesIns_Inst_Sbox_12_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L9_U1 ( .a ({new_AGEMA_signal_8868, new_AGEMA_signal_8867, SubBytesIns_Inst_Sbox_12_M52}), .b ({new_AGEMA_signal_9278, new_AGEMA_signal_9277, SubBytesIns_Inst_Sbox_12_M53}), .c ({new_AGEMA_signal_9652, new_AGEMA_signal_9651, SubBytesIns_Inst_Sbox_12_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L10_U1 ( .a ({new_AGEMA_signal_9278, new_AGEMA_signal_9277, SubBytesIns_Inst_Sbox_12_M53}), .b ({new_AGEMA_signal_9286, new_AGEMA_signal_9285, SubBytesIns_Inst_Sbox_12_L4}), .c ({new_AGEMA_signal_9654, new_AGEMA_signal_9653, SubBytesIns_Inst_Sbox_12_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L11_U1 ( .a ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, SubBytesIns_Inst_Sbox_12_M60}), .b ({new_AGEMA_signal_9282, new_AGEMA_signal_9281, SubBytesIns_Inst_Sbox_12_L2}), .c ({new_AGEMA_signal_9656, new_AGEMA_signal_9655, SubBytesIns_Inst_Sbox_12_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L12_U1 ( .a ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, SubBytesIns_Inst_Sbox_12_M48}), .b ({new_AGEMA_signal_8396, new_AGEMA_signal_8395, SubBytesIns_Inst_Sbox_12_M51}), .c ({new_AGEMA_signal_8884, new_AGEMA_signal_8883, SubBytesIns_Inst_Sbox_12_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L13_U1 ( .a ({new_AGEMA_signal_8394, new_AGEMA_signal_8393, SubBytesIns_Inst_Sbox_12_M50}), .b ({new_AGEMA_signal_9646, new_AGEMA_signal_9645, SubBytesIns_Inst_Sbox_12_L0}), .c ({new_AGEMA_signal_10070, new_AGEMA_signal_10069, SubBytesIns_Inst_Sbox_12_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L14_U1 ( .a ({new_AGEMA_signal_8868, new_AGEMA_signal_8867, SubBytesIns_Inst_Sbox_12_M52}), .b ({new_AGEMA_signal_8876, new_AGEMA_signal_8875, SubBytesIns_Inst_Sbox_12_M61}), .c ({new_AGEMA_signal_9290, new_AGEMA_signal_9289, SubBytesIns_Inst_Sbox_12_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L15_U1 ( .a ({new_AGEMA_signal_8872, new_AGEMA_signal_8871, SubBytesIns_Inst_Sbox_12_M55}), .b ({new_AGEMA_signal_8880, new_AGEMA_signal_8879, SubBytesIns_Inst_Sbox_12_L1}), .c ({new_AGEMA_signal_9292, new_AGEMA_signal_9291, SubBytesIns_Inst_Sbox_12_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L16_U1 ( .a ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, SubBytesIns_Inst_Sbox_12_M56}), .b ({new_AGEMA_signal_9646, new_AGEMA_signal_9645, SubBytesIns_Inst_Sbox_12_L0}), .c ({new_AGEMA_signal_10072, new_AGEMA_signal_10071, SubBytesIns_Inst_Sbox_12_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L17_U1 ( .a ({new_AGEMA_signal_8400, new_AGEMA_signal_8399, SubBytesIns_Inst_Sbox_12_M57}), .b ({new_AGEMA_signal_8880, new_AGEMA_signal_8879, SubBytesIns_Inst_Sbox_12_L1}), .c ({new_AGEMA_signal_9294, new_AGEMA_signal_9293, SubBytesIns_Inst_Sbox_12_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L18_U1 ( .a ({new_AGEMA_signal_8874, new_AGEMA_signal_8873, SubBytesIns_Inst_Sbox_12_M58}), .b ({new_AGEMA_signal_8882, new_AGEMA_signal_8881, SubBytesIns_Inst_Sbox_12_L8}), .c ({new_AGEMA_signal_9296, new_AGEMA_signal_9295, SubBytesIns_Inst_Sbox_12_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L19_U1 ( .a ({new_AGEMA_signal_8878, new_AGEMA_signal_8877, SubBytesIns_Inst_Sbox_12_M63}), .b ({new_AGEMA_signal_9286, new_AGEMA_signal_9285, SubBytesIns_Inst_Sbox_12_L4}), .c ({new_AGEMA_signal_9658, new_AGEMA_signal_9657, SubBytesIns_Inst_Sbox_12_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L20_U1 ( .a ({new_AGEMA_signal_9646, new_AGEMA_signal_9645, SubBytesIns_Inst_Sbox_12_L0}), .b ({new_AGEMA_signal_8880, new_AGEMA_signal_8879, SubBytesIns_Inst_Sbox_12_L1}), .c ({new_AGEMA_signal_10074, new_AGEMA_signal_10073, SubBytesIns_Inst_Sbox_12_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L21_U1 ( .a ({new_AGEMA_signal_8880, new_AGEMA_signal_8879, SubBytesIns_Inst_Sbox_12_L1}), .b ({new_AGEMA_signal_9650, new_AGEMA_signal_9649, SubBytesIns_Inst_Sbox_12_L7}), .c ({new_AGEMA_signal_10076, new_AGEMA_signal_10075, SubBytesIns_Inst_Sbox_12_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L22_U1 ( .a ({new_AGEMA_signal_9284, new_AGEMA_signal_9283, SubBytesIns_Inst_Sbox_12_L3}), .b ({new_AGEMA_signal_8884, new_AGEMA_signal_8883, SubBytesIns_Inst_Sbox_12_L12}), .c ({new_AGEMA_signal_9660, new_AGEMA_signal_9659, SubBytesIns_Inst_Sbox_12_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L23_U1 ( .a ({new_AGEMA_signal_9296, new_AGEMA_signal_9295, SubBytesIns_Inst_Sbox_12_L18}), .b ({new_AGEMA_signal_9282, new_AGEMA_signal_9281, SubBytesIns_Inst_Sbox_12_L2}), .c ({new_AGEMA_signal_9662, new_AGEMA_signal_9661, SubBytesIns_Inst_Sbox_12_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L24_U1 ( .a ({new_AGEMA_signal_9292, new_AGEMA_signal_9291, SubBytesIns_Inst_Sbox_12_L15}), .b ({new_AGEMA_signal_9652, new_AGEMA_signal_9651, SubBytesIns_Inst_Sbox_12_L9}), .c ({new_AGEMA_signal_10078, new_AGEMA_signal_10077, SubBytesIns_Inst_Sbox_12_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L25_U1 ( .a ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_9654, new_AGEMA_signal_9653, SubBytesIns_Inst_Sbox_12_L10}), .c ({new_AGEMA_signal_10080, new_AGEMA_signal_10079, SubBytesIns_Inst_Sbox_12_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L26_U1 ( .a ({new_AGEMA_signal_9650, new_AGEMA_signal_9649, SubBytesIns_Inst_Sbox_12_L7}), .b ({new_AGEMA_signal_9652, new_AGEMA_signal_9651, SubBytesIns_Inst_Sbox_12_L9}), .c ({new_AGEMA_signal_10082, new_AGEMA_signal_10081, SubBytesIns_Inst_Sbox_12_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L27_U1 ( .a ({new_AGEMA_signal_8882, new_AGEMA_signal_8881, SubBytesIns_Inst_Sbox_12_L8}), .b ({new_AGEMA_signal_9654, new_AGEMA_signal_9653, SubBytesIns_Inst_Sbox_12_L10}), .c ({new_AGEMA_signal_10084, new_AGEMA_signal_10083, SubBytesIns_Inst_Sbox_12_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L28_U1 ( .a ({new_AGEMA_signal_9656, new_AGEMA_signal_9655, SubBytesIns_Inst_Sbox_12_L11}), .b ({new_AGEMA_signal_9290, new_AGEMA_signal_9289, SubBytesIns_Inst_Sbox_12_L14}), .c ({new_AGEMA_signal_10086, new_AGEMA_signal_10085, SubBytesIns_Inst_Sbox_12_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L29_U1 ( .a ({new_AGEMA_signal_9656, new_AGEMA_signal_9655, SubBytesIns_Inst_Sbox_12_L11}), .b ({new_AGEMA_signal_9294, new_AGEMA_signal_9293, SubBytesIns_Inst_Sbox_12_L17}), .c ({new_AGEMA_signal_10088, new_AGEMA_signal_10087, SubBytesIns_Inst_Sbox_12_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S0_U1 ( .a ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_10078, new_AGEMA_signal_10077, SubBytesIns_Inst_Sbox_12_L24}), .c ({new_AGEMA_signal_10390, new_AGEMA_signal_10389, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S1_U1 ( .a ({new_AGEMA_signal_10072, new_AGEMA_signal_10071, SubBytesIns_Inst_Sbox_12_L16}), .b ({new_AGEMA_signal_10082, new_AGEMA_signal_10081, SubBytesIns_Inst_Sbox_12_L26}), .c ({new_AGEMA_signal_10392, new_AGEMA_signal_10391, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S2_U1 ( .a ({new_AGEMA_signal_9658, new_AGEMA_signal_9657, SubBytesIns_Inst_Sbox_12_L19}), .b ({new_AGEMA_signal_10086, new_AGEMA_signal_10085, SubBytesIns_Inst_Sbox_12_L28}), .c ({new_AGEMA_signal_10394, new_AGEMA_signal_10393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S3_U1 ( .a ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_10076, new_AGEMA_signal_10075, SubBytesIns_Inst_Sbox_12_L21}), .c ({new_AGEMA_signal_10396, new_AGEMA_signal_10395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S4_U1 ( .a ({new_AGEMA_signal_10074, new_AGEMA_signal_10073, SubBytesIns_Inst_Sbox_12_L20}), .b ({new_AGEMA_signal_9660, new_AGEMA_signal_9659, SubBytesIns_Inst_Sbox_12_L22}), .c ({new_AGEMA_signal_10398, new_AGEMA_signal_10397, MixColumnsInput[67]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S5_U1 ( .a ({new_AGEMA_signal_10080, new_AGEMA_signal_10079, SubBytesIns_Inst_Sbox_12_L25}), .b ({new_AGEMA_signal_10088, new_AGEMA_signal_10087, SubBytesIns_Inst_Sbox_12_L29}), .c ({new_AGEMA_signal_10400, new_AGEMA_signal_10399, MixColumnsInput[66]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S6_U1 ( .a ({new_AGEMA_signal_10070, new_AGEMA_signal_10069, SubBytesIns_Inst_Sbox_12_L13}), .b ({new_AGEMA_signal_10084, new_AGEMA_signal_10083, SubBytesIns_Inst_Sbox_12_L27}), .c ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S7_U1 ( .a ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_9662, new_AGEMA_signal_9661, SubBytesIns_Inst_Sbox_12_L23}), .c ({new_AGEMA_signal_10090, new_AGEMA_signal_10089, MixColumnsInput[64]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M46_U1 ( .a ({new_AGEMA_signal_8412, new_AGEMA_signal_8411, SubBytesIns_Inst_Sbox_13_M44}), .b ({new_AGEMA_signal_5990, new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_13_T6}), .clk (clk), .r ({Fresh[1664], Fresh[1663], Fresh[1662]}), .c ({new_AGEMA_signal_8888, new_AGEMA_signal_8887, SubBytesIns_Inst_Sbox_13_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M47_U1 ( .a ({new_AGEMA_signal_7980, new_AGEMA_signal_7979, SubBytesIns_Inst_Sbox_13_M40}), .b ({new_AGEMA_signal_6480, new_AGEMA_signal_6479, SubBytesIns_Inst_Sbox_13_T8}), .clk (clk), .r ({Fresh[1667], Fresh[1666], Fresh[1665]}), .c ({new_AGEMA_signal_8414, new_AGEMA_signal_8413, SubBytesIns_Inst_Sbox_13_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M48_U1 ( .a ({new_AGEMA_signal_7978, new_AGEMA_signal_7977, SubBytesIns_Inst_Sbox_13_M39}), .b ({ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .clk (clk), .r ({Fresh[1670], Fresh[1669], Fresh[1668]}), .c ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, SubBytesIns_Inst_Sbox_13_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M49_U1 ( .a ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, SubBytesIns_Inst_Sbox_13_M43}), .b ({new_AGEMA_signal_5998, new_AGEMA_signal_5997, SubBytesIns_Inst_Sbox_13_T16}), .clk (clk), .r ({Fresh[1673], Fresh[1672], Fresh[1671]}), .c ({new_AGEMA_signal_8890, new_AGEMA_signal_8889, SubBytesIns_Inst_Sbox_13_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M50_U1 ( .a ({new_AGEMA_signal_7976, new_AGEMA_signal_7975, SubBytesIns_Inst_Sbox_13_M38}), .b ({new_AGEMA_signal_5992, new_AGEMA_signal_5991, SubBytesIns_Inst_Sbox_13_T9}), .clk (clk), .r ({Fresh[1676], Fresh[1675], Fresh[1674]}), .c ({new_AGEMA_signal_8418, new_AGEMA_signal_8417, SubBytesIns_Inst_Sbox_13_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M51_U1 ( .a ({new_AGEMA_signal_7974, new_AGEMA_signal_7973, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_6486, new_AGEMA_signal_6485, SubBytesIns_Inst_Sbox_13_T17}), .clk (clk), .r ({Fresh[1679], Fresh[1678], Fresh[1677]}), .c ({new_AGEMA_signal_8420, new_AGEMA_signal_8419, SubBytesIns_Inst_Sbox_13_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M52_U1 ( .a ({new_AGEMA_signal_8408, new_AGEMA_signal_8407, SubBytesIns_Inst_Sbox_13_M42}), .b ({new_AGEMA_signal_5996, new_AGEMA_signal_5995, SubBytesIns_Inst_Sbox_13_T15}), .clk (clk), .r ({Fresh[1682], Fresh[1681], Fresh[1680]}), .c ({new_AGEMA_signal_8892, new_AGEMA_signal_8891, SubBytesIns_Inst_Sbox_13_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M53_U1 ( .a ({new_AGEMA_signal_8886, new_AGEMA_signal_8885, SubBytesIns_Inst_Sbox_13_M45}), .b ({new_AGEMA_signal_6004, new_AGEMA_signal_6003, SubBytesIns_Inst_Sbox_13_T27}), .clk (clk), .r ({Fresh[1685], Fresh[1684], Fresh[1683]}), .c ({new_AGEMA_signal_9298, new_AGEMA_signal_9297, SubBytesIns_Inst_Sbox_13_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M54_U1 ( .a ({new_AGEMA_signal_8406, new_AGEMA_signal_8405, SubBytesIns_Inst_Sbox_13_M41}), .b ({new_AGEMA_signal_6482, new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_13_T10}), .clk (clk), .r ({Fresh[1688], Fresh[1687], Fresh[1686]}), .c ({new_AGEMA_signal_8894, new_AGEMA_signal_8893, SubBytesIns_Inst_Sbox_13_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M55_U1 ( .a ({new_AGEMA_signal_8412, new_AGEMA_signal_8411, SubBytesIns_Inst_Sbox_13_M44}), .b ({new_AGEMA_signal_5994, new_AGEMA_signal_5993, SubBytesIns_Inst_Sbox_13_T13}), .clk (clk), .r ({Fresh[1691], Fresh[1690], Fresh[1689]}), .c ({new_AGEMA_signal_8896, new_AGEMA_signal_8895, SubBytesIns_Inst_Sbox_13_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M56_U1 ( .a ({new_AGEMA_signal_7980, new_AGEMA_signal_7979, SubBytesIns_Inst_Sbox_13_M40}), .b ({new_AGEMA_signal_6490, new_AGEMA_signal_6489, SubBytesIns_Inst_Sbox_13_T23}), .clk (clk), .r ({Fresh[1694], Fresh[1693], Fresh[1692]}), .c ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, SubBytesIns_Inst_Sbox_13_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M57_U1 ( .a ({new_AGEMA_signal_7978, new_AGEMA_signal_7977, SubBytesIns_Inst_Sbox_13_M39}), .b ({new_AGEMA_signal_6000, new_AGEMA_signal_5999, SubBytesIns_Inst_Sbox_13_T19}), .clk (clk), .r ({Fresh[1697], Fresh[1696], Fresh[1695]}), .c ({new_AGEMA_signal_8424, new_AGEMA_signal_8423, SubBytesIns_Inst_Sbox_13_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M58_U1 ( .a ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, SubBytesIns_Inst_Sbox_13_M43}), .b ({new_AGEMA_signal_5662, new_AGEMA_signal_5661, SubBytesIns_Inst_Sbox_13_T3}), .clk (clk), .r ({Fresh[1700], Fresh[1699], Fresh[1698]}), .c ({new_AGEMA_signal_8898, new_AGEMA_signal_8897, SubBytesIns_Inst_Sbox_13_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M59_U1 ( .a ({new_AGEMA_signal_7976, new_AGEMA_signal_7975, SubBytesIns_Inst_Sbox_13_M38}), .b ({new_AGEMA_signal_6002, new_AGEMA_signal_6001, SubBytesIns_Inst_Sbox_13_T22}), .clk (clk), .r ({Fresh[1703], Fresh[1702], Fresh[1701]}), .c ({new_AGEMA_signal_8426, new_AGEMA_signal_8425, SubBytesIns_Inst_Sbox_13_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M60_U1 ( .a ({new_AGEMA_signal_7974, new_AGEMA_signal_7973, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_6488, new_AGEMA_signal_6487, SubBytesIns_Inst_Sbox_13_T20}), .clk (clk), .r ({Fresh[1706], Fresh[1705], Fresh[1704]}), .c ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, SubBytesIns_Inst_Sbox_13_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M61_U1 ( .a ({new_AGEMA_signal_8408, new_AGEMA_signal_8407, SubBytesIns_Inst_Sbox_13_M42}), .b ({new_AGEMA_signal_5658, new_AGEMA_signal_5657, SubBytesIns_Inst_Sbox_13_T1}), .clk (clk), .r ({Fresh[1709], Fresh[1708], Fresh[1707]}), .c ({new_AGEMA_signal_8900, new_AGEMA_signal_8899, SubBytesIns_Inst_Sbox_13_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M62_U1 ( .a ({new_AGEMA_signal_8886, new_AGEMA_signal_8885, SubBytesIns_Inst_Sbox_13_M45}), .b ({new_AGEMA_signal_5664, new_AGEMA_signal_5663, SubBytesIns_Inst_Sbox_13_T4}), .clk (clk), .r ({Fresh[1712], Fresh[1711], Fresh[1710]}), .c ({new_AGEMA_signal_9300, new_AGEMA_signal_9299, SubBytesIns_Inst_Sbox_13_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M63_U1 ( .a ({new_AGEMA_signal_8406, new_AGEMA_signal_8405, SubBytesIns_Inst_Sbox_13_M41}), .b ({new_AGEMA_signal_5660, new_AGEMA_signal_5659, SubBytesIns_Inst_Sbox_13_T2}), .clk (clk), .r ({Fresh[1715], Fresh[1714], Fresh[1713]}), .c ({new_AGEMA_signal_8902, new_AGEMA_signal_8901, SubBytesIns_Inst_Sbox_13_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L0_U1 ( .a ({new_AGEMA_signal_8900, new_AGEMA_signal_8899, SubBytesIns_Inst_Sbox_13_M61}), .b ({new_AGEMA_signal_9300, new_AGEMA_signal_9299, SubBytesIns_Inst_Sbox_13_M62}), .c ({new_AGEMA_signal_9664, new_AGEMA_signal_9663, SubBytesIns_Inst_Sbox_13_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L1_U1 ( .a ({new_AGEMA_signal_8418, new_AGEMA_signal_8417, SubBytesIns_Inst_Sbox_13_M50}), .b ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, SubBytesIns_Inst_Sbox_13_M56}), .c ({new_AGEMA_signal_8904, new_AGEMA_signal_8903, SubBytesIns_Inst_Sbox_13_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L2_U1 ( .a ({new_AGEMA_signal_8888, new_AGEMA_signal_8887, SubBytesIns_Inst_Sbox_13_M46}), .b ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, SubBytesIns_Inst_Sbox_13_M48}), .c ({new_AGEMA_signal_9302, new_AGEMA_signal_9301, SubBytesIns_Inst_Sbox_13_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L3_U1 ( .a ({new_AGEMA_signal_8414, new_AGEMA_signal_8413, SubBytesIns_Inst_Sbox_13_M47}), .b ({new_AGEMA_signal_8896, new_AGEMA_signal_8895, SubBytesIns_Inst_Sbox_13_M55}), .c ({new_AGEMA_signal_9304, new_AGEMA_signal_9303, SubBytesIns_Inst_Sbox_13_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L4_U1 ( .a ({new_AGEMA_signal_8894, new_AGEMA_signal_8893, SubBytesIns_Inst_Sbox_13_M54}), .b ({new_AGEMA_signal_8898, new_AGEMA_signal_8897, SubBytesIns_Inst_Sbox_13_M58}), .c ({new_AGEMA_signal_9306, new_AGEMA_signal_9305, SubBytesIns_Inst_Sbox_13_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L5_U1 ( .a ({new_AGEMA_signal_8890, new_AGEMA_signal_8889, SubBytesIns_Inst_Sbox_13_M49}), .b ({new_AGEMA_signal_8900, new_AGEMA_signal_8899, SubBytesIns_Inst_Sbox_13_M61}), .c ({new_AGEMA_signal_9308, new_AGEMA_signal_9307, SubBytesIns_Inst_Sbox_13_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L6_U1 ( .a ({new_AGEMA_signal_9300, new_AGEMA_signal_9299, SubBytesIns_Inst_Sbox_13_M62}), .b ({new_AGEMA_signal_9308, new_AGEMA_signal_9307, SubBytesIns_Inst_Sbox_13_L5}), .c ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, SubBytesIns_Inst_Sbox_13_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L7_U1 ( .a ({new_AGEMA_signal_8888, new_AGEMA_signal_8887, SubBytesIns_Inst_Sbox_13_M46}), .b ({new_AGEMA_signal_9304, new_AGEMA_signal_9303, SubBytesIns_Inst_Sbox_13_L3}), .c ({new_AGEMA_signal_9668, new_AGEMA_signal_9667, SubBytesIns_Inst_Sbox_13_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L8_U1 ( .a ({new_AGEMA_signal_8420, new_AGEMA_signal_8419, SubBytesIns_Inst_Sbox_13_M51}), .b ({new_AGEMA_signal_8426, new_AGEMA_signal_8425, SubBytesIns_Inst_Sbox_13_M59}), .c ({new_AGEMA_signal_8906, new_AGEMA_signal_8905, SubBytesIns_Inst_Sbox_13_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L9_U1 ( .a ({new_AGEMA_signal_8892, new_AGEMA_signal_8891, SubBytesIns_Inst_Sbox_13_M52}), .b ({new_AGEMA_signal_9298, new_AGEMA_signal_9297, SubBytesIns_Inst_Sbox_13_M53}), .c ({new_AGEMA_signal_9670, new_AGEMA_signal_9669, SubBytesIns_Inst_Sbox_13_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L10_U1 ( .a ({new_AGEMA_signal_9298, new_AGEMA_signal_9297, SubBytesIns_Inst_Sbox_13_M53}), .b ({new_AGEMA_signal_9306, new_AGEMA_signal_9305, SubBytesIns_Inst_Sbox_13_L4}), .c ({new_AGEMA_signal_9672, new_AGEMA_signal_9671, SubBytesIns_Inst_Sbox_13_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L11_U1 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, SubBytesIns_Inst_Sbox_13_M60}), .b ({new_AGEMA_signal_9302, new_AGEMA_signal_9301, SubBytesIns_Inst_Sbox_13_L2}), .c ({new_AGEMA_signal_9674, new_AGEMA_signal_9673, SubBytesIns_Inst_Sbox_13_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L12_U1 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, SubBytesIns_Inst_Sbox_13_M48}), .b ({new_AGEMA_signal_8420, new_AGEMA_signal_8419, SubBytesIns_Inst_Sbox_13_M51}), .c ({new_AGEMA_signal_8908, new_AGEMA_signal_8907, SubBytesIns_Inst_Sbox_13_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L13_U1 ( .a ({new_AGEMA_signal_8418, new_AGEMA_signal_8417, SubBytesIns_Inst_Sbox_13_M50}), .b ({new_AGEMA_signal_9664, new_AGEMA_signal_9663, SubBytesIns_Inst_Sbox_13_L0}), .c ({new_AGEMA_signal_10092, new_AGEMA_signal_10091, SubBytesIns_Inst_Sbox_13_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L14_U1 ( .a ({new_AGEMA_signal_8892, new_AGEMA_signal_8891, SubBytesIns_Inst_Sbox_13_M52}), .b ({new_AGEMA_signal_8900, new_AGEMA_signal_8899, SubBytesIns_Inst_Sbox_13_M61}), .c ({new_AGEMA_signal_9310, new_AGEMA_signal_9309, SubBytesIns_Inst_Sbox_13_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L15_U1 ( .a ({new_AGEMA_signal_8896, new_AGEMA_signal_8895, SubBytesIns_Inst_Sbox_13_M55}), .b ({new_AGEMA_signal_8904, new_AGEMA_signal_8903, SubBytesIns_Inst_Sbox_13_L1}), .c ({new_AGEMA_signal_9312, new_AGEMA_signal_9311, SubBytesIns_Inst_Sbox_13_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L16_U1 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, SubBytesIns_Inst_Sbox_13_M56}), .b ({new_AGEMA_signal_9664, new_AGEMA_signal_9663, SubBytesIns_Inst_Sbox_13_L0}), .c ({new_AGEMA_signal_10094, new_AGEMA_signal_10093, SubBytesIns_Inst_Sbox_13_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L17_U1 ( .a ({new_AGEMA_signal_8424, new_AGEMA_signal_8423, SubBytesIns_Inst_Sbox_13_M57}), .b ({new_AGEMA_signal_8904, new_AGEMA_signal_8903, SubBytesIns_Inst_Sbox_13_L1}), .c ({new_AGEMA_signal_9314, new_AGEMA_signal_9313, SubBytesIns_Inst_Sbox_13_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L18_U1 ( .a ({new_AGEMA_signal_8898, new_AGEMA_signal_8897, SubBytesIns_Inst_Sbox_13_M58}), .b ({new_AGEMA_signal_8906, new_AGEMA_signal_8905, SubBytesIns_Inst_Sbox_13_L8}), .c ({new_AGEMA_signal_9316, new_AGEMA_signal_9315, SubBytesIns_Inst_Sbox_13_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L19_U1 ( .a ({new_AGEMA_signal_8902, new_AGEMA_signal_8901, SubBytesIns_Inst_Sbox_13_M63}), .b ({new_AGEMA_signal_9306, new_AGEMA_signal_9305, SubBytesIns_Inst_Sbox_13_L4}), .c ({new_AGEMA_signal_9676, new_AGEMA_signal_9675, SubBytesIns_Inst_Sbox_13_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L20_U1 ( .a ({new_AGEMA_signal_9664, new_AGEMA_signal_9663, SubBytesIns_Inst_Sbox_13_L0}), .b ({new_AGEMA_signal_8904, new_AGEMA_signal_8903, SubBytesIns_Inst_Sbox_13_L1}), .c ({new_AGEMA_signal_10096, new_AGEMA_signal_10095, SubBytesIns_Inst_Sbox_13_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L21_U1 ( .a ({new_AGEMA_signal_8904, new_AGEMA_signal_8903, SubBytesIns_Inst_Sbox_13_L1}), .b ({new_AGEMA_signal_9668, new_AGEMA_signal_9667, SubBytesIns_Inst_Sbox_13_L7}), .c ({new_AGEMA_signal_10098, new_AGEMA_signal_10097, SubBytesIns_Inst_Sbox_13_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L22_U1 ( .a ({new_AGEMA_signal_9304, new_AGEMA_signal_9303, SubBytesIns_Inst_Sbox_13_L3}), .b ({new_AGEMA_signal_8908, new_AGEMA_signal_8907, SubBytesIns_Inst_Sbox_13_L12}), .c ({new_AGEMA_signal_9678, new_AGEMA_signal_9677, SubBytesIns_Inst_Sbox_13_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L23_U1 ( .a ({new_AGEMA_signal_9316, new_AGEMA_signal_9315, SubBytesIns_Inst_Sbox_13_L18}), .b ({new_AGEMA_signal_9302, new_AGEMA_signal_9301, SubBytesIns_Inst_Sbox_13_L2}), .c ({new_AGEMA_signal_9680, new_AGEMA_signal_9679, SubBytesIns_Inst_Sbox_13_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L24_U1 ( .a ({new_AGEMA_signal_9312, new_AGEMA_signal_9311, SubBytesIns_Inst_Sbox_13_L15}), .b ({new_AGEMA_signal_9670, new_AGEMA_signal_9669, SubBytesIns_Inst_Sbox_13_L9}), .c ({new_AGEMA_signal_10100, new_AGEMA_signal_10099, SubBytesIns_Inst_Sbox_13_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L25_U1 ( .a ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_9672, new_AGEMA_signal_9671, SubBytesIns_Inst_Sbox_13_L10}), .c ({new_AGEMA_signal_10102, new_AGEMA_signal_10101, SubBytesIns_Inst_Sbox_13_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L26_U1 ( .a ({new_AGEMA_signal_9668, new_AGEMA_signal_9667, SubBytesIns_Inst_Sbox_13_L7}), .b ({new_AGEMA_signal_9670, new_AGEMA_signal_9669, SubBytesIns_Inst_Sbox_13_L9}), .c ({new_AGEMA_signal_10104, new_AGEMA_signal_10103, SubBytesIns_Inst_Sbox_13_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L27_U1 ( .a ({new_AGEMA_signal_8906, new_AGEMA_signal_8905, SubBytesIns_Inst_Sbox_13_L8}), .b ({new_AGEMA_signal_9672, new_AGEMA_signal_9671, SubBytesIns_Inst_Sbox_13_L10}), .c ({new_AGEMA_signal_10106, new_AGEMA_signal_10105, SubBytesIns_Inst_Sbox_13_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L28_U1 ( .a ({new_AGEMA_signal_9674, new_AGEMA_signal_9673, SubBytesIns_Inst_Sbox_13_L11}), .b ({new_AGEMA_signal_9310, new_AGEMA_signal_9309, SubBytesIns_Inst_Sbox_13_L14}), .c ({new_AGEMA_signal_10108, new_AGEMA_signal_10107, SubBytesIns_Inst_Sbox_13_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L29_U1 ( .a ({new_AGEMA_signal_9674, new_AGEMA_signal_9673, SubBytesIns_Inst_Sbox_13_L11}), .b ({new_AGEMA_signal_9314, new_AGEMA_signal_9313, SubBytesIns_Inst_Sbox_13_L17}), .c ({new_AGEMA_signal_10110, new_AGEMA_signal_10109, SubBytesIns_Inst_Sbox_13_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S0_U1 ( .a ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_10100, new_AGEMA_signal_10099, SubBytesIns_Inst_Sbox_13_L24}), .c ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S1_U1 ( .a ({new_AGEMA_signal_10094, new_AGEMA_signal_10093, SubBytesIns_Inst_Sbox_13_L16}), .b ({new_AGEMA_signal_10104, new_AGEMA_signal_10103, SubBytesIns_Inst_Sbox_13_L26}), .c ({new_AGEMA_signal_10406, new_AGEMA_signal_10405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S2_U1 ( .a ({new_AGEMA_signal_9676, new_AGEMA_signal_9675, SubBytesIns_Inst_Sbox_13_L19}), .b ({new_AGEMA_signal_10108, new_AGEMA_signal_10107, SubBytesIns_Inst_Sbox_13_L28}), .c ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S3_U1 ( .a ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_10098, new_AGEMA_signal_10097, SubBytesIns_Inst_Sbox_13_L21}), .c ({new_AGEMA_signal_10410, new_AGEMA_signal_10409, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S4_U1 ( .a ({new_AGEMA_signal_10096, new_AGEMA_signal_10095, SubBytesIns_Inst_Sbox_13_L20}), .b ({new_AGEMA_signal_9678, new_AGEMA_signal_9677, SubBytesIns_Inst_Sbox_13_L22}), .c ({new_AGEMA_signal_10412, new_AGEMA_signal_10411, MixColumnsInput[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S5_U1 ( .a ({new_AGEMA_signal_10102, new_AGEMA_signal_10101, SubBytesIns_Inst_Sbox_13_L25}), .b ({new_AGEMA_signal_10110, new_AGEMA_signal_10109, SubBytesIns_Inst_Sbox_13_L29}), .c ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, MixColumnsInput[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S6_U1 ( .a ({new_AGEMA_signal_10092, new_AGEMA_signal_10091, SubBytesIns_Inst_Sbox_13_L13}), .b ({new_AGEMA_signal_10106, new_AGEMA_signal_10105, SubBytesIns_Inst_Sbox_13_L27}), .c ({new_AGEMA_signal_10416, new_AGEMA_signal_10415, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S7_U1 ( .a ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_9680, new_AGEMA_signal_9679, SubBytesIns_Inst_Sbox_13_L23}), .c ({new_AGEMA_signal_10112, new_AGEMA_signal_10111, MixColumnsInput[40]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M46_U1 ( .a ({new_AGEMA_signal_8436, new_AGEMA_signal_8435, SubBytesIns_Inst_Sbox_14_M44}), .b ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, SubBytesIns_Inst_Sbox_14_T6}), .clk (clk), .r ({Fresh[1718], Fresh[1717], Fresh[1716]}), .c ({new_AGEMA_signal_8912, new_AGEMA_signal_8911, SubBytesIns_Inst_Sbox_14_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M47_U1 ( .a ({new_AGEMA_signal_7988, new_AGEMA_signal_7987, SubBytesIns_Inst_Sbox_14_M40}), .b ({new_AGEMA_signal_6506, new_AGEMA_signal_6505, SubBytesIns_Inst_Sbox_14_T8}), .clk (clk), .r ({Fresh[1721], Fresh[1720], Fresh[1719]}), .c ({new_AGEMA_signal_8438, new_AGEMA_signal_8437, SubBytesIns_Inst_Sbox_14_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M48_U1 ( .a ({new_AGEMA_signal_7986, new_AGEMA_signal_7985, SubBytesIns_Inst_Sbox_14_M39}), .b ({ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .clk (clk), .r ({Fresh[1724], Fresh[1723], Fresh[1722]}), .c ({new_AGEMA_signal_8440, new_AGEMA_signal_8439, SubBytesIns_Inst_Sbox_14_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M49_U1 ( .a ({new_AGEMA_signal_8434, new_AGEMA_signal_8433, SubBytesIns_Inst_Sbox_14_M43}), .b ({new_AGEMA_signal_6014, new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_14_T16}), .clk (clk), .r ({Fresh[1727], Fresh[1726], Fresh[1725]}), .c ({new_AGEMA_signal_8914, new_AGEMA_signal_8913, SubBytesIns_Inst_Sbox_14_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M50_U1 ( .a ({new_AGEMA_signal_7984, new_AGEMA_signal_7983, SubBytesIns_Inst_Sbox_14_M38}), .b ({new_AGEMA_signal_6008, new_AGEMA_signal_6007, SubBytesIns_Inst_Sbox_14_T9}), .clk (clk), .r ({Fresh[1730], Fresh[1729], Fresh[1728]}), .c ({new_AGEMA_signal_8442, new_AGEMA_signal_8441, SubBytesIns_Inst_Sbox_14_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M51_U1 ( .a ({new_AGEMA_signal_7982, new_AGEMA_signal_7981, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_6512, new_AGEMA_signal_6511, SubBytesIns_Inst_Sbox_14_T17}), .clk (clk), .r ({Fresh[1733], Fresh[1732], Fresh[1731]}), .c ({new_AGEMA_signal_8444, new_AGEMA_signal_8443, SubBytesIns_Inst_Sbox_14_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M52_U1 ( .a ({new_AGEMA_signal_8432, new_AGEMA_signal_8431, SubBytesIns_Inst_Sbox_14_M42}), .b ({new_AGEMA_signal_6012, new_AGEMA_signal_6011, SubBytesIns_Inst_Sbox_14_T15}), .clk (clk), .r ({Fresh[1736], Fresh[1735], Fresh[1734]}), .c ({new_AGEMA_signal_8916, new_AGEMA_signal_8915, SubBytesIns_Inst_Sbox_14_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M53_U1 ( .a ({new_AGEMA_signal_8910, new_AGEMA_signal_8909, SubBytesIns_Inst_Sbox_14_M45}), .b ({new_AGEMA_signal_6020, new_AGEMA_signal_6019, SubBytesIns_Inst_Sbox_14_T27}), .clk (clk), .r ({Fresh[1739], Fresh[1738], Fresh[1737]}), .c ({new_AGEMA_signal_9318, new_AGEMA_signal_9317, SubBytesIns_Inst_Sbox_14_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M54_U1 ( .a ({new_AGEMA_signal_8430, new_AGEMA_signal_8429, SubBytesIns_Inst_Sbox_14_M41}), .b ({new_AGEMA_signal_6508, new_AGEMA_signal_6507, SubBytesIns_Inst_Sbox_14_T10}), .clk (clk), .r ({Fresh[1742], Fresh[1741], Fresh[1740]}), .c ({new_AGEMA_signal_8918, new_AGEMA_signal_8917, SubBytesIns_Inst_Sbox_14_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M55_U1 ( .a ({new_AGEMA_signal_8436, new_AGEMA_signal_8435, SubBytesIns_Inst_Sbox_14_M44}), .b ({new_AGEMA_signal_6010, new_AGEMA_signal_6009, SubBytesIns_Inst_Sbox_14_T13}), .clk (clk), .r ({Fresh[1745], Fresh[1744], Fresh[1743]}), .c ({new_AGEMA_signal_8920, new_AGEMA_signal_8919, SubBytesIns_Inst_Sbox_14_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M56_U1 ( .a ({new_AGEMA_signal_7988, new_AGEMA_signal_7987, SubBytesIns_Inst_Sbox_14_M40}), .b ({new_AGEMA_signal_6516, new_AGEMA_signal_6515, SubBytesIns_Inst_Sbox_14_T23}), .clk (clk), .r ({Fresh[1748], Fresh[1747], Fresh[1746]}), .c ({new_AGEMA_signal_8446, new_AGEMA_signal_8445, SubBytesIns_Inst_Sbox_14_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M57_U1 ( .a ({new_AGEMA_signal_7986, new_AGEMA_signal_7985, SubBytesIns_Inst_Sbox_14_M39}), .b ({new_AGEMA_signal_6016, new_AGEMA_signal_6015, SubBytesIns_Inst_Sbox_14_T19}), .clk (clk), .r ({Fresh[1751], Fresh[1750], Fresh[1749]}), .c ({new_AGEMA_signal_8448, new_AGEMA_signal_8447, SubBytesIns_Inst_Sbox_14_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M58_U1 ( .a ({new_AGEMA_signal_8434, new_AGEMA_signal_8433, SubBytesIns_Inst_Sbox_14_M43}), .b ({new_AGEMA_signal_5682, new_AGEMA_signal_5681, SubBytesIns_Inst_Sbox_14_T3}), .clk (clk), .r ({Fresh[1754], Fresh[1753], Fresh[1752]}), .c ({new_AGEMA_signal_8922, new_AGEMA_signal_8921, SubBytesIns_Inst_Sbox_14_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M59_U1 ( .a ({new_AGEMA_signal_7984, new_AGEMA_signal_7983, SubBytesIns_Inst_Sbox_14_M38}), .b ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, SubBytesIns_Inst_Sbox_14_T22}), .clk (clk), .r ({Fresh[1757], Fresh[1756], Fresh[1755]}), .c ({new_AGEMA_signal_8450, new_AGEMA_signal_8449, SubBytesIns_Inst_Sbox_14_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M60_U1 ( .a ({new_AGEMA_signal_7982, new_AGEMA_signal_7981, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_6514, new_AGEMA_signal_6513, SubBytesIns_Inst_Sbox_14_T20}), .clk (clk), .r ({Fresh[1760], Fresh[1759], Fresh[1758]}), .c ({new_AGEMA_signal_8452, new_AGEMA_signal_8451, SubBytesIns_Inst_Sbox_14_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M61_U1 ( .a ({new_AGEMA_signal_8432, new_AGEMA_signal_8431, SubBytesIns_Inst_Sbox_14_M42}), .b ({new_AGEMA_signal_5678, new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_14_T1}), .clk (clk), .r ({Fresh[1763], Fresh[1762], Fresh[1761]}), .c ({new_AGEMA_signal_8924, new_AGEMA_signal_8923, SubBytesIns_Inst_Sbox_14_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M62_U1 ( .a ({new_AGEMA_signal_8910, new_AGEMA_signal_8909, SubBytesIns_Inst_Sbox_14_M45}), .b ({new_AGEMA_signal_5684, new_AGEMA_signal_5683, SubBytesIns_Inst_Sbox_14_T4}), .clk (clk), .r ({Fresh[1766], Fresh[1765], Fresh[1764]}), .c ({new_AGEMA_signal_9320, new_AGEMA_signal_9319, SubBytesIns_Inst_Sbox_14_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M63_U1 ( .a ({new_AGEMA_signal_8430, new_AGEMA_signal_8429, SubBytesIns_Inst_Sbox_14_M41}), .b ({new_AGEMA_signal_5680, new_AGEMA_signal_5679, SubBytesIns_Inst_Sbox_14_T2}), .clk (clk), .r ({Fresh[1769], Fresh[1768], Fresh[1767]}), .c ({new_AGEMA_signal_8926, new_AGEMA_signal_8925, SubBytesIns_Inst_Sbox_14_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L0_U1 ( .a ({new_AGEMA_signal_8924, new_AGEMA_signal_8923, SubBytesIns_Inst_Sbox_14_M61}), .b ({new_AGEMA_signal_9320, new_AGEMA_signal_9319, SubBytesIns_Inst_Sbox_14_M62}), .c ({new_AGEMA_signal_9682, new_AGEMA_signal_9681, SubBytesIns_Inst_Sbox_14_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L1_U1 ( .a ({new_AGEMA_signal_8442, new_AGEMA_signal_8441, SubBytesIns_Inst_Sbox_14_M50}), .b ({new_AGEMA_signal_8446, new_AGEMA_signal_8445, SubBytesIns_Inst_Sbox_14_M56}), .c ({new_AGEMA_signal_8928, new_AGEMA_signal_8927, SubBytesIns_Inst_Sbox_14_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L2_U1 ( .a ({new_AGEMA_signal_8912, new_AGEMA_signal_8911, SubBytesIns_Inst_Sbox_14_M46}), .b ({new_AGEMA_signal_8440, new_AGEMA_signal_8439, SubBytesIns_Inst_Sbox_14_M48}), .c ({new_AGEMA_signal_9322, new_AGEMA_signal_9321, SubBytesIns_Inst_Sbox_14_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L3_U1 ( .a ({new_AGEMA_signal_8438, new_AGEMA_signal_8437, SubBytesIns_Inst_Sbox_14_M47}), .b ({new_AGEMA_signal_8920, new_AGEMA_signal_8919, SubBytesIns_Inst_Sbox_14_M55}), .c ({new_AGEMA_signal_9324, new_AGEMA_signal_9323, SubBytesIns_Inst_Sbox_14_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L4_U1 ( .a ({new_AGEMA_signal_8918, new_AGEMA_signal_8917, SubBytesIns_Inst_Sbox_14_M54}), .b ({new_AGEMA_signal_8922, new_AGEMA_signal_8921, SubBytesIns_Inst_Sbox_14_M58}), .c ({new_AGEMA_signal_9326, new_AGEMA_signal_9325, SubBytesIns_Inst_Sbox_14_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L5_U1 ( .a ({new_AGEMA_signal_8914, new_AGEMA_signal_8913, SubBytesIns_Inst_Sbox_14_M49}), .b ({new_AGEMA_signal_8924, new_AGEMA_signal_8923, SubBytesIns_Inst_Sbox_14_M61}), .c ({new_AGEMA_signal_9328, new_AGEMA_signal_9327, SubBytesIns_Inst_Sbox_14_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L6_U1 ( .a ({new_AGEMA_signal_9320, new_AGEMA_signal_9319, SubBytesIns_Inst_Sbox_14_M62}), .b ({new_AGEMA_signal_9328, new_AGEMA_signal_9327, SubBytesIns_Inst_Sbox_14_L5}), .c ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, SubBytesIns_Inst_Sbox_14_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L7_U1 ( .a ({new_AGEMA_signal_8912, new_AGEMA_signal_8911, SubBytesIns_Inst_Sbox_14_M46}), .b ({new_AGEMA_signal_9324, new_AGEMA_signal_9323, SubBytesIns_Inst_Sbox_14_L3}), .c ({new_AGEMA_signal_9686, new_AGEMA_signal_9685, SubBytesIns_Inst_Sbox_14_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L8_U1 ( .a ({new_AGEMA_signal_8444, new_AGEMA_signal_8443, SubBytesIns_Inst_Sbox_14_M51}), .b ({new_AGEMA_signal_8450, new_AGEMA_signal_8449, SubBytesIns_Inst_Sbox_14_M59}), .c ({new_AGEMA_signal_8930, new_AGEMA_signal_8929, SubBytesIns_Inst_Sbox_14_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L9_U1 ( .a ({new_AGEMA_signal_8916, new_AGEMA_signal_8915, SubBytesIns_Inst_Sbox_14_M52}), .b ({new_AGEMA_signal_9318, new_AGEMA_signal_9317, SubBytesIns_Inst_Sbox_14_M53}), .c ({new_AGEMA_signal_9688, new_AGEMA_signal_9687, SubBytesIns_Inst_Sbox_14_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L10_U1 ( .a ({new_AGEMA_signal_9318, new_AGEMA_signal_9317, SubBytesIns_Inst_Sbox_14_M53}), .b ({new_AGEMA_signal_9326, new_AGEMA_signal_9325, SubBytesIns_Inst_Sbox_14_L4}), .c ({new_AGEMA_signal_9690, new_AGEMA_signal_9689, SubBytesIns_Inst_Sbox_14_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L11_U1 ( .a ({new_AGEMA_signal_8452, new_AGEMA_signal_8451, SubBytesIns_Inst_Sbox_14_M60}), .b ({new_AGEMA_signal_9322, new_AGEMA_signal_9321, SubBytesIns_Inst_Sbox_14_L2}), .c ({new_AGEMA_signal_9692, new_AGEMA_signal_9691, SubBytesIns_Inst_Sbox_14_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L12_U1 ( .a ({new_AGEMA_signal_8440, new_AGEMA_signal_8439, SubBytesIns_Inst_Sbox_14_M48}), .b ({new_AGEMA_signal_8444, new_AGEMA_signal_8443, SubBytesIns_Inst_Sbox_14_M51}), .c ({new_AGEMA_signal_8932, new_AGEMA_signal_8931, SubBytesIns_Inst_Sbox_14_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L13_U1 ( .a ({new_AGEMA_signal_8442, new_AGEMA_signal_8441, SubBytesIns_Inst_Sbox_14_M50}), .b ({new_AGEMA_signal_9682, new_AGEMA_signal_9681, SubBytesIns_Inst_Sbox_14_L0}), .c ({new_AGEMA_signal_10114, new_AGEMA_signal_10113, SubBytesIns_Inst_Sbox_14_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L14_U1 ( .a ({new_AGEMA_signal_8916, new_AGEMA_signal_8915, SubBytesIns_Inst_Sbox_14_M52}), .b ({new_AGEMA_signal_8924, new_AGEMA_signal_8923, SubBytesIns_Inst_Sbox_14_M61}), .c ({new_AGEMA_signal_9330, new_AGEMA_signal_9329, SubBytesIns_Inst_Sbox_14_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L15_U1 ( .a ({new_AGEMA_signal_8920, new_AGEMA_signal_8919, SubBytesIns_Inst_Sbox_14_M55}), .b ({new_AGEMA_signal_8928, new_AGEMA_signal_8927, SubBytesIns_Inst_Sbox_14_L1}), .c ({new_AGEMA_signal_9332, new_AGEMA_signal_9331, SubBytesIns_Inst_Sbox_14_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L16_U1 ( .a ({new_AGEMA_signal_8446, new_AGEMA_signal_8445, SubBytesIns_Inst_Sbox_14_M56}), .b ({new_AGEMA_signal_9682, new_AGEMA_signal_9681, SubBytesIns_Inst_Sbox_14_L0}), .c ({new_AGEMA_signal_10116, new_AGEMA_signal_10115, SubBytesIns_Inst_Sbox_14_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L17_U1 ( .a ({new_AGEMA_signal_8448, new_AGEMA_signal_8447, SubBytesIns_Inst_Sbox_14_M57}), .b ({new_AGEMA_signal_8928, new_AGEMA_signal_8927, SubBytesIns_Inst_Sbox_14_L1}), .c ({new_AGEMA_signal_9334, new_AGEMA_signal_9333, SubBytesIns_Inst_Sbox_14_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L18_U1 ( .a ({new_AGEMA_signal_8922, new_AGEMA_signal_8921, SubBytesIns_Inst_Sbox_14_M58}), .b ({new_AGEMA_signal_8930, new_AGEMA_signal_8929, SubBytesIns_Inst_Sbox_14_L8}), .c ({new_AGEMA_signal_9336, new_AGEMA_signal_9335, SubBytesIns_Inst_Sbox_14_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L19_U1 ( .a ({new_AGEMA_signal_8926, new_AGEMA_signal_8925, SubBytesIns_Inst_Sbox_14_M63}), .b ({new_AGEMA_signal_9326, new_AGEMA_signal_9325, SubBytesIns_Inst_Sbox_14_L4}), .c ({new_AGEMA_signal_9694, new_AGEMA_signal_9693, SubBytesIns_Inst_Sbox_14_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L20_U1 ( .a ({new_AGEMA_signal_9682, new_AGEMA_signal_9681, SubBytesIns_Inst_Sbox_14_L0}), .b ({new_AGEMA_signal_8928, new_AGEMA_signal_8927, SubBytesIns_Inst_Sbox_14_L1}), .c ({new_AGEMA_signal_10118, new_AGEMA_signal_10117, SubBytesIns_Inst_Sbox_14_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L21_U1 ( .a ({new_AGEMA_signal_8928, new_AGEMA_signal_8927, SubBytesIns_Inst_Sbox_14_L1}), .b ({new_AGEMA_signal_9686, new_AGEMA_signal_9685, SubBytesIns_Inst_Sbox_14_L7}), .c ({new_AGEMA_signal_10120, new_AGEMA_signal_10119, SubBytesIns_Inst_Sbox_14_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L22_U1 ( .a ({new_AGEMA_signal_9324, new_AGEMA_signal_9323, SubBytesIns_Inst_Sbox_14_L3}), .b ({new_AGEMA_signal_8932, new_AGEMA_signal_8931, SubBytesIns_Inst_Sbox_14_L12}), .c ({new_AGEMA_signal_9696, new_AGEMA_signal_9695, SubBytesIns_Inst_Sbox_14_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L23_U1 ( .a ({new_AGEMA_signal_9336, new_AGEMA_signal_9335, SubBytesIns_Inst_Sbox_14_L18}), .b ({new_AGEMA_signal_9322, new_AGEMA_signal_9321, SubBytesIns_Inst_Sbox_14_L2}), .c ({new_AGEMA_signal_9698, new_AGEMA_signal_9697, SubBytesIns_Inst_Sbox_14_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L24_U1 ( .a ({new_AGEMA_signal_9332, new_AGEMA_signal_9331, SubBytesIns_Inst_Sbox_14_L15}), .b ({new_AGEMA_signal_9688, new_AGEMA_signal_9687, SubBytesIns_Inst_Sbox_14_L9}), .c ({new_AGEMA_signal_10122, new_AGEMA_signal_10121, SubBytesIns_Inst_Sbox_14_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L25_U1 ( .a ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_9690, new_AGEMA_signal_9689, SubBytesIns_Inst_Sbox_14_L10}), .c ({new_AGEMA_signal_10124, new_AGEMA_signal_10123, SubBytesIns_Inst_Sbox_14_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L26_U1 ( .a ({new_AGEMA_signal_9686, new_AGEMA_signal_9685, SubBytesIns_Inst_Sbox_14_L7}), .b ({new_AGEMA_signal_9688, new_AGEMA_signal_9687, SubBytesIns_Inst_Sbox_14_L9}), .c ({new_AGEMA_signal_10126, new_AGEMA_signal_10125, SubBytesIns_Inst_Sbox_14_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L27_U1 ( .a ({new_AGEMA_signal_8930, new_AGEMA_signal_8929, SubBytesIns_Inst_Sbox_14_L8}), .b ({new_AGEMA_signal_9690, new_AGEMA_signal_9689, SubBytesIns_Inst_Sbox_14_L10}), .c ({new_AGEMA_signal_10128, new_AGEMA_signal_10127, SubBytesIns_Inst_Sbox_14_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L28_U1 ( .a ({new_AGEMA_signal_9692, new_AGEMA_signal_9691, SubBytesIns_Inst_Sbox_14_L11}), .b ({new_AGEMA_signal_9330, new_AGEMA_signal_9329, SubBytesIns_Inst_Sbox_14_L14}), .c ({new_AGEMA_signal_10130, new_AGEMA_signal_10129, SubBytesIns_Inst_Sbox_14_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L29_U1 ( .a ({new_AGEMA_signal_9692, new_AGEMA_signal_9691, SubBytesIns_Inst_Sbox_14_L11}), .b ({new_AGEMA_signal_9334, new_AGEMA_signal_9333, SubBytesIns_Inst_Sbox_14_L17}), .c ({new_AGEMA_signal_10132, new_AGEMA_signal_10131, SubBytesIns_Inst_Sbox_14_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S0_U1 ( .a ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_10122, new_AGEMA_signal_10121, SubBytesIns_Inst_Sbox_14_L24}), .c ({new_AGEMA_signal_10418, new_AGEMA_signal_10417, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S1_U1 ( .a ({new_AGEMA_signal_10116, new_AGEMA_signal_10115, SubBytesIns_Inst_Sbox_14_L16}), .b ({new_AGEMA_signal_10126, new_AGEMA_signal_10125, SubBytesIns_Inst_Sbox_14_L26}), .c ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S2_U1 ( .a ({new_AGEMA_signal_9694, new_AGEMA_signal_9693, SubBytesIns_Inst_Sbox_14_L19}), .b ({new_AGEMA_signal_10130, new_AGEMA_signal_10129, SubBytesIns_Inst_Sbox_14_L28}), .c ({new_AGEMA_signal_10422, new_AGEMA_signal_10421, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S3_U1 ( .a ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_10120, new_AGEMA_signal_10119, SubBytesIns_Inst_Sbox_14_L21}), .c ({new_AGEMA_signal_10424, new_AGEMA_signal_10423, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S4_U1 ( .a ({new_AGEMA_signal_10118, new_AGEMA_signal_10117, SubBytesIns_Inst_Sbox_14_L20}), .b ({new_AGEMA_signal_9696, new_AGEMA_signal_9695, SubBytesIns_Inst_Sbox_14_L22}), .c ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, MixColumnsInput[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S5_U1 ( .a ({new_AGEMA_signal_10124, new_AGEMA_signal_10123, SubBytesIns_Inst_Sbox_14_L25}), .b ({new_AGEMA_signal_10132, new_AGEMA_signal_10131, SubBytesIns_Inst_Sbox_14_L29}), .c ({new_AGEMA_signal_10428, new_AGEMA_signal_10427, MixColumnsInput[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S6_U1 ( .a ({new_AGEMA_signal_10114, new_AGEMA_signal_10113, SubBytesIns_Inst_Sbox_14_L13}), .b ({new_AGEMA_signal_10128, new_AGEMA_signal_10127, SubBytesIns_Inst_Sbox_14_L27}), .c ({new_AGEMA_signal_10430, new_AGEMA_signal_10429, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S7_U1 ( .a ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_9698, new_AGEMA_signal_9697, SubBytesIns_Inst_Sbox_14_L23}), .c ({new_AGEMA_signal_10134, new_AGEMA_signal_10133, MixColumnsInput[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M46_U1 ( .a ({new_AGEMA_signal_8460, new_AGEMA_signal_8459, SubBytesIns_Inst_Sbox_15_M44}), .b ({new_AGEMA_signal_6022, new_AGEMA_signal_6021, SubBytesIns_Inst_Sbox_15_T6}), .clk (clk), .r ({Fresh[1772], Fresh[1771], Fresh[1770]}), .c ({new_AGEMA_signal_8936, new_AGEMA_signal_8935, SubBytesIns_Inst_Sbox_15_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M47_U1 ( .a ({new_AGEMA_signal_7996, new_AGEMA_signal_7995, SubBytesIns_Inst_Sbox_15_M40}), .b ({new_AGEMA_signal_6532, new_AGEMA_signal_6531, SubBytesIns_Inst_Sbox_15_T8}), .clk (clk), .r ({Fresh[1775], Fresh[1774], Fresh[1773]}), .c ({new_AGEMA_signal_8462, new_AGEMA_signal_8461, SubBytesIns_Inst_Sbox_15_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M48_U1 ( .a ({new_AGEMA_signal_7994, new_AGEMA_signal_7993, SubBytesIns_Inst_Sbox_15_M39}), .b ({ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .clk (clk), .r ({Fresh[1778], Fresh[1777], Fresh[1776]}), .c ({new_AGEMA_signal_8464, new_AGEMA_signal_8463, SubBytesIns_Inst_Sbox_15_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M49_U1 ( .a ({new_AGEMA_signal_8458, new_AGEMA_signal_8457, SubBytesIns_Inst_Sbox_15_M43}), .b ({new_AGEMA_signal_6030, new_AGEMA_signal_6029, SubBytesIns_Inst_Sbox_15_T16}), .clk (clk), .r ({Fresh[1781], Fresh[1780], Fresh[1779]}), .c ({new_AGEMA_signal_8938, new_AGEMA_signal_8937, SubBytesIns_Inst_Sbox_15_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M50_U1 ( .a ({new_AGEMA_signal_7992, new_AGEMA_signal_7991, SubBytesIns_Inst_Sbox_15_M38}), .b ({new_AGEMA_signal_6024, new_AGEMA_signal_6023, SubBytesIns_Inst_Sbox_15_T9}), .clk (clk), .r ({Fresh[1784], Fresh[1783], Fresh[1782]}), .c ({new_AGEMA_signal_8466, new_AGEMA_signal_8465, SubBytesIns_Inst_Sbox_15_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M51_U1 ( .a ({new_AGEMA_signal_7990, new_AGEMA_signal_7989, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_6538, new_AGEMA_signal_6537, SubBytesIns_Inst_Sbox_15_T17}), .clk (clk), .r ({Fresh[1787], Fresh[1786], Fresh[1785]}), .c ({new_AGEMA_signal_8468, new_AGEMA_signal_8467, SubBytesIns_Inst_Sbox_15_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M52_U1 ( .a ({new_AGEMA_signal_8456, new_AGEMA_signal_8455, SubBytesIns_Inst_Sbox_15_M42}), .b ({new_AGEMA_signal_6028, new_AGEMA_signal_6027, SubBytesIns_Inst_Sbox_15_T15}), .clk (clk), .r ({Fresh[1790], Fresh[1789], Fresh[1788]}), .c ({new_AGEMA_signal_8940, new_AGEMA_signal_8939, SubBytesIns_Inst_Sbox_15_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M53_U1 ( .a ({new_AGEMA_signal_8934, new_AGEMA_signal_8933, SubBytesIns_Inst_Sbox_15_M45}), .b ({new_AGEMA_signal_6036, new_AGEMA_signal_6035, SubBytesIns_Inst_Sbox_15_T27}), .clk (clk), .r ({Fresh[1793], Fresh[1792], Fresh[1791]}), .c ({new_AGEMA_signal_9338, new_AGEMA_signal_9337, SubBytesIns_Inst_Sbox_15_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M54_U1 ( .a ({new_AGEMA_signal_8454, new_AGEMA_signal_8453, SubBytesIns_Inst_Sbox_15_M41}), .b ({new_AGEMA_signal_6534, new_AGEMA_signal_6533, SubBytesIns_Inst_Sbox_15_T10}), .clk (clk), .r ({Fresh[1796], Fresh[1795], Fresh[1794]}), .c ({new_AGEMA_signal_8942, new_AGEMA_signal_8941, SubBytesIns_Inst_Sbox_15_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M55_U1 ( .a ({new_AGEMA_signal_8460, new_AGEMA_signal_8459, SubBytesIns_Inst_Sbox_15_M44}), .b ({new_AGEMA_signal_6026, new_AGEMA_signal_6025, SubBytesIns_Inst_Sbox_15_T13}), .clk (clk), .r ({Fresh[1799], Fresh[1798], Fresh[1797]}), .c ({new_AGEMA_signal_8944, new_AGEMA_signal_8943, SubBytesIns_Inst_Sbox_15_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M56_U1 ( .a ({new_AGEMA_signal_7996, new_AGEMA_signal_7995, SubBytesIns_Inst_Sbox_15_M40}), .b ({new_AGEMA_signal_6542, new_AGEMA_signal_6541, SubBytesIns_Inst_Sbox_15_T23}), .clk (clk), .r ({Fresh[1802], Fresh[1801], Fresh[1800]}), .c ({new_AGEMA_signal_8470, new_AGEMA_signal_8469, SubBytesIns_Inst_Sbox_15_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M57_U1 ( .a ({new_AGEMA_signal_7994, new_AGEMA_signal_7993, SubBytesIns_Inst_Sbox_15_M39}), .b ({new_AGEMA_signal_6032, new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_15_T19}), .clk (clk), .r ({Fresh[1805], Fresh[1804], Fresh[1803]}), .c ({new_AGEMA_signal_8472, new_AGEMA_signal_8471, SubBytesIns_Inst_Sbox_15_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M58_U1 ( .a ({new_AGEMA_signal_8458, new_AGEMA_signal_8457, SubBytesIns_Inst_Sbox_15_M43}), .b ({new_AGEMA_signal_5702, new_AGEMA_signal_5701, SubBytesIns_Inst_Sbox_15_T3}), .clk (clk), .r ({Fresh[1808], Fresh[1807], Fresh[1806]}), .c ({new_AGEMA_signal_8946, new_AGEMA_signal_8945, SubBytesIns_Inst_Sbox_15_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M59_U1 ( .a ({new_AGEMA_signal_7992, new_AGEMA_signal_7991, SubBytesIns_Inst_Sbox_15_M38}), .b ({new_AGEMA_signal_6034, new_AGEMA_signal_6033, SubBytesIns_Inst_Sbox_15_T22}), .clk (clk), .r ({Fresh[1811], Fresh[1810], Fresh[1809]}), .c ({new_AGEMA_signal_8474, new_AGEMA_signal_8473, SubBytesIns_Inst_Sbox_15_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M60_U1 ( .a ({new_AGEMA_signal_7990, new_AGEMA_signal_7989, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_6540, new_AGEMA_signal_6539, SubBytesIns_Inst_Sbox_15_T20}), .clk (clk), .r ({Fresh[1814], Fresh[1813], Fresh[1812]}), .c ({new_AGEMA_signal_8476, new_AGEMA_signal_8475, SubBytesIns_Inst_Sbox_15_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M61_U1 ( .a ({new_AGEMA_signal_8456, new_AGEMA_signal_8455, SubBytesIns_Inst_Sbox_15_M42}), .b ({new_AGEMA_signal_5698, new_AGEMA_signal_5697, SubBytesIns_Inst_Sbox_15_T1}), .clk (clk), .r ({Fresh[1817], Fresh[1816], Fresh[1815]}), .c ({new_AGEMA_signal_8948, new_AGEMA_signal_8947, SubBytesIns_Inst_Sbox_15_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M62_U1 ( .a ({new_AGEMA_signal_8934, new_AGEMA_signal_8933, SubBytesIns_Inst_Sbox_15_M45}), .b ({new_AGEMA_signal_5704, new_AGEMA_signal_5703, SubBytesIns_Inst_Sbox_15_T4}), .clk (clk), .r ({Fresh[1820], Fresh[1819], Fresh[1818]}), .c ({new_AGEMA_signal_9340, new_AGEMA_signal_9339, SubBytesIns_Inst_Sbox_15_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M63_U1 ( .a ({new_AGEMA_signal_8454, new_AGEMA_signal_8453, SubBytesIns_Inst_Sbox_15_M41}), .b ({new_AGEMA_signal_5700, new_AGEMA_signal_5699, SubBytesIns_Inst_Sbox_15_T2}), .clk (clk), .r ({Fresh[1823], Fresh[1822], Fresh[1821]}), .c ({new_AGEMA_signal_8950, new_AGEMA_signal_8949, SubBytesIns_Inst_Sbox_15_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L0_U1 ( .a ({new_AGEMA_signal_8948, new_AGEMA_signal_8947, SubBytesIns_Inst_Sbox_15_M61}), .b ({new_AGEMA_signal_9340, new_AGEMA_signal_9339, SubBytesIns_Inst_Sbox_15_M62}), .c ({new_AGEMA_signal_9700, new_AGEMA_signal_9699, SubBytesIns_Inst_Sbox_15_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L1_U1 ( .a ({new_AGEMA_signal_8466, new_AGEMA_signal_8465, SubBytesIns_Inst_Sbox_15_M50}), .b ({new_AGEMA_signal_8470, new_AGEMA_signal_8469, SubBytesIns_Inst_Sbox_15_M56}), .c ({new_AGEMA_signal_8952, new_AGEMA_signal_8951, SubBytesIns_Inst_Sbox_15_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L2_U1 ( .a ({new_AGEMA_signal_8936, new_AGEMA_signal_8935, SubBytesIns_Inst_Sbox_15_M46}), .b ({new_AGEMA_signal_8464, new_AGEMA_signal_8463, SubBytesIns_Inst_Sbox_15_M48}), .c ({new_AGEMA_signal_9342, new_AGEMA_signal_9341, SubBytesIns_Inst_Sbox_15_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L3_U1 ( .a ({new_AGEMA_signal_8462, new_AGEMA_signal_8461, SubBytesIns_Inst_Sbox_15_M47}), .b ({new_AGEMA_signal_8944, new_AGEMA_signal_8943, SubBytesIns_Inst_Sbox_15_M55}), .c ({new_AGEMA_signal_9344, new_AGEMA_signal_9343, SubBytesIns_Inst_Sbox_15_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L4_U1 ( .a ({new_AGEMA_signal_8942, new_AGEMA_signal_8941, SubBytesIns_Inst_Sbox_15_M54}), .b ({new_AGEMA_signal_8946, new_AGEMA_signal_8945, SubBytesIns_Inst_Sbox_15_M58}), .c ({new_AGEMA_signal_9346, new_AGEMA_signal_9345, SubBytesIns_Inst_Sbox_15_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L5_U1 ( .a ({new_AGEMA_signal_8938, new_AGEMA_signal_8937, SubBytesIns_Inst_Sbox_15_M49}), .b ({new_AGEMA_signal_8948, new_AGEMA_signal_8947, SubBytesIns_Inst_Sbox_15_M61}), .c ({new_AGEMA_signal_9348, new_AGEMA_signal_9347, SubBytesIns_Inst_Sbox_15_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L6_U1 ( .a ({new_AGEMA_signal_9340, new_AGEMA_signal_9339, SubBytesIns_Inst_Sbox_15_M62}), .b ({new_AGEMA_signal_9348, new_AGEMA_signal_9347, SubBytesIns_Inst_Sbox_15_L5}), .c ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, SubBytesIns_Inst_Sbox_15_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L7_U1 ( .a ({new_AGEMA_signal_8936, new_AGEMA_signal_8935, SubBytesIns_Inst_Sbox_15_M46}), .b ({new_AGEMA_signal_9344, new_AGEMA_signal_9343, SubBytesIns_Inst_Sbox_15_L3}), .c ({new_AGEMA_signal_9704, new_AGEMA_signal_9703, SubBytesIns_Inst_Sbox_15_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L8_U1 ( .a ({new_AGEMA_signal_8468, new_AGEMA_signal_8467, SubBytesIns_Inst_Sbox_15_M51}), .b ({new_AGEMA_signal_8474, new_AGEMA_signal_8473, SubBytesIns_Inst_Sbox_15_M59}), .c ({new_AGEMA_signal_8954, new_AGEMA_signal_8953, SubBytesIns_Inst_Sbox_15_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L9_U1 ( .a ({new_AGEMA_signal_8940, new_AGEMA_signal_8939, SubBytesIns_Inst_Sbox_15_M52}), .b ({new_AGEMA_signal_9338, new_AGEMA_signal_9337, SubBytesIns_Inst_Sbox_15_M53}), .c ({new_AGEMA_signal_9706, new_AGEMA_signal_9705, SubBytesIns_Inst_Sbox_15_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L10_U1 ( .a ({new_AGEMA_signal_9338, new_AGEMA_signal_9337, SubBytesIns_Inst_Sbox_15_M53}), .b ({new_AGEMA_signal_9346, new_AGEMA_signal_9345, SubBytesIns_Inst_Sbox_15_L4}), .c ({new_AGEMA_signal_9708, new_AGEMA_signal_9707, SubBytesIns_Inst_Sbox_15_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L11_U1 ( .a ({new_AGEMA_signal_8476, new_AGEMA_signal_8475, SubBytesIns_Inst_Sbox_15_M60}), .b ({new_AGEMA_signal_9342, new_AGEMA_signal_9341, SubBytesIns_Inst_Sbox_15_L2}), .c ({new_AGEMA_signal_9710, new_AGEMA_signal_9709, SubBytesIns_Inst_Sbox_15_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L12_U1 ( .a ({new_AGEMA_signal_8464, new_AGEMA_signal_8463, SubBytesIns_Inst_Sbox_15_M48}), .b ({new_AGEMA_signal_8468, new_AGEMA_signal_8467, SubBytesIns_Inst_Sbox_15_M51}), .c ({new_AGEMA_signal_8956, new_AGEMA_signal_8955, SubBytesIns_Inst_Sbox_15_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L13_U1 ( .a ({new_AGEMA_signal_8466, new_AGEMA_signal_8465, SubBytesIns_Inst_Sbox_15_M50}), .b ({new_AGEMA_signal_9700, new_AGEMA_signal_9699, SubBytesIns_Inst_Sbox_15_L0}), .c ({new_AGEMA_signal_10136, new_AGEMA_signal_10135, SubBytesIns_Inst_Sbox_15_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L14_U1 ( .a ({new_AGEMA_signal_8940, new_AGEMA_signal_8939, SubBytesIns_Inst_Sbox_15_M52}), .b ({new_AGEMA_signal_8948, new_AGEMA_signal_8947, SubBytesIns_Inst_Sbox_15_M61}), .c ({new_AGEMA_signal_9350, new_AGEMA_signal_9349, SubBytesIns_Inst_Sbox_15_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L15_U1 ( .a ({new_AGEMA_signal_8944, new_AGEMA_signal_8943, SubBytesIns_Inst_Sbox_15_M55}), .b ({new_AGEMA_signal_8952, new_AGEMA_signal_8951, SubBytesIns_Inst_Sbox_15_L1}), .c ({new_AGEMA_signal_9352, new_AGEMA_signal_9351, SubBytesIns_Inst_Sbox_15_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L16_U1 ( .a ({new_AGEMA_signal_8470, new_AGEMA_signal_8469, SubBytesIns_Inst_Sbox_15_M56}), .b ({new_AGEMA_signal_9700, new_AGEMA_signal_9699, SubBytesIns_Inst_Sbox_15_L0}), .c ({new_AGEMA_signal_10138, new_AGEMA_signal_10137, SubBytesIns_Inst_Sbox_15_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L17_U1 ( .a ({new_AGEMA_signal_8472, new_AGEMA_signal_8471, SubBytesIns_Inst_Sbox_15_M57}), .b ({new_AGEMA_signal_8952, new_AGEMA_signal_8951, SubBytesIns_Inst_Sbox_15_L1}), .c ({new_AGEMA_signal_9354, new_AGEMA_signal_9353, SubBytesIns_Inst_Sbox_15_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L18_U1 ( .a ({new_AGEMA_signal_8946, new_AGEMA_signal_8945, SubBytesIns_Inst_Sbox_15_M58}), .b ({new_AGEMA_signal_8954, new_AGEMA_signal_8953, SubBytesIns_Inst_Sbox_15_L8}), .c ({new_AGEMA_signal_9356, new_AGEMA_signal_9355, SubBytesIns_Inst_Sbox_15_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L19_U1 ( .a ({new_AGEMA_signal_8950, new_AGEMA_signal_8949, SubBytesIns_Inst_Sbox_15_M63}), .b ({new_AGEMA_signal_9346, new_AGEMA_signal_9345, SubBytesIns_Inst_Sbox_15_L4}), .c ({new_AGEMA_signal_9712, new_AGEMA_signal_9711, SubBytesIns_Inst_Sbox_15_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L20_U1 ( .a ({new_AGEMA_signal_9700, new_AGEMA_signal_9699, SubBytesIns_Inst_Sbox_15_L0}), .b ({new_AGEMA_signal_8952, new_AGEMA_signal_8951, SubBytesIns_Inst_Sbox_15_L1}), .c ({new_AGEMA_signal_10140, new_AGEMA_signal_10139, SubBytesIns_Inst_Sbox_15_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L21_U1 ( .a ({new_AGEMA_signal_8952, new_AGEMA_signal_8951, SubBytesIns_Inst_Sbox_15_L1}), .b ({new_AGEMA_signal_9704, new_AGEMA_signal_9703, SubBytesIns_Inst_Sbox_15_L7}), .c ({new_AGEMA_signal_10142, new_AGEMA_signal_10141, SubBytesIns_Inst_Sbox_15_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L22_U1 ( .a ({new_AGEMA_signal_9344, new_AGEMA_signal_9343, SubBytesIns_Inst_Sbox_15_L3}), .b ({new_AGEMA_signal_8956, new_AGEMA_signal_8955, SubBytesIns_Inst_Sbox_15_L12}), .c ({new_AGEMA_signal_9714, new_AGEMA_signal_9713, SubBytesIns_Inst_Sbox_15_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L23_U1 ( .a ({new_AGEMA_signal_9356, new_AGEMA_signal_9355, SubBytesIns_Inst_Sbox_15_L18}), .b ({new_AGEMA_signal_9342, new_AGEMA_signal_9341, SubBytesIns_Inst_Sbox_15_L2}), .c ({new_AGEMA_signal_9716, new_AGEMA_signal_9715, SubBytesIns_Inst_Sbox_15_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L24_U1 ( .a ({new_AGEMA_signal_9352, new_AGEMA_signal_9351, SubBytesIns_Inst_Sbox_15_L15}), .b ({new_AGEMA_signal_9706, new_AGEMA_signal_9705, SubBytesIns_Inst_Sbox_15_L9}), .c ({new_AGEMA_signal_10144, new_AGEMA_signal_10143, SubBytesIns_Inst_Sbox_15_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L25_U1 ( .a ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_9708, new_AGEMA_signal_9707, SubBytesIns_Inst_Sbox_15_L10}), .c ({new_AGEMA_signal_10146, new_AGEMA_signal_10145, SubBytesIns_Inst_Sbox_15_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L26_U1 ( .a ({new_AGEMA_signal_9704, new_AGEMA_signal_9703, SubBytesIns_Inst_Sbox_15_L7}), .b ({new_AGEMA_signal_9706, new_AGEMA_signal_9705, SubBytesIns_Inst_Sbox_15_L9}), .c ({new_AGEMA_signal_10148, new_AGEMA_signal_10147, SubBytesIns_Inst_Sbox_15_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L27_U1 ( .a ({new_AGEMA_signal_8954, new_AGEMA_signal_8953, SubBytesIns_Inst_Sbox_15_L8}), .b ({new_AGEMA_signal_9708, new_AGEMA_signal_9707, SubBytesIns_Inst_Sbox_15_L10}), .c ({new_AGEMA_signal_10150, new_AGEMA_signal_10149, SubBytesIns_Inst_Sbox_15_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L28_U1 ( .a ({new_AGEMA_signal_9710, new_AGEMA_signal_9709, SubBytesIns_Inst_Sbox_15_L11}), .b ({new_AGEMA_signal_9350, new_AGEMA_signal_9349, SubBytesIns_Inst_Sbox_15_L14}), .c ({new_AGEMA_signal_10152, new_AGEMA_signal_10151, SubBytesIns_Inst_Sbox_15_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L29_U1 ( .a ({new_AGEMA_signal_9710, new_AGEMA_signal_9709, SubBytesIns_Inst_Sbox_15_L11}), .b ({new_AGEMA_signal_9354, new_AGEMA_signal_9353, SubBytesIns_Inst_Sbox_15_L17}), .c ({new_AGEMA_signal_10154, new_AGEMA_signal_10153, SubBytesIns_Inst_Sbox_15_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S0_U1 ( .a ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_10144, new_AGEMA_signal_10143, SubBytesIns_Inst_Sbox_15_L24}), .c ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S1_U1 ( .a ({new_AGEMA_signal_10138, new_AGEMA_signal_10137, SubBytesIns_Inst_Sbox_15_L16}), .b ({new_AGEMA_signal_10148, new_AGEMA_signal_10147, SubBytesIns_Inst_Sbox_15_L26}), .c ({new_AGEMA_signal_10434, new_AGEMA_signal_10433, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S2_U1 ( .a ({new_AGEMA_signal_9712, new_AGEMA_signal_9711, SubBytesIns_Inst_Sbox_15_L19}), .b ({new_AGEMA_signal_10152, new_AGEMA_signal_10151, SubBytesIns_Inst_Sbox_15_L28}), .c ({new_AGEMA_signal_10436, new_AGEMA_signal_10435, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S3_U1 ( .a ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_10142, new_AGEMA_signal_10141, SubBytesIns_Inst_Sbox_15_L21}), .c ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S4_U1 ( .a ({new_AGEMA_signal_10140, new_AGEMA_signal_10139, SubBytesIns_Inst_Sbox_15_L20}), .b ({new_AGEMA_signal_9714, new_AGEMA_signal_9713, SubBytesIns_Inst_Sbox_15_L22}), .c ({new_AGEMA_signal_10440, new_AGEMA_signal_10439, MixColumnsInput[123]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S5_U1 ( .a ({new_AGEMA_signal_10146, new_AGEMA_signal_10145, SubBytesIns_Inst_Sbox_15_L25}), .b ({new_AGEMA_signal_10154, new_AGEMA_signal_10153, SubBytesIns_Inst_Sbox_15_L29}), .c ({new_AGEMA_signal_10442, new_AGEMA_signal_10441, MixColumnsInput[122]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S6_U1 ( .a ({new_AGEMA_signal_10136, new_AGEMA_signal_10135, SubBytesIns_Inst_Sbox_15_L13}), .b ({new_AGEMA_signal_10150, new_AGEMA_signal_10149, SubBytesIns_Inst_Sbox_15_L27}), .c ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S7_U1 ( .a ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_9716, new_AGEMA_signal_9715, SubBytesIns_Inst_Sbox_15_L23}), .c ({new_AGEMA_signal_10156, new_AGEMA_signal_10155, MixColumnsInput[120]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U96 ( .a ({new_AGEMA_signal_11390, new_AGEMA_signal_11389, MixColumnsIns_MixOneColumnInst_0_n64}), .b ({new_AGEMA_signal_10374, new_AGEMA_signal_10373, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .c ({new_AGEMA_signal_11992, new_AGEMA_signal_11991, MixColumnsOutput[105]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U95 ( .a ({new_AGEMA_signal_10984, new_AGEMA_signal_10983, MixColumnsIns_MixOneColumnInst_0_n63}), .b ({new_AGEMA_signal_10976, new_AGEMA_signal_10975, MixColumnsIns_MixOneColumnInst_0_n62}), .c ({new_AGEMA_signal_11390, new_AGEMA_signal_11389, MixColumnsIns_MixOneColumnInst_0_n64}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U94 ( .a ({new_AGEMA_signal_10942, new_AGEMA_signal_10941, MixColumnsIns_MixOneColumnInst_0_n61}), .b ({new_AGEMA_signal_10540, new_AGEMA_signal_10539, MixColumnsIns_MixOneColumnInst_0_n60}), .c ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, MixColumnsOutput[104]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U93 ( .a ({new_AGEMA_signal_10560, new_AGEMA_signal_10559, MixColumnsIns_MixOneColumnInst_0_n59}), .b ({new_AGEMA_signal_10046, new_AGEMA_signal_10045, MixColumnsInput[112]}), .c ({new_AGEMA_signal_10942, new_AGEMA_signal_10941, MixColumnsIns_MixOneColumnInst_0_n61}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U92 ( .a ({new_AGEMA_signal_10944, new_AGEMA_signal_10943, MixColumnsIns_MixOneColumnInst_0_n58}), .b ({new_AGEMA_signal_10522, new_AGEMA_signal_10521, MixColumnsIns_MixOneColumnInst_0_n57}), .c ({new_AGEMA_signal_11394, new_AGEMA_signal_11393, MixColumnsOutput[103]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U91 ( .a ({new_AGEMA_signal_10544, new_AGEMA_signal_10543, MixColumnsIns_MixOneColumnInst_0_n56}), .b ({new_AGEMA_signal_10292, new_AGEMA_signal_10291, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .c ({new_AGEMA_signal_10944, new_AGEMA_signal_10943, MixColumnsIns_MixOneColumnInst_0_n58}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U90 ( .a ({new_AGEMA_signal_10946, new_AGEMA_signal_10945, MixColumnsIns_MixOneColumnInst_0_n55}), .b ({new_AGEMA_signal_10524, new_AGEMA_signal_10523, MixColumnsIns_MixOneColumnInst_0_n54}), .c ({new_AGEMA_signal_11396, new_AGEMA_signal_11395, MixColumnsOutput[102]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U89 ( .a ({new_AGEMA_signal_10548, new_AGEMA_signal_10547, MixColumnsIns_MixOneColumnInst_0_n53}), .b ({new_AGEMA_signal_10294, new_AGEMA_signal_10293, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .c ({new_AGEMA_signal_10946, new_AGEMA_signal_10945, MixColumnsIns_MixOneColumnInst_0_n55}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U88 ( .a ({new_AGEMA_signal_10948, new_AGEMA_signal_10947, MixColumnsIns_MixOneColumnInst_0_n52}), .b ({new_AGEMA_signal_10526, new_AGEMA_signal_10525, MixColumnsIns_MixOneColumnInst_0_n51}), .c ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, MixColumnsOutput[101]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U87 ( .a ({new_AGEMA_signal_10552, new_AGEMA_signal_10551, MixColumnsIns_MixOneColumnInst_0_n50}), .b ({new_AGEMA_signal_10296, new_AGEMA_signal_10295, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .c ({new_AGEMA_signal_10948, new_AGEMA_signal_10947, MixColumnsIns_MixOneColumnInst_0_n52}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U86 ( .a ({new_AGEMA_signal_11400, new_AGEMA_signal_11399, MixColumnsIns_MixOneColumnInst_0_n49}), .b ({new_AGEMA_signal_10958, new_AGEMA_signal_10957, MixColumnsIns_MixOneColumnInst_0_n48}), .c ({new_AGEMA_signal_11994, new_AGEMA_signal_11993, MixColumnsOutput[100]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U85 ( .a ({new_AGEMA_signal_10996, new_AGEMA_signal_10995, MixColumnsIns_MixOneColumnInst_0_n47}), .b ({new_AGEMA_signal_10298, new_AGEMA_signal_10297, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .c ({new_AGEMA_signal_11400, new_AGEMA_signal_11399, MixColumnsIns_MixOneColumnInst_0_n49}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U84 ( .a ({new_AGEMA_signal_11402, new_AGEMA_signal_11401, MixColumnsIns_MixOneColumnInst_0_n46}), .b ({new_AGEMA_signal_10960, new_AGEMA_signal_10959, MixColumnsIns_MixOneColumnInst_0_n45}), .c ({new_AGEMA_signal_11996, new_AGEMA_signal_11995, MixColumnsOutput[99]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U83 ( .a ({new_AGEMA_signal_11000, new_AGEMA_signal_10999, MixColumnsIns_MixOneColumnInst_0_n44}), .b ({new_AGEMA_signal_10300, new_AGEMA_signal_10299, MixColumnsInput[107]}), .c ({new_AGEMA_signal_11402, new_AGEMA_signal_11401, MixColumnsIns_MixOneColumnInst_0_n46}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U82 ( .a ({new_AGEMA_signal_10950, new_AGEMA_signal_10949, MixColumnsIns_MixOneColumnInst_0_n43}), .b ({new_AGEMA_signal_10522, new_AGEMA_signal_10521, MixColumnsIns_MixOneColumnInst_0_n57}), .c ({new_AGEMA_signal_11404, new_AGEMA_signal_11403, MixColumnsOutput[127]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U81 ( .a ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_10434, new_AGEMA_signal_10433, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .c ({new_AGEMA_signal_10522, new_AGEMA_signal_10521, MixColumnsIns_MixOneColumnInst_0_n57}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U80 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_10530, new_AGEMA_signal_10529, MixColumnsIns_MixOneColumnInst_0_n42}), .c ({new_AGEMA_signal_10950, new_AGEMA_signal_10949, MixColumnsIns_MixOneColumnInst_0_n43}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U79 ( .a ({new_AGEMA_signal_10952, new_AGEMA_signal_10951, MixColumnsIns_MixOneColumnInst_0_n41}), .b ({new_AGEMA_signal_10524, new_AGEMA_signal_10523, MixColumnsIns_MixOneColumnInst_0_n54}), .c ({new_AGEMA_signal_11406, new_AGEMA_signal_11405, MixColumnsOutput[126]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U78 ( .a ({new_AGEMA_signal_10364, new_AGEMA_signal_10363, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .b ({new_AGEMA_signal_10436, new_AGEMA_signal_10435, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .c ({new_AGEMA_signal_10524, new_AGEMA_signal_10523, MixColumnsIns_MixOneColumnInst_0_n54}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U77 ( .a ({new_AGEMA_signal_10224, new_AGEMA_signal_10223, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .b ({new_AGEMA_signal_10532, new_AGEMA_signal_10531, MixColumnsIns_MixOneColumnInst_0_n40}), .c ({new_AGEMA_signal_10952, new_AGEMA_signal_10951, MixColumnsIns_MixOneColumnInst_0_n41}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U76 ( .a ({new_AGEMA_signal_10954, new_AGEMA_signal_10953, MixColumnsIns_MixOneColumnInst_0_n39}), .b ({new_AGEMA_signal_10528, new_AGEMA_signal_10527, MixColumnsIns_MixOneColumnInst_0_n38}), .c ({new_AGEMA_signal_11408, new_AGEMA_signal_11407, MixColumnsOutput[98]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U75 ( .a ({new_AGEMA_signal_10556, new_AGEMA_signal_10555, MixColumnsIns_MixOneColumnInst_0_n37}), .b ({new_AGEMA_signal_10302, new_AGEMA_signal_10301, MixColumnsInput[106]}), .c ({new_AGEMA_signal_10954, new_AGEMA_signal_10953, MixColumnsIns_MixOneColumnInst_0_n39}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U74 ( .a ({new_AGEMA_signal_10956, new_AGEMA_signal_10955, MixColumnsIns_MixOneColumnInst_0_n36}), .b ({new_AGEMA_signal_10526, new_AGEMA_signal_10525, MixColumnsIns_MixOneColumnInst_0_n51}), .c ({new_AGEMA_signal_11410, new_AGEMA_signal_11409, MixColumnsOutput[125]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U73 ( .a ({new_AGEMA_signal_10366, new_AGEMA_signal_10365, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .b ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .c ({new_AGEMA_signal_10526, new_AGEMA_signal_10525, MixColumnsIns_MixOneColumnInst_0_n51}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U72 ( .a ({new_AGEMA_signal_10226, new_AGEMA_signal_10225, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .b ({new_AGEMA_signal_10534, new_AGEMA_signal_10533, MixColumnsIns_MixOneColumnInst_0_n35}), .c ({new_AGEMA_signal_10956, new_AGEMA_signal_10955, MixColumnsIns_MixOneColumnInst_0_n36}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U71 ( .a ({new_AGEMA_signal_11412, new_AGEMA_signal_11411, MixColumnsIns_MixOneColumnInst_0_n34}), .b ({new_AGEMA_signal_10958, new_AGEMA_signal_10957, MixColumnsIns_MixOneColumnInst_0_n48}), .c ({new_AGEMA_signal_11998, new_AGEMA_signal_11997, MixColumnsOutput[124]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U70 ( .a ({new_AGEMA_signal_10368, new_AGEMA_signal_10367, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .b ({new_AGEMA_signal_10562, new_AGEMA_signal_10561, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]}), .c ({new_AGEMA_signal_10958, new_AGEMA_signal_10957, MixColumnsIns_MixOneColumnInst_0_n48}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U69 ( .a ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .b ({new_AGEMA_signal_10972, new_AGEMA_signal_10971, MixColumnsIns_MixOneColumnInst_0_n33}), .c ({new_AGEMA_signal_11412, new_AGEMA_signal_11411, MixColumnsIns_MixOneColumnInst_0_n34}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U68 ( .a ({new_AGEMA_signal_11414, new_AGEMA_signal_11413, MixColumnsIns_MixOneColumnInst_0_n32}), .b ({new_AGEMA_signal_10960, new_AGEMA_signal_10959, MixColumnsIns_MixOneColumnInst_0_n45}), .c ({new_AGEMA_signal_12000, new_AGEMA_signal_11999, MixColumnsOutput[123]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U67 ( .a ({new_AGEMA_signal_10370, new_AGEMA_signal_10369, MixColumnsInput[115]}), .b ({new_AGEMA_signal_10564, new_AGEMA_signal_10563, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]}), .c ({new_AGEMA_signal_10960, new_AGEMA_signal_10959, MixColumnsIns_MixOneColumnInst_0_n45}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U66 ( .a ({new_AGEMA_signal_10230, new_AGEMA_signal_10229, MixColumnsInput[99]}), .b ({new_AGEMA_signal_10978, new_AGEMA_signal_10977, MixColumnsIns_MixOneColumnInst_0_n31}), .c ({new_AGEMA_signal_11414, new_AGEMA_signal_11413, MixColumnsIns_MixOneColumnInst_0_n32}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U65 ( .a ({new_AGEMA_signal_10962, new_AGEMA_signal_10961, MixColumnsIns_MixOneColumnInst_0_n30}), .b ({new_AGEMA_signal_10528, new_AGEMA_signal_10527, MixColumnsIns_MixOneColumnInst_0_n38}), .c ({new_AGEMA_signal_11416, new_AGEMA_signal_11415, MixColumnsOutput[122]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U64 ( .a ({new_AGEMA_signal_10372, new_AGEMA_signal_10371, MixColumnsInput[114]}), .b ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .c ({new_AGEMA_signal_10528, new_AGEMA_signal_10527, MixColumnsIns_MixOneColumnInst_0_n38}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U63 ( .a ({new_AGEMA_signal_10232, new_AGEMA_signal_10231, MixColumnsInput[98]}), .b ({new_AGEMA_signal_10536, new_AGEMA_signal_10535, MixColumnsIns_MixOneColumnInst_0_n29}), .c ({new_AGEMA_signal_10962, new_AGEMA_signal_10961, MixColumnsIns_MixOneColumnInst_0_n30}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U62 ( .a ({new_AGEMA_signal_11418, new_AGEMA_signal_11417, MixColumnsIns_MixOneColumnInst_0_n28}), .b ({new_AGEMA_signal_10974, new_AGEMA_signal_10973, MixColumnsIns_MixOneColumnInst_0_n27}), .c ({new_AGEMA_signal_12002, new_AGEMA_signal_12001, MixColumnsOutput[121]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U61 ( .a ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .b ({new_AGEMA_signal_10982, new_AGEMA_signal_10981, MixColumnsIns_MixOneColumnInst_0_n26}), .c ({new_AGEMA_signal_11418, new_AGEMA_signal_11417, MixColumnsIns_MixOneColumnInst_0_n28}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U60 ( .a ({new_AGEMA_signal_10964, new_AGEMA_signal_10963, MixColumnsIns_MixOneColumnInst_0_n25}), .b ({new_AGEMA_signal_10538, new_AGEMA_signal_10537, MixColumnsIns_MixOneColumnInst_0_n24}), .c ({new_AGEMA_signal_11420, new_AGEMA_signal_11419, MixColumnsOutput[120]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U59 ( .a ({new_AGEMA_signal_10558, new_AGEMA_signal_10557, MixColumnsIns_MixOneColumnInst_0_n23}), .b ({new_AGEMA_signal_9826, new_AGEMA_signal_9825, MixColumnsInput[96]}), .c ({new_AGEMA_signal_10964, new_AGEMA_signal_10963, MixColumnsIns_MixOneColumnInst_0_n25}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U58 ( .a ({new_AGEMA_signal_10966, new_AGEMA_signal_10965, MixColumnsIns_MixOneColumnInst_0_n22}), .b ({new_AGEMA_signal_10530, new_AGEMA_signal_10529, MixColumnsIns_MixOneColumnInst_0_n42}), .c ({new_AGEMA_signal_11422, new_AGEMA_signal_11421, MixColumnsOutput[119]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U57 ( .a ({new_AGEMA_signal_10292, new_AGEMA_signal_10291, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_10364, new_AGEMA_signal_10363, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .c ({new_AGEMA_signal_10530, new_AGEMA_signal_10529, MixColumnsIns_MixOneColumnInst_0_n42}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U56 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_10542, new_AGEMA_signal_10541, MixColumnsIns_MixOneColumnInst_0_n21}), .c ({new_AGEMA_signal_10966, new_AGEMA_signal_10965, MixColumnsIns_MixOneColumnInst_0_n22}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U55 ( .a ({new_AGEMA_signal_10968, new_AGEMA_signal_10967, MixColumnsIns_MixOneColumnInst_0_n20}), .b ({new_AGEMA_signal_10532, new_AGEMA_signal_10531, MixColumnsIns_MixOneColumnInst_0_n40}), .c ({new_AGEMA_signal_11424, new_AGEMA_signal_11423, MixColumnsOutput[118]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U54 ( .a ({new_AGEMA_signal_10294, new_AGEMA_signal_10293, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .b ({new_AGEMA_signal_10366, new_AGEMA_signal_10365, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .c ({new_AGEMA_signal_10532, new_AGEMA_signal_10531, MixColumnsIns_MixOneColumnInst_0_n40}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U53 ( .a ({new_AGEMA_signal_10434, new_AGEMA_signal_10433, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .b ({new_AGEMA_signal_10546, new_AGEMA_signal_10545, MixColumnsIns_MixOneColumnInst_0_n19}), .c ({new_AGEMA_signal_10968, new_AGEMA_signal_10967, MixColumnsIns_MixOneColumnInst_0_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U52 ( .a ({new_AGEMA_signal_10970, new_AGEMA_signal_10969, MixColumnsIns_MixOneColumnInst_0_n18}), .b ({new_AGEMA_signal_10534, new_AGEMA_signal_10533, MixColumnsIns_MixOneColumnInst_0_n35}), .c ({new_AGEMA_signal_11426, new_AGEMA_signal_11425, MixColumnsOutput[117]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U51 ( .a ({new_AGEMA_signal_10296, new_AGEMA_signal_10295, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .b ({new_AGEMA_signal_10368, new_AGEMA_signal_10367, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .c ({new_AGEMA_signal_10534, new_AGEMA_signal_10533, MixColumnsIns_MixOneColumnInst_0_n35}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U50 ( .a ({new_AGEMA_signal_10436, new_AGEMA_signal_10435, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .b ({new_AGEMA_signal_10550, new_AGEMA_signal_10549, MixColumnsIns_MixOneColumnInst_0_n17}), .c ({new_AGEMA_signal_10970, new_AGEMA_signal_10969, MixColumnsIns_MixOneColumnInst_0_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U49 ( .a ({new_AGEMA_signal_11428, new_AGEMA_signal_11427, MixColumnsIns_MixOneColumnInst_0_n16}), .b ({new_AGEMA_signal_10972, new_AGEMA_signal_10971, MixColumnsIns_MixOneColumnInst_0_n33}), .c ({new_AGEMA_signal_12004, new_AGEMA_signal_12003, MixColumnsOutput[116]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U48 ( .a ({new_AGEMA_signal_10298, new_AGEMA_signal_10297, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .b ({new_AGEMA_signal_10568, new_AGEMA_signal_10567, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]}), .c ({new_AGEMA_signal_10972, new_AGEMA_signal_10971, MixColumnsIns_MixOneColumnInst_0_n33}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U47 ( .a ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .b ({new_AGEMA_signal_10994, new_AGEMA_signal_10993, MixColumnsIns_MixOneColumnInst_0_n15}), .c ({new_AGEMA_signal_11428, new_AGEMA_signal_11427, MixColumnsIns_MixOneColumnInst_0_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U46 ( .a ({new_AGEMA_signal_11430, new_AGEMA_signal_11429, MixColumnsIns_MixOneColumnInst_0_n14}), .b ({new_AGEMA_signal_10974, new_AGEMA_signal_10973, MixColumnsIns_MixOneColumnInst_0_n27}), .c ({new_AGEMA_signal_12006, new_AGEMA_signal_12005, MixColumnsOutput[97]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U45 ( .a ({new_AGEMA_signal_10374, new_AGEMA_signal_10373, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .b ({new_AGEMA_signal_10566, new_AGEMA_signal_10565, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]}), .c ({new_AGEMA_signal_10974, new_AGEMA_signal_10973, MixColumnsIns_MixOneColumnInst_0_n27}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U44 ( .a ({new_AGEMA_signal_10304, new_AGEMA_signal_10303, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .b ({new_AGEMA_signal_10976, new_AGEMA_signal_10975, MixColumnsIns_MixOneColumnInst_0_n62}), .c ({new_AGEMA_signal_11430, new_AGEMA_signal_11429, MixColumnsIns_MixOneColumnInst_0_n14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U43 ( .a ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .b ({new_AGEMA_signal_10584, new_AGEMA_signal_10583, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]}), .c ({new_AGEMA_signal_10976, new_AGEMA_signal_10975, MixColumnsIns_MixOneColumnInst_0_n62}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U42 ( .a ({new_AGEMA_signal_11432, new_AGEMA_signal_11431, MixColumnsIns_MixOneColumnInst_0_n13}), .b ({new_AGEMA_signal_10978, new_AGEMA_signal_10977, MixColumnsIns_MixOneColumnInst_0_n31}), .c ({new_AGEMA_signal_12008, new_AGEMA_signal_12007, MixColumnsOutput[115]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U41 ( .a ({new_AGEMA_signal_10300, new_AGEMA_signal_10299, MixColumnsInput[107]}), .b ({new_AGEMA_signal_10570, new_AGEMA_signal_10569, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]}), .c ({new_AGEMA_signal_10978, new_AGEMA_signal_10977, MixColumnsIns_MixOneColumnInst_0_n31}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U40 ( .a ({new_AGEMA_signal_10440, new_AGEMA_signal_10439, MixColumnsInput[123]}), .b ({new_AGEMA_signal_10998, new_AGEMA_signal_10997, MixColumnsIns_MixOneColumnInst_0_n12}), .c ({new_AGEMA_signal_11432, new_AGEMA_signal_11431, MixColumnsIns_MixOneColumnInst_0_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U39 ( .a ({new_AGEMA_signal_10980, new_AGEMA_signal_10979, MixColumnsIns_MixOneColumnInst_0_n11}), .b ({new_AGEMA_signal_10536, new_AGEMA_signal_10535, MixColumnsIns_MixOneColumnInst_0_n29}), .c ({new_AGEMA_signal_11434, new_AGEMA_signal_11433, MixColumnsOutput[114]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U38 ( .a ({new_AGEMA_signal_10302, new_AGEMA_signal_10301, MixColumnsInput[106]}), .b ({new_AGEMA_signal_10374, new_AGEMA_signal_10373, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .c ({new_AGEMA_signal_10536, new_AGEMA_signal_10535, MixColumnsIns_MixOneColumnInst_0_n29}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U37 ( .a ({new_AGEMA_signal_10442, new_AGEMA_signal_10441, MixColumnsInput[122]}), .b ({new_AGEMA_signal_10554, new_AGEMA_signal_10553, MixColumnsIns_MixOneColumnInst_0_n10}), .c ({new_AGEMA_signal_10980, new_AGEMA_signal_10979, MixColumnsIns_MixOneColumnInst_0_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U36 ( .a ({new_AGEMA_signal_11436, new_AGEMA_signal_11435, MixColumnsIns_MixOneColumnInst_0_n9}), .b ({new_AGEMA_signal_10982, new_AGEMA_signal_10981, MixColumnsIns_MixOneColumnInst_0_n26}), .c ({new_AGEMA_signal_12010, new_AGEMA_signal_12009, MixColumnsOutput[113]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U35 ( .a ({new_AGEMA_signal_10572, new_AGEMA_signal_10571, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]}), .b ({new_AGEMA_signal_10304, new_AGEMA_signal_10303, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .c ({new_AGEMA_signal_10982, new_AGEMA_signal_10981, MixColumnsIns_MixOneColumnInst_0_n26}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U34 ( .a ({new_AGEMA_signal_10984, new_AGEMA_signal_10983, MixColumnsIns_MixOneColumnInst_0_n63}), .b ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .c ({new_AGEMA_signal_11436, new_AGEMA_signal_11435, MixColumnsIns_MixOneColumnInst_0_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U33 ( .a ({new_AGEMA_signal_10578, new_AGEMA_signal_10577, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]}), .b ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .c ({new_AGEMA_signal_10984, new_AGEMA_signal_10983, MixColumnsIns_MixOneColumnInst_0_n63}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U32 ( .a ({new_AGEMA_signal_10986, new_AGEMA_signal_10985, MixColumnsIns_MixOneColumnInst_0_n8}), .b ({new_AGEMA_signal_10538, new_AGEMA_signal_10537, MixColumnsIns_MixOneColumnInst_0_n24}), .c ({new_AGEMA_signal_11438, new_AGEMA_signal_11437, MixColumnsOutput[112]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U31 ( .a ({new_AGEMA_signal_9936, new_AGEMA_signal_9935, MixColumnsInput[104]}), .b ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .c ({new_AGEMA_signal_10538, new_AGEMA_signal_10537, MixColumnsIns_MixOneColumnInst_0_n24}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U30 ( .a ({new_AGEMA_signal_10156, new_AGEMA_signal_10155, MixColumnsInput[120]}), .b ({new_AGEMA_signal_10540, new_AGEMA_signal_10539, MixColumnsIns_MixOneColumnInst_0_n60}), .c ({new_AGEMA_signal_10986, new_AGEMA_signal_10985, MixColumnsIns_MixOneColumnInst_0_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U29 ( .a ({new_AGEMA_signal_10292, new_AGEMA_signal_10291, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_9826, new_AGEMA_signal_9825, MixColumnsInput[96]}), .c ({new_AGEMA_signal_10540, new_AGEMA_signal_10539, MixColumnsIns_MixOneColumnInst_0_n60}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U28 ( .a ({new_AGEMA_signal_10988, new_AGEMA_signal_10987, MixColumnsIns_MixOneColumnInst_0_n7}), .b ({new_AGEMA_signal_10542, new_AGEMA_signal_10541, MixColumnsIns_MixOneColumnInst_0_n21}), .c ({new_AGEMA_signal_11440, new_AGEMA_signal_11439, MixColumnsOutput[111]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U27 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_10294, new_AGEMA_signal_10293, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .c ({new_AGEMA_signal_10542, new_AGEMA_signal_10541, MixColumnsIns_MixOneColumnInst_0_n21}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U26 ( .a ({new_AGEMA_signal_10544, new_AGEMA_signal_10543, MixColumnsIns_MixOneColumnInst_0_n56}), .b ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .c ({new_AGEMA_signal_10988, new_AGEMA_signal_10987, MixColumnsIns_MixOneColumnInst_0_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U25 ( .a ({new_AGEMA_signal_10224, new_AGEMA_signal_10223, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .b ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .c ({new_AGEMA_signal_10544, new_AGEMA_signal_10543, MixColumnsIns_MixOneColumnInst_0_n56}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U24 ( .a ({new_AGEMA_signal_10990, new_AGEMA_signal_10989, MixColumnsIns_MixOneColumnInst_0_n6}), .b ({new_AGEMA_signal_10546, new_AGEMA_signal_10545, MixColumnsIns_MixOneColumnInst_0_n19}), .c ({new_AGEMA_signal_11442, new_AGEMA_signal_11441, MixColumnsOutput[110]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U23 ( .a ({new_AGEMA_signal_10224, new_AGEMA_signal_10223, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .b ({new_AGEMA_signal_10296, new_AGEMA_signal_10295, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .c ({new_AGEMA_signal_10546, new_AGEMA_signal_10545, MixColumnsIns_MixOneColumnInst_0_n19}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U22 ( .a ({new_AGEMA_signal_10548, new_AGEMA_signal_10547, MixColumnsIns_MixOneColumnInst_0_n53}), .b ({new_AGEMA_signal_10364, new_AGEMA_signal_10363, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .c ({new_AGEMA_signal_10990, new_AGEMA_signal_10989, MixColumnsIns_MixOneColumnInst_0_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U21 ( .a ({new_AGEMA_signal_10226, new_AGEMA_signal_10225, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .b ({new_AGEMA_signal_10434, new_AGEMA_signal_10433, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .c ({new_AGEMA_signal_10548, new_AGEMA_signal_10547, MixColumnsIns_MixOneColumnInst_0_n53}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U20 ( .a ({new_AGEMA_signal_10992, new_AGEMA_signal_10991, MixColumnsIns_MixOneColumnInst_0_n5}), .b ({new_AGEMA_signal_10550, new_AGEMA_signal_10549, MixColumnsIns_MixOneColumnInst_0_n17}), .c ({new_AGEMA_signal_11444, new_AGEMA_signal_11443, MixColumnsOutput[109]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U19 ( .a ({new_AGEMA_signal_10226, new_AGEMA_signal_10225, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .b ({new_AGEMA_signal_10298, new_AGEMA_signal_10297, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .c ({new_AGEMA_signal_10550, new_AGEMA_signal_10549, MixColumnsIns_MixOneColumnInst_0_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U18 ( .a ({new_AGEMA_signal_10552, new_AGEMA_signal_10551, MixColumnsIns_MixOneColumnInst_0_n50}), .b ({new_AGEMA_signal_10366, new_AGEMA_signal_10365, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .c ({new_AGEMA_signal_10992, new_AGEMA_signal_10991, MixColumnsIns_MixOneColumnInst_0_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U17 ( .a ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .b ({new_AGEMA_signal_10436, new_AGEMA_signal_10435, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .c ({new_AGEMA_signal_10552, new_AGEMA_signal_10551, MixColumnsIns_MixOneColumnInst_0_n50}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U16 ( .a ({new_AGEMA_signal_11446, new_AGEMA_signal_11445, MixColumnsIns_MixOneColumnInst_0_n4}), .b ({new_AGEMA_signal_10994, new_AGEMA_signal_10993, MixColumnsIns_MixOneColumnInst_0_n15}), .c ({new_AGEMA_signal_12012, new_AGEMA_signal_12011, MixColumnsOutput[108]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U15 ( .a ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .b ({new_AGEMA_signal_10574, new_AGEMA_signal_10573, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]}), .c ({new_AGEMA_signal_10994, new_AGEMA_signal_10993, MixColumnsIns_MixOneColumnInst_0_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U14 ( .a ({new_AGEMA_signal_10996, new_AGEMA_signal_10995, MixColumnsIns_MixOneColumnInst_0_n47}), .b ({new_AGEMA_signal_10368, new_AGEMA_signal_10367, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .c ({new_AGEMA_signal_11446, new_AGEMA_signal_11445, MixColumnsIns_MixOneColumnInst_0_n4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U13 ( .a ({new_AGEMA_signal_10580, new_AGEMA_signal_10579, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]}), .b ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .c ({new_AGEMA_signal_10996, new_AGEMA_signal_10995, MixColumnsIns_MixOneColumnInst_0_n47}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U12 ( .a ({new_AGEMA_signal_11448, new_AGEMA_signal_11447, MixColumnsIns_MixOneColumnInst_0_n3}), .b ({new_AGEMA_signal_10998, new_AGEMA_signal_10997, MixColumnsIns_MixOneColumnInst_0_n12}), .c ({new_AGEMA_signal_12014, new_AGEMA_signal_12013, MixColumnsOutput[107]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U11 ( .a ({new_AGEMA_signal_10230, new_AGEMA_signal_10229, MixColumnsInput[99]}), .b ({new_AGEMA_signal_10576, new_AGEMA_signal_10575, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]}), .c ({new_AGEMA_signal_10998, new_AGEMA_signal_10997, MixColumnsIns_MixOneColumnInst_0_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U10 ( .a ({new_AGEMA_signal_11000, new_AGEMA_signal_10999, MixColumnsIns_MixOneColumnInst_0_n44}), .b ({new_AGEMA_signal_10370, new_AGEMA_signal_10369, MixColumnsInput[115]}), .c ({new_AGEMA_signal_11448, new_AGEMA_signal_11447, MixColumnsIns_MixOneColumnInst_0_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U9 ( .a ({new_AGEMA_signal_10582, new_AGEMA_signal_10581, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]}), .b ({new_AGEMA_signal_10440, new_AGEMA_signal_10439, MixColumnsInput[123]}), .c ({new_AGEMA_signal_11000, new_AGEMA_signal_10999, MixColumnsIns_MixOneColumnInst_0_n44}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U8 ( .a ({new_AGEMA_signal_11002, new_AGEMA_signal_11001, MixColumnsIns_MixOneColumnInst_0_n2}), .b ({new_AGEMA_signal_10554, new_AGEMA_signal_10553, MixColumnsIns_MixOneColumnInst_0_n10}), .c ({new_AGEMA_signal_11450, new_AGEMA_signal_11449, MixColumnsOutput[106]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U7 ( .a ({new_AGEMA_signal_10232, new_AGEMA_signal_10231, MixColumnsInput[98]}), .b ({new_AGEMA_signal_10304, new_AGEMA_signal_10303, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .c ({new_AGEMA_signal_10554, new_AGEMA_signal_10553, MixColumnsIns_MixOneColumnInst_0_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U6 ( .a ({new_AGEMA_signal_10556, new_AGEMA_signal_10555, MixColumnsIns_MixOneColumnInst_0_n37}), .b ({new_AGEMA_signal_10372, new_AGEMA_signal_10371, MixColumnsInput[114]}), .c ({new_AGEMA_signal_11002, new_AGEMA_signal_11001, MixColumnsIns_MixOneColumnInst_0_n2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U5 ( .a ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .b ({new_AGEMA_signal_10442, new_AGEMA_signal_10441, MixColumnsInput[122]}), .c ({new_AGEMA_signal_10556, new_AGEMA_signal_10555, MixColumnsIns_MixOneColumnInst_0_n37}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U4 ( .a ({new_AGEMA_signal_11004, new_AGEMA_signal_11003, MixColumnsIns_MixOneColumnInst_0_n1}), .b ({new_AGEMA_signal_9936, new_AGEMA_signal_9935, MixColumnsInput[104]}), .c ({new_AGEMA_signal_11452, new_AGEMA_signal_11451, MixColumnsOutput[96]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U3 ( .a ({new_AGEMA_signal_10560, new_AGEMA_signal_10559, MixColumnsIns_MixOneColumnInst_0_n59}), .b ({new_AGEMA_signal_10558, new_AGEMA_signal_10557, MixColumnsIns_MixOneColumnInst_0_n23}), .c ({new_AGEMA_signal_11004, new_AGEMA_signal_11003, MixColumnsIns_MixOneColumnInst_0_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U2 ( .a ({new_AGEMA_signal_10046, new_AGEMA_signal_10045, MixColumnsInput[112]}), .b ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .c ({new_AGEMA_signal_10558, new_AGEMA_signal_10557, MixColumnsIns_MixOneColumnInst_0_n23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U1 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_10156, new_AGEMA_signal_10155, MixColumnsInput[120]}), .c ({new_AGEMA_signal_10560, new_AGEMA_signal_10559, MixColumnsIns_MixOneColumnInst_0_n59}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_10440, new_AGEMA_signal_10439, MixColumnsInput[123]}), .c ({new_AGEMA_signal_10562, new_AGEMA_signal_10561, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_10442, new_AGEMA_signal_10441, MixColumnsInput[122]}), .c ({new_AGEMA_signal_10564, new_AGEMA_signal_10563, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_10156, new_AGEMA_signal_10155, MixColumnsInput[120]}), .c ({new_AGEMA_signal_10566, new_AGEMA_signal_10565, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_10370, new_AGEMA_signal_10369, MixColumnsInput[115]}), .c ({new_AGEMA_signal_10568, new_AGEMA_signal_10567, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_10372, new_AGEMA_signal_10371, MixColumnsInput[114]}), .c ({new_AGEMA_signal_10570, new_AGEMA_signal_10569, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_10046, new_AGEMA_signal_10045, MixColumnsInput[112]}), .c ({new_AGEMA_signal_10572, new_AGEMA_signal_10571, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_10292, new_AGEMA_signal_10291, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_10300, new_AGEMA_signal_10299, MixColumnsInput[107]}), .c ({new_AGEMA_signal_10574, new_AGEMA_signal_10573, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_10292, new_AGEMA_signal_10291, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_10302, new_AGEMA_signal_10301, MixColumnsInput[106]}), .c ({new_AGEMA_signal_10576, new_AGEMA_signal_10575, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_10292, new_AGEMA_signal_10291, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_9936, new_AGEMA_signal_9935, MixColumnsInput[104]}), .c ({new_AGEMA_signal_10578, new_AGEMA_signal_10577, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_10230, new_AGEMA_signal_10229, MixColumnsInput[99]}), .c ({new_AGEMA_signal_10580, new_AGEMA_signal_10579, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_10232, new_AGEMA_signal_10231, MixColumnsInput[98]}), .c ({new_AGEMA_signal_10582, new_AGEMA_signal_10581, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_9826, new_AGEMA_signal_9825, MixColumnsInput[96]}), .c ({new_AGEMA_signal_10584, new_AGEMA_signal_10583, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U96 ( .a ({new_AGEMA_signal_11454, new_AGEMA_signal_11453, MixColumnsIns_MixOneColumnInst_1_n64}), .b ({new_AGEMA_signal_10318, new_AGEMA_signal_10317, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .c ({new_AGEMA_signal_12016, new_AGEMA_signal_12015, MixColumnsOutput[73]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U95 ( .a ({new_AGEMA_signal_11048, new_AGEMA_signal_11047, MixColumnsIns_MixOneColumnInst_1_n63}), .b ({new_AGEMA_signal_11040, new_AGEMA_signal_11039, MixColumnsIns_MixOneColumnInst_1_n62}), .c ({new_AGEMA_signal_11454, new_AGEMA_signal_11453, MixColumnsIns_MixOneColumnInst_1_n64}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U94 ( .a ({new_AGEMA_signal_11006, new_AGEMA_signal_11005, MixColumnsIns_MixOneColumnInst_1_n61}), .b ({new_AGEMA_signal_10604, new_AGEMA_signal_10603, MixColumnsIns_MixOneColumnInst_1_n60}), .c ({new_AGEMA_signal_11456, new_AGEMA_signal_11455, MixColumnsOutput[72]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U93 ( .a ({new_AGEMA_signal_10624, new_AGEMA_signal_10623, MixColumnsIns_MixOneColumnInst_1_n59}), .b ({new_AGEMA_signal_9958, new_AGEMA_signal_9957, MixColumnsInput[80]}), .c ({new_AGEMA_signal_11006, new_AGEMA_signal_11005, MixColumnsIns_MixOneColumnInst_1_n61}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U92 ( .a ({new_AGEMA_signal_11008, new_AGEMA_signal_11007, MixColumnsIns_MixOneColumnInst_1_n58}), .b ({new_AGEMA_signal_10586, new_AGEMA_signal_10585, MixColumnsIns_MixOneColumnInst_1_n57}), .c ({new_AGEMA_signal_11458, new_AGEMA_signal_11457, MixColumnsOutput[71]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U91 ( .a ({new_AGEMA_signal_10608, new_AGEMA_signal_10607, MixColumnsIns_MixOneColumnInst_1_n56}), .b ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .c ({new_AGEMA_signal_11008, new_AGEMA_signal_11007, MixColumnsIns_MixOneColumnInst_1_n58}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U90 ( .a ({new_AGEMA_signal_11010, new_AGEMA_signal_11009, MixColumnsIns_MixOneColumnInst_1_n55}), .b ({new_AGEMA_signal_10588, new_AGEMA_signal_10587, MixColumnsIns_MixOneColumnInst_1_n54}), .c ({new_AGEMA_signal_11460, new_AGEMA_signal_11459, MixColumnsOutput[70]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U89 ( .a ({new_AGEMA_signal_10612, new_AGEMA_signal_10611, MixColumnsIns_MixOneColumnInst_1_n53}), .b ({new_AGEMA_signal_10238, new_AGEMA_signal_10237, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .c ({new_AGEMA_signal_11010, new_AGEMA_signal_11009, MixColumnsIns_MixOneColumnInst_1_n55}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U88 ( .a ({new_AGEMA_signal_11012, new_AGEMA_signal_11011, MixColumnsIns_MixOneColumnInst_1_n52}), .b ({new_AGEMA_signal_10590, new_AGEMA_signal_10589, MixColumnsIns_MixOneColumnInst_1_n51}), .c ({new_AGEMA_signal_11462, new_AGEMA_signal_11461, MixColumnsOutput[69]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U87 ( .a ({new_AGEMA_signal_10616, new_AGEMA_signal_10615, MixColumnsIns_MixOneColumnInst_1_n50}), .b ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .c ({new_AGEMA_signal_11012, new_AGEMA_signal_11011, MixColumnsIns_MixOneColumnInst_1_n52}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U86 ( .a ({new_AGEMA_signal_11464, new_AGEMA_signal_11463, MixColumnsIns_MixOneColumnInst_1_n49}), .b ({new_AGEMA_signal_11022, new_AGEMA_signal_11021, MixColumnsIns_MixOneColumnInst_1_n48}), .c ({new_AGEMA_signal_12018, new_AGEMA_signal_12017, MixColumnsOutput[68]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U85 ( .a ({new_AGEMA_signal_11060, new_AGEMA_signal_11059, MixColumnsIns_MixOneColumnInst_1_n47}), .b ({new_AGEMA_signal_10242, new_AGEMA_signal_10241, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .c ({new_AGEMA_signal_11464, new_AGEMA_signal_11463, MixColumnsIns_MixOneColumnInst_1_n49}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U84 ( .a ({new_AGEMA_signal_11466, new_AGEMA_signal_11465, MixColumnsIns_MixOneColumnInst_1_n46}), .b ({new_AGEMA_signal_11024, new_AGEMA_signal_11023, MixColumnsIns_MixOneColumnInst_1_n45}), .c ({new_AGEMA_signal_12020, new_AGEMA_signal_12019, MixColumnsOutput[67]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U83 ( .a ({new_AGEMA_signal_11064, new_AGEMA_signal_11063, MixColumnsIns_MixOneColumnInst_1_n44}), .b ({new_AGEMA_signal_10244, new_AGEMA_signal_10243, MixColumnsInput[75]}), .c ({new_AGEMA_signal_11466, new_AGEMA_signal_11465, MixColumnsIns_MixOneColumnInst_1_n46}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U82 ( .a ({new_AGEMA_signal_11014, new_AGEMA_signal_11013, MixColumnsIns_MixOneColumnInst_1_n43}), .b ({new_AGEMA_signal_10586, new_AGEMA_signal_10585, MixColumnsIns_MixOneColumnInst_1_n57}), .c ({new_AGEMA_signal_11468, new_AGEMA_signal_11467, MixColumnsOutput[95]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U81 ( .a ({new_AGEMA_signal_10306, new_AGEMA_signal_10305, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_10378, new_AGEMA_signal_10377, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .c ({new_AGEMA_signal_10586, new_AGEMA_signal_10585, MixColumnsIns_MixOneColumnInst_1_n57}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U80 ( .a ({new_AGEMA_signal_10390, new_AGEMA_signal_10389, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_10594, new_AGEMA_signal_10593, MixColumnsIns_MixOneColumnInst_1_n42}), .c ({new_AGEMA_signal_11014, new_AGEMA_signal_11013, MixColumnsIns_MixOneColumnInst_1_n43}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U79 ( .a ({new_AGEMA_signal_11016, new_AGEMA_signal_11015, MixColumnsIns_MixOneColumnInst_1_n41}), .b ({new_AGEMA_signal_10588, new_AGEMA_signal_10587, MixColumnsIns_MixOneColumnInst_1_n54}), .c ({new_AGEMA_signal_11470, new_AGEMA_signal_11469, MixColumnsOutput[94]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U78 ( .a ({new_AGEMA_signal_10308, new_AGEMA_signal_10307, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .b ({new_AGEMA_signal_10380, new_AGEMA_signal_10379, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .c ({new_AGEMA_signal_10588, new_AGEMA_signal_10587, MixColumnsIns_MixOneColumnInst_1_n54}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U77 ( .a ({new_AGEMA_signal_10392, new_AGEMA_signal_10391, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .b ({new_AGEMA_signal_10596, new_AGEMA_signal_10595, MixColumnsIns_MixOneColumnInst_1_n40}), .c ({new_AGEMA_signal_11016, new_AGEMA_signal_11015, MixColumnsIns_MixOneColumnInst_1_n41}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U76 ( .a ({new_AGEMA_signal_11018, new_AGEMA_signal_11017, MixColumnsIns_MixOneColumnInst_1_n39}), .b ({new_AGEMA_signal_10592, new_AGEMA_signal_10591, MixColumnsIns_MixOneColumnInst_1_n38}), .c ({new_AGEMA_signal_11472, new_AGEMA_signal_11471, MixColumnsOutput[66]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U75 ( .a ({new_AGEMA_signal_10620, new_AGEMA_signal_10619, MixColumnsIns_MixOneColumnInst_1_n37}), .b ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, MixColumnsInput[74]}), .c ({new_AGEMA_signal_11018, new_AGEMA_signal_11017, MixColumnsIns_MixOneColumnInst_1_n39}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U74 ( .a ({new_AGEMA_signal_11020, new_AGEMA_signal_11019, MixColumnsIns_MixOneColumnInst_1_n36}), .b ({new_AGEMA_signal_10590, new_AGEMA_signal_10589, MixColumnsIns_MixOneColumnInst_1_n51}), .c ({new_AGEMA_signal_11474, new_AGEMA_signal_11473, MixColumnsOutput[93]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U73 ( .a ({new_AGEMA_signal_10310, new_AGEMA_signal_10309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .b ({new_AGEMA_signal_10382, new_AGEMA_signal_10381, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .c ({new_AGEMA_signal_10590, new_AGEMA_signal_10589, MixColumnsIns_MixOneColumnInst_1_n51}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U72 ( .a ({new_AGEMA_signal_10394, new_AGEMA_signal_10393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .b ({new_AGEMA_signal_10598, new_AGEMA_signal_10597, MixColumnsIns_MixOneColumnInst_1_n35}), .c ({new_AGEMA_signal_11020, new_AGEMA_signal_11019, MixColumnsIns_MixOneColumnInst_1_n36}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U71 ( .a ({new_AGEMA_signal_11476, new_AGEMA_signal_11475, MixColumnsIns_MixOneColumnInst_1_n34}), .b ({new_AGEMA_signal_11022, new_AGEMA_signal_11021, MixColumnsIns_MixOneColumnInst_1_n48}), .c ({new_AGEMA_signal_12022, new_AGEMA_signal_12021, MixColumnsOutput[92]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U70 ( .a ({new_AGEMA_signal_10312, new_AGEMA_signal_10311, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .b ({new_AGEMA_signal_10626, new_AGEMA_signal_10625, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]}), .c ({new_AGEMA_signal_11022, new_AGEMA_signal_11021, MixColumnsIns_MixOneColumnInst_1_n48}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U69 ( .a ({new_AGEMA_signal_10396, new_AGEMA_signal_10395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .b ({new_AGEMA_signal_11036, new_AGEMA_signal_11035, MixColumnsIns_MixOneColumnInst_1_n33}), .c ({new_AGEMA_signal_11476, new_AGEMA_signal_11475, MixColumnsIns_MixOneColumnInst_1_n34}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U68 ( .a ({new_AGEMA_signal_11478, new_AGEMA_signal_11477, MixColumnsIns_MixOneColumnInst_1_n32}), .b ({new_AGEMA_signal_11024, new_AGEMA_signal_11023, MixColumnsIns_MixOneColumnInst_1_n45}), .c ({new_AGEMA_signal_12024, new_AGEMA_signal_12023, MixColumnsOutput[91]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U67 ( .a ({new_AGEMA_signal_10314, new_AGEMA_signal_10313, MixColumnsInput[83]}), .b ({new_AGEMA_signal_10628, new_AGEMA_signal_10627, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]}), .c ({new_AGEMA_signal_11024, new_AGEMA_signal_11023, MixColumnsIns_MixOneColumnInst_1_n45}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U66 ( .a ({new_AGEMA_signal_10398, new_AGEMA_signal_10397, MixColumnsInput[67]}), .b ({new_AGEMA_signal_11042, new_AGEMA_signal_11041, MixColumnsIns_MixOneColumnInst_1_n31}), .c ({new_AGEMA_signal_11478, new_AGEMA_signal_11477, MixColumnsIns_MixOneColumnInst_1_n32}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U65 ( .a ({new_AGEMA_signal_11026, new_AGEMA_signal_11025, MixColumnsIns_MixOneColumnInst_1_n30}), .b ({new_AGEMA_signal_10592, new_AGEMA_signal_10591, MixColumnsIns_MixOneColumnInst_1_n38}), .c ({new_AGEMA_signal_11480, new_AGEMA_signal_11479, MixColumnsOutput[90]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U64 ( .a ({new_AGEMA_signal_10316, new_AGEMA_signal_10315, MixColumnsInput[82]}), .b ({new_AGEMA_signal_10388, new_AGEMA_signal_10387, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .c ({new_AGEMA_signal_10592, new_AGEMA_signal_10591, MixColumnsIns_MixOneColumnInst_1_n38}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U63 ( .a ({new_AGEMA_signal_10400, new_AGEMA_signal_10399, MixColumnsInput[66]}), .b ({new_AGEMA_signal_10600, new_AGEMA_signal_10599, MixColumnsIns_MixOneColumnInst_1_n29}), .c ({new_AGEMA_signal_11026, new_AGEMA_signal_11025, MixColumnsIns_MixOneColumnInst_1_n30}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U62 ( .a ({new_AGEMA_signal_11482, new_AGEMA_signal_11481, MixColumnsIns_MixOneColumnInst_1_n28}), .b ({new_AGEMA_signal_11038, new_AGEMA_signal_11037, MixColumnsIns_MixOneColumnInst_1_n27}), .c ({new_AGEMA_signal_12026, new_AGEMA_signal_12025, MixColumnsOutput[89]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U61 ( .a ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .b ({new_AGEMA_signal_11046, new_AGEMA_signal_11045, MixColumnsIns_MixOneColumnInst_1_n26}), .c ({new_AGEMA_signal_11482, new_AGEMA_signal_11481, MixColumnsIns_MixOneColumnInst_1_n28}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U60 ( .a ({new_AGEMA_signal_11028, new_AGEMA_signal_11027, MixColumnsIns_MixOneColumnInst_1_n25}), .b ({new_AGEMA_signal_10602, new_AGEMA_signal_10601, MixColumnsIns_MixOneColumnInst_1_n24}), .c ({new_AGEMA_signal_11484, new_AGEMA_signal_11483, MixColumnsOutput[88]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U59 ( .a ({new_AGEMA_signal_10622, new_AGEMA_signal_10621, MixColumnsIns_MixOneColumnInst_1_n23}), .b ({new_AGEMA_signal_10090, new_AGEMA_signal_10089, MixColumnsInput[64]}), .c ({new_AGEMA_signal_11028, new_AGEMA_signal_11027, MixColumnsIns_MixOneColumnInst_1_n25}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U58 ( .a ({new_AGEMA_signal_11030, new_AGEMA_signal_11029, MixColumnsIns_MixOneColumnInst_1_n22}), .b ({new_AGEMA_signal_10594, new_AGEMA_signal_10593, MixColumnsIns_MixOneColumnInst_1_n42}), .c ({new_AGEMA_signal_11486, new_AGEMA_signal_11485, MixColumnsOutput[87]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U57 ( .a ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_10308, new_AGEMA_signal_10307, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .c ({new_AGEMA_signal_10594, new_AGEMA_signal_10593, MixColumnsIns_MixOneColumnInst_1_n42}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U56 ( .a ({new_AGEMA_signal_10376, new_AGEMA_signal_10375, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_10606, new_AGEMA_signal_10605, MixColumnsIns_MixOneColumnInst_1_n21}), .c ({new_AGEMA_signal_11030, new_AGEMA_signal_11029, MixColumnsIns_MixOneColumnInst_1_n22}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U55 ( .a ({new_AGEMA_signal_11032, new_AGEMA_signal_11031, MixColumnsIns_MixOneColumnInst_1_n20}), .b ({new_AGEMA_signal_10596, new_AGEMA_signal_10595, MixColumnsIns_MixOneColumnInst_1_n40}), .c ({new_AGEMA_signal_11488, new_AGEMA_signal_11487, MixColumnsOutput[86]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U54 ( .a ({new_AGEMA_signal_10238, new_AGEMA_signal_10237, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .b ({new_AGEMA_signal_10310, new_AGEMA_signal_10309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .c ({new_AGEMA_signal_10596, new_AGEMA_signal_10595, MixColumnsIns_MixOneColumnInst_1_n40}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U53 ( .a ({new_AGEMA_signal_10378, new_AGEMA_signal_10377, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .b ({new_AGEMA_signal_10610, new_AGEMA_signal_10609, MixColumnsIns_MixOneColumnInst_1_n19}), .c ({new_AGEMA_signal_11032, new_AGEMA_signal_11031, MixColumnsIns_MixOneColumnInst_1_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U52 ( .a ({new_AGEMA_signal_11034, new_AGEMA_signal_11033, MixColumnsIns_MixOneColumnInst_1_n18}), .b ({new_AGEMA_signal_10598, new_AGEMA_signal_10597, MixColumnsIns_MixOneColumnInst_1_n35}), .c ({new_AGEMA_signal_11490, new_AGEMA_signal_11489, MixColumnsOutput[85]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U51 ( .a ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .b ({new_AGEMA_signal_10312, new_AGEMA_signal_10311, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .c ({new_AGEMA_signal_10598, new_AGEMA_signal_10597, MixColumnsIns_MixOneColumnInst_1_n35}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U50 ( .a ({new_AGEMA_signal_10380, new_AGEMA_signal_10379, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .b ({new_AGEMA_signal_10614, new_AGEMA_signal_10613, MixColumnsIns_MixOneColumnInst_1_n17}), .c ({new_AGEMA_signal_11034, new_AGEMA_signal_11033, MixColumnsIns_MixOneColumnInst_1_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U49 ( .a ({new_AGEMA_signal_11492, new_AGEMA_signal_11491, MixColumnsIns_MixOneColumnInst_1_n16}), .b ({new_AGEMA_signal_11036, new_AGEMA_signal_11035, MixColumnsIns_MixOneColumnInst_1_n33}), .c ({new_AGEMA_signal_12028, new_AGEMA_signal_12027, MixColumnsOutput[84]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U48 ( .a ({new_AGEMA_signal_10242, new_AGEMA_signal_10241, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .b ({new_AGEMA_signal_10632, new_AGEMA_signal_10631, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]}), .c ({new_AGEMA_signal_11036, new_AGEMA_signal_11035, MixColumnsIns_MixOneColumnInst_1_n33}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U47 ( .a ({new_AGEMA_signal_10382, new_AGEMA_signal_10381, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .b ({new_AGEMA_signal_11058, new_AGEMA_signal_11057, MixColumnsIns_MixOneColumnInst_1_n15}), .c ({new_AGEMA_signal_11492, new_AGEMA_signal_11491, MixColumnsIns_MixOneColumnInst_1_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U46 ( .a ({new_AGEMA_signal_11494, new_AGEMA_signal_11493, MixColumnsIns_MixOneColumnInst_1_n14}), .b ({new_AGEMA_signal_11038, new_AGEMA_signal_11037, MixColumnsIns_MixOneColumnInst_1_n27}), .c ({new_AGEMA_signal_12030, new_AGEMA_signal_12029, MixColumnsOutput[65]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U45 ( .a ({new_AGEMA_signal_10318, new_AGEMA_signal_10317, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .b ({new_AGEMA_signal_10630, new_AGEMA_signal_10629, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]}), .c ({new_AGEMA_signal_11038, new_AGEMA_signal_11037, MixColumnsIns_MixOneColumnInst_1_n27}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U44 ( .a ({new_AGEMA_signal_10248, new_AGEMA_signal_10247, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .b ({new_AGEMA_signal_11040, new_AGEMA_signal_11039, MixColumnsIns_MixOneColumnInst_1_n62}), .c ({new_AGEMA_signal_11494, new_AGEMA_signal_11493, MixColumnsIns_MixOneColumnInst_1_n14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U43 ( .a ({new_AGEMA_signal_10388, new_AGEMA_signal_10387, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .b ({new_AGEMA_signal_10648, new_AGEMA_signal_10647, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]}), .c ({new_AGEMA_signal_11040, new_AGEMA_signal_11039, MixColumnsIns_MixOneColumnInst_1_n62}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U42 ( .a ({new_AGEMA_signal_11496, new_AGEMA_signal_11495, MixColumnsIns_MixOneColumnInst_1_n13}), .b ({new_AGEMA_signal_11042, new_AGEMA_signal_11041, MixColumnsIns_MixOneColumnInst_1_n31}), .c ({new_AGEMA_signal_12032, new_AGEMA_signal_12031, MixColumnsOutput[83]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U41 ( .a ({new_AGEMA_signal_10244, new_AGEMA_signal_10243, MixColumnsInput[75]}), .b ({new_AGEMA_signal_10634, new_AGEMA_signal_10633, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]}), .c ({new_AGEMA_signal_11042, new_AGEMA_signal_11041, MixColumnsIns_MixOneColumnInst_1_n31}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U40 ( .a ({new_AGEMA_signal_10384, new_AGEMA_signal_10383, MixColumnsInput[91]}), .b ({new_AGEMA_signal_11062, new_AGEMA_signal_11061, MixColumnsIns_MixOneColumnInst_1_n12}), .c ({new_AGEMA_signal_11496, new_AGEMA_signal_11495, MixColumnsIns_MixOneColumnInst_1_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U39 ( .a ({new_AGEMA_signal_11044, new_AGEMA_signal_11043, MixColumnsIns_MixOneColumnInst_1_n11}), .b ({new_AGEMA_signal_10600, new_AGEMA_signal_10599, MixColumnsIns_MixOneColumnInst_1_n29}), .c ({new_AGEMA_signal_11498, new_AGEMA_signal_11497, MixColumnsOutput[82]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U38 ( .a ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, MixColumnsInput[74]}), .b ({new_AGEMA_signal_10318, new_AGEMA_signal_10317, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .c ({new_AGEMA_signal_10600, new_AGEMA_signal_10599, MixColumnsIns_MixOneColumnInst_1_n29}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U37 ( .a ({new_AGEMA_signal_10386, new_AGEMA_signal_10385, MixColumnsInput[90]}), .b ({new_AGEMA_signal_10618, new_AGEMA_signal_10617, MixColumnsIns_MixOneColumnInst_1_n10}), .c ({new_AGEMA_signal_11044, new_AGEMA_signal_11043, MixColumnsIns_MixOneColumnInst_1_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U36 ( .a ({new_AGEMA_signal_11500, new_AGEMA_signal_11499, MixColumnsIns_MixOneColumnInst_1_n9}), .b ({new_AGEMA_signal_11046, new_AGEMA_signal_11045, MixColumnsIns_MixOneColumnInst_1_n26}), .c ({new_AGEMA_signal_12034, new_AGEMA_signal_12033, MixColumnsOutput[81]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U35 ( .a ({new_AGEMA_signal_10636, new_AGEMA_signal_10635, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]}), .b ({new_AGEMA_signal_10248, new_AGEMA_signal_10247, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .c ({new_AGEMA_signal_11046, new_AGEMA_signal_11045, MixColumnsIns_MixOneColumnInst_1_n26}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U34 ( .a ({new_AGEMA_signal_11048, new_AGEMA_signal_11047, MixColumnsIns_MixOneColumnInst_1_n63}), .b ({new_AGEMA_signal_10388, new_AGEMA_signal_10387, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .c ({new_AGEMA_signal_11500, new_AGEMA_signal_11499, MixColumnsIns_MixOneColumnInst_1_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U33 ( .a ({new_AGEMA_signal_10642, new_AGEMA_signal_10641, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]}), .b ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .c ({new_AGEMA_signal_11048, new_AGEMA_signal_11047, MixColumnsIns_MixOneColumnInst_1_n63}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U32 ( .a ({new_AGEMA_signal_11050, new_AGEMA_signal_11049, MixColumnsIns_MixOneColumnInst_1_n8}), .b ({new_AGEMA_signal_10602, new_AGEMA_signal_10601, MixColumnsIns_MixOneColumnInst_1_n24}), .c ({new_AGEMA_signal_11502, new_AGEMA_signal_11501, MixColumnsOutput[80]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U31 ( .a ({new_AGEMA_signal_9848, new_AGEMA_signal_9847, MixColumnsInput[72]}), .b ({new_AGEMA_signal_10306, new_AGEMA_signal_10305, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .c ({new_AGEMA_signal_10602, new_AGEMA_signal_10601, MixColumnsIns_MixOneColumnInst_1_n24}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U30 ( .a ({new_AGEMA_signal_10068, new_AGEMA_signal_10067, MixColumnsInput[88]}), .b ({new_AGEMA_signal_10604, new_AGEMA_signal_10603, MixColumnsIns_MixOneColumnInst_1_n60}), .c ({new_AGEMA_signal_11050, new_AGEMA_signal_11049, MixColumnsIns_MixOneColumnInst_1_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U29 ( .a ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_10090, new_AGEMA_signal_10089, MixColumnsInput[64]}), .c ({new_AGEMA_signal_10604, new_AGEMA_signal_10603, MixColumnsIns_MixOneColumnInst_1_n60}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U28 ( .a ({new_AGEMA_signal_11052, new_AGEMA_signal_11051, MixColumnsIns_MixOneColumnInst_1_n7}), .b ({new_AGEMA_signal_10606, new_AGEMA_signal_10605, MixColumnsIns_MixOneColumnInst_1_n21}), .c ({new_AGEMA_signal_11504, new_AGEMA_signal_11503, MixColumnsOutput[79]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U27 ( .a ({new_AGEMA_signal_10390, new_AGEMA_signal_10389, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_10238, new_AGEMA_signal_10237, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .c ({new_AGEMA_signal_10606, new_AGEMA_signal_10605, MixColumnsIns_MixOneColumnInst_1_n21}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U26 ( .a ({new_AGEMA_signal_10608, new_AGEMA_signal_10607, MixColumnsIns_MixOneColumnInst_1_n56}), .b ({new_AGEMA_signal_10306, new_AGEMA_signal_10305, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .c ({new_AGEMA_signal_11052, new_AGEMA_signal_11051, MixColumnsIns_MixOneColumnInst_1_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U25 ( .a ({new_AGEMA_signal_10392, new_AGEMA_signal_10391, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .b ({new_AGEMA_signal_10376, new_AGEMA_signal_10375, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .c ({new_AGEMA_signal_10608, new_AGEMA_signal_10607, MixColumnsIns_MixOneColumnInst_1_n56}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U24 ( .a ({new_AGEMA_signal_11054, new_AGEMA_signal_11053, MixColumnsIns_MixOneColumnInst_1_n6}), .b ({new_AGEMA_signal_10610, new_AGEMA_signal_10609, MixColumnsIns_MixOneColumnInst_1_n19}), .c ({new_AGEMA_signal_11506, new_AGEMA_signal_11505, MixColumnsOutput[78]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U23 ( .a ({new_AGEMA_signal_10392, new_AGEMA_signal_10391, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .b ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .c ({new_AGEMA_signal_10610, new_AGEMA_signal_10609, MixColumnsIns_MixOneColumnInst_1_n19}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U22 ( .a ({new_AGEMA_signal_10612, new_AGEMA_signal_10611, MixColumnsIns_MixOneColumnInst_1_n53}), .b ({new_AGEMA_signal_10308, new_AGEMA_signal_10307, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .c ({new_AGEMA_signal_11054, new_AGEMA_signal_11053, MixColumnsIns_MixOneColumnInst_1_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U21 ( .a ({new_AGEMA_signal_10394, new_AGEMA_signal_10393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .b ({new_AGEMA_signal_10378, new_AGEMA_signal_10377, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .c ({new_AGEMA_signal_10612, new_AGEMA_signal_10611, MixColumnsIns_MixOneColumnInst_1_n53}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U20 ( .a ({new_AGEMA_signal_11056, new_AGEMA_signal_11055, MixColumnsIns_MixOneColumnInst_1_n5}), .b ({new_AGEMA_signal_10614, new_AGEMA_signal_10613, MixColumnsIns_MixOneColumnInst_1_n17}), .c ({new_AGEMA_signal_11508, new_AGEMA_signal_11507, MixColumnsOutput[77]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U19 ( .a ({new_AGEMA_signal_10394, new_AGEMA_signal_10393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .b ({new_AGEMA_signal_10242, new_AGEMA_signal_10241, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .c ({new_AGEMA_signal_10614, new_AGEMA_signal_10613, MixColumnsIns_MixOneColumnInst_1_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U18 ( .a ({new_AGEMA_signal_10616, new_AGEMA_signal_10615, MixColumnsIns_MixOneColumnInst_1_n50}), .b ({new_AGEMA_signal_10310, new_AGEMA_signal_10309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .c ({new_AGEMA_signal_11056, new_AGEMA_signal_11055, MixColumnsIns_MixOneColumnInst_1_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U17 ( .a ({new_AGEMA_signal_10396, new_AGEMA_signal_10395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .b ({new_AGEMA_signal_10380, new_AGEMA_signal_10379, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .c ({new_AGEMA_signal_10616, new_AGEMA_signal_10615, MixColumnsIns_MixOneColumnInst_1_n50}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U16 ( .a ({new_AGEMA_signal_11510, new_AGEMA_signal_11509, MixColumnsIns_MixOneColumnInst_1_n4}), .b ({new_AGEMA_signal_11058, new_AGEMA_signal_11057, MixColumnsIns_MixOneColumnInst_1_n15}), .c ({new_AGEMA_signal_12036, new_AGEMA_signal_12035, MixColumnsOutput[76]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U15 ( .a ({new_AGEMA_signal_10396, new_AGEMA_signal_10395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .b ({new_AGEMA_signal_10638, new_AGEMA_signal_10637, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]}), .c ({new_AGEMA_signal_11058, new_AGEMA_signal_11057, MixColumnsIns_MixOneColumnInst_1_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U14 ( .a ({new_AGEMA_signal_11060, new_AGEMA_signal_11059, MixColumnsIns_MixOneColumnInst_1_n47}), .b ({new_AGEMA_signal_10312, new_AGEMA_signal_10311, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .c ({new_AGEMA_signal_11510, new_AGEMA_signal_11509, MixColumnsIns_MixOneColumnInst_1_n4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U13 ( .a ({new_AGEMA_signal_10644, new_AGEMA_signal_10643, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]}), .b ({new_AGEMA_signal_10382, new_AGEMA_signal_10381, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .c ({new_AGEMA_signal_11060, new_AGEMA_signal_11059, MixColumnsIns_MixOneColumnInst_1_n47}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U12 ( .a ({new_AGEMA_signal_11512, new_AGEMA_signal_11511, MixColumnsIns_MixOneColumnInst_1_n3}), .b ({new_AGEMA_signal_11062, new_AGEMA_signal_11061, MixColumnsIns_MixOneColumnInst_1_n12}), .c ({new_AGEMA_signal_12038, new_AGEMA_signal_12037, MixColumnsOutput[75]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U11 ( .a ({new_AGEMA_signal_10398, new_AGEMA_signal_10397, MixColumnsInput[67]}), .b ({new_AGEMA_signal_10640, new_AGEMA_signal_10639, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]}), .c ({new_AGEMA_signal_11062, new_AGEMA_signal_11061, MixColumnsIns_MixOneColumnInst_1_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U10 ( .a ({new_AGEMA_signal_11064, new_AGEMA_signal_11063, MixColumnsIns_MixOneColumnInst_1_n44}), .b ({new_AGEMA_signal_10314, new_AGEMA_signal_10313, MixColumnsInput[83]}), .c ({new_AGEMA_signal_11512, new_AGEMA_signal_11511, MixColumnsIns_MixOneColumnInst_1_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U9 ( .a ({new_AGEMA_signal_10646, new_AGEMA_signal_10645, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]}), .b ({new_AGEMA_signal_10384, new_AGEMA_signal_10383, MixColumnsInput[91]}), .c ({new_AGEMA_signal_11064, new_AGEMA_signal_11063, MixColumnsIns_MixOneColumnInst_1_n44}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U8 ( .a ({new_AGEMA_signal_11066, new_AGEMA_signal_11065, MixColumnsIns_MixOneColumnInst_1_n2}), .b ({new_AGEMA_signal_10618, new_AGEMA_signal_10617, MixColumnsIns_MixOneColumnInst_1_n10}), .c ({new_AGEMA_signal_11514, new_AGEMA_signal_11513, MixColumnsOutput[74]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U7 ( .a ({new_AGEMA_signal_10400, new_AGEMA_signal_10399, MixColumnsInput[66]}), .b ({new_AGEMA_signal_10248, new_AGEMA_signal_10247, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .c ({new_AGEMA_signal_10618, new_AGEMA_signal_10617, MixColumnsIns_MixOneColumnInst_1_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U6 ( .a ({new_AGEMA_signal_10620, new_AGEMA_signal_10619, MixColumnsIns_MixOneColumnInst_1_n37}), .b ({new_AGEMA_signal_10316, new_AGEMA_signal_10315, MixColumnsInput[82]}), .c ({new_AGEMA_signal_11066, new_AGEMA_signal_11065, MixColumnsIns_MixOneColumnInst_1_n2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U5 ( .a ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .b ({new_AGEMA_signal_10386, new_AGEMA_signal_10385, MixColumnsInput[90]}), .c ({new_AGEMA_signal_10620, new_AGEMA_signal_10619, MixColumnsIns_MixOneColumnInst_1_n37}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U4 ( .a ({new_AGEMA_signal_11068, new_AGEMA_signal_11067, MixColumnsIns_MixOneColumnInst_1_n1}), .b ({new_AGEMA_signal_9848, new_AGEMA_signal_9847, MixColumnsInput[72]}), .c ({new_AGEMA_signal_11516, new_AGEMA_signal_11515, MixColumnsOutput[64]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U3 ( .a ({new_AGEMA_signal_10624, new_AGEMA_signal_10623, MixColumnsIns_MixOneColumnInst_1_n59}), .b ({new_AGEMA_signal_10622, new_AGEMA_signal_10621, MixColumnsIns_MixOneColumnInst_1_n23}), .c ({new_AGEMA_signal_11068, new_AGEMA_signal_11067, MixColumnsIns_MixOneColumnInst_1_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U2 ( .a ({new_AGEMA_signal_9958, new_AGEMA_signal_9957, MixColumnsInput[80]}), .b ({new_AGEMA_signal_10376, new_AGEMA_signal_10375, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .c ({new_AGEMA_signal_10622, new_AGEMA_signal_10621, MixColumnsIns_MixOneColumnInst_1_n23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U1 ( .a ({new_AGEMA_signal_10390, new_AGEMA_signal_10389, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_10068, new_AGEMA_signal_10067, MixColumnsInput[88]}), .c ({new_AGEMA_signal_10624, new_AGEMA_signal_10623, MixColumnsIns_MixOneColumnInst_1_n59}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_10376, new_AGEMA_signal_10375, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_10384, new_AGEMA_signal_10383, MixColumnsInput[91]}), .c ({new_AGEMA_signal_10626, new_AGEMA_signal_10625, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_10376, new_AGEMA_signal_10375, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_10386, new_AGEMA_signal_10385, MixColumnsInput[90]}), .c ({new_AGEMA_signal_10628, new_AGEMA_signal_10627, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_10376, new_AGEMA_signal_10375, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_10068, new_AGEMA_signal_10067, MixColumnsInput[88]}), .c ({new_AGEMA_signal_10630, new_AGEMA_signal_10629, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_10306, new_AGEMA_signal_10305, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_10314, new_AGEMA_signal_10313, MixColumnsInput[83]}), .c ({new_AGEMA_signal_10632, new_AGEMA_signal_10631, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_10306, new_AGEMA_signal_10305, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_10316, new_AGEMA_signal_10315, MixColumnsInput[82]}), .c ({new_AGEMA_signal_10634, new_AGEMA_signal_10633, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_10306, new_AGEMA_signal_10305, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_9958, new_AGEMA_signal_9957, MixColumnsInput[80]}), .c ({new_AGEMA_signal_10636, new_AGEMA_signal_10635, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_10244, new_AGEMA_signal_10243, MixColumnsInput[75]}), .c ({new_AGEMA_signal_10638, new_AGEMA_signal_10637, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, MixColumnsInput[74]}), .c ({new_AGEMA_signal_10640, new_AGEMA_signal_10639, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_9848, new_AGEMA_signal_9847, MixColumnsInput[72]}), .c ({new_AGEMA_signal_10642, new_AGEMA_signal_10641, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_10390, new_AGEMA_signal_10389, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_10398, new_AGEMA_signal_10397, MixColumnsInput[67]}), .c ({new_AGEMA_signal_10644, new_AGEMA_signal_10643, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_10390, new_AGEMA_signal_10389, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_10400, new_AGEMA_signal_10399, MixColumnsInput[66]}), .c ({new_AGEMA_signal_10646, new_AGEMA_signal_10645, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_10390, new_AGEMA_signal_10389, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_10090, new_AGEMA_signal_10089, MixColumnsInput[64]}), .c ({new_AGEMA_signal_10648, new_AGEMA_signal_10647, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U96 ( .a ({new_AGEMA_signal_11518, new_AGEMA_signal_11517, MixColumnsIns_MixOneColumnInst_2_n64}), .b ({new_AGEMA_signal_10262, new_AGEMA_signal_10261, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .c ({new_AGEMA_signal_12040, new_AGEMA_signal_12039, MixColumnsOutput[41]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U95 ( .a ({new_AGEMA_signal_11112, new_AGEMA_signal_11111, MixColumnsIns_MixOneColumnInst_2_n63}), .b ({new_AGEMA_signal_11104, new_AGEMA_signal_11103, MixColumnsIns_MixOneColumnInst_2_n62}), .c ({new_AGEMA_signal_11518, new_AGEMA_signal_11517, MixColumnsIns_MixOneColumnInst_2_n64}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U94 ( .a ({new_AGEMA_signal_11070, new_AGEMA_signal_11069, MixColumnsIns_MixOneColumnInst_2_n61}), .b ({new_AGEMA_signal_10668, new_AGEMA_signal_10667, MixColumnsIns_MixOneColumnInst_2_n60}), .c ({new_AGEMA_signal_11520, new_AGEMA_signal_11519, MixColumnsOutput[40]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U93 ( .a ({new_AGEMA_signal_10688, new_AGEMA_signal_10687, MixColumnsIns_MixOneColumnInst_2_n59}), .b ({new_AGEMA_signal_9870, new_AGEMA_signal_9869, MixColumnsInput[48]}), .c ({new_AGEMA_signal_11070, new_AGEMA_signal_11069, MixColumnsIns_MixOneColumnInst_2_n61}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U92 ( .a ({new_AGEMA_signal_11072, new_AGEMA_signal_11071, MixColumnsIns_MixOneColumnInst_2_n58}), .b ({new_AGEMA_signal_10650, new_AGEMA_signal_10649, MixColumnsIns_MixOneColumnInst_2_n57}), .c ({new_AGEMA_signal_11522, new_AGEMA_signal_11521, MixColumnsOutput[39]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U91 ( .a ({new_AGEMA_signal_10672, new_AGEMA_signal_10671, MixColumnsIns_MixOneColumnInst_2_n56}), .b ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .c ({new_AGEMA_signal_11072, new_AGEMA_signal_11071, MixColumnsIns_MixOneColumnInst_2_n58}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U90 ( .a ({new_AGEMA_signal_11074, new_AGEMA_signal_11073, MixColumnsIns_MixOneColumnInst_2_n55}), .b ({new_AGEMA_signal_10652, new_AGEMA_signal_10651, MixColumnsIns_MixOneColumnInst_2_n54}), .c ({new_AGEMA_signal_11524, new_AGEMA_signal_11523, MixColumnsOutput[38]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U89 ( .a ({new_AGEMA_signal_10676, new_AGEMA_signal_10675, MixColumnsIns_MixOneColumnInst_2_n53}), .b ({new_AGEMA_signal_10406, new_AGEMA_signal_10405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .c ({new_AGEMA_signal_11074, new_AGEMA_signal_11073, MixColumnsIns_MixOneColumnInst_2_n55}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U88 ( .a ({new_AGEMA_signal_11076, new_AGEMA_signal_11075, MixColumnsIns_MixOneColumnInst_2_n52}), .b ({new_AGEMA_signal_10654, new_AGEMA_signal_10653, MixColumnsIns_MixOneColumnInst_2_n51}), .c ({new_AGEMA_signal_11526, new_AGEMA_signal_11525, MixColumnsOutput[37]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U87 ( .a ({new_AGEMA_signal_10680, new_AGEMA_signal_10679, MixColumnsIns_MixOneColumnInst_2_n50}), .b ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .c ({new_AGEMA_signal_11076, new_AGEMA_signal_11075, MixColumnsIns_MixOneColumnInst_2_n52}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U86 ( .a ({new_AGEMA_signal_11528, new_AGEMA_signal_11527, MixColumnsIns_MixOneColumnInst_2_n49}), .b ({new_AGEMA_signal_11086, new_AGEMA_signal_11085, MixColumnsIns_MixOneColumnInst_2_n48}), .c ({new_AGEMA_signal_12042, new_AGEMA_signal_12041, MixColumnsOutput[36]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U85 ( .a ({new_AGEMA_signal_11124, new_AGEMA_signal_11123, MixColumnsIns_MixOneColumnInst_2_n47}), .b ({new_AGEMA_signal_10410, new_AGEMA_signal_10409, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .c ({new_AGEMA_signal_11528, new_AGEMA_signal_11527, MixColumnsIns_MixOneColumnInst_2_n49}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U84 ( .a ({new_AGEMA_signal_11530, new_AGEMA_signal_11529, MixColumnsIns_MixOneColumnInst_2_n46}), .b ({new_AGEMA_signal_11088, new_AGEMA_signal_11087, MixColumnsIns_MixOneColumnInst_2_n45}), .c ({new_AGEMA_signal_12044, new_AGEMA_signal_12043, MixColumnsOutput[35]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U83 ( .a ({new_AGEMA_signal_11128, new_AGEMA_signal_11127, MixColumnsIns_MixOneColumnInst_2_n44}), .b ({new_AGEMA_signal_10412, new_AGEMA_signal_10411, MixColumnsInput[43]}), .c ({new_AGEMA_signal_11530, new_AGEMA_signal_11529, MixColumnsIns_MixOneColumnInst_2_n46}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U82 ( .a ({new_AGEMA_signal_11078, new_AGEMA_signal_11077, MixColumnsIns_MixOneColumnInst_2_n43}), .b ({new_AGEMA_signal_10650, new_AGEMA_signal_10649, MixColumnsIns_MixOneColumnInst_2_n57}), .c ({new_AGEMA_signal_11532, new_AGEMA_signal_11531, MixColumnsOutput[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U81 ( .a ({new_AGEMA_signal_10250, new_AGEMA_signal_10249, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_10322, new_AGEMA_signal_10321, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .c ({new_AGEMA_signal_10650, new_AGEMA_signal_10649, MixColumnsIns_MixOneColumnInst_2_n57}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U80 ( .a ({new_AGEMA_signal_10334, new_AGEMA_signal_10333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_10658, new_AGEMA_signal_10657, MixColumnsIns_MixOneColumnInst_2_n42}), .c ({new_AGEMA_signal_11078, new_AGEMA_signal_11077, MixColumnsIns_MixOneColumnInst_2_n43}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U79 ( .a ({new_AGEMA_signal_11080, new_AGEMA_signal_11079, MixColumnsIns_MixOneColumnInst_2_n41}), .b ({new_AGEMA_signal_10652, new_AGEMA_signal_10651, MixColumnsIns_MixOneColumnInst_2_n54}), .c ({new_AGEMA_signal_11534, new_AGEMA_signal_11533, MixColumnsOutput[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U78 ( .a ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .b ({new_AGEMA_signal_10324, new_AGEMA_signal_10323, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .c ({new_AGEMA_signal_10652, new_AGEMA_signal_10651, MixColumnsIns_MixOneColumnInst_2_n54}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U77 ( .a ({new_AGEMA_signal_10336, new_AGEMA_signal_10335, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .b ({new_AGEMA_signal_10660, new_AGEMA_signal_10659, MixColumnsIns_MixOneColumnInst_2_n40}), .c ({new_AGEMA_signal_11080, new_AGEMA_signal_11079, MixColumnsIns_MixOneColumnInst_2_n41}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U76 ( .a ({new_AGEMA_signal_11082, new_AGEMA_signal_11081, MixColumnsIns_MixOneColumnInst_2_n39}), .b ({new_AGEMA_signal_10656, new_AGEMA_signal_10655, MixColumnsIns_MixOneColumnInst_2_n38}), .c ({new_AGEMA_signal_11536, new_AGEMA_signal_11535, MixColumnsOutput[34]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U75 ( .a ({new_AGEMA_signal_10684, new_AGEMA_signal_10683, MixColumnsIns_MixOneColumnInst_2_n37}), .b ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, MixColumnsInput[42]}), .c ({new_AGEMA_signal_11082, new_AGEMA_signal_11081, MixColumnsIns_MixOneColumnInst_2_n39}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U74 ( .a ({new_AGEMA_signal_11084, new_AGEMA_signal_11083, MixColumnsIns_MixOneColumnInst_2_n36}), .b ({new_AGEMA_signal_10654, new_AGEMA_signal_10653, MixColumnsIns_MixOneColumnInst_2_n51}), .c ({new_AGEMA_signal_11538, new_AGEMA_signal_11537, MixColumnsOutput[61]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U73 ( .a ({new_AGEMA_signal_10254, new_AGEMA_signal_10253, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .b ({new_AGEMA_signal_10326, new_AGEMA_signal_10325, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .c ({new_AGEMA_signal_10654, new_AGEMA_signal_10653, MixColumnsIns_MixOneColumnInst_2_n51}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U72 ( .a ({new_AGEMA_signal_10338, new_AGEMA_signal_10337, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .b ({new_AGEMA_signal_10662, new_AGEMA_signal_10661, MixColumnsIns_MixOneColumnInst_2_n35}), .c ({new_AGEMA_signal_11084, new_AGEMA_signal_11083, MixColumnsIns_MixOneColumnInst_2_n36}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U71 ( .a ({new_AGEMA_signal_11540, new_AGEMA_signal_11539, MixColumnsIns_MixOneColumnInst_2_n34}), .b ({new_AGEMA_signal_11086, new_AGEMA_signal_11085, MixColumnsIns_MixOneColumnInst_2_n48}), .c ({new_AGEMA_signal_12046, new_AGEMA_signal_12045, MixColumnsOutput[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U70 ( .a ({new_AGEMA_signal_10256, new_AGEMA_signal_10255, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .b ({new_AGEMA_signal_10690, new_AGEMA_signal_10689, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]}), .c ({new_AGEMA_signal_11086, new_AGEMA_signal_11085, MixColumnsIns_MixOneColumnInst_2_n48}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U69 ( .a ({new_AGEMA_signal_10340, new_AGEMA_signal_10339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .b ({new_AGEMA_signal_11100, new_AGEMA_signal_11099, MixColumnsIns_MixOneColumnInst_2_n33}), .c ({new_AGEMA_signal_11540, new_AGEMA_signal_11539, MixColumnsIns_MixOneColumnInst_2_n34}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U68 ( .a ({new_AGEMA_signal_11542, new_AGEMA_signal_11541, MixColumnsIns_MixOneColumnInst_2_n32}), .b ({new_AGEMA_signal_11088, new_AGEMA_signal_11087, MixColumnsIns_MixOneColumnInst_2_n45}), .c ({new_AGEMA_signal_12048, new_AGEMA_signal_12047, MixColumnsOutput[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U67 ( .a ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, MixColumnsInput[51]}), .b ({new_AGEMA_signal_10692, new_AGEMA_signal_10691, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]}), .c ({new_AGEMA_signal_11088, new_AGEMA_signal_11087, MixColumnsIns_MixOneColumnInst_2_n45}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U66 ( .a ({new_AGEMA_signal_10342, new_AGEMA_signal_10341, MixColumnsInput[35]}), .b ({new_AGEMA_signal_11106, new_AGEMA_signal_11105, MixColumnsIns_MixOneColumnInst_2_n31}), .c ({new_AGEMA_signal_11542, new_AGEMA_signal_11541, MixColumnsIns_MixOneColumnInst_2_n32}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U65 ( .a ({new_AGEMA_signal_11090, new_AGEMA_signal_11089, MixColumnsIns_MixOneColumnInst_2_n30}), .b ({new_AGEMA_signal_10656, new_AGEMA_signal_10655, MixColumnsIns_MixOneColumnInst_2_n38}), .c ({new_AGEMA_signal_11544, new_AGEMA_signal_11543, MixColumnsOutput[58]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U64 ( .a ({new_AGEMA_signal_10260, new_AGEMA_signal_10259, MixColumnsInput[50]}), .b ({new_AGEMA_signal_10332, new_AGEMA_signal_10331, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .c ({new_AGEMA_signal_10656, new_AGEMA_signal_10655, MixColumnsIns_MixOneColumnInst_2_n38}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U63 ( .a ({new_AGEMA_signal_10344, new_AGEMA_signal_10343, MixColumnsInput[34]}), .b ({new_AGEMA_signal_10664, new_AGEMA_signal_10663, MixColumnsIns_MixOneColumnInst_2_n29}), .c ({new_AGEMA_signal_11090, new_AGEMA_signal_11089, MixColumnsIns_MixOneColumnInst_2_n30}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U62 ( .a ({new_AGEMA_signal_11546, new_AGEMA_signal_11545, MixColumnsIns_MixOneColumnInst_2_n28}), .b ({new_AGEMA_signal_11102, new_AGEMA_signal_11101, MixColumnsIns_MixOneColumnInst_2_n27}), .c ({new_AGEMA_signal_12050, new_AGEMA_signal_12049, MixColumnsOutput[57]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U61 ( .a ({new_AGEMA_signal_10346, new_AGEMA_signal_10345, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .b ({new_AGEMA_signal_11110, new_AGEMA_signal_11109, MixColumnsIns_MixOneColumnInst_2_n26}), .c ({new_AGEMA_signal_11546, new_AGEMA_signal_11545, MixColumnsIns_MixOneColumnInst_2_n28}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U60 ( .a ({new_AGEMA_signal_11092, new_AGEMA_signal_11091, MixColumnsIns_MixOneColumnInst_2_n25}), .b ({new_AGEMA_signal_10666, new_AGEMA_signal_10665, MixColumnsIns_MixOneColumnInst_2_n24}), .c ({new_AGEMA_signal_11548, new_AGEMA_signal_11547, MixColumnsOutput[56]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U59 ( .a ({new_AGEMA_signal_10686, new_AGEMA_signal_10685, MixColumnsIns_MixOneColumnInst_2_n23}), .b ({new_AGEMA_signal_10002, new_AGEMA_signal_10001, MixColumnsInput[32]}), .c ({new_AGEMA_signal_11092, new_AGEMA_signal_11091, MixColumnsIns_MixOneColumnInst_2_n25}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U58 ( .a ({new_AGEMA_signal_11094, new_AGEMA_signal_11093, MixColumnsIns_MixOneColumnInst_2_n22}), .b ({new_AGEMA_signal_10658, new_AGEMA_signal_10657, MixColumnsIns_MixOneColumnInst_2_n42}), .c ({new_AGEMA_signal_11550, new_AGEMA_signal_11549, MixColumnsOutput[55]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U57 ( .a ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .c ({new_AGEMA_signal_10658, new_AGEMA_signal_10657, MixColumnsIns_MixOneColumnInst_2_n42}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U56 ( .a ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_10670, new_AGEMA_signal_10669, MixColumnsIns_MixOneColumnInst_2_n21}), .c ({new_AGEMA_signal_11094, new_AGEMA_signal_11093, MixColumnsIns_MixOneColumnInst_2_n22}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U55 ( .a ({new_AGEMA_signal_11096, new_AGEMA_signal_11095, MixColumnsIns_MixOneColumnInst_2_n20}), .b ({new_AGEMA_signal_10660, new_AGEMA_signal_10659, MixColumnsIns_MixOneColumnInst_2_n40}), .c ({new_AGEMA_signal_11552, new_AGEMA_signal_11551, MixColumnsOutput[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U54 ( .a ({new_AGEMA_signal_10406, new_AGEMA_signal_10405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .b ({new_AGEMA_signal_10254, new_AGEMA_signal_10253, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .c ({new_AGEMA_signal_10660, new_AGEMA_signal_10659, MixColumnsIns_MixOneColumnInst_2_n40}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U53 ( .a ({new_AGEMA_signal_10322, new_AGEMA_signal_10321, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .b ({new_AGEMA_signal_10674, new_AGEMA_signal_10673, MixColumnsIns_MixOneColumnInst_2_n19}), .c ({new_AGEMA_signal_11096, new_AGEMA_signal_11095, MixColumnsIns_MixOneColumnInst_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U52 ( .a ({new_AGEMA_signal_11098, new_AGEMA_signal_11097, MixColumnsIns_MixOneColumnInst_2_n18}), .b ({new_AGEMA_signal_10662, new_AGEMA_signal_10661, MixColumnsIns_MixOneColumnInst_2_n35}), .c ({new_AGEMA_signal_11554, new_AGEMA_signal_11553, MixColumnsOutput[53]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U51 ( .a ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .b ({new_AGEMA_signal_10256, new_AGEMA_signal_10255, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .c ({new_AGEMA_signal_10662, new_AGEMA_signal_10661, MixColumnsIns_MixOneColumnInst_2_n35}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U50 ( .a ({new_AGEMA_signal_10324, new_AGEMA_signal_10323, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .b ({new_AGEMA_signal_10678, new_AGEMA_signal_10677, MixColumnsIns_MixOneColumnInst_2_n17}), .c ({new_AGEMA_signal_11098, new_AGEMA_signal_11097, MixColumnsIns_MixOneColumnInst_2_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U49 ( .a ({new_AGEMA_signal_11556, new_AGEMA_signal_11555, MixColumnsIns_MixOneColumnInst_2_n16}), .b ({new_AGEMA_signal_11100, new_AGEMA_signal_11099, MixColumnsIns_MixOneColumnInst_2_n33}), .c ({new_AGEMA_signal_12052, new_AGEMA_signal_12051, MixColumnsOutput[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U48 ( .a ({new_AGEMA_signal_10410, new_AGEMA_signal_10409, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .b ({new_AGEMA_signal_10696, new_AGEMA_signal_10695, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]}), .c ({new_AGEMA_signal_11100, new_AGEMA_signal_11099, MixColumnsIns_MixOneColumnInst_2_n33}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U47 ( .a ({new_AGEMA_signal_10326, new_AGEMA_signal_10325, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .b ({new_AGEMA_signal_11122, new_AGEMA_signal_11121, MixColumnsIns_MixOneColumnInst_2_n15}), .c ({new_AGEMA_signal_11556, new_AGEMA_signal_11555, MixColumnsIns_MixOneColumnInst_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U46 ( .a ({new_AGEMA_signal_11558, new_AGEMA_signal_11557, MixColumnsIns_MixOneColumnInst_2_n14}), .b ({new_AGEMA_signal_11102, new_AGEMA_signal_11101, MixColumnsIns_MixOneColumnInst_2_n27}), .c ({new_AGEMA_signal_12054, new_AGEMA_signal_12053, MixColumnsOutput[33]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U45 ( .a ({new_AGEMA_signal_10262, new_AGEMA_signal_10261, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .b ({new_AGEMA_signal_10694, new_AGEMA_signal_10693, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]}), .c ({new_AGEMA_signal_11102, new_AGEMA_signal_11101, MixColumnsIns_MixOneColumnInst_2_n27}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U44 ( .a ({new_AGEMA_signal_10416, new_AGEMA_signal_10415, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .b ({new_AGEMA_signal_11104, new_AGEMA_signal_11103, MixColumnsIns_MixOneColumnInst_2_n62}), .c ({new_AGEMA_signal_11558, new_AGEMA_signal_11557, MixColumnsIns_MixOneColumnInst_2_n14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U43 ( .a ({new_AGEMA_signal_10332, new_AGEMA_signal_10331, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .b ({new_AGEMA_signal_10712, new_AGEMA_signal_10711, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]}), .c ({new_AGEMA_signal_11104, new_AGEMA_signal_11103, MixColumnsIns_MixOneColumnInst_2_n62}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U42 ( .a ({new_AGEMA_signal_11560, new_AGEMA_signal_11559, MixColumnsIns_MixOneColumnInst_2_n13}), .b ({new_AGEMA_signal_11106, new_AGEMA_signal_11105, MixColumnsIns_MixOneColumnInst_2_n31}), .c ({new_AGEMA_signal_12056, new_AGEMA_signal_12055, MixColumnsOutput[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U41 ( .a ({new_AGEMA_signal_10412, new_AGEMA_signal_10411, MixColumnsInput[43]}), .b ({new_AGEMA_signal_10698, new_AGEMA_signal_10697, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]}), .c ({new_AGEMA_signal_11106, new_AGEMA_signal_11105, MixColumnsIns_MixOneColumnInst_2_n31}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U40 ( .a ({new_AGEMA_signal_10328, new_AGEMA_signal_10327, MixColumnsInput[59]}), .b ({new_AGEMA_signal_11126, new_AGEMA_signal_11125, MixColumnsIns_MixOneColumnInst_2_n12}), .c ({new_AGEMA_signal_11560, new_AGEMA_signal_11559, MixColumnsIns_MixOneColumnInst_2_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U39 ( .a ({new_AGEMA_signal_11108, new_AGEMA_signal_11107, MixColumnsIns_MixOneColumnInst_2_n11}), .b ({new_AGEMA_signal_10664, new_AGEMA_signal_10663, MixColumnsIns_MixOneColumnInst_2_n29}), .c ({new_AGEMA_signal_11562, new_AGEMA_signal_11561, MixColumnsOutput[50]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U38 ( .a ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, MixColumnsInput[42]}), .b ({new_AGEMA_signal_10262, new_AGEMA_signal_10261, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .c ({new_AGEMA_signal_10664, new_AGEMA_signal_10663, MixColumnsIns_MixOneColumnInst_2_n29}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U37 ( .a ({new_AGEMA_signal_10330, new_AGEMA_signal_10329, MixColumnsInput[58]}), .b ({new_AGEMA_signal_10682, new_AGEMA_signal_10681, MixColumnsIns_MixOneColumnInst_2_n10}), .c ({new_AGEMA_signal_11108, new_AGEMA_signal_11107, MixColumnsIns_MixOneColumnInst_2_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U36 ( .a ({new_AGEMA_signal_11564, new_AGEMA_signal_11563, MixColumnsIns_MixOneColumnInst_2_n9}), .b ({new_AGEMA_signal_11110, new_AGEMA_signal_11109, MixColumnsIns_MixOneColumnInst_2_n26}), .c ({new_AGEMA_signal_12058, new_AGEMA_signal_12057, MixColumnsOutput[49]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U35 ( .a ({new_AGEMA_signal_10700, new_AGEMA_signal_10699, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]}), .b ({new_AGEMA_signal_10416, new_AGEMA_signal_10415, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .c ({new_AGEMA_signal_11110, new_AGEMA_signal_11109, MixColumnsIns_MixOneColumnInst_2_n26}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U34 ( .a ({new_AGEMA_signal_11112, new_AGEMA_signal_11111, MixColumnsIns_MixOneColumnInst_2_n63}), .b ({new_AGEMA_signal_10332, new_AGEMA_signal_10331, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .c ({new_AGEMA_signal_11564, new_AGEMA_signal_11563, MixColumnsIns_MixOneColumnInst_2_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U33 ( .a ({new_AGEMA_signal_10706, new_AGEMA_signal_10705, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]}), .b ({new_AGEMA_signal_10346, new_AGEMA_signal_10345, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .c ({new_AGEMA_signal_11112, new_AGEMA_signal_11111, MixColumnsIns_MixOneColumnInst_2_n63}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U32 ( .a ({new_AGEMA_signal_11114, new_AGEMA_signal_11113, MixColumnsIns_MixOneColumnInst_2_n8}), .b ({new_AGEMA_signal_10666, new_AGEMA_signal_10665, MixColumnsIns_MixOneColumnInst_2_n24}), .c ({new_AGEMA_signal_11566, new_AGEMA_signal_11565, MixColumnsOutput[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U31 ( .a ({new_AGEMA_signal_10112, new_AGEMA_signal_10111, MixColumnsInput[40]}), .b ({new_AGEMA_signal_10250, new_AGEMA_signal_10249, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .c ({new_AGEMA_signal_10666, new_AGEMA_signal_10665, MixColumnsIns_MixOneColumnInst_2_n24}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U30 ( .a ({new_AGEMA_signal_9980, new_AGEMA_signal_9979, MixColumnsInput[56]}), .b ({new_AGEMA_signal_10668, new_AGEMA_signal_10667, MixColumnsIns_MixOneColumnInst_2_n60}), .c ({new_AGEMA_signal_11114, new_AGEMA_signal_11113, MixColumnsIns_MixOneColumnInst_2_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U29 ( .a ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_10002, new_AGEMA_signal_10001, MixColumnsInput[32]}), .c ({new_AGEMA_signal_10668, new_AGEMA_signal_10667, MixColumnsIns_MixOneColumnInst_2_n60}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U28 ( .a ({new_AGEMA_signal_11116, new_AGEMA_signal_11115, MixColumnsIns_MixOneColumnInst_2_n7}), .b ({new_AGEMA_signal_10670, new_AGEMA_signal_10669, MixColumnsIns_MixOneColumnInst_2_n21}), .c ({new_AGEMA_signal_11568, new_AGEMA_signal_11567, MixColumnsOutput[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U27 ( .a ({new_AGEMA_signal_10334, new_AGEMA_signal_10333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_10406, new_AGEMA_signal_10405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .c ({new_AGEMA_signal_10670, new_AGEMA_signal_10669, MixColumnsIns_MixOneColumnInst_2_n21}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U26 ( .a ({new_AGEMA_signal_10672, new_AGEMA_signal_10671, MixColumnsIns_MixOneColumnInst_2_n56}), .b ({new_AGEMA_signal_10250, new_AGEMA_signal_10249, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .c ({new_AGEMA_signal_11116, new_AGEMA_signal_11115, MixColumnsIns_MixOneColumnInst_2_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U25 ( .a ({new_AGEMA_signal_10336, new_AGEMA_signal_10335, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .b ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .c ({new_AGEMA_signal_10672, new_AGEMA_signal_10671, MixColumnsIns_MixOneColumnInst_2_n56}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U24 ( .a ({new_AGEMA_signal_11118, new_AGEMA_signal_11117, MixColumnsIns_MixOneColumnInst_2_n6}), .b ({new_AGEMA_signal_10674, new_AGEMA_signal_10673, MixColumnsIns_MixOneColumnInst_2_n19}), .c ({new_AGEMA_signal_11570, new_AGEMA_signal_11569, MixColumnsOutput[46]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U23 ( .a ({new_AGEMA_signal_10336, new_AGEMA_signal_10335, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .b ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .c ({new_AGEMA_signal_10674, new_AGEMA_signal_10673, MixColumnsIns_MixOneColumnInst_2_n19}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U22 ( .a ({new_AGEMA_signal_10676, new_AGEMA_signal_10675, MixColumnsIns_MixOneColumnInst_2_n53}), .b ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .c ({new_AGEMA_signal_11118, new_AGEMA_signal_11117, MixColumnsIns_MixOneColumnInst_2_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U21 ( .a ({new_AGEMA_signal_10338, new_AGEMA_signal_10337, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .b ({new_AGEMA_signal_10322, new_AGEMA_signal_10321, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .c ({new_AGEMA_signal_10676, new_AGEMA_signal_10675, MixColumnsIns_MixOneColumnInst_2_n53}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U20 ( .a ({new_AGEMA_signal_11120, new_AGEMA_signal_11119, MixColumnsIns_MixOneColumnInst_2_n5}), .b ({new_AGEMA_signal_10678, new_AGEMA_signal_10677, MixColumnsIns_MixOneColumnInst_2_n17}), .c ({new_AGEMA_signal_11572, new_AGEMA_signal_11571, MixColumnsOutput[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U19 ( .a ({new_AGEMA_signal_10338, new_AGEMA_signal_10337, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .b ({new_AGEMA_signal_10410, new_AGEMA_signal_10409, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .c ({new_AGEMA_signal_10678, new_AGEMA_signal_10677, MixColumnsIns_MixOneColumnInst_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U18 ( .a ({new_AGEMA_signal_10680, new_AGEMA_signal_10679, MixColumnsIns_MixOneColumnInst_2_n50}), .b ({new_AGEMA_signal_10254, new_AGEMA_signal_10253, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .c ({new_AGEMA_signal_11120, new_AGEMA_signal_11119, MixColumnsIns_MixOneColumnInst_2_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U17 ( .a ({new_AGEMA_signal_10340, new_AGEMA_signal_10339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .b ({new_AGEMA_signal_10324, new_AGEMA_signal_10323, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .c ({new_AGEMA_signal_10680, new_AGEMA_signal_10679, MixColumnsIns_MixOneColumnInst_2_n50}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U16 ( .a ({new_AGEMA_signal_11574, new_AGEMA_signal_11573, MixColumnsIns_MixOneColumnInst_2_n4}), .b ({new_AGEMA_signal_11122, new_AGEMA_signal_11121, MixColumnsIns_MixOneColumnInst_2_n15}), .c ({new_AGEMA_signal_12060, new_AGEMA_signal_12059, MixColumnsOutput[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U15 ( .a ({new_AGEMA_signal_10340, new_AGEMA_signal_10339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .b ({new_AGEMA_signal_10702, new_AGEMA_signal_10701, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]}), .c ({new_AGEMA_signal_11122, new_AGEMA_signal_11121, MixColumnsIns_MixOneColumnInst_2_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U14 ( .a ({new_AGEMA_signal_11124, new_AGEMA_signal_11123, MixColumnsIns_MixOneColumnInst_2_n47}), .b ({new_AGEMA_signal_10256, new_AGEMA_signal_10255, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .c ({new_AGEMA_signal_11574, new_AGEMA_signal_11573, MixColumnsIns_MixOneColumnInst_2_n4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U13 ( .a ({new_AGEMA_signal_10708, new_AGEMA_signal_10707, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]}), .b ({new_AGEMA_signal_10326, new_AGEMA_signal_10325, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .c ({new_AGEMA_signal_11124, new_AGEMA_signal_11123, MixColumnsIns_MixOneColumnInst_2_n47}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U12 ( .a ({new_AGEMA_signal_11576, new_AGEMA_signal_11575, MixColumnsIns_MixOneColumnInst_2_n3}), .b ({new_AGEMA_signal_11126, new_AGEMA_signal_11125, MixColumnsIns_MixOneColumnInst_2_n12}), .c ({new_AGEMA_signal_12062, new_AGEMA_signal_12061, MixColumnsOutput[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U11 ( .a ({new_AGEMA_signal_10342, new_AGEMA_signal_10341, MixColumnsInput[35]}), .b ({new_AGEMA_signal_10704, new_AGEMA_signal_10703, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]}), .c ({new_AGEMA_signal_11126, new_AGEMA_signal_11125, MixColumnsIns_MixOneColumnInst_2_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U10 ( .a ({new_AGEMA_signal_11128, new_AGEMA_signal_11127, MixColumnsIns_MixOneColumnInst_2_n44}), .b ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, MixColumnsInput[51]}), .c ({new_AGEMA_signal_11576, new_AGEMA_signal_11575, MixColumnsIns_MixOneColumnInst_2_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U9 ( .a ({new_AGEMA_signal_10710, new_AGEMA_signal_10709, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]}), .b ({new_AGEMA_signal_10328, new_AGEMA_signal_10327, MixColumnsInput[59]}), .c ({new_AGEMA_signal_11128, new_AGEMA_signal_11127, MixColumnsIns_MixOneColumnInst_2_n44}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U8 ( .a ({new_AGEMA_signal_11130, new_AGEMA_signal_11129, MixColumnsIns_MixOneColumnInst_2_n2}), .b ({new_AGEMA_signal_10682, new_AGEMA_signal_10681, MixColumnsIns_MixOneColumnInst_2_n10}), .c ({new_AGEMA_signal_11578, new_AGEMA_signal_11577, MixColumnsOutput[42]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U7 ( .a ({new_AGEMA_signal_10344, new_AGEMA_signal_10343, MixColumnsInput[34]}), .b ({new_AGEMA_signal_10416, new_AGEMA_signal_10415, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .c ({new_AGEMA_signal_10682, new_AGEMA_signal_10681, MixColumnsIns_MixOneColumnInst_2_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U6 ( .a ({new_AGEMA_signal_10684, new_AGEMA_signal_10683, MixColumnsIns_MixOneColumnInst_2_n37}), .b ({new_AGEMA_signal_10260, new_AGEMA_signal_10259, MixColumnsInput[50]}), .c ({new_AGEMA_signal_11130, new_AGEMA_signal_11129, MixColumnsIns_MixOneColumnInst_2_n2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U5 ( .a ({new_AGEMA_signal_10346, new_AGEMA_signal_10345, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .b ({new_AGEMA_signal_10330, new_AGEMA_signal_10329, MixColumnsInput[58]}), .c ({new_AGEMA_signal_10684, new_AGEMA_signal_10683, MixColumnsIns_MixOneColumnInst_2_n37}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U4 ( .a ({new_AGEMA_signal_11132, new_AGEMA_signal_11131, MixColumnsIns_MixOneColumnInst_2_n1}), .b ({new_AGEMA_signal_10112, new_AGEMA_signal_10111, MixColumnsInput[40]}), .c ({new_AGEMA_signal_11580, new_AGEMA_signal_11579, MixColumnsOutput[32]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U3 ( .a ({new_AGEMA_signal_10688, new_AGEMA_signal_10687, MixColumnsIns_MixOneColumnInst_2_n59}), .b ({new_AGEMA_signal_10686, new_AGEMA_signal_10685, MixColumnsIns_MixOneColumnInst_2_n23}), .c ({new_AGEMA_signal_11132, new_AGEMA_signal_11131, MixColumnsIns_MixOneColumnInst_2_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U2 ( .a ({new_AGEMA_signal_9870, new_AGEMA_signal_9869, MixColumnsInput[48]}), .b ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .c ({new_AGEMA_signal_10686, new_AGEMA_signal_10685, MixColumnsIns_MixOneColumnInst_2_n23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U1 ( .a ({new_AGEMA_signal_10334, new_AGEMA_signal_10333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_9980, new_AGEMA_signal_9979, MixColumnsInput[56]}), .c ({new_AGEMA_signal_10688, new_AGEMA_signal_10687, MixColumnsIns_MixOneColumnInst_2_n59}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_10328, new_AGEMA_signal_10327, MixColumnsInput[59]}), .c ({new_AGEMA_signal_10690, new_AGEMA_signal_10689, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_10330, new_AGEMA_signal_10329, MixColumnsInput[58]}), .c ({new_AGEMA_signal_10692, new_AGEMA_signal_10691, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_9980, new_AGEMA_signal_9979, MixColumnsInput[56]}), .c ({new_AGEMA_signal_10694, new_AGEMA_signal_10693, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_10250, new_AGEMA_signal_10249, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, MixColumnsInput[51]}), .c ({new_AGEMA_signal_10696, new_AGEMA_signal_10695, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_10250, new_AGEMA_signal_10249, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_10260, new_AGEMA_signal_10259, MixColumnsInput[50]}), .c ({new_AGEMA_signal_10698, new_AGEMA_signal_10697, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_10250, new_AGEMA_signal_10249, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_9870, new_AGEMA_signal_9869, MixColumnsInput[48]}), .c ({new_AGEMA_signal_10700, new_AGEMA_signal_10699, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_10412, new_AGEMA_signal_10411, MixColumnsInput[43]}), .c ({new_AGEMA_signal_10702, new_AGEMA_signal_10701, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, MixColumnsInput[42]}), .c ({new_AGEMA_signal_10704, new_AGEMA_signal_10703, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_10112, new_AGEMA_signal_10111, MixColumnsInput[40]}), .c ({new_AGEMA_signal_10706, new_AGEMA_signal_10705, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_10334, new_AGEMA_signal_10333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_10342, new_AGEMA_signal_10341, MixColumnsInput[35]}), .c ({new_AGEMA_signal_10708, new_AGEMA_signal_10707, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_10334, new_AGEMA_signal_10333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_10344, new_AGEMA_signal_10343, MixColumnsInput[34]}), .c ({new_AGEMA_signal_10710, new_AGEMA_signal_10709, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_10334, new_AGEMA_signal_10333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_10002, new_AGEMA_signal_10001, MixColumnsInput[32]}), .c ({new_AGEMA_signal_10712, new_AGEMA_signal_10711, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U96 ( .a ({new_AGEMA_signal_11582, new_AGEMA_signal_11581, MixColumnsIns_MixOneColumnInst_3_n64}), .b ({new_AGEMA_signal_10430, new_AGEMA_signal_10429, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .c ({new_AGEMA_signal_12064, new_AGEMA_signal_12063, MixColumnsOutput[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U95 ( .a ({new_AGEMA_signal_11176, new_AGEMA_signal_11175, MixColumnsIns_MixOneColumnInst_3_n63}), .b ({new_AGEMA_signal_11168, new_AGEMA_signal_11167, MixColumnsIns_MixOneColumnInst_3_n62}), .c ({new_AGEMA_signal_11582, new_AGEMA_signal_11581, MixColumnsIns_MixOneColumnInst_3_n64}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U94 ( .a ({new_AGEMA_signal_11134, new_AGEMA_signal_11133, MixColumnsIns_MixOneColumnInst_3_n61}), .b ({new_AGEMA_signal_10732, new_AGEMA_signal_10731, MixColumnsIns_MixOneColumnInst_3_n60}), .c ({new_AGEMA_signal_11584, new_AGEMA_signal_11583, MixColumnsOutput[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U93 ( .a ({new_AGEMA_signal_10752, new_AGEMA_signal_10751, MixColumnsIns_MixOneColumnInst_3_n59}), .b ({new_AGEMA_signal_10134, new_AGEMA_signal_10133, MixColumnsInput[16]}), .c ({new_AGEMA_signal_11134, new_AGEMA_signal_11133, MixColumnsIns_MixOneColumnInst_3_n61}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U92 ( .a ({new_AGEMA_signal_11136, new_AGEMA_signal_11135, MixColumnsIns_MixOneColumnInst_3_n58}), .b ({new_AGEMA_signal_10714, new_AGEMA_signal_10713, MixColumnsIns_MixOneColumnInst_3_n57}), .c ({new_AGEMA_signal_11586, new_AGEMA_signal_11585, MixColumnsOutput[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U91 ( .a ({new_AGEMA_signal_10736, new_AGEMA_signal_10735, MixColumnsIns_MixOneColumnInst_3_n56}), .b ({new_AGEMA_signal_10348, new_AGEMA_signal_10347, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .c ({new_AGEMA_signal_11136, new_AGEMA_signal_11135, MixColumnsIns_MixOneColumnInst_3_n58}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U90 ( .a ({new_AGEMA_signal_11138, new_AGEMA_signal_11137, MixColumnsIns_MixOneColumnInst_3_n55}), .b ({new_AGEMA_signal_10716, new_AGEMA_signal_10715, MixColumnsIns_MixOneColumnInst_3_n54}), .c ({new_AGEMA_signal_11588, new_AGEMA_signal_11587, MixColumnsOutput[6]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U89 ( .a ({new_AGEMA_signal_10740, new_AGEMA_signal_10739, MixColumnsIns_MixOneColumnInst_3_n53}), .b ({new_AGEMA_signal_10350, new_AGEMA_signal_10349, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .c ({new_AGEMA_signal_11138, new_AGEMA_signal_11137, MixColumnsIns_MixOneColumnInst_3_n55}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U88 ( .a ({new_AGEMA_signal_11140, new_AGEMA_signal_11139, MixColumnsIns_MixOneColumnInst_3_n52}), .b ({new_AGEMA_signal_10718, new_AGEMA_signal_10717, MixColumnsIns_MixOneColumnInst_3_n51}), .c ({new_AGEMA_signal_11590, new_AGEMA_signal_11589, MixColumnsOutput[5]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U87 ( .a ({new_AGEMA_signal_10744, new_AGEMA_signal_10743, MixColumnsIns_MixOneColumnInst_3_n50}), .b ({new_AGEMA_signal_10352, new_AGEMA_signal_10351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .c ({new_AGEMA_signal_11140, new_AGEMA_signal_11139, MixColumnsIns_MixOneColumnInst_3_n52}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U86 ( .a ({new_AGEMA_signal_11592, new_AGEMA_signal_11591, MixColumnsIns_MixOneColumnInst_3_n49}), .b ({new_AGEMA_signal_11150, new_AGEMA_signal_11149, MixColumnsIns_MixOneColumnInst_3_n48}), .c ({new_AGEMA_signal_12066, new_AGEMA_signal_12065, MixColumnsOutput[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U85 ( .a ({new_AGEMA_signal_11188, new_AGEMA_signal_11187, MixColumnsIns_MixOneColumnInst_3_n47}), .b ({new_AGEMA_signal_10354, new_AGEMA_signal_10353, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .c ({new_AGEMA_signal_11592, new_AGEMA_signal_11591, MixColumnsIns_MixOneColumnInst_3_n49}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U84 ( .a ({new_AGEMA_signal_11594, new_AGEMA_signal_11593, MixColumnsIns_MixOneColumnInst_3_n46}), .b ({new_AGEMA_signal_11152, new_AGEMA_signal_11151, MixColumnsIns_MixOneColumnInst_3_n45}), .c ({new_AGEMA_signal_12068, new_AGEMA_signal_12067, MixColumnsOutput[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U83 ( .a ({new_AGEMA_signal_11192, new_AGEMA_signal_11191, MixColumnsIns_MixOneColumnInst_3_n44}), .b ({new_AGEMA_signal_10356, new_AGEMA_signal_10355, MixColumnsInput[11]}), .c ({new_AGEMA_signal_11594, new_AGEMA_signal_11593, MixColumnsIns_MixOneColumnInst_3_n46}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U82 ( .a ({new_AGEMA_signal_11142, new_AGEMA_signal_11141, MixColumnsIns_MixOneColumnInst_3_n43}), .b ({new_AGEMA_signal_10714, new_AGEMA_signal_10713, MixColumnsIns_MixOneColumnInst_3_n57}), .c ({new_AGEMA_signal_11596, new_AGEMA_signal_11595, MixColumnsOutput[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U81 ( .a ({new_AGEMA_signal_10418, new_AGEMA_signal_10417, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_10266, new_AGEMA_signal_10265, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .c ({new_AGEMA_signal_10714, new_AGEMA_signal_10713, MixColumnsIns_MixOneColumnInst_3_n57}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U80 ( .a ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_10722, new_AGEMA_signal_10721, MixColumnsIns_MixOneColumnInst_3_n42}), .c ({new_AGEMA_signal_11142, new_AGEMA_signal_11141, MixColumnsIns_MixOneColumnInst_3_n43}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U79 ( .a ({new_AGEMA_signal_11144, new_AGEMA_signal_11143, MixColumnsIns_MixOneColumnInst_3_n41}), .b ({new_AGEMA_signal_10716, new_AGEMA_signal_10715, MixColumnsIns_MixOneColumnInst_3_n54}), .c ({new_AGEMA_signal_11598, new_AGEMA_signal_11597, MixColumnsOutput[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U78 ( .a ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .b ({new_AGEMA_signal_10268, new_AGEMA_signal_10267, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .c ({new_AGEMA_signal_10716, new_AGEMA_signal_10715, MixColumnsIns_MixOneColumnInst_3_n54}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U77 ( .a ({new_AGEMA_signal_10280, new_AGEMA_signal_10279, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .b ({new_AGEMA_signal_10724, new_AGEMA_signal_10723, MixColumnsIns_MixOneColumnInst_3_n40}), .c ({new_AGEMA_signal_11144, new_AGEMA_signal_11143, MixColumnsIns_MixOneColumnInst_3_n41}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U76 ( .a ({new_AGEMA_signal_11146, new_AGEMA_signal_11145, MixColumnsIns_MixOneColumnInst_3_n39}), .b ({new_AGEMA_signal_10720, new_AGEMA_signal_10719, MixColumnsIns_MixOneColumnInst_3_n38}), .c ({new_AGEMA_signal_11600, new_AGEMA_signal_11599, MixColumnsOutput[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U75 ( .a ({new_AGEMA_signal_10748, new_AGEMA_signal_10747, MixColumnsIns_MixOneColumnInst_3_n37}), .b ({new_AGEMA_signal_10358, new_AGEMA_signal_10357, MixColumnsInput[10]}), .c ({new_AGEMA_signal_11146, new_AGEMA_signal_11145, MixColumnsIns_MixOneColumnInst_3_n39}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U74 ( .a ({new_AGEMA_signal_11148, new_AGEMA_signal_11147, MixColumnsIns_MixOneColumnInst_3_n36}), .b ({new_AGEMA_signal_10718, new_AGEMA_signal_10717, MixColumnsIns_MixOneColumnInst_3_n51}), .c ({new_AGEMA_signal_11602, new_AGEMA_signal_11601, MixColumnsOutput[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U73 ( .a ({new_AGEMA_signal_10422, new_AGEMA_signal_10421, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .b ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .c ({new_AGEMA_signal_10718, new_AGEMA_signal_10717, MixColumnsIns_MixOneColumnInst_3_n51}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U72 ( .a ({new_AGEMA_signal_10282, new_AGEMA_signal_10281, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .b ({new_AGEMA_signal_10726, new_AGEMA_signal_10725, MixColumnsIns_MixOneColumnInst_3_n35}), .c ({new_AGEMA_signal_11148, new_AGEMA_signal_11147, MixColumnsIns_MixOneColumnInst_3_n36}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U71 ( .a ({new_AGEMA_signal_11604, new_AGEMA_signal_11603, MixColumnsIns_MixOneColumnInst_3_n34}), .b ({new_AGEMA_signal_11150, new_AGEMA_signal_11149, MixColumnsIns_MixOneColumnInst_3_n48}), .c ({new_AGEMA_signal_12070, new_AGEMA_signal_12069, MixColumnsOutput[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U70 ( .a ({new_AGEMA_signal_10424, new_AGEMA_signal_10423, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .b ({new_AGEMA_signal_10754, new_AGEMA_signal_10753, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]}), .c ({new_AGEMA_signal_11150, new_AGEMA_signal_11149, MixColumnsIns_MixOneColumnInst_3_n48}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U69 ( .a ({new_AGEMA_signal_10284, new_AGEMA_signal_10283, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .b ({new_AGEMA_signal_11164, new_AGEMA_signal_11163, MixColumnsIns_MixOneColumnInst_3_n33}), .c ({new_AGEMA_signal_11604, new_AGEMA_signal_11603, MixColumnsIns_MixOneColumnInst_3_n34}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U68 ( .a ({new_AGEMA_signal_11606, new_AGEMA_signal_11605, MixColumnsIns_MixOneColumnInst_3_n32}), .b ({new_AGEMA_signal_11152, new_AGEMA_signal_11151, MixColumnsIns_MixOneColumnInst_3_n45}), .c ({new_AGEMA_signal_12072, new_AGEMA_signal_12071, MixColumnsOutput[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U67 ( .a ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, MixColumnsInput[19]}), .b ({new_AGEMA_signal_10756, new_AGEMA_signal_10755, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]}), .c ({new_AGEMA_signal_11152, new_AGEMA_signal_11151, MixColumnsIns_MixOneColumnInst_3_n45}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U66 ( .a ({new_AGEMA_signal_10286, new_AGEMA_signal_10285, MixColumnsInput[3]}), .b ({new_AGEMA_signal_11170, new_AGEMA_signal_11169, MixColumnsIns_MixOneColumnInst_3_n31}), .c ({new_AGEMA_signal_11606, new_AGEMA_signal_11605, MixColumnsIns_MixOneColumnInst_3_n32}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U65 ( .a ({new_AGEMA_signal_11154, new_AGEMA_signal_11153, MixColumnsIns_MixOneColumnInst_3_n30}), .b ({new_AGEMA_signal_10720, new_AGEMA_signal_10719, MixColumnsIns_MixOneColumnInst_3_n38}), .c ({new_AGEMA_signal_11608, new_AGEMA_signal_11607, MixColumnsOutput[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U64 ( .a ({new_AGEMA_signal_10428, new_AGEMA_signal_10427, MixColumnsInput[18]}), .b ({new_AGEMA_signal_10276, new_AGEMA_signal_10275, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .c ({new_AGEMA_signal_10720, new_AGEMA_signal_10719, MixColumnsIns_MixOneColumnInst_3_n38}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U63 ( .a ({new_AGEMA_signal_10288, new_AGEMA_signal_10287, MixColumnsInput[2]}), .b ({new_AGEMA_signal_10728, new_AGEMA_signal_10727, MixColumnsIns_MixOneColumnInst_3_n29}), .c ({new_AGEMA_signal_11154, new_AGEMA_signal_11153, MixColumnsIns_MixOneColumnInst_3_n30}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U62 ( .a ({new_AGEMA_signal_11610, new_AGEMA_signal_11609, MixColumnsIns_MixOneColumnInst_3_n28}), .b ({new_AGEMA_signal_11166, new_AGEMA_signal_11165, MixColumnsIns_MixOneColumnInst_3_n27}), .c ({new_AGEMA_signal_12074, new_AGEMA_signal_12073, MixColumnsOutput[25]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U61 ( .a ({new_AGEMA_signal_10290, new_AGEMA_signal_10289, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .b ({new_AGEMA_signal_11174, new_AGEMA_signal_11173, MixColumnsIns_MixOneColumnInst_3_n26}), .c ({new_AGEMA_signal_11610, new_AGEMA_signal_11609, MixColumnsIns_MixOneColumnInst_3_n28}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U60 ( .a ({new_AGEMA_signal_11156, new_AGEMA_signal_11155, MixColumnsIns_MixOneColumnInst_3_n25}), .b ({new_AGEMA_signal_10730, new_AGEMA_signal_10729, MixColumnsIns_MixOneColumnInst_3_n24}), .c ({new_AGEMA_signal_11612, new_AGEMA_signal_11611, MixColumnsOutput[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U59 ( .a ({new_AGEMA_signal_10750, new_AGEMA_signal_10749, MixColumnsIns_MixOneColumnInst_3_n23}), .b ({new_AGEMA_signal_9914, new_AGEMA_signal_9913, MixColumnsInput[0]}), .c ({new_AGEMA_signal_11156, new_AGEMA_signal_11155, MixColumnsIns_MixOneColumnInst_3_n25}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U58 ( .a ({new_AGEMA_signal_11158, new_AGEMA_signal_11157, MixColumnsIns_MixOneColumnInst_3_n22}), .b ({new_AGEMA_signal_10722, new_AGEMA_signal_10721, MixColumnsIns_MixOneColumnInst_3_n42}), .c ({new_AGEMA_signal_11614, new_AGEMA_signal_11613, MixColumnsOutput[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U57 ( .a ({new_AGEMA_signal_10348, new_AGEMA_signal_10347, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .c ({new_AGEMA_signal_10722, new_AGEMA_signal_10721, MixColumnsIns_MixOneColumnInst_3_n42}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U56 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_10734, new_AGEMA_signal_10733, MixColumnsIns_MixOneColumnInst_3_n21}), .c ({new_AGEMA_signal_11158, new_AGEMA_signal_11157, MixColumnsIns_MixOneColumnInst_3_n22}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U55 ( .a ({new_AGEMA_signal_11160, new_AGEMA_signal_11159, MixColumnsIns_MixOneColumnInst_3_n20}), .b ({new_AGEMA_signal_10724, new_AGEMA_signal_10723, MixColumnsIns_MixOneColumnInst_3_n40}), .c ({new_AGEMA_signal_11616, new_AGEMA_signal_11615, MixColumnsOutput[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U54 ( .a ({new_AGEMA_signal_10350, new_AGEMA_signal_10349, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .b ({new_AGEMA_signal_10422, new_AGEMA_signal_10421, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .c ({new_AGEMA_signal_10724, new_AGEMA_signal_10723, MixColumnsIns_MixOneColumnInst_3_n40}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U53 ( .a ({new_AGEMA_signal_10266, new_AGEMA_signal_10265, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .b ({new_AGEMA_signal_10738, new_AGEMA_signal_10737, MixColumnsIns_MixOneColumnInst_3_n19}), .c ({new_AGEMA_signal_11160, new_AGEMA_signal_11159, MixColumnsIns_MixOneColumnInst_3_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U52 ( .a ({new_AGEMA_signal_11162, new_AGEMA_signal_11161, MixColumnsIns_MixOneColumnInst_3_n18}), .b ({new_AGEMA_signal_10726, new_AGEMA_signal_10725, MixColumnsIns_MixOneColumnInst_3_n35}), .c ({new_AGEMA_signal_11618, new_AGEMA_signal_11617, MixColumnsOutput[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U51 ( .a ({new_AGEMA_signal_10352, new_AGEMA_signal_10351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .b ({new_AGEMA_signal_10424, new_AGEMA_signal_10423, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .c ({new_AGEMA_signal_10726, new_AGEMA_signal_10725, MixColumnsIns_MixOneColumnInst_3_n35}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U50 ( .a ({new_AGEMA_signal_10268, new_AGEMA_signal_10267, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .b ({new_AGEMA_signal_10742, new_AGEMA_signal_10741, MixColumnsIns_MixOneColumnInst_3_n17}), .c ({new_AGEMA_signal_11162, new_AGEMA_signal_11161, MixColumnsIns_MixOneColumnInst_3_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U49 ( .a ({new_AGEMA_signal_11620, new_AGEMA_signal_11619, MixColumnsIns_MixOneColumnInst_3_n16}), .b ({new_AGEMA_signal_11164, new_AGEMA_signal_11163, MixColumnsIns_MixOneColumnInst_3_n33}), .c ({new_AGEMA_signal_12076, new_AGEMA_signal_12075, MixColumnsOutput[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U48 ( .a ({new_AGEMA_signal_10354, new_AGEMA_signal_10353, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .b ({new_AGEMA_signal_10760, new_AGEMA_signal_10759, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]}), .c ({new_AGEMA_signal_11164, new_AGEMA_signal_11163, MixColumnsIns_MixOneColumnInst_3_n33}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U47 ( .a ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .b ({new_AGEMA_signal_11186, new_AGEMA_signal_11185, MixColumnsIns_MixOneColumnInst_3_n15}), .c ({new_AGEMA_signal_11620, new_AGEMA_signal_11619, MixColumnsIns_MixOneColumnInst_3_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U46 ( .a ({new_AGEMA_signal_11622, new_AGEMA_signal_11621, MixColumnsIns_MixOneColumnInst_3_n14}), .b ({new_AGEMA_signal_11166, new_AGEMA_signal_11165, MixColumnsIns_MixOneColumnInst_3_n27}), .c ({new_AGEMA_signal_12078, new_AGEMA_signal_12077, MixColumnsOutput[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U45 ( .a ({new_AGEMA_signal_10430, new_AGEMA_signal_10429, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .b ({new_AGEMA_signal_10758, new_AGEMA_signal_10757, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]}), .c ({new_AGEMA_signal_11166, new_AGEMA_signal_11165, MixColumnsIns_MixOneColumnInst_3_n27}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U44 ( .a ({new_AGEMA_signal_10360, new_AGEMA_signal_10359, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .b ({new_AGEMA_signal_11168, new_AGEMA_signal_11167, MixColumnsIns_MixOneColumnInst_3_n62}), .c ({new_AGEMA_signal_11622, new_AGEMA_signal_11621, MixColumnsIns_MixOneColumnInst_3_n14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U43 ( .a ({new_AGEMA_signal_10276, new_AGEMA_signal_10275, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .b ({new_AGEMA_signal_10776, new_AGEMA_signal_10775, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]}), .c ({new_AGEMA_signal_11168, new_AGEMA_signal_11167, MixColumnsIns_MixOneColumnInst_3_n62}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U42 ( .a ({new_AGEMA_signal_11624, new_AGEMA_signal_11623, MixColumnsIns_MixOneColumnInst_3_n13}), .b ({new_AGEMA_signal_11170, new_AGEMA_signal_11169, MixColumnsIns_MixOneColumnInst_3_n31}), .c ({new_AGEMA_signal_12080, new_AGEMA_signal_12079, MixColumnsOutput[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U41 ( .a ({new_AGEMA_signal_10356, new_AGEMA_signal_10355, MixColumnsInput[11]}), .b ({new_AGEMA_signal_10762, new_AGEMA_signal_10761, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]}), .c ({new_AGEMA_signal_11170, new_AGEMA_signal_11169, MixColumnsIns_MixOneColumnInst_3_n31}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U40 ( .a ({new_AGEMA_signal_10272, new_AGEMA_signal_10271, MixColumnsInput[27]}), .b ({new_AGEMA_signal_11190, new_AGEMA_signal_11189, MixColumnsIns_MixOneColumnInst_3_n12}), .c ({new_AGEMA_signal_11624, new_AGEMA_signal_11623, MixColumnsIns_MixOneColumnInst_3_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U39 ( .a ({new_AGEMA_signal_11172, new_AGEMA_signal_11171, MixColumnsIns_MixOneColumnInst_3_n11}), .b ({new_AGEMA_signal_10728, new_AGEMA_signal_10727, MixColumnsIns_MixOneColumnInst_3_n29}), .c ({new_AGEMA_signal_11626, new_AGEMA_signal_11625, MixColumnsOutput[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U38 ( .a ({new_AGEMA_signal_10358, new_AGEMA_signal_10357, MixColumnsInput[10]}), .b ({new_AGEMA_signal_10430, new_AGEMA_signal_10429, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .c ({new_AGEMA_signal_10728, new_AGEMA_signal_10727, MixColumnsIns_MixOneColumnInst_3_n29}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U37 ( .a ({new_AGEMA_signal_10274, new_AGEMA_signal_10273, MixColumnsInput[26]}), .b ({new_AGEMA_signal_10746, new_AGEMA_signal_10745, MixColumnsIns_MixOneColumnInst_3_n10}), .c ({new_AGEMA_signal_11172, new_AGEMA_signal_11171, MixColumnsIns_MixOneColumnInst_3_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U36 ( .a ({new_AGEMA_signal_11628, new_AGEMA_signal_11627, MixColumnsIns_MixOneColumnInst_3_n9}), .b ({new_AGEMA_signal_11174, new_AGEMA_signal_11173, MixColumnsIns_MixOneColumnInst_3_n26}), .c ({new_AGEMA_signal_12082, new_AGEMA_signal_12081, MixColumnsOutput[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U35 ( .a ({new_AGEMA_signal_10764, new_AGEMA_signal_10763, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]}), .b ({new_AGEMA_signal_10360, new_AGEMA_signal_10359, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .c ({new_AGEMA_signal_11174, new_AGEMA_signal_11173, MixColumnsIns_MixOneColumnInst_3_n26}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U34 ( .a ({new_AGEMA_signal_11176, new_AGEMA_signal_11175, MixColumnsIns_MixOneColumnInst_3_n63}), .b ({new_AGEMA_signal_10276, new_AGEMA_signal_10275, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .c ({new_AGEMA_signal_11628, new_AGEMA_signal_11627, MixColumnsIns_MixOneColumnInst_3_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U33 ( .a ({new_AGEMA_signal_10770, new_AGEMA_signal_10769, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]}), .b ({new_AGEMA_signal_10290, new_AGEMA_signal_10289, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .c ({new_AGEMA_signal_11176, new_AGEMA_signal_11175, MixColumnsIns_MixOneColumnInst_3_n63}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U32 ( .a ({new_AGEMA_signal_11178, new_AGEMA_signal_11177, MixColumnsIns_MixOneColumnInst_3_n8}), .b ({new_AGEMA_signal_10730, new_AGEMA_signal_10729, MixColumnsIns_MixOneColumnInst_3_n24}), .c ({new_AGEMA_signal_11630, new_AGEMA_signal_11629, MixColumnsOutput[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U31 ( .a ({new_AGEMA_signal_10024, new_AGEMA_signal_10023, MixColumnsInput[8]}), .b ({new_AGEMA_signal_10418, new_AGEMA_signal_10417, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .c ({new_AGEMA_signal_10730, new_AGEMA_signal_10729, MixColumnsIns_MixOneColumnInst_3_n24}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U30 ( .a ({new_AGEMA_signal_9892, new_AGEMA_signal_9891, MixColumnsInput[24]}), .b ({new_AGEMA_signal_10732, new_AGEMA_signal_10731, MixColumnsIns_MixOneColumnInst_3_n60}), .c ({new_AGEMA_signal_11178, new_AGEMA_signal_11177, MixColumnsIns_MixOneColumnInst_3_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U29 ( .a ({new_AGEMA_signal_10348, new_AGEMA_signal_10347, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_9914, new_AGEMA_signal_9913, MixColumnsInput[0]}), .c ({new_AGEMA_signal_10732, new_AGEMA_signal_10731, MixColumnsIns_MixOneColumnInst_3_n60}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U28 ( .a ({new_AGEMA_signal_11180, new_AGEMA_signal_11179, MixColumnsIns_MixOneColumnInst_3_n7}), .b ({new_AGEMA_signal_10734, new_AGEMA_signal_10733, MixColumnsIns_MixOneColumnInst_3_n21}), .c ({new_AGEMA_signal_11632, new_AGEMA_signal_11631, MixColumnsOutput[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U27 ( .a ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_10350, new_AGEMA_signal_10349, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .c ({new_AGEMA_signal_10734, new_AGEMA_signal_10733, MixColumnsIns_MixOneColumnInst_3_n21}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U26 ( .a ({new_AGEMA_signal_10736, new_AGEMA_signal_10735, MixColumnsIns_MixOneColumnInst_3_n56}), .b ({new_AGEMA_signal_10418, new_AGEMA_signal_10417, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .c ({new_AGEMA_signal_11180, new_AGEMA_signal_11179, MixColumnsIns_MixOneColumnInst_3_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U25 ( .a ({new_AGEMA_signal_10280, new_AGEMA_signal_10279, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .b ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .c ({new_AGEMA_signal_10736, new_AGEMA_signal_10735, MixColumnsIns_MixOneColumnInst_3_n56}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U24 ( .a ({new_AGEMA_signal_11182, new_AGEMA_signal_11181, MixColumnsIns_MixOneColumnInst_3_n6}), .b ({new_AGEMA_signal_10738, new_AGEMA_signal_10737, MixColumnsIns_MixOneColumnInst_3_n19}), .c ({new_AGEMA_signal_11634, new_AGEMA_signal_11633, MixColumnsOutput[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U23 ( .a ({new_AGEMA_signal_10280, new_AGEMA_signal_10279, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .b ({new_AGEMA_signal_10352, new_AGEMA_signal_10351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .c ({new_AGEMA_signal_10738, new_AGEMA_signal_10737, MixColumnsIns_MixOneColumnInst_3_n19}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U22 ( .a ({new_AGEMA_signal_10740, new_AGEMA_signal_10739, MixColumnsIns_MixOneColumnInst_3_n53}), .b ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .c ({new_AGEMA_signal_11182, new_AGEMA_signal_11181, MixColumnsIns_MixOneColumnInst_3_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U21 ( .a ({new_AGEMA_signal_10282, new_AGEMA_signal_10281, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .b ({new_AGEMA_signal_10266, new_AGEMA_signal_10265, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .c ({new_AGEMA_signal_10740, new_AGEMA_signal_10739, MixColumnsIns_MixOneColumnInst_3_n53}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U20 ( .a ({new_AGEMA_signal_11184, new_AGEMA_signal_11183, MixColumnsIns_MixOneColumnInst_3_n5}), .b ({new_AGEMA_signal_10742, new_AGEMA_signal_10741, MixColumnsIns_MixOneColumnInst_3_n17}), .c ({new_AGEMA_signal_11636, new_AGEMA_signal_11635, MixColumnsOutput[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U19 ( .a ({new_AGEMA_signal_10282, new_AGEMA_signal_10281, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .b ({new_AGEMA_signal_10354, new_AGEMA_signal_10353, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .c ({new_AGEMA_signal_10742, new_AGEMA_signal_10741, MixColumnsIns_MixOneColumnInst_3_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U18 ( .a ({new_AGEMA_signal_10744, new_AGEMA_signal_10743, MixColumnsIns_MixOneColumnInst_3_n50}), .b ({new_AGEMA_signal_10422, new_AGEMA_signal_10421, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .c ({new_AGEMA_signal_11184, new_AGEMA_signal_11183, MixColumnsIns_MixOneColumnInst_3_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U17 ( .a ({new_AGEMA_signal_10284, new_AGEMA_signal_10283, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .b ({new_AGEMA_signal_10268, new_AGEMA_signal_10267, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .c ({new_AGEMA_signal_10744, new_AGEMA_signal_10743, MixColumnsIns_MixOneColumnInst_3_n50}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U16 ( .a ({new_AGEMA_signal_11638, new_AGEMA_signal_11637, MixColumnsIns_MixOneColumnInst_3_n4}), .b ({new_AGEMA_signal_11186, new_AGEMA_signal_11185, MixColumnsIns_MixOneColumnInst_3_n15}), .c ({new_AGEMA_signal_12084, new_AGEMA_signal_12083, MixColumnsOutput[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U15 ( .a ({new_AGEMA_signal_10284, new_AGEMA_signal_10283, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .b ({new_AGEMA_signal_10766, new_AGEMA_signal_10765, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]}), .c ({new_AGEMA_signal_11186, new_AGEMA_signal_11185, MixColumnsIns_MixOneColumnInst_3_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U14 ( .a ({new_AGEMA_signal_11188, new_AGEMA_signal_11187, MixColumnsIns_MixOneColumnInst_3_n47}), .b ({new_AGEMA_signal_10424, new_AGEMA_signal_10423, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .c ({new_AGEMA_signal_11638, new_AGEMA_signal_11637, MixColumnsIns_MixOneColumnInst_3_n4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U13 ( .a ({new_AGEMA_signal_10772, new_AGEMA_signal_10771, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]}), .b ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .c ({new_AGEMA_signal_11188, new_AGEMA_signal_11187, MixColumnsIns_MixOneColumnInst_3_n47}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U12 ( .a ({new_AGEMA_signal_11640, new_AGEMA_signal_11639, MixColumnsIns_MixOneColumnInst_3_n3}), .b ({new_AGEMA_signal_11190, new_AGEMA_signal_11189, MixColumnsIns_MixOneColumnInst_3_n12}), .c ({new_AGEMA_signal_12086, new_AGEMA_signal_12085, MixColumnsOutput[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U11 ( .a ({new_AGEMA_signal_10286, new_AGEMA_signal_10285, MixColumnsInput[3]}), .b ({new_AGEMA_signal_10768, new_AGEMA_signal_10767, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]}), .c ({new_AGEMA_signal_11190, new_AGEMA_signal_11189, MixColumnsIns_MixOneColumnInst_3_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U10 ( .a ({new_AGEMA_signal_11192, new_AGEMA_signal_11191, MixColumnsIns_MixOneColumnInst_3_n44}), .b ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, MixColumnsInput[19]}), .c ({new_AGEMA_signal_11640, new_AGEMA_signal_11639, MixColumnsIns_MixOneColumnInst_3_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U9 ( .a ({new_AGEMA_signal_10774, new_AGEMA_signal_10773, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]}), .b ({new_AGEMA_signal_10272, new_AGEMA_signal_10271, MixColumnsInput[27]}), .c ({new_AGEMA_signal_11192, new_AGEMA_signal_11191, MixColumnsIns_MixOneColumnInst_3_n44}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U8 ( .a ({new_AGEMA_signal_11194, new_AGEMA_signal_11193, MixColumnsIns_MixOneColumnInst_3_n2}), .b ({new_AGEMA_signal_10746, new_AGEMA_signal_10745, MixColumnsIns_MixOneColumnInst_3_n10}), .c ({new_AGEMA_signal_11642, new_AGEMA_signal_11641, MixColumnsOutput[10]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U7 ( .a ({new_AGEMA_signal_10288, new_AGEMA_signal_10287, MixColumnsInput[2]}), .b ({new_AGEMA_signal_10360, new_AGEMA_signal_10359, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .c ({new_AGEMA_signal_10746, new_AGEMA_signal_10745, MixColumnsIns_MixOneColumnInst_3_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U6 ( .a ({new_AGEMA_signal_10748, new_AGEMA_signal_10747, MixColumnsIns_MixOneColumnInst_3_n37}), .b ({new_AGEMA_signal_10428, new_AGEMA_signal_10427, MixColumnsInput[18]}), .c ({new_AGEMA_signal_11194, new_AGEMA_signal_11193, MixColumnsIns_MixOneColumnInst_3_n2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U5 ( .a ({new_AGEMA_signal_10290, new_AGEMA_signal_10289, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .b ({new_AGEMA_signal_10274, new_AGEMA_signal_10273, MixColumnsInput[26]}), .c ({new_AGEMA_signal_10748, new_AGEMA_signal_10747, MixColumnsIns_MixOneColumnInst_3_n37}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U4 ( .a ({new_AGEMA_signal_11196, new_AGEMA_signal_11195, MixColumnsIns_MixOneColumnInst_3_n1}), .b ({new_AGEMA_signal_10024, new_AGEMA_signal_10023, MixColumnsInput[8]}), .c ({new_AGEMA_signal_11644, new_AGEMA_signal_11643, MixColumnsOutput[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U3 ( .a ({new_AGEMA_signal_10752, new_AGEMA_signal_10751, MixColumnsIns_MixOneColumnInst_3_n59}), .b ({new_AGEMA_signal_10750, new_AGEMA_signal_10749, MixColumnsIns_MixOneColumnInst_3_n23}), .c ({new_AGEMA_signal_11196, new_AGEMA_signal_11195, MixColumnsIns_MixOneColumnInst_3_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U2 ( .a ({new_AGEMA_signal_10134, new_AGEMA_signal_10133, MixColumnsInput[16]}), .b ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .c ({new_AGEMA_signal_10750, new_AGEMA_signal_10749, MixColumnsIns_MixOneColumnInst_3_n23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U1 ( .a ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_9892, new_AGEMA_signal_9891, MixColumnsInput[24]}), .c ({new_AGEMA_signal_10752, new_AGEMA_signal_10751, MixColumnsIns_MixOneColumnInst_3_n59}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_10272, new_AGEMA_signal_10271, MixColumnsInput[27]}), .c ({new_AGEMA_signal_10754, new_AGEMA_signal_10753, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_10274, new_AGEMA_signal_10273, MixColumnsInput[26]}), .c ({new_AGEMA_signal_10756, new_AGEMA_signal_10755, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_9892, new_AGEMA_signal_9891, MixColumnsInput[24]}), .c ({new_AGEMA_signal_10758, new_AGEMA_signal_10757, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_10418, new_AGEMA_signal_10417, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, MixColumnsInput[19]}), .c ({new_AGEMA_signal_10760, new_AGEMA_signal_10759, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_10418, new_AGEMA_signal_10417, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_10428, new_AGEMA_signal_10427, MixColumnsInput[18]}), .c ({new_AGEMA_signal_10762, new_AGEMA_signal_10761, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_10418, new_AGEMA_signal_10417, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_10134, new_AGEMA_signal_10133, MixColumnsInput[16]}), .c ({new_AGEMA_signal_10764, new_AGEMA_signal_10763, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_10348, new_AGEMA_signal_10347, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_10356, new_AGEMA_signal_10355, MixColumnsInput[11]}), .c ({new_AGEMA_signal_10766, new_AGEMA_signal_10765, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_10348, new_AGEMA_signal_10347, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_10358, new_AGEMA_signal_10357, MixColumnsInput[10]}), .c ({new_AGEMA_signal_10768, new_AGEMA_signal_10767, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_10348, new_AGEMA_signal_10347, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_10024, new_AGEMA_signal_10023, MixColumnsInput[8]}), .c ({new_AGEMA_signal_10770, new_AGEMA_signal_10769, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_10286, new_AGEMA_signal_10285, MixColumnsInput[3]}), .c ({new_AGEMA_signal_10772, new_AGEMA_signal_10771, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_10288, new_AGEMA_signal_10287, MixColumnsInput[2]}), .c ({new_AGEMA_signal_10774, new_AGEMA_signal_10773, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_9914, new_AGEMA_signal_9913, MixColumnsInput[0]}), .c ({new_AGEMA_signal_10776, new_AGEMA_signal_10775, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11388, new_AGEMA_signal_11387, KeyExpansionOutput[0]}), .a ({key_s2[0], key_s1[0], key_s0[0]}), .c ({new_AGEMA_signal_11648, new_AGEMA_signal_11647, KeyReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11812, new_AGEMA_signal_11811, KeyExpansionOutput[1]}), .a ({key_s2[1], key_s1[1], key_s0[1]}), .c ({new_AGEMA_signal_12090, new_AGEMA_signal_12089, KeyReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11790, new_AGEMA_signal_11789, KeyExpansionOutput[2]}), .a ({key_s2[2], key_s1[2], key_s0[2]}), .c ({new_AGEMA_signal_12094, new_AGEMA_signal_12093, KeyReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11784, new_AGEMA_signal_11783, KeyExpansionOutput[3]}), .a ({key_s2[3], key_s1[3], key_s0[3]}), .c ({new_AGEMA_signal_12098, new_AGEMA_signal_12097, KeyReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11782, new_AGEMA_signal_11781, KeyExpansionOutput[4]}), .a ({key_s2[4], key_s1[4], key_s0[4]}), .c ({new_AGEMA_signal_12102, new_AGEMA_signal_12101, KeyReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11780, new_AGEMA_signal_11779, KeyExpansionOutput[5]}), .a ({key_s2[5], key_s1[5], key_s0[5]}), .c ({new_AGEMA_signal_12106, new_AGEMA_signal_12105, KeyReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11778, new_AGEMA_signal_11777, KeyExpansionOutput[6]}), .a ({key_s2[6], key_s1[6], key_s0[6]}), .c ({new_AGEMA_signal_12110, new_AGEMA_signal_12109, KeyReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11776, new_AGEMA_signal_11775, KeyExpansionOutput[7]}), .a ({key_s2[7], key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_12114, new_AGEMA_signal_12113, KeyReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11326, new_AGEMA_signal_11325, KeyExpansionOutput[8]}), .a ({key_s2[8], key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_11652, new_AGEMA_signal_11651, KeyReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11774, new_AGEMA_signal_11773, KeyExpansionOutput[9]}), .a ({key_s2[9], key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_12118, new_AGEMA_signal_12117, KeyReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11830, new_AGEMA_signal_11829, KeyExpansionOutput[10]}), .a ({key_s2[10], key_s1[10], key_s0[10]}), .c ({new_AGEMA_signal_12122, new_AGEMA_signal_12121, KeyReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11828, new_AGEMA_signal_11827, KeyExpansionOutput[11]}), .a ({key_s2[11], key_s1[11], key_s0[11]}), .c ({new_AGEMA_signal_12126, new_AGEMA_signal_12125, KeyReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11826, new_AGEMA_signal_11825, KeyExpansionOutput[12]}), .a ({key_s2[12], key_s1[12], key_s0[12]}), .c ({new_AGEMA_signal_12130, new_AGEMA_signal_12129, KeyReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11824, new_AGEMA_signal_11823, KeyExpansionOutput[13]}), .a ({key_s2[13], key_s1[13], key_s0[13]}), .c ({new_AGEMA_signal_12134, new_AGEMA_signal_12133, KeyReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11822, new_AGEMA_signal_11821, KeyExpansionOutput[14]}), .a ({key_s2[14], key_s1[14], key_s0[14]}), .c ({new_AGEMA_signal_12138, new_AGEMA_signal_12137, KeyReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11820, new_AGEMA_signal_11819, KeyExpansionOutput[15]}), .a ({key_s2[15], key_s1[15], key_s0[15]}), .c ({new_AGEMA_signal_12142, new_AGEMA_signal_12141, KeyReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11374, new_AGEMA_signal_11373, KeyExpansionOutput[16]}), .a ({key_s2[16], key_s1[16], key_s0[16]}), .c ({new_AGEMA_signal_11656, new_AGEMA_signal_11655, KeyReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11818, new_AGEMA_signal_11817, KeyExpansionOutput[17]}), .a ({key_s2[17], key_s1[17], key_s0[17]}), .c ({new_AGEMA_signal_12146, new_AGEMA_signal_12145, KeyReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11816, new_AGEMA_signal_11815, KeyExpansionOutput[18]}), .a ({key_s2[18], key_s1[18], key_s0[18]}), .c ({new_AGEMA_signal_12150, new_AGEMA_signal_12149, KeyReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11814, new_AGEMA_signal_11813, KeyExpansionOutput[19]}), .a ({key_s2[19], key_s1[19], key_s0[19]}), .c ({new_AGEMA_signal_12154, new_AGEMA_signal_12153, KeyReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11810, new_AGEMA_signal_11809, KeyExpansionOutput[20]}), .a ({key_s2[20], key_s1[20], key_s0[20]}), .c ({new_AGEMA_signal_12158, new_AGEMA_signal_12157, KeyReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11808, new_AGEMA_signal_11807, KeyExpansionOutput[21]}), .a ({key_s2[21], key_s1[21], key_s0[21]}), .c ({new_AGEMA_signal_12162, new_AGEMA_signal_12161, KeyReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11806, new_AGEMA_signal_11805, KeyExpansionOutput[22]}), .a ({key_s2[22], key_s1[22], key_s0[22]}), .c ({new_AGEMA_signal_12166, new_AGEMA_signal_12165, KeyReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11804, new_AGEMA_signal_11803, KeyExpansionOutput[23]}), .a ({key_s2[23], key_s1[23], key_s0[23]}), .c ({new_AGEMA_signal_12170, new_AGEMA_signal_12169, KeyReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11802, new_AGEMA_signal_11801, KeyExpansionOutput[24]}), .a ({key_s2[24], key_s1[24], key_s0[24]}), .c ({new_AGEMA_signal_12174, new_AGEMA_signal_12173, KeyReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12216, new_AGEMA_signal_12215, KeyExpansionOutput[25]}), .a ({key_s2[25], key_s1[25], key_s0[25]}), .c ({new_AGEMA_signal_12636, new_AGEMA_signal_12635, KeyReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12214, new_AGEMA_signal_12213, KeyExpansionOutput[26]}), .a ({key_s2[26], key_s1[26], key_s0[26]}), .c ({new_AGEMA_signal_12640, new_AGEMA_signal_12639, KeyReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12212, new_AGEMA_signal_12211, KeyExpansionOutput[27]}), .a ({key_s2[27], key_s1[27], key_s0[27]}), .c ({new_AGEMA_signal_12644, new_AGEMA_signal_12643, KeyReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12210, new_AGEMA_signal_12209, KeyExpansionOutput[28]}), .a ({key_s2[28], key_s1[28], key_s0[28]}), .c ({new_AGEMA_signal_12648, new_AGEMA_signal_12647, KeyReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12208, new_AGEMA_signal_12207, KeyExpansionOutput[29]}), .a ({key_s2[29], key_s1[29], key_s0[29]}), .c ({new_AGEMA_signal_12652, new_AGEMA_signal_12651, KeyReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12206, new_AGEMA_signal_12205, KeyExpansionOutput[30]}), .a ({key_s2[30], key_s1[30], key_s0[30]}), .c ({new_AGEMA_signal_12656, new_AGEMA_signal_12655, KeyReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12204, new_AGEMA_signal_12203, KeyExpansionOutput[31]}), .a ({key_s2[31], key_s1[31], key_s0[31]}), .c ({new_AGEMA_signal_12660, new_AGEMA_signal_12659, KeyReg_Inst_ff_SDE_31_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10940, new_AGEMA_signal_10939, KeyExpansionOutput[32]}), .a ({key_s2[32], key_s1[32], key_s0[32]}), .c ({new_AGEMA_signal_11200, new_AGEMA_signal_11199, KeyReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11366, new_AGEMA_signal_11365, KeyExpansionOutput[33]}), .a ({key_s2[33], key_s1[33], key_s0[33]}), .c ({new_AGEMA_signal_11660, new_AGEMA_signal_11659, KeyReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11344, new_AGEMA_signal_11343, KeyExpansionOutput[34]}), .a ({key_s2[34], key_s1[34], key_s0[34]}), .c ({new_AGEMA_signal_11664, new_AGEMA_signal_11663, KeyReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11338, new_AGEMA_signal_11337, KeyExpansionOutput[35]}), .a ({key_s2[35], key_s1[35], key_s0[35]}), .c ({new_AGEMA_signal_11668, new_AGEMA_signal_11667, KeyReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11336, new_AGEMA_signal_11335, KeyExpansionOutput[36]}), .a ({key_s2[36], key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_11672, new_AGEMA_signal_11671, KeyReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11334, new_AGEMA_signal_11333, KeyExpansionOutput[37]}), .a ({key_s2[37], key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_11676, new_AGEMA_signal_11675, KeyReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11332, new_AGEMA_signal_11331, KeyExpansionOutput[38]}), .a ({key_s2[38], key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_11680, new_AGEMA_signal_11679, KeyReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11330, new_AGEMA_signal_11329, KeyExpansionOutput[39]}), .a ({key_s2[39], key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_11684, new_AGEMA_signal_11683, KeyReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10880, new_AGEMA_signal_10879, KeyExpansionOutput[40]}), .a ({key_s2[40], key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_11204, new_AGEMA_signal_11203, KeyReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11328, new_AGEMA_signal_11327, KeyExpansionOutput[41]}), .a ({key_s2[41], key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_11688, new_AGEMA_signal_11687, KeyReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, KeyExpansionOutput[42]}), .a ({key_s2[42], key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_11692, new_AGEMA_signal_11691, KeyReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11384, new_AGEMA_signal_11383, KeyExpansionOutput[43]}), .a ({key_s2[43], key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_11696, new_AGEMA_signal_11695, KeyReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11382, new_AGEMA_signal_11381, KeyExpansionOutput[44]}), .a ({key_s2[44], key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_11700, new_AGEMA_signal_11699, KeyReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, KeyExpansionOutput[45]}), .a ({key_s2[45], key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_11704, new_AGEMA_signal_11703, KeyReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11378, new_AGEMA_signal_11377, KeyExpansionOutput[46]}), .a ({key_s2[46], key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_11708, new_AGEMA_signal_11707, KeyReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11376, new_AGEMA_signal_11375, KeyExpansionOutput[47]}), .a ({key_s2[47], key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_11712, new_AGEMA_signal_11711, KeyReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10912, new_AGEMA_signal_10911, KeyExpansionOutput[48]}), .a ({key_s2[48], key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_11208, new_AGEMA_signal_11207, KeyReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11372, new_AGEMA_signal_11371, KeyExpansionOutput[49]}), .a ({key_s2[49], key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_11716, new_AGEMA_signal_11715, KeyReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11370, new_AGEMA_signal_11369, KeyExpansionOutput[50]}), .a ({key_s2[50], key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_11720, new_AGEMA_signal_11719, KeyReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11368, new_AGEMA_signal_11367, KeyExpansionOutput[51]}), .a ({key_s2[51], key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_11724, new_AGEMA_signal_11723, KeyReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11364, new_AGEMA_signal_11363, KeyExpansionOutput[52]}), .a ({key_s2[52], key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_11728, new_AGEMA_signal_11727, KeyReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11362, new_AGEMA_signal_11361, KeyExpansionOutput[53]}), .a ({key_s2[53], key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_11732, new_AGEMA_signal_11731, KeyReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11360, new_AGEMA_signal_11359, KeyExpansionOutput[54]}), .a ({key_s2[54], key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_11736, new_AGEMA_signal_11735, KeyReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11358, new_AGEMA_signal_11357, KeyExpansionOutput[55]}), .a ({key_s2[55], key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_11740, new_AGEMA_signal_11739, KeyReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11356, new_AGEMA_signal_11355, KeyExpansionOutput[56]}), .a ({key_s2[56], key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_11744, new_AGEMA_signal_11743, KeyReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11800, new_AGEMA_signal_11799, KeyExpansionOutput[57]}), .a ({key_s2[57], key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_12178, new_AGEMA_signal_12177, KeyReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11798, new_AGEMA_signal_11797, KeyExpansionOutput[58]}), .a ({key_s2[58], key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_12182, new_AGEMA_signal_12181, KeyReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11796, new_AGEMA_signal_11795, KeyExpansionOutput[59]}), .a ({key_s2[59], key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_12186, new_AGEMA_signal_12185, KeyReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11794, new_AGEMA_signal_11793, KeyExpansionOutput[60]}), .a ({key_s2[60], key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_12190, new_AGEMA_signal_12189, KeyReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11792, new_AGEMA_signal_11791, KeyExpansionOutput[61]}), .a ({key_s2[61], key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_12194, new_AGEMA_signal_12193, KeyReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11788, new_AGEMA_signal_11787, KeyExpansionOutput[62]}), .a ({key_s2[62], key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_12198, new_AGEMA_signal_12197, KeyReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11786, new_AGEMA_signal_11785, KeyExpansionOutput[63]}), .a ({key_s2[63], key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_12202, new_AGEMA_signal_12201, KeyReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10506, new_AGEMA_signal_10505, KeyExpansionOutput[64]}), .a ({key_s2[64], key_s1[64], key_s0[64]}), .c ({new_AGEMA_signal_10780, new_AGEMA_signal_10779, KeyReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10904, new_AGEMA_signal_10903, KeyExpansionOutput[65]}), .a ({key_s2[65], key_s1[65], key_s0[65]}), .c ({new_AGEMA_signal_11212, new_AGEMA_signal_11211, KeyReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10892, new_AGEMA_signal_10891, KeyExpansionOutput[66]}), .a ({key_s2[66], key_s1[66], key_s0[66]}), .c ({new_AGEMA_signal_11216, new_AGEMA_signal_11215, KeyReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10890, new_AGEMA_signal_10889, KeyExpansionOutput[67]}), .a ({key_s2[67], key_s1[67], key_s0[67]}), .c ({new_AGEMA_signal_11220, new_AGEMA_signal_11219, KeyReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10888, new_AGEMA_signal_10887, KeyExpansionOutput[68]}), .a ({key_s2[68], key_s1[68], key_s0[68]}), .c ({new_AGEMA_signal_11224, new_AGEMA_signal_11223, KeyReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10886, new_AGEMA_signal_10885, KeyExpansionOutput[69]}), .a ({key_s2[69], key_s1[69], key_s0[69]}), .c ({new_AGEMA_signal_11228, new_AGEMA_signal_11227, KeyReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10884, new_AGEMA_signal_10883, KeyExpansionOutput[70]}), .a ({key_s2[70], key_s1[70], key_s0[70]}), .c ({new_AGEMA_signal_11232, new_AGEMA_signal_11231, KeyReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10882, new_AGEMA_signal_10881, KeyExpansionOutput[71]}), .a ({key_s2[71], key_s1[71], key_s0[71]}), .c ({new_AGEMA_signal_11236, new_AGEMA_signal_11235, KeyReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10458, new_AGEMA_signal_10457, KeyExpansionOutput[72]}), .a ({key_s2[72], key_s1[72], key_s0[72]}), .c ({new_AGEMA_signal_10784, new_AGEMA_signal_10783, KeyReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10878, new_AGEMA_signal_10877, KeyExpansionOutput[73]}), .a ({key_s2[73], key_s1[73], key_s0[73]}), .c ({new_AGEMA_signal_11240, new_AGEMA_signal_11239, KeyReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10938, new_AGEMA_signal_10937, KeyExpansionOutput[74]}), .a ({key_s2[74], key_s1[74], key_s0[74]}), .c ({new_AGEMA_signal_11244, new_AGEMA_signal_11243, KeyReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10936, new_AGEMA_signal_10935, KeyExpansionOutput[75]}), .a ({key_s2[75], key_s1[75], key_s0[75]}), .c ({new_AGEMA_signal_11248, new_AGEMA_signal_11247, KeyReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10920, new_AGEMA_signal_10919, KeyExpansionOutput[76]}), .a ({key_s2[76], key_s1[76], key_s0[76]}), .c ({new_AGEMA_signal_11252, new_AGEMA_signal_11251, KeyReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10918, new_AGEMA_signal_10917, KeyExpansionOutput[77]}), .a ({key_s2[77], key_s1[77], key_s0[77]}), .c ({new_AGEMA_signal_11256, new_AGEMA_signal_11255, KeyReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10916, new_AGEMA_signal_10915, KeyExpansionOutput[78]}), .a ({key_s2[78], key_s1[78], key_s0[78]}), .c ({new_AGEMA_signal_11260, new_AGEMA_signal_11259, KeyReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10914, new_AGEMA_signal_10913, KeyExpansionOutput[79]}), .a ({key_s2[79], key_s1[79], key_s0[79]}), .c ({new_AGEMA_signal_11264, new_AGEMA_signal_11263, KeyReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10466, new_AGEMA_signal_10465, KeyExpansionOutput[80]}), .a ({key_s2[80], key_s1[80], key_s0[80]}), .c ({new_AGEMA_signal_10788, new_AGEMA_signal_10787, KeyReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10910, new_AGEMA_signal_10909, KeyExpansionOutput[81]}), .a ({key_s2[81], key_s1[81], key_s0[81]}), .c ({new_AGEMA_signal_11268, new_AGEMA_signal_11267, KeyReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10908, new_AGEMA_signal_10907, KeyExpansionOutput[82]}), .a ({key_s2[82], key_s1[82], key_s0[82]}), .c ({new_AGEMA_signal_11272, new_AGEMA_signal_11271, KeyReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10906, new_AGEMA_signal_10905, KeyExpansionOutput[83]}), .a ({key_s2[83], key_s1[83], key_s0[83]}), .c ({new_AGEMA_signal_11276, new_AGEMA_signal_11275, KeyReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10902, new_AGEMA_signal_10901, KeyExpansionOutput[84]}), .a ({key_s2[84], key_s1[84], key_s0[84]}), .c ({new_AGEMA_signal_11280, new_AGEMA_signal_11279, KeyReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10900, new_AGEMA_signal_10899, KeyExpansionOutput[85]}), .a ({key_s2[85], key_s1[85], key_s0[85]}), .c ({new_AGEMA_signal_11284, new_AGEMA_signal_11283, KeyReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10898, new_AGEMA_signal_10897, KeyExpansionOutput[86]}), .a ({key_s2[86], key_s1[86], key_s0[86]}), .c ({new_AGEMA_signal_11288, new_AGEMA_signal_11287, KeyReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10896, new_AGEMA_signal_10895, KeyExpansionOutput[87]}), .a ({key_s2[87], key_s1[87], key_s0[87]}), .c ({new_AGEMA_signal_11292, new_AGEMA_signal_11291, KeyReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10894, new_AGEMA_signal_10893, KeyExpansionOutput[88]}), .a ({key_s2[88], key_s1[88], key_s0[88]}), .c ({new_AGEMA_signal_11296, new_AGEMA_signal_11295, KeyReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11354, new_AGEMA_signal_11353, KeyExpansionOutput[89]}), .a ({key_s2[89], key_s1[89], key_s0[89]}), .c ({new_AGEMA_signal_11748, new_AGEMA_signal_11747, KeyReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11352, new_AGEMA_signal_11351, KeyExpansionOutput[90]}), .a ({key_s2[90], key_s1[90], key_s0[90]}), .c ({new_AGEMA_signal_11752, new_AGEMA_signal_11751, KeyReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11350, new_AGEMA_signal_11349, KeyExpansionOutput[91]}), .a ({key_s2[91], key_s1[91], key_s0[91]}), .c ({new_AGEMA_signal_11756, new_AGEMA_signal_11755, KeyReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11348, new_AGEMA_signal_11347, KeyExpansionOutput[92]}), .a ({key_s2[92], key_s1[92], key_s0[92]}), .c ({new_AGEMA_signal_11760, new_AGEMA_signal_11759, KeyReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11346, new_AGEMA_signal_11345, KeyExpansionOutput[93]}), .a ({key_s2[93], key_s1[93], key_s0[93]}), .c ({new_AGEMA_signal_11764, new_AGEMA_signal_11763, KeyReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11342, new_AGEMA_signal_11341, KeyExpansionOutput[94]}), .a ({key_s2[94], key_s1[94], key_s0[94]}), .c ({new_AGEMA_signal_11768, new_AGEMA_signal_11767, KeyReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_11340, new_AGEMA_signal_11339, KeyExpansionOutput[95]}), .a ({key_s2[95], key_s1[95], key_s0[95]}), .c ({new_AGEMA_signal_11772, new_AGEMA_signal_11771, KeyReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10162, new_AGEMA_signal_10161, KeyExpansionOutput[96]}), .a ({key_s2[96], key_s1[96], key_s0[96]}), .c ({new_AGEMA_signal_10448, new_AGEMA_signal_10447, KeyReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10464, new_AGEMA_signal_10463, KeyExpansionOutput[97]}), .a ({key_s2[97], key_s1[97], key_s0[97]}), .c ({new_AGEMA_signal_10792, new_AGEMA_signal_10791, KeyReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, KeyExpansionOutput[98]}), .a ({key_s2[98], key_s1[98], key_s0[98]}), .c ({new_AGEMA_signal_10796, new_AGEMA_signal_10795, KeyReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10460, new_AGEMA_signal_10459, KeyExpansionOutput[99]}), .a ({key_s2[99], key_s1[99], key_s0[99]}), .c ({new_AGEMA_signal_10800, new_AGEMA_signal_10799, KeyReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10504, new_AGEMA_signal_10503, KeyExpansionOutput[100]}), .a ({key_s2[100], key_s1[100], key_s0[100]}), .c ({new_AGEMA_signal_10804, new_AGEMA_signal_10803, KeyReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10502, new_AGEMA_signal_10501, KeyExpansionOutput[101]}), .a ({key_s2[101], key_s1[101], key_s0[101]}), .c ({new_AGEMA_signal_10808, new_AGEMA_signal_10807, KeyReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10500, new_AGEMA_signal_10499, KeyExpansionOutput[102]}), .a ({key_s2[102], key_s1[102], key_s0[102]}), .c ({new_AGEMA_signal_10812, new_AGEMA_signal_10811, KeyReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10498, new_AGEMA_signal_10497, KeyExpansionOutput[103]}), .a ({key_s2[103], key_s1[103], key_s0[103]}), .c ({new_AGEMA_signal_10816, new_AGEMA_signal_10815, KeyReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10160, new_AGEMA_signal_10159, KeyExpansionOutput[104]}), .a ({key_s2[104], key_s1[104], key_s0[104]}), .c ({new_AGEMA_signal_10452, new_AGEMA_signal_10451, KeyReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10496, new_AGEMA_signal_10495, KeyExpansionOutput[105]}), .a ({key_s2[105], key_s1[105], key_s0[105]}), .c ({new_AGEMA_signal_10820, new_AGEMA_signal_10819, KeyReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10494, new_AGEMA_signal_10493, KeyExpansionOutput[106]}), .a ({key_s2[106], key_s1[106], key_s0[106]}), .c ({new_AGEMA_signal_10824, new_AGEMA_signal_10823, KeyReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10492, new_AGEMA_signal_10491, KeyExpansionOutput[107]}), .a ({key_s2[107], key_s1[107], key_s0[107]}), .c ({new_AGEMA_signal_10828, new_AGEMA_signal_10827, KeyReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10490, new_AGEMA_signal_10489, KeyExpansionOutput[108]}), .a ({key_s2[108], key_s1[108], key_s0[108]}), .c ({new_AGEMA_signal_10832, new_AGEMA_signal_10831, KeyReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10488, new_AGEMA_signal_10487, KeyExpansionOutput[109]}), .a ({key_s2[109], key_s1[109], key_s0[109]}), .c ({new_AGEMA_signal_10836, new_AGEMA_signal_10835, KeyReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10486, new_AGEMA_signal_10485, KeyExpansionOutput[110]}), .a ({key_s2[110], key_s1[110], key_s0[110]}), .c ({new_AGEMA_signal_10840, new_AGEMA_signal_10839, KeyReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10484, new_AGEMA_signal_10483, KeyExpansionOutput[111]}), .a ({key_s2[111], key_s1[111], key_s0[111]}), .c ({new_AGEMA_signal_10844, new_AGEMA_signal_10843, KeyReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10158, new_AGEMA_signal_10157, KeyExpansionOutput[112]}), .a ({key_s2[112], key_s1[112], key_s0[112]}), .c ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, KeyReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10482, new_AGEMA_signal_10481, KeyExpansionOutput[113]}), .a ({key_s2[113], key_s1[113], key_s0[113]}), .c ({new_AGEMA_signal_10848, new_AGEMA_signal_10847, KeyReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10480, new_AGEMA_signal_10479, KeyExpansionOutput[114]}), .a ({key_s2[114], key_s1[114], key_s0[114]}), .c ({new_AGEMA_signal_10852, new_AGEMA_signal_10851, KeyReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10478, new_AGEMA_signal_10477, KeyExpansionOutput[115]}), .a ({key_s2[115], key_s1[115], key_s0[115]}), .c ({new_AGEMA_signal_10856, new_AGEMA_signal_10855, KeyReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10476, new_AGEMA_signal_10475, KeyExpansionOutput[116]}), .a ({key_s2[116], key_s1[116], key_s0[116]}), .c ({new_AGEMA_signal_10860, new_AGEMA_signal_10859, KeyReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10474, new_AGEMA_signal_10473, KeyExpansionOutput[117]}), .a ({key_s2[117], key_s1[117], key_s0[117]}), .c ({new_AGEMA_signal_10864, new_AGEMA_signal_10863, KeyReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10472, new_AGEMA_signal_10471, KeyExpansionOutput[118]}), .a ({key_s2[118], key_s1[118], key_s0[118]}), .c ({new_AGEMA_signal_10868, new_AGEMA_signal_10867, KeyReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10470, new_AGEMA_signal_10469, KeyExpansionOutput[119]}), .a ({key_s2[119], key_s1[119], key_s0[119]}), .c ({new_AGEMA_signal_10872, new_AGEMA_signal_10871, KeyReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, KeyExpansionOutput[120]}), .a ({key_s2[120], key_s1[120], key_s0[120]}), .c ({new_AGEMA_signal_10876, new_AGEMA_signal_10875, KeyReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10934, new_AGEMA_signal_10933, KeyExpansionOutput[121]}), .a ({key_s2[121], key_s1[121], key_s0[121]}), .c ({new_AGEMA_signal_11300, new_AGEMA_signal_11299, KeyReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10932, new_AGEMA_signal_10931, KeyExpansionOutput[122]}), .a ({key_s2[122], key_s1[122], key_s0[122]}), .c ({new_AGEMA_signal_11304, new_AGEMA_signal_11303, KeyReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10930, new_AGEMA_signal_10929, KeyExpansionOutput[123]}), .a ({key_s2[123], key_s1[123], key_s0[123]}), .c ({new_AGEMA_signal_11308, new_AGEMA_signal_11307, KeyReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10928, new_AGEMA_signal_10927, KeyExpansionOutput[124]}), .a ({key_s2[124], key_s1[124], key_s0[124]}), .c ({new_AGEMA_signal_11312, new_AGEMA_signal_11311, KeyReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10926, new_AGEMA_signal_10925, KeyExpansionOutput[125]}), .a ({key_s2[125], key_s1[125], key_s0[125]}), .c ({new_AGEMA_signal_11316, new_AGEMA_signal_11315, KeyReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10924, new_AGEMA_signal_10923, KeyExpansionOutput[126]}), .a ({key_s2[126], key_s1[126], key_s0[126]}), .c ({new_AGEMA_signal_11320, new_AGEMA_signal_11319, KeyReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_10922, new_AGEMA_signal_10921, KeyExpansionOutput[127]}), .a ({key_s2[127], key_s1[127], key_s0[127]}), .c ({new_AGEMA_signal_11324, new_AGEMA_signal_11323, KeyReg_Inst_ff_SDE_127_next_state}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U128 ( .a ({new_AGEMA_signal_5314, new_AGEMA_signal_5313, RoundKey[9]}), .b ({new_AGEMA_signal_11328, new_AGEMA_signal_11327, KeyExpansionOutput[41]}), .c ({new_AGEMA_signal_11774, new_AGEMA_signal_11773, KeyExpansionOutput[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U127 ( .a ({new_AGEMA_signal_5248, new_AGEMA_signal_5247, RoundKey[8]}), .b ({new_AGEMA_signal_10880, new_AGEMA_signal_10879, KeyExpansionOutput[40]}), .c ({new_AGEMA_signal_11326, new_AGEMA_signal_11325, KeyExpansionOutput[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U126 ( .a ({new_AGEMA_signal_5182, new_AGEMA_signal_5181, RoundKey[7]}), .b ({new_AGEMA_signal_11330, new_AGEMA_signal_11329, KeyExpansionOutput[39]}), .c ({new_AGEMA_signal_11776, new_AGEMA_signal_11775, KeyExpansionOutput[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U125 ( .a ({new_AGEMA_signal_5116, new_AGEMA_signal_5115, RoundKey[6]}), .b ({new_AGEMA_signal_11332, new_AGEMA_signal_11331, KeyExpansionOutput[38]}), .c ({new_AGEMA_signal_11778, new_AGEMA_signal_11777, KeyExpansionOutput[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U124 ( .a ({new_AGEMA_signal_5050, new_AGEMA_signal_5049, RoundKey[5]}), .b ({new_AGEMA_signal_11334, new_AGEMA_signal_11333, KeyExpansionOutput[37]}), .c ({new_AGEMA_signal_11780, new_AGEMA_signal_11779, KeyExpansionOutput[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U123 ( .a ({new_AGEMA_signal_4984, new_AGEMA_signal_4983, RoundKey[4]}), .b ({new_AGEMA_signal_11336, new_AGEMA_signal_11335, KeyExpansionOutput[36]}), .c ({new_AGEMA_signal_11782, new_AGEMA_signal_11781, KeyExpansionOutput[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U122 ( .a ({new_AGEMA_signal_4930, new_AGEMA_signal_4929, RoundKey[41]}), .b ({new_AGEMA_signal_10878, new_AGEMA_signal_10877, KeyExpansionOutput[73]}), .c ({new_AGEMA_signal_11328, new_AGEMA_signal_11327, KeyExpansionOutput[41]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U121 ( .a ({new_AGEMA_signal_5140, new_AGEMA_signal_5139, RoundKey[73]}), .b ({new_AGEMA_signal_10496, new_AGEMA_signal_10495, KeyExpansionOutput[105]}), .c ({new_AGEMA_signal_10878, new_AGEMA_signal_10877, KeyExpansionOutput[73]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U120 ( .a ({new_AGEMA_signal_4924, new_AGEMA_signal_4923, RoundKey[40]}), .b ({new_AGEMA_signal_10458, new_AGEMA_signal_10457, KeyExpansionOutput[72]}), .c ({new_AGEMA_signal_10880, new_AGEMA_signal_10879, KeyExpansionOutput[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U119 ( .a ({new_AGEMA_signal_5134, new_AGEMA_signal_5133, RoundKey[72]}), .b ({new_AGEMA_signal_10160, new_AGEMA_signal_10159, KeyExpansionOutput[104]}), .c ({new_AGEMA_signal_10458, new_AGEMA_signal_10457, KeyExpansionOutput[72]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U118 ( .a ({new_AGEMA_signal_4918, new_AGEMA_signal_4917, RoundKey[3]}), .b ({new_AGEMA_signal_11338, new_AGEMA_signal_11337, KeyExpansionOutput[35]}), .c ({new_AGEMA_signal_11784, new_AGEMA_signal_11783, KeyExpansionOutput[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U117 ( .a ({new_AGEMA_signal_4912, new_AGEMA_signal_4911, RoundKey[39]}), .b ({new_AGEMA_signal_10882, new_AGEMA_signal_10881, KeyExpansionOutput[71]}), .c ({new_AGEMA_signal_11330, new_AGEMA_signal_11329, KeyExpansionOutput[39]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U116 ( .a ({new_AGEMA_signal_5128, new_AGEMA_signal_5127, RoundKey[71]}), .b ({new_AGEMA_signal_10498, new_AGEMA_signal_10497, KeyExpansionOutput[103]}), .c ({new_AGEMA_signal_10882, new_AGEMA_signal_10881, KeyExpansionOutput[71]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U115 ( .a ({new_AGEMA_signal_4906, new_AGEMA_signal_4905, RoundKey[38]}), .b ({new_AGEMA_signal_10884, new_AGEMA_signal_10883, KeyExpansionOutput[70]}), .c ({new_AGEMA_signal_11332, new_AGEMA_signal_11331, KeyExpansionOutput[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U114 ( .a ({new_AGEMA_signal_5122, new_AGEMA_signal_5121, RoundKey[70]}), .b ({new_AGEMA_signal_10500, new_AGEMA_signal_10499, KeyExpansionOutput[102]}), .c ({new_AGEMA_signal_10884, new_AGEMA_signal_10883, KeyExpansionOutput[70]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U113 ( .a ({new_AGEMA_signal_4900, new_AGEMA_signal_4899, RoundKey[37]}), .b ({new_AGEMA_signal_10886, new_AGEMA_signal_10885, KeyExpansionOutput[69]}), .c ({new_AGEMA_signal_11334, new_AGEMA_signal_11333, KeyExpansionOutput[37]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U112 ( .a ({new_AGEMA_signal_5110, new_AGEMA_signal_5109, RoundKey[69]}), .b ({new_AGEMA_signal_10502, new_AGEMA_signal_10501, KeyExpansionOutput[101]}), .c ({new_AGEMA_signal_10886, new_AGEMA_signal_10885, KeyExpansionOutput[69]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U111 ( .a ({new_AGEMA_signal_4894, new_AGEMA_signal_4893, RoundKey[36]}), .b ({new_AGEMA_signal_10888, new_AGEMA_signal_10887, KeyExpansionOutput[68]}), .c ({new_AGEMA_signal_11336, new_AGEMA_signal_11335, KeyExpansionOutput[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U110 ( .a ({new_AGEMA_signal_5104, new_AGEMA_signal_5103, RoundKey[68]}), .b ({new_AGEMA_signal_10504, new_AGEMA_signal_10503, KeyExpansionOutput[100]}), .c ({new_AGEMA_signal_10888, new_AGEMA_signal_10887, KeyExpansionOutput[68]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U109 ( .a ({new_AGEMA_signal_4888, new_AGEMA_signal_4887, RoundKey[35]}), .b ({new_AGEMA_signal_10890, new_AGEMA_signal_10889, KeyExpansionOutput[67]}), .c ({new_AGEMA_signal_11338, new_AGEMA_signal_11337, KeyExpansionOutput[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U108 ( .a ({new_AGEMA_signal_5098, new_AGEMA_signal_5097, RoundKey[67]}), .b ({new_AGEMA_signal_10460, new_AGEMA_signal_10459, KeyExpansionOutput[99]}), .c ({new_AGEMA_signal_10890, new_AGEMA_signal_10889, KeyExpansionOutput[67]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U107 ( .a ({new_AGEMA_signal_5308, new_AGEMA_signal_5307, RoundKey[99]}), .b ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_10460, new_AGEMA_signal_10459, KeyExpansionOutput[99]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U106 ( .a ({new_AGEMA_signal_4864, new_AGEMA_signal_4863, RoundKey[31]}), .b ({new_AGEMA_signal_11786, new_AGEMA_signal_11785, KeyExpansionOutput[63]}), .c ({new_AGEMA_signal_12204, new_AGEMA_signal_12203, KeyExpansionOutput[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U105 ( .a ({new_AGEMA_signal_5074, new_AGEMA_signal_5073, RoundKey[63]}), .b ({new_AGEMA_signal_11340, new_AGEMA_signal_11339, KeyExpansionOutput[95]}), .c ({new_AGEMA_signal_11786, new_AGEMA_signal_11785, KeyExpansionOutput[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U104 ( .a ({new_AGEMA_signal_5284, new_AGEMA_signal_5283, RoundKey[95]}), .b ({new_AGEMA_signal_10922, new_AGEMA_signal_10921, KeyExpansionOutput[127]}), .c ({new_AGEMA_signal_11340, new_AGEMA_signal_11339, KeyExpansionOutput[95]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U103 ( .a ({new_AGEMA_signal_4858, new_AGEMA_signal_4857, RoundKey[30]}), .b ({new_AGEMA_signal_11788, new_AGEMA_signal_11787, KeyExpansionOutput[62]}), .c ({new_AGEMA_signal_12206, new_AGEMA_signal_12205, KeyExpansionOutput[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U102 ( .a ({new_AGEMA_signal_5068, new_AGEMA_signal_5067, RoundKey[62]}), .b ({new_AGEMA_signal_11342, new_AGEMA_signal_11341, KeyExpansionOutput[94]}), .c ({new_AGEMA_signal_11788, new_AGEMA_signal_11787, KeyExpansionOutput[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U101 ( .a ({new_AGEMA_signal_5278, new_AGEMA_signal_5277, RoundKey[94]}), .b ({new_AGEMA_signal_10924, new_AGEMA_signal_10923, KeyExpansionOutput[126]}), .c ({new_AGEMA_signal_11342, new_AGEMA_signal_11341, KeyExpansionOutput[94]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U100 ( .a ({new_AGEMA_signal_4852, new_AGEMA_signal_4851, RoundKey[2]}), .b ({new_AGEMA_signal_11344, new_AGEMA_signal_11343, KeyExpansionOutput[34]}), .c ({new_AGEMA_signal_11790, new_AGEMA_signal_11789, KeyExpansionOutput[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U99 ( .a ({new_AGEMA_signal_4882, new_AGEMA_signal_4881, RoundKey[34]}), .b ({new_AGEMA_signal_10892, new_AGEMA_signal_10891, KeyExpansionOutput[66]}), .c ({new_AGEMA_signal_11344, new_AGEMA_signal_11343, KeyExpansionOutput[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U98 ( .a ({new_AGEMA_signal_5092, new_AGEMA_signal_5091, RoundKey[66]}), .b ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, KeyExpansionOutput[98]}), .c ({new_AGEMA_signal_10892, new_AGEMA_signal_10891, KeyExpansionOutput[66]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U97 ( .a ({new_AGEMA_signal_5302, new_AGEMA_signal_5301, RoundKey[98]}), .b ({new_AGEMA_signal_10218, new_AGEMA_signal_10217, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, KeyExpansionOutput[98]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U96 ( .a ({new_AGEMA_signal_4846, new_AGEMA_signal_4845, RoundKey[29]}), .b ({new_AGEMA_signal_11792, new_AGEMA_signal_11791, KeyExpansionOutput[61]}), .c ({new_AGEMA_signal_12208, new_AGEMA_signal_12207, KeyExpansionOutput[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U95 ( .a ({new_AGEMA_signal_5062, new_AGEMA_signal_5061, RoundKey[61]}), .b ({new_AGEMA_signal_11346, new_AGEMA_signal_11345, KeyExpansionOutput[93]}), .c ({new_AGEMA_signal_11792, new_AGEMA_signal_11791, KeyExpansionOutput[61]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U94 ( .a ({new_AGEMA_signal_5272, new_AGEMA_signal_5271, RoundKey[93]}), .b ({new_AGEMA_signal_10926, new_AGEMA_signal_10925, KeyExpansionOutput[125]}), .c ({new_AGEMA_signal_11346, new_AGEMA_signal_11345, KeyExpansionOutput[93]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U93 ( .a ({new_AGEMA_signal_4840, new_AGEMA_signal_4839, RoundKey[28]}), .b ({new_AGEMA_signal_11794, new_AGEMA_signal_11793, KeyExpansionOutput[60]}), .c ({new_AGEMA_signal_12210, new_AGEMA_signal_12209, KeyExpansionOutput[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U92 ( .a ({new_AGEMA_signal_5056, new_AGEMA_signal_5055, RoundKey[60]}), .b ({new_AGEMA_signal_11348, new_AGEMA_signal_11347, KeyExpansionOutput[92]}), .c ({new_AGEMA_signal_11794, new_AGEMA_signal_11793, KeyExpansionOutput[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U91 ( .a ({new_AGEMA_signal_5266, new_AGEMA_signal_5265, RoundKey[92]}), .b ({new_AGEMA_signal_10928, new_AGEMA_signal_10927, KeyExpansionOutput[124]}), .c ({new_AGEMA_signal_11348, new_AGEMA_signal_11347, KeyExpansionOutput[92]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U90 ( .a ({new_AGEMA_signal_4834, new_AGEMA_signal_4833, RoundKey[27]}), .b ({new_AGEMA_signal_11796, new_AGEMA_signal_11795, KeyExpansionOutput[59]}), .c ({new_AGEMA_signal_12212, new_AGEMA_signal_12211, KeyExpansionOutput[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U89 ( .a ({new_AGEMA_signal_5044, new_AGEMA_signal_5043, RoundKey[59]}), .b ({new_AGEMA_signal_11350, new_AGEMA_signal_11349, KeyExpansionOutput[91]}), .c ({new_AGEMA_signal_11796, new_AGEMA_signal_11795, KeyExpansionOutput[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U88 ( .a ({new_AGEMA_signal_5260, new_AGEMA_signal_5259, RoundKey[91]}), .b ({new_AGEMA_signal_10930, new_AGEMA_signal_10929, KeyExpansionOutput[123]}), .c ({new_AGEMA_signal_11350, new_AGEMA_signal_11349, KeyExpansionOutput[91]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U87 ( .a ({new_AGEMA_signal_4828, new_AGEMA_signal_4827, RoundKey[26]}), .b ({new_AGEMA_signal_11798, new_AGEMA_signal_11797, KeyExpansionOutput[58]}), .c ({new_AGEMA_signal_12214, new_AGEMA_signal_12213, KeyExpansionOutput[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U86 ( .a ({new_AGEMA_signal_5038, new_AGEMA_signal_5037, RoundKey[58]}), .b ({new_AGEMA_signal_11352, new_AGEMA_signal_11351, KeyExpansionOutput[90]}), .c ({new_AGEMA_signal_11798, new_AGEMA_signal_11797, KeyExpansionOutput[58]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U85 ( .a ({new_AGEMA_signal_5254, new_AGEMA_signal_5253, RoundKey[90]}), .b ({new_AGEMA_signal_10932, new_AGEMA_signal_10931, KeyExpansionOutput[122]}), .c ({new_AGEMA_signal_11352, new_AGEMA_signal_11351, KeyExpansionOutput[90]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U84 ( .a ({new_AGEMA_signal_4822, new_AGEMA_signal_4821, RoundKey[25]}), .b ({new_AGEMA_signal_11800, new_AGEMA_signal_11799, KeyExpansionOutput[57]}), .c ({new_AGEMA_signal_12216, new_AGEMA_signal_12215, KeyExpansionOutput[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U83 ( .a ({new_AGEMA_signal_5032, new_AGEMA_signal_5031, RoundKey[57]}), .b ({new_AGEMA_signal_11354, new_AGEMA_signal_11353, KeyExpansionOutput[89]}), .c ({new_AGEMA_signal_11800, new_AGEMA_signal_11799, KeyExpansionOutput[57]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U82 ( .a ({new_AGEMA_signal_5242, new_AGEMA_signal_5241, RoundKey[89]}), .b ({new_AGEMA_signal_10934, new_AGEMA_signal_10933, KeyExpansionOutput[121]}), .c ({new_AGEMA_signal_11354, new_AGEMA_signal_11353, KeyExpansionOutput[89]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U81 ( .a ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, RoundKey[24]}), .b ({new_AGEMA_signal_11356, new_AGEMA_signal_11355, KeyExpansionOutput[56]}), .c ({new_AGEMA_signal_11802, new_AGEMA_signal_11801, KeyExpansionOutput[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U80 ( .a ({new_AGEMA_signal_5026, new_AGEMA_signal_5025, RoundKey[56]}), .b ({new_AGEMA_signal_10894, new_AGEMA_signal_10893, KeyExpansionOutput[88]}), .c ({new_AGEMA_signal_11356, new_AGEMA_signal_11355, KeyExpansionOutput[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U79 ( .a ({new_AGEMA_signal_5236, new_AGEMA_signal_5235, RoundKey[88]}), .b ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, KeyExpansionOutput[120]}), .c ({new_AGEMA_signal_10894, new_AGEMA_signal_10893, KeyExpansionOutput[88]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U78 ( .a ({new_AGEMA_signal_4810, new_AGEMA_signal_4809, RoundKey[23]}), .b ({new_AGEMA_signal_11358, new_AGEMA_signal_11357, KeyExpansionOutput[55]}), .c ({new_AGEMA_signal_11804, new_AGEMA_signal_11803, KeyExpansionOutput[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U77 ( .a ({new_AGEMA_signal_5020, new_AGEMA_signal_5019, RoundKey[55]}), .b ({new_AGEMA_signal_10896, new_AGEMA_signal_10895, KeyExpansionOutput[87]}), .c ({new_AGEMA_signal_11358, new_AGEMA_signal_11357, KeyExpansionOutput[55]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U76 ( .a ({new_AGEMA_signal_5230, new_AGEMA_signal_5229, RoundKey[87]}), .b ({new_AGEMA_signal_10470, new_AGEMA_signal_10469, KeyExpansionOutput[119]}), .c ({new_AGEMA_signal_10896, new_AGEMA_signal_10895, KeyExpansionOutput[87]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U75 ( .a ({new_AGEMA_signal_4804, new_AGEMA_signal_4803, RoundKey[22]}), .b ({new_AGEMA_signal_11360, new_AGEMA_signal_11359, KeyExpansionOutput[54]}), .c ({new_AGEMA_signal_11806, new_AGEMA_signal_11805, KeyExpansionOutput[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U74 ( .a ({new_AGEMA_signal_5014, new_AGEMA_signal_5013, RoundKey[54]}), .b ({new_AGEMA_signal_10898, new_AGEMA_signal_10897, KeyExpansionOutput[86]}), .c ({new_AGEMA_signal_11360, new_AGEMA_signal_11359, KeyExpansionOutput[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U73 ( .a ({new_AGEMA_signal_5224, new_AGEMA_signal_5223, RoundKey[86]}), .b ({new_AGEMA_signal_10472, new_AGEMA_signal_10471, KeyExpansionOutput[118]}), .c ({new_AGEMA_signal_10898, new_AGEMA_signal_10897, KeyExpansionOutput[86]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U72 ( .a ({new_AGEMA_signal_4798, new_AGEMA_signal_4797, RoundKey[21]}), .b ({new_AGEMA_signal_11362, new_AGEMA_signal_11361, KeyExpansionOutput[53]}), .c ({new_AGEMA_signal_11808, new_AGEMA_signal_11807, KeyExpansionOutput[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U71 ( .a ({new_AGEMA_signal_5008, new_AGEMA_signal_5007, RoundKey[53]}), .b ({new_AGEMA_signal_10900, new_AGEMA_signal_10899, KeyExpansionOutput[85]}), .c ({new_AGEMA_signal_11362, new_AGEMA_signal_11361, KeyExpansionOutput[53]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U70 ( .a ({new_AGEMA_signal_5218, new_AGEMA_signal_5217, RoundKey[85]}), .b ({new_AGEMA_signal_10474, new_AGEMA_signal_10473, KeyExpansionOutput[117]}), .c ({new_AGEMA_signal_10900, new_AGEMA_signal_10899, KeyExpansionOutput[85]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U69 ( .a ({new_AGEMA_signal_4792, new_AGEMA_signal_4791, RoundKey[20]}), .b ({new_AGEMA_signal_11364, new_AGEMA_signal_11363, KeyExpansionOutput[52]}), .c ({new_AGEMA_signal_11810, new_AGEMA_signal_11809, KeyExpansionOutput[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U68 ( .a ({new_AGEMA_signal_5002, new_AGEMA_signal_5001, RoundKey[52]}), .b ({new_AGEMA_signal_10902, new_AGEMA_signal_10901, KeyExpansionOutput[84]}), .c ({new_AGEMA_signal_11364, new_AGEMA_signal_11363, KeyExpansionOutput[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U67 ( .a ({new_AGEMA_signal_5212, new_AGEMA_signal_5211, RoundKey[84]}), .b ({new_AGEMA_signal_10476, new_AGEMA_signal_10475, KeyExpansionOutput[116]}), .c ({new_AGEMA_signal_10902, new_AGEMA_signal_10901, KeyExpansionOutput[84]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U66 ( .a ({new_AGEMA_signal_4786, new_AGEMA_signal_4785, RoundKey[1]}), .b ({new_AGEMA_signal_11366, new_AGEMA_signal_11365, KeyExpansionOutput[33]}), .c ({new_AGEMA_signal_11812, new_AGEMA_signal_11811, KeyExpansionOutput[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U65 ( .a ({new_AGEMA_signal_4876, new_AGEMA_signal_4875, RoundKey[33]}), .b ({new_AGEMA_signal_10904, new_AGEMA_signal_10903, KeyExpansionOutput[65]}), .c ({new_AGEMA_signal_11366, new_AGEMA_signal_11365, KeyExpansionOutput[33]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U64 ( .a ({new_AGEMA_signal_5086, new_AGEMA_signal_5085, RoundKey[65]}), .b ({new_AGEMA_signal_10464, new_AGEMA_signal_10463, KeyExpansionOutput[97]}), .c ({new_AGEMA_signal_10904, new_AGEMA_signal_10903, KeyExpansionOutput[65]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U63 ( .a ({new_AGEMA_signal_5296, new_AGEMA_signal_5295, RoundKey[97]}), .b ({new_AGEMA_signal_10220, new_AGEMA_signal_10219, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_10464, new_AGEMA_signal_10463, KeyExpansionOutput[97]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U62 ( .a ({new_AGEMA_signal_4780, new_AGEMA_signal_4779, RoundKey[19]}), .b ({new_AGEMA_signal_11368, new_AGEMA_signal_11367, KeyExpansionOutput[51]}), .c ({new_AGEMA_signal_11814, new_AGEMA_signal_11813, KeyExpansionOutput[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U61 ( .a ({new_AGEMA_signal_4996, new_AGEMA_signal_4995, RoundKey[51]}), .b ({new_AGEMA_signal_10906, new_AGEMA_signal_10905, KeyExpansionOutput[83]}), .c ({new_AGEMA_signal_11368, new_AGEMA_signal_11367, KeyExpansionOutput[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U60 ( .a ({new_AGEMA_signal_5206, new_AGEMA_signal_5205, RoundKey[83]}), .b ({new_AGEMA_signal_10478, new_AGEMA_signal_10477, KeyExpansionOutput[115]}), .c ({new_AGEMA_signal_10906, new_AGEMA_signal_10905, KeyExpansionOutput[83]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U59 ( .a ({new_AGEMA_signal_4774, new_AGEMA_signal_4773, RoundKey[18]}), .b ({new_AGEMA_signal_11370, new_AGEMA_signal_11369, KeyExpansionOutput[50]}), .c ({new_AGEMA_signal_11816, new_AGEMA_signal_11815, KeyExpansionOutput[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U58 ( .a ({new_AGEMA_signal_4990, new_AGEMA_signal_4989, RoundKey[50]}), .b ({new_AGEMA_signal_10908, new_AGEMA_signal_10907, KeyExpansionOutput[82]}), .c ({new_AGEMA_signal_11370, new_AGEMA_signal_11369, KeyExpansionOutput[50]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U57 ( .a ({new_AGEMA_signal_5200, new_AGEMA_signal_5199, RoundKey[82]}), .b ({new_AGEMA_signal_10480, new_AGEMA_signal_10479, KeyExpansionOutput[114]}), .c ({new_AGEMA_signal_10908, new_AGEMA_signal_10907, KeyExpansionOutput[82]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U56 ( .a ({new_AGEMA_signal_4768, new_AGEMA_signal_4767, RoundKey[17]}), .b ({new_AGEMA_signal_11372, new_AGEMA_signal_11371, KeyExpansionOutput[49]}), .c ({new_AGEMA_signal_11818, new_AGEMA_signal_11817, KeyExpansionOutput[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U55 ( .a ({new_AGEMA_signal_4978, new_AGEMA_signal_4977, RoundKey[49]}), .b ({new_AGEMA_signal_10910, new_AGEMA_signal_10909, KeyExpansionOutput[81]}), .c ({new_AGEMA_signal_11372, new_AGEMA_signal_11371, KeyExpansionOutput[49]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U54 ( .a ({new_AGEMA_signal_5194, new_AGEMA_signal_5193, RoundKey[81]}), .b ({new_AGEMA_signal_10482, new_AGEMA_signal_10481, KeyExpansionOutput[113]}), .c ({new_AGEMA_signal_10910, new_AGEMA_signal_10909, KeyExpansionOutput[81]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U53 ( .a ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, RoundKey[16]}), .b ({new_AGEMA_signal_10912, new_AGEMA_signal_10911, KeyExpansionOutput[48]}), .c ({new_AGEMA_signal_11374, new_AGEMA_signal_11373, KeyExpansionOutput[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U52 ( .a ({new_AGEMA_signal_4972, new_AGEMA_signal_4971, RoundKey[48]}), .b ({new_AGEMA_signal_10466, new_AGEMA_signal_10465, KeyExpansionOutput[80]}), .c ({new_AGEMA_signal_10912, new_AGEMA_signal_10911, KeyExpansionOutput[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U51 ( .a ({new_AGEMA_signal_5188, new_AGEMA_signal_5187, RoundKey[80]}), .b ({new_AGEMA_signal_10158, new_AGEMA_signal_10157, KeyExpansionOutput[112]}), .c ({new_AGEMA_signal_10466, new_AGEMA_signal_10465, KeyExpansionOutput[80]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U50 ( .a ({new_AGEMA_signal_4756, new_AGEMA_signal_4755, RoundKey[15]}), .b ({new_AGEMA_signal_11376, new_AGEMA_signal_11375, KeyExpansionOutput[47]}), .c ({new_AGEMA_signal_11820, new_AGEMA_signal_11819, KeyExpansionOutput[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U49 ( .a ({new_AGEMA_signal_4966, new_AGEMA_signal_4965, RoundKey[47]}), .b ({new_AGEMA_signal_10914, new_AGEMA_signal_10913, KeyExpansionOutput[79]}), .c ({new_AGEMA_signal_11376, new_AGEMA_signal_11375, KeyExpansionOutput[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U48 ( .a ({new_AGEMA_signal_5176, new_AGEMA_signal_5175, RoundKey[79]}), .b ({new_AGEMA_signal_10484, new_AGEMA_signal_10483, KeyExpansionOutput[111]}), .c ({new_AGEMA_signal_10914, new_AGEMA_signal_10913, KeyExpansionOutput[79]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U47 ( .a ({new_AGEMA_signal_4750, new_AGEMA_signal_4749, RoundKey[14]}), .b ({new_AGEMA_signal_11378, new_AGEMA_signal_11377, KeyExpansionOutput[46]}), .c ({new_AGEMA_signal_11822, new_AGEMA_signal_11821, KeyExpansionOutput[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U46 ( .a ({new_AGEMA_signal_4960, new_AGEMA_signal_4959, RoundKey[46]}), .b ({new_AGEMA_signal_10916, new_AGEMA_signal_10915, KeyExpansionOutput[78]}), .c ({new_AGEMA_signal_11378, new_AGEMA_signal_11377, KeyExpansionOutput[46]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U45 ( .a ({new_AGEMA_signal_5170, new_AGEMA_signal_5169, RoundKey[78]}), .b ({new_AGEMA_signal_10486, new_AGEMA_signal_10485, KeyExpansionOutput[110]}), .c ({new_AGEMA_signal_10916, new_AGEMA_signal_10915, KeyExpansionOutput[78]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U44 ( .a ({new_AGEMA_signal_4744, new_AGEMA_signal_4743, RoundKey[13]}), .b ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, KeyExpansionOutput[45]}), .c ({new_AGEMA_signal_11824, new_AGEMA_signal_11823, KeyExpansionOutput[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U43 ( .a ({new_AGEMA_signal_4954, new_AGEMA_signal_4953, RoundKey[45]}), .b ({new_AGEMA_signal_10918, new_AGEMA_signal_10917, KeyExpansionOutput[77]}), .c ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, KeyExpansionOutput[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U42 ( .a ({new_AGEMA_signal_5164, new_AGEMA_signal_5163, RoundKey[77]}), .b ({new_AGEMA_signal_10488, new_AGEMA_signal_10487, KeyExpansionOutput[109]}), .c ({new_AGEMA_signal_10918, new_AGEMA_signal_10917, KeyExpansionOutput[77]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U41 ( .a ({new_AGEMA_signal_4738, new_AGEMA_signal_4737, RoundKey[12]}), .b ({new_AGEMA_signal_11382, new_AGEMA_signal_11381, KeyExpansionOutput[44]}), .c ({new_AGEMA_signal_11826, new_AGEMA_signal_11825, KeyExpansionOutput[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U40 ( .a ({new_AGEMA_signal_4948, new_AGEMA_signal_4947, RoundKey[44]}), .b ({new_AGEMA_signal_10920, new_AGEMA_signal_10919, KeyExpansionOutput[76]}), .c ({new_AGEMA_signal_11382, new_AGEMA_signal_11381, KeyExpansionOutput[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U39 ( .a ({new_AGEMA_signal_5158, new_AGEMA_signal_5157, RoundKey[76]}), .b ({new_AGEMA_signal_10490, new_AGEMA_signal_10489, KeyExpansionOutput[108]}), .c ({new_AGEMA_signal_10920, new_AGEMA_signal_10919, KeyExpansionOutput[76]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U38 ( .a ({new_AGEMA_signal_4732, new_AGEMA_signal_4731, RoundKey[127]}), .b ({new_AGEMA_signal_10508, new_AGEMA_signal_10507, KeyExpansionIns_tmp[31]}), .c ({new_AGEMA_signal_10922, new_AGEMA_signal_10921, KeyExpansionOutput[127]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U37 ( .a ({new_AGEMA_signal_4726, new_AGEMA_signal_4725, RoundKey[126]}), .b ({new_AGEMA_signal_10510, new_AGEMA_signal_10509, KeyExpansionIns_tmp[30]}), .c ({new_AGEMA_signal_10924, new_AGEMA_signal_10923, KeyExpansionOutput[126]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U36 ( .a ({new_AGEMA_signal_4720, new_AGEMA_signal_4719, RoundKey[125]}), .b ({new_AGEMA_signal_10512, new_AGEMA_signal_10511, KeyExpansionIns_tmp[29]}), .c ({new_AGEMA_signal_10926, new_AGEMA_signal_10925, KeyExpansionOutput[125]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U35 ( .a ({new_AGEMA_signal_4714, new_AGEMA_signal_4713, RoundKey[124]}), .b ({new_AGEMA_signal_10514, new_AGEMA_signal_10513, KeyExpansionIns_tmp[28]}), .c ({new_AGEMA_signal_10928, new_AGEMA_signal_10927, KeyExpansionOutput[124]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U34 ( .a ({new_AGEMA_signal_4708, new_AGEMA_signal_4707, RoundKey[123]}), .b ({new_AGEMA_signal_10516, new_AGEMA_signal_10515, KeyExpansionIns_tmp[27]}), .c ({new_AGEMA_signal_10930, new_AGEMA_signal_10929, KeyExpansionOutput[123]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U33 ( .a ({new_AGEMA_signal_4702, new_AGEMA_signal_4701, RoundKey[122]}), .b ({new_AGEMA_signal_10518, new_AGEMA_signal_10517, KeyExpansionIns_tmp[26]}), .c ({new_AGEMA_signal_10932, new_AGEMA_signal_10931, KeyExpansionOutput[122]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U32 ( .a ({new_AGEMA_signal_4696, new_AGEMA_signal_4695, RoundKey[121]}), .b ({new_AGEMA_signal_10520, new_AGEMA_signal_10519, KeyExpansionIns_tmp[25]}), .c ({new_AGEMA_signal_10934, new_AGEMA_signal_10933, KeyExpansionOutput[121]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U31 ( .a ({new_AGEMA_signal_4690, new_AGEMA_signal_4689, RoundKey[120]}), .b ({new_AGEMA_signal_10164, new_AGEMA_signal_10163, KeyExpansionIns_tmp[24]}), .c ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, KeyExpansionOutput[120]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U30 ( .a ({new_AGEMA_signal_4684, new_AGEMA_signal_4683, RoundKey[11]}), .b ({new_AGEMA_signal_11384, new_AGEMA_signal_11383, KeyExpansionOutput[43]}), .c ({new_AGEMA_signal_11828, new_AGEMA_signal_11827, KeyExpansionOutput[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U29 ( .a ({new_AGEMA_signal_4942, new_AGEMA_signal_4941, RoundKey[43]}), .b ({new_AGEMA_signal_10936, new_AGEMA_signal_10935, KeyExpansionOutput[75]}), .c ({new_AGEMA_signal_11384, new_AGEMA_signal_11383, KeyExpansionOutput[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U28 ( .a ({new_AGEMA_signal_5152, new_AGEMA_signal_5151, RoundKey[75]}), .b ({new_AGEMA_signal_10492, new_AGEMA_signal_10491, KeyExpansionOutput[107]}), .c ({new_AGEMA_signal_10936, new_AGEMA_signal_10935, KeyExpansionOutput[75]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U27 ( .a ({new_AGEMA_signal_4678, new_AGEMA_signal_4677, RoundKey[119]}), .b ({new_AGEMA_signal_10180, new_AGEMA_signal_10179, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_10470, new_AGEMA_signal_10469, KeyExpansionOutput[119]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U26 ( .a ({new_AGEMA_signal_4672, new_AGEMA_signal_4671, RoundKey[118]}), .b ({new_AGEMA_signal_10182, new_AGEMA_signal_10181, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_10472, new_AGEMA_signal_10471, KeyExpansionOutput[118]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U25 ( .a ({new_AGEMA_signal_4666, new_AGEMA_signal_4665, RoundKey[117]}), .b ({new_AGEMA_signal_10184, new_AGEMA_signal_10183, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_10474, new_AGEMA_signal_10473, KeyExpansionOutput[117]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U24 ( .a ({new_AGEMA_signal_4660, new_AGEMA_signal_4659, RoundKey[116]}), .b ({new_AGEMA_signal_10186, new_AGEMA_signal_10185, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_10476, new_AGEMA_signal_10475, KeyExpansionOutput[116]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U23 ( .a ({new_AGEMA_signal_4654, new_AGEMA_signal_4653, RoundKey[115]}), .b ({new_AGEMA_signal_10188, new_AGEMA_signal_10187, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_10478, new_AGEMA_signal_10477, KeyExpansionOutput[115]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U22 ( .a ({new_AGEMA_signal_4648, new_AGEMA_signal_4647, RoundKey[114]}), .b ({new_AGEMA_signal_10190, new_AGEMA_signal_10189, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_10480, new_AGEMA_signal_10479, KeyExpansionOutput[114]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U21 ( .a ({new_AGEMA_signal_4642, new_AGEMA_signal_4641, RoundKey[113]}), .b ({new_AGEMA_signal_10192, new_AGEMA_signal_10191, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_10482, new_AGEMA_signal_10481, KeyExpansionOutput[113]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U20 ( .a ({new_AGEMA_signal_4636, new_AGEMA_signal_4635, RoundKey[112]}), .b ({new_AGEMA_signal_9760, new_AGEMA_signal_9759, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_10158, new_AGEMA_signal_10157, KeyExpansionOutput[112]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U19 ( .a ({new_AGEMA_signal_4630, new_AGEMA_signal_4629, RoundKey[111]}), .b ({new_AGEMA_signal_10194, new_AGEMA_signal_10193, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_10484, new_AGEMA_signal_10483, KeyExpansionOutput[111]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U18 ( .a ({new_AGEMA_signal_4624, new_AGEMA_signal_4623, RoundKey[110]}), .b ({new_AGEMA_signal_10196, new_AGEMA_signal_10195, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_10486, new_AGEMA_signal_10485, KeyExpansionOutput[110]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U17 ( .a ({new_AGEMA_signal_4618, new_AGEMA_signal_4617, RoundKey[10]}), .b ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, KeyExpansionOutput[42]}), .c ({new_AGEMA_signal_11830, new_AGEMA_signal_11829, KeyExpansionOutput[10]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U16 ( .a ({new_AGEMA_signal_4936, new_AGEMA_signal_4935, RoundKey[42]}), .b ({new_AGEMA_signal_10938, new_AGEMA_signal_10937, KeyExpansionOutput[74]}), .c ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, KeyExpansionOutput[42]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U15 ( .a ({new_AGEMA_signal_5146, new_AGEMA_signal_5145, RoundKey[74]}), .b ({new_AGEMA_signal_10494, new_AGEMA_signal_10493, KeyExpansionOutput[106]}), .c ({new_AGEMA_signal_10938, new_AGEMA_signal_10937, KeyExpansionOutput[74]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U14 ( .a ({new_AGEMA_signal_4612, new_AGEMA_signal_4611, RoundKey[109]}), .b ({new_AGEMA_signal_10198, new_AGEMA_signal_10197, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_10488, new_AGEMA_signal_10487, KeyExpansionOutput[109]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U13 ( .a ({new_AGEMA_signal_4606, new_AGEMA_signal_4605, RoundKey[108]}), .b ({new_AGEMA_signal_10200, new_AGEMA_signal_10199, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_10490, new_AGEMA_signal_10489, KeyExpansionOutput[108]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U12 ( .a ({new_AGEMA_signal_4600, new_AGEMA_signal_4599, RoundKey[107]}), .b ({new_AGEMA_signal_10202, new_AGEMA_signal_10201, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_10492, new_AGEMA_signal_10491, KeyExpansionOutput[107]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U11 ( .a ({new_AGEMA_signal_4594, new_AGEMA_signal_4593, RoundKey[106]}), .b ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_10494, new_AGEMA_signal_10493, KeyExpansionOutput[106]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U10 ( .a ({new_AGEMA_signal_4588, new_AGEMA_signal_4587, RoundKey[105]}), .b ({new_AGEMA_signal_10206, new_AGEMA_signal_10205, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_10496, new_AGEMA_signal_10495, KeyExpansionOutput[105]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U9 ( .a ({new_AGEMA_signal_4582, new_AGEMA_signal_4581, RoundKey[104]}), .b ({new_AGEMA_signal_9782, new_AGEMA_signal_9781, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_10160, new_AGEMA_signal_10159, KeyExpansionOutput[104]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U8 ( .a ({new_AGEMA_signal_4576, new_AGEMA_signal_4575, RoundKey[103]}), .b ({new_AGEMA_signal_10208, new_AGEMA_signal_10207, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_10498, new_AGEMA_signal_10497, KeyExpansionOutput[103]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U7 ( .a ({new_AGEMA_signal_4570, new_AGEMA_signal_4569, RoundKey[102]}), .b ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_10500, new_AGEMA_signal_10499, KeyExpansionOutput[102]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U6 ( .a ({new_AGEMA_signal_4564, new_AGEMA_signal_4563, RoundKey[101]}), .b ({new_AGEMA_signal_10212, new_AGEMA_signal_10211, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_10502, new_AGEMA_signal_10501, KeyExpansionOutput[101]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U5 ( .a ({new_AGEMA_signal_4558, new_AGEMA_signal_4557, RoundKey[100]}), .b ({new_AGEMA_signal_10214, new_AGEMA_signal_10213, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_10504, new_AGEMA_signal_10503, KeyExpansionOutput[100]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U4 ( .a ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, RoundKey[0]}), .b ({new_AGEMA_signal_10940, new_AGEMA_signal_10939, KeyExpansionOutput[32]}), .c ({new_AGEMA_signal_11388, new_AGEMA_signal_11387, KeyExpansionOutput[0]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U3 ( .a ({new_AGEMA_signal_4870, new_AGEMA_signal_4869, RoundKey[32]}), .b ({new_AGEMA_signal_10506, new_AGEMA_signal_10505, KeyExpansionOutput[64]}), .c ({new_AGEMA_signal_10940, new_AGEMA_signal_10939, KeyExpansionOutput[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U2 ( .a ({new_AGEMA_signal_5080, new_AGEMA_signal_5079, RoundKey[64]}), .b ({new_AGEMA_signal_10162, new_AGEMA_signal_10161, KeyExpansionOutput[96]}), .c ({new_AGEMA_signal_10506, new_AGEMA_signal_10505, KeyExpansionOutput[64]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U1 ( .a ({new_AGEMA_signal_5290, new_AGEMA_signal_5289, RoundKey[96]}), .b ({new_AGEMA_signal_9804, new_AGEMA_signal_9803, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_10162, new_AGEMA_signal_10161, KeyExpansionOutput[96]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U8 ( .a ({new_AGEMA_signal_10166, new_AGEMA_signal_10165, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_}), .b ({1'b0, 1'b0, n283}), .c ({new_AGEMA_signal_10508, new_AGEMA_signal_10507, KeyExpansionIns_tmp[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U7 ( .a ({new_AGEMA_signal_10168, new_AGEMA_signal_10167, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_}), .b ({1'b0, 1'b0, n285}), .c ({new_AGEMA_signal_10510, new_AGEMA_signal_10509, KeyExpansionIns_tmp[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U6 ( .a ({new_AGEMA_signal_10170, new_AGEMA_signal_10169, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_}), .b ({1'b0, 1'b0, Rcon[5]}), .c ({new_AGEMA_signal_10512, new_AGEMA_signal_10511, KeyExpansionIns_tmp[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U5 ( .a ({new_AGEMA_signal_10172, new_AGEMA_signal_10171, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_}), .b ({1'b0, 1'b0, Rcon[4]}), .c ({new_AGEMA_signal_10514, new_AGEMA_signal_10513, KeyExpansionIns_tmp[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U4 ( .a ({new_AGEMA_signal_10174, new_AGEMA_signal_10173, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_}), .b ({1'b0, 1'b0, Rcon[3]}), .c ({new_AGEMA_signal_10516, new_AGEMA_signal_10515, KeyExpansionIns_tmp[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U3 ( .a ({new_AGEMA_signal_10176, new_AGEMA_signal_10175, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_}), .b ({1'b0, 1'b0, Rcon[2]}), .c ({new_AGEMA_signal_10518, new_AGEMA_signal_10517, KeyExpansionIns_tmp[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U2 ( .a ({new_AGEMA_signal_10178, new_AGEMA_signal_10177, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_}), .b ({1'b0, 1'b0, Rcon[1]}), .c ({new_AGEMA_signal_10520, new_AGEMA_signal_10519, KeyExpansionIns_tmp[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U1 ( .a ({new_AGEMA_signal_9738, new_AGEMA_signal_9737, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_}), .b ({1'b0, 1'b0, Rcon[0]}), .c ({new_AGEMA_signal_10164, new_AGEMA_signal_10163, KeyExpansionIns_tmp[24]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M46_U1 ( .a ({new_AGEMA_signal_8004, new_AGEMA_signal_8003, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .clk (clk), .r ({Fresh[1826], Fresh[1825], Fresh[1824]}), .c ({new_AGEMA_signal_8480, new_AGEMA_signal_8479, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M47_U1 ( .a ({new_AGEMA_signal_7844, new_AGEMA_signal_7843, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_6038, new_AGEMA_signal_6037, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8}), .clk (clk), .r ({Fresh[1829], Fresh[1828], Fresh[1827]}), .c ({new_AGEMA_signal_8006, new_AGEMA_signal_8005, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M48_U1 ( .a ({new_AGEMA_signal_7842, new_AGEMA_signal_7841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, RoundKey[16]}), .clk (clk), .r ({Fresh[1832], Fresh[1831], Fresh[1830]}), .c ({new_AGEMA_signal_8008, new_AGEMA_signal_8007, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M49_U1 ( .a ({new_AGEMA_signal_8002, new_AGEMA_signal_8001, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_5726, new_AGEMA_signal_5725, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .clk (clk), .r ({Fresh[1835], Fresh[1834], Fresh[1833]}), .c ({new_AGEMA_signal_8482, new_AGEMA_signal_8481, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M50_U1 ( .a ({new_AGEMA_signal_7840, new_AGEMA_signal_7839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_5720, new_AGEMA_signal_5719, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}), .clk (clk), .r ({Fresh[1838], Fresh[1837], Fresh[1836]}), .c ({new_AGEMA_signal_8010, new_AGEMA_signal_8009, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M51_U1 ( .a ({new_AGEMA_signal_7838, new_AGEMA_signal_7837, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_6044, new_AGEMA_signal_6043, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}), .clk (clk), .r ({Fresh[1841], Fresh[1840], Fresh[1839]}), .c ({new_AGEMA_signal_8012, new_AGEMA_signal_8011, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M52_U1 ( .a ({new_AGEMA_signal_8000, new_AGEMA_signal_7999, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_5724, new_AGEMA_signal_5723, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15}), .clk (clk), .r ({Fresh[1844], Fresh[1843], Fresh[1842]}), .c ({new_AGEMA_signal_8484, new_AGEMA_signal_8483, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M53_U1 ( .a ({new_AGEMA_signal_8478, new_AGEMA_signal_8477, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_5732, new_AGEMA_signal_5731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27}), .clk (clk), .r ({Fresh[1847], Fresh[1846], Fresh[1845]}), .c ({new_AGEMA_signal_8958, new_AGEMA_signal_8957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M54_U1 ( .a ({new_AGEMA_signal_7998, new_AGEMA_signal_7997, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_6040, new_AGEMA_signal_6039, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}), .clk (clk), .r ({Fresh[1850], Fresh[1849], Fresh[1848]}), .c ({new_AGEMA_signal_8486, new_AGEMA_signal_8485, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M55_U1 ( .a ({new_AGEMA_signal_8004, new_AGEMA_signal_8003, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_5722, new_AGEMA_signal_5721, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13}), .clk (clk), .r ({Fresh[1853], Fresh[1852], Fresh[1851]}), .c ({new_AGEMA_signal_8488, new_AGEMA_signal_8487, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M56_U1 ( .a ({new_AGEMA_signal_7844, new_AGEMA_signal_7843, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_6048, new_AGEMA_signal_6047, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23}), .clk (clk), .r ({Fresh[1856], Fresh[1855], Fresh[1854]}), .c ({new_AGEMA_signal_8014, new_AGEMA_signal_8013, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M57_U1 ( .a ({new_AGEMA_signal_7842, new_AGEMA_signal_7841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_5728, new_AGEMA_signal_5727, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}), .clk (clk), .r ({Fresh[1859], Fresh[1858], Fresh[1857]}), .c ({new_AGEMA_signal_8016, new_AGEMA_signal_8015, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M58_U1 ( .a ({new_AGEMA_signal_8002, new_AGEMA_signal_8001, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_5322, new_AGEMA_signal_5321, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .clk (clk), .r ({Fresh[1862], Fresh[1861], Fresh[1860]}), .c ({new_AGEMA_signal_8490, new_AGEMA_signal_8489, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M59_U1 ( .a ({new_AGEMA_signal_7840, new_AGEMA_signal_7839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_5730, new_AGEMA_signal_5729, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}), .clk (clk), .r ({Fresh[1865], Fresh[1864], Fresh[1863]}), .c ({new_AGEMA_signal_8018, new_AGEMA_signal_8017, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M60_U1 ( .a ({new_AGEMA_signal_7838, new_AGEMA_signal_7837, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_6046, new_AGEMA_signal_6045, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}), .clk (clk), .r ({Fresh[1868], Fresh[1867], Fresh[1866]}), .c ({new_AGEMA_signal_8020, new_AGEMA_signal_8019, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M61_U1 ( .a ({new_AGEMA_signal_8000, new_AGEMA_signal_7999, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_5318, new_AGEMA_signal_5317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .clk (clk), .r ({Fresh[1871], Fresh[1870], Fresh[1869]}), .c ({new_AGEMA_signal_8492, new_AGEMA_signal_8491, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M62_U1 ( .a ({new_AGEMA_signal_8478, new_AGEMA_signal_8477, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_5324, new_AGEMA_signal_5323, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}), .clk (clk), .r ({Fresh[1874], Fresh[1873], Fresh[1872]}), .c ({new_AGEMA_signal_8960, new_AGEMA_signal_8959, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M63_U1 ( .a ({new_AGEMA_signal_7998, new_AGEMA_signal_7997, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_5320, new_AGEMA_signal_5319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .clk (clk), .r ({Fresh[1877], Fresh[1876], Fresh[1875]}), .c ({new_AGEMA_signal_8494, new_AGEMA_signal_8493, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L0_U1 ( .a ({new_AGEMA_signal_8492, new_AGEMA_signal_8491, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}), .b ({new_AGEMA_signal_8960, new_AGEMA_signal_8959, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62}), .c ({new_AGEMA_signal_9358, new_AGEMA_signal_9357, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L1_U1 ( .a ({new_AGEMA_signal_8010, new_AGEMA_signal_8009, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_8014, new_AGEMA_signal_8013, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56}), .c ({new_AGEMA_signal_8496, new_AGEMA_signal_8495, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L2_U1 ( .a ({new_AGEMA_signal_8480, new_AGEMA_signal_8479, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_8008, new_AGEMA_signal_8007, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48}), .c ({new_AGEMA_signal_8962, new_AGEMA_signal_8961, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L3_U1 ( .a ({new_AGEMA_signal_8006, new_AGEMA_signal_8005, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47}), .b ({new_AGEMA_signal_8488, new_AGEMA_signal_8487, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55}), .c ({new_AGEMA_signal_8964, new_AGEMA_signal_8963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L4_U1 ( .a ({new_AGEMA_signal_8486, new_AGEMA_signal_8485, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54}), .b ({new_AGEMA_signal_8490, new_AGEMA_signal_8489, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58}), .c ({new_AGEMA_signal_8966, new_AGEMA_signal_8965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L5_U1 ( .a ({new_AGEMA_signal_8482, new_AGEMA_signal_8481, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49}), .b ({new_AGEMA_signal_8492, new_AGEMA_signal_8491, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_8968, new_AGEMA_signal_8967, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L6_U1 ( .a ({new_AGEMA_signal_8960, new_AGEMA_signal_8959, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62}), .b ({new_AGEMA_signal_8968, new_AGEMA_signal_8967, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5}), .c ({new_AGEMA_signal_9360, new_AGEMA_signal_9359, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L7_U1 ( .a ({new_AGEMA_signal_8480, new_AGEMA_signal_8479, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_8964, new_AGEMA_signal_8963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3}), .c ({new_AGEMA_signal_9362, new_AGEMA_signal_9361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L8_U1 ( .a ({new_AGEMA_signal_8012, new_AGEMA_signal_8011, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51}), .b ({new_AGEMA_signal_8018, new_AGEMA_signal_8017, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59}), .c ({new_AGEMA_signal_8498, new_AGEMA_signal_8497, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L9_U1 ( .a ({new_AGEMA_signal_8484, new_AGEMA_signal_8483, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_8958, new_AGEMA_signal_8957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53}), .c ({new_AGEMA_signal_9364, new_AGEMA_signal_9363, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L10_U1 ( .a ({new_AGEMA_signal_8958, new_AGEMA_signal_8957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53}), .b ({new_AGEMA_signal_8966, new_AGEMA_signal_8965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_9366, new_AGEMA_signal_9365, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L11_U1 ( .a ({new_AGEMA_signal_8020, new_AGEMA_signal_8019, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60}), .b ({new_AGEMA_signal_8962, new_AGEMA_signal_8961, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_9368, new_AGEMA_signal_9367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L12_U1 ( .a ({new_AGEMA_signal_8008, new_AGEMA_signal_8007, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48}), .b ({new_AGEMA_signal_8012, new_AGEMA_signal_8011, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51}), .c ({new_AGEMA_signal_8500, new_AGEMA_signal_8499, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L13_U1 ( .a ({new_AGEMA_signal_8010, new_AGEMA_signal_8009, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_9358, new_AGEMA_signal_9357, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_9718, new_AGEMA_signal_9717, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L14_U1 ( .a ({new_AGEMA_signal_8484, new_AGEMA_signal_8483, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_8492, new_AGEMA_signal_8491, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_8970, new_AGEMA_signal_8969, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L15_U1 ( .a ({new_AGEMA_signal_8488, new_AGEMA_signal_8487, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55}), .b ({new_AGEMA_signal_8496, new_AGEMA_signal_8495, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_8972, new_AGEMA_signal_8971, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L16_U1 ( .a ({new_AGEMA_signal_8014, new_AGEMA_signal_8013, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56}), .b ({new_AGEMA_signal_9358, new_AGEMA_signal_9357, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_9720, new_AGEMA_signal_9719, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L17_U1 ( .a ({new_AGEMA_signal_8016, new_AGEMA_signal_8015, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57}), .b ({new_AGEMA_signal_8496, new_AGEMA_signal_8495, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_8974, new_AGEMA_signal_8973, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L18_U1 ( .a ({new_AGEMA_signal_8490, new_AGEMA_signal_8489, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58}), .b ({new_AGEMA_signal_8498, new_AGEMA_signal_8497, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8}), .c ({new_AGEMA_signal_8976, new_AGEMA_signal_8975, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L19_U1 ( .a ({new_AGEMA_signal_8494, new_AGEMA_signal_8493, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63}), .b ({new_AGEMA_signal_8966, new_AGEMA_signal_8965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_9370, new_AGEMA_signal_9369, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L20_U1 ( .a ({new_AGEMA_signal_9358, new_AGEMA_signal_9357, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}), .b ({new_AGEMA_signal_8496, new_AGEMA_signal_8495, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_9722, new_AGEMA_signal_9721, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L21_U1 ( .a ({new_AGEMA_signal_8496, new_AGEMA_signal_8495, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .b ({new_AGEMA_signal_9362, new_AGEMA_signal_9361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7}), .c ({new_AGEMA_signal_9724, new_AGEMA_signal_9723, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L22_U1 ( .a ({new_AGEMA_signal_8964, new_AGEMA_signal_8963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3}), .b ({new_AGEMA_signal_8500, new_AGEMA_signal_8499, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12}), .c ({new_AGEMA_signal_9372, new_AGEMA_signal_9371, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L23_U1 ( .a ({new_AGEMA_signal_8976, new_AGEMA_signal_8975, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18}), .b ({new_AGEMA_signal_8962, new_AGEMA_signal_8961, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_9374, new_AGEMA_signal_9373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L24_U1 ( .a ({new_AGEMA_signal_8972, new_AGEMA_signal_8971, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15}), .b ({new_AGEMA_signal_9364, new_AGEMA_signal_9363, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_9726, new_AGEMA_signal_9725, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L25_U1 ( .a ({new_AGEMA_signal_9360, new_AGEMA_signal_9359, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_9366, new_AGEMA_signal_9365, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_9728, new_AGEMA_signal_9727, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L26_U1 ( .a ({new_AGEMA_signal_9362, new_AGEMA_signal_9361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7}), .b ({new_AGEMA_signal_9364, new_AGEMA_signal_9363, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_9730, new_AGEMA_signal_9729, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L27_U1 ( .a ({new_AGEMA_signal_8498, new_AGEMA_signal_8497, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8}), .b ({new_AGEMA_signal_9366, new_AGEMA_signal_9365, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_9732, new_AGEMA_signal_9731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L28_U1 ( .a ({new_AGEMA_signal_9368, new_AGEMA_signal_9367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_8970, new_AGEMA_signal_8969, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14}), .c ({new_AGEMA_signal_9734, new_AGEMA_signal_9733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L29_U1 ( .a ({new_AGEMA_signal_9368, new_AGEMA_signal_9367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_8974, new_AGEMA_signal_8973, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17}), .c ({new_AGEMA_signal_9736, new_AGEMA_signal_9735, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S0_U1 ( .a ({new_AGEMA_signal_9360, new_AGEMA_signal_9359, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_9726, new_AGEMA_signal_9725, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24}), .c ({new_AGEMA_signal_10166, new_AGEMA_signal_10165, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S1_U1 ( .a ({new_AGEMA_signal_9720, new_AGEMA_signal_9719, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16}), .b ({new_AGEMA_signal_9730, new_AGEMA_signal_9729, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26}), .c ({new_AGEMA_signal_10168, new_AGEMA_signal_10167, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S2_U1 ( .a ({new_AGEMA_signal_9370, new_AGEMA_signal_9369, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19}), .b ({new_AGEMA_signal_9734, new_AGEMA_signal_9733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28}), .c ({new_AGEMA_signal_10170, new_AGEMA_signal_10169, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S3_U1 ( .a ({new_AGEMA_signal_9360, new_AGEMA_signal_9359, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_9724, new_AGEMA_signal_9723, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21}), .c ({new_AGEMA_signal_10172, new_AGEMA_signal_10171, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S4_U1 ( .a ({new_AGEMA_signal_9722, new_AGEMA_signal_9721, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20}), .b ({new_AGEMA_signal_9372, new_AGEMA_signal_9371, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22}), .c ({new_AGEMA_signal_10174, new_AGEMA_signal_10173, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S5_U1 ( .a ({new_AGEMA_signal_9728, new_AGEMA_signal_9727, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25}), .b ({new_AGEMA_signal_9736, new_AGEMA_signal_9735, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29}), .c ({new_AGEMA_signal_10176, new_AGEMA_signal_10175, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S6_U1 ( .a ({new_AGEMA_signal_9718, new_AGEMA_signal_9717, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13}), .b ({new_AGEMA_signal_9732, new_AGEMA_signal_9731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27}), .c ({new_AGEMA_signal_10178, new_AGEMA_signal_10177, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S7_U1 ( .a ({new_AGEMA_signal_9360, new_AGEMA_signal_9359, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_9374, new_AGEMA_signal_9373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23}), .c ({new_AGEMA_signal_9738, new_AGEMA_signal_9737, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M46_U1 ( .a ({new_AGEMA_signal_8028, new_AGEMA_signal_8027, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_5734, new_AGEMA_signal_5733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .clk (clk), .r ({Fresh[1880], Fresh[1879], Fresh[1878]}), .c ({new_AGEMA_signal_8504, new_AGEMA_signal_8503, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M47_U1 ( .a ({new_AGEMA_signal_7852, new_AGEMA_signal_7851, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_6064, new_AGEMA_signal_6063, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8}), .clk (clk), .r ({Fresh[1883], Fresh[1882], Fresh[1881]}), .c ({new_AGEMA_signal_8030, new_AGEMA_signal_8029, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M48_U1 ( .a ({new_AGEMA_signal_7850, new_AGEMA_signal_7849, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_5248, new_AGEMA_signal_5247, RoundKey[8]}), .clk (clk), .r ({Fresh[1886], Fresh[1885], Fresh[1884]}), .c ({new_AGEMA_signal_8032, new_AGEMA_signal_8031, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M49_U1 ( .a ({new_AGEMA_signal_8026, new_AGEMA_signal_8025, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .clk (clk), .r ({Fresh[1889], Fresh[1888], Fresh[1887]}), .c ({new_AGEMA_signal_8506, new_AGEMA_signal_8505, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M50_U1 ( .a ({new_AGEMA_signal_7848, new_AGEMA_signal_7847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_5736, new_AGEMA_signal_5735, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}), .clk (clk), .r ({Fresh[1892], Fresh[1891], Fresh[1890]}), .c ({new_AGEMA_signal_8034, new_AGEMA_signal_8033, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M51_U1 ( .a ({new_AGEMA_signal_7846, new_AGEMA_signal_7845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_6070, new_AGEMA_signal_6069, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}), .clk (clk), .r ({Fresh[1895], Fresh[1894], Fresh[1893]}), .c ({new_AGEMA_signal_8036, new_AGEMA_signal_8035, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M52_U1 ( .a ({new_AGEMA_signal_8024, new_AGEMA_signal_8023, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_5740, new_AGEMA_signal_5739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15}), .clk (clk), .r ({Fresh[1898], Fresh[1897], Fresh[1896]}), .c ({new_AGEMA_signal_8508, new_AGEMA_signal_8507, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M53_U1 ( .a ({new_AGEMA_signal_8502, new_AGEMA_signal_8501, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27}), .clk (clk), .r ({Fresh[1901], Fresh[1900], Fresh[1899]}), .c ({new_AGEMA_signal_8978, new_AGEMA_signal_8977, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M54_U1 ( .a ({new_AGEMA_signal_8022, new_AGEMA_signal_8021, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_6066, new_AGEMA_signal_6065, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}), .clk (clk), .r ({Fresh[1904], Fresh[1903], Fresh[1902]}), .c ({new_AGEMA_signal_8510, new_AGEMA_signal_8509, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M55_U1 ( .a ({new_AGEMA_signal_8028, new_AGEMA_signal_8027, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_5738, new_AGEMA_signal_5737, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13}), .clk (clk), .r ({Fresh[1907], Fresh[1906], Fresh[1905]}), .c ({new_AGEMA_signal_8512, new_AGEMA_signal_8511, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M56_U1 ( .a ({new_AGEMA_signal_7852, new_AGEMA_signal_7851, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_6074, new_AGEMA_signal_6073, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23}), .clk (clk), .r ({Fresh[1910], Fresh[1909], Fresh[1908]}), .c ({new_AGEMA_signal_8038, new_AGEMA_signal_8037, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M57_U1 ( .a ({new_AGEMA_signal_7850, new_AGEMA_signal_7849, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_5744, new_AGEMA_signal_5743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}), .clk (clk), .r ({Fresh[1913], Fresh[1912], Fresh[1911]}), .c ({new_AGEMA_signal_8040, new_AGEMA_signal_8039, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M58_U1 ( .a ({new_AGEMA_signal_8026, new_AGEMA_signal_8025, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_5342, new_AGEMA_signal_5341, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .clk (clk), .r ({Fresh[1916], Fresh[1915], Fresh[1914]}), .c ({new_AGEMA_signal_8514, new_AGEMA_signal_8513, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M59_U1 ( .a ({new_AGEMA_signal_7848, new_AGEMA_signal_7847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_5746, new_AGEMA_signal_5745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}), .clk (clk), .r ({Fresh[1919], Fresh[1918], Fresh[1917]}), .c ({new_AGEMA_signal_8042, new_AGEMA_signal_8041, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M60_U1 ( .a ({new_AGEMA_signal_7846, new_AGEMA_signal_7845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_6072, new_AGEMA_signal_6071, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}), .clk (clk), .r ({Fresh[1922], Fresh[1921], Fresh[1920]}), .c ({new_AGEMA_signal_8044, new_AGEMA_signal_8043, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M61_U1 ( .a ({new_AGEMA_signal_8024, new_AGEMA_signal_8023, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_5338, new_AGEMA_signal_5337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .clk (clk), .r ({Fresh[1925], Fresh[1924], Fresh[1923]}), .c ({new_AGEMA_signal_8516, new_AGEMA_signal_8515, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M62_U1 ( .a ({new_AGEMA_signal_8502, new_AGEMA_signal_8501, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_5344, new_AGEMA_signal_5343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}), .clk (clk), .r ({Fresh[1928], Fresh[1927], Fresh[1926]}), .c ({new_AGEMA_signal_8980, new_AGEMA_signal_8979, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M63_U1 ( .a ({new_AGEMA_signal_8022, new_AGEMA_signal_8021, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_5340, new_AGEMA_signal_5339, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .clk (clk), .r ({Fresh[1931], Fresh[1930], Fresh[1929]}), .c ({new_AGEMA_signal_8518, new_AGEMA_signal_8517, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L0_U1 ( .a ({new_AGEMA_signal_8516, new_AGEMA_signal_8515, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}), .b ({new_AGEMA_signal_8980, new_AGEMA_signal_8979, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62}), .c ({new_AGEMA_signal_9376, new_AGEMA_signal_9375, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L1_U1 ( .a ({new_AGEMA_signal_8034, new_AGEMA_signal_8033, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_8038, new_AGEMA_signal_8037, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56}), .c ({new_AGEMA_signal_8520, new_AGEMA_signal_8519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L2_U1 ( .a ({new_AGEMA_signal_8504, new_AGEMA_signal_8503, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_8032, new_AGEMA_signal_8031, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48}), .c ({new_AGEMA_signal_8982, new_AGEMA_signal_8981, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L3_U1 ( .a ({new_AGEMA_signal_8030, new_AGEMA_signal_8029, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47}), .b ({new_AGEMA_signal_8512, new_AGEMA_signal_8511, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55}), .c ({new_AGEMA_signal_8984, new_AGEMA_signal_8983, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L4_U1 ( .a ({new_AGEMA_signal_8510, new_AGEMA_signal_8509, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54}), .b ({new_AGEMA_signal_8514, new_AGEMA_signal_8513, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58}), .c ({new_AGEMA_signal_8986, new_AGEMA_signal_8985, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L5_U1 ( .a ({new_AGEMA_signal_8506, new_AGEMA_signal_8505, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49}), .b ({new_AGEMA_signal_8516, new_AGEMA_signal_8515, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_8988, new_AGEMA_signal_8987, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L6_U1 ( .a ({new_AGEMA_signal_8980, new_AGEMA_signal_8979, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62}), .b ({new_AGEMA_signal_8988, new_AGEMA_signal_8987, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5}), .c ({new_AGEMA_signal_9378, new_AGEMA_signal_9377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L7_U1 ( .a ({new_AGEMA_signal_8504, new_AGEMA_signal_8503, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_8984, new_AGEMA_signal_8983, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3}), .c ({new_AGEMA_signal_9380, new_AGEMA_signal_9379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L8_U1 ( .a ({new_AGEMA_signal_8036, new_AGEMA_signal_8035, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51}), .b ({new_AGEMA_signal_8042, new_AGEMA_signal_8041, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59}), .c ({new_AGEMA_signal_8522, new_AGEMA_signal_8521, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L9_U1 ( .a ({new_AGEMA_signal_8508, new_AGEMA_signal_8507, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_8978, new_AGEMA_signal_8977, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53}), .c ({new_AGEMA_signal_9382, new_AGEMA_signal_9381, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L10_U1 ( .a ({new_AGEMA_signal_8978, new_AGEMA_signal_8977, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53}), .b ({new_AGEMA_signal_8986, new_AGEMA_signal_8985, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_9384, new_AGEMA_signal_9383, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L11_U1 ( .a ({new_AGEMA_signal_8044, new_AGEMA_signal_8043, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60}), .b ({new_AGEMA_signal_8982, new_AGEMA_signal_8981, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_9386, new_AGEMA_signal_9385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L12_U1 ( .a ({new_AGEMA_signal_8032, new_AGEMA_signal_8031, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48}), .b ({new_AGEMA_signal_8036, new_AGEMA_signal_8035, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51}), .c ({new_AGEMA_signal_8524, new_AGEMA_signal_8523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L13_U1 ( .a ({new_AGEMA_signal_8034, new_AGEMA_signal_8033, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_9376, new_AGEMA_signal_9375, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_9740, new_AGEMA_signal_9739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L14_U1 ( .a ({new_AGEMA_signal_8508, new_AGEMA_signal_8507, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_8516, new_AGEMA_signal_8515, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_8990, new_AGEMA_signal_8989, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L15_U1 ( .a ({new_AGEMA_signal_8512, new_AGEMA_signal_8511, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55}), .b ({new_AGEMA_signal_8520, new_AGEMA_signal_8519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_8992, new_AGEMA_signal_8991, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L16_U1 ( .a ({new_AGEMA_signal_8038, new_AGEMA_signal_8037, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56}), .b ({new_AGEMA_signal_9376, new_AGEMA_signal_9375, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_9742, new_AGEMA_signal_9741, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L17_U1 ( .a ({new_AGEMA_signal_8040, new_AGEMA_signal_8039, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57}), .b ({new_AGEMA_signal_8520, new_AGEMA_signal_8519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_8994, new_AGEMA_signal_8993, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L18_U1 ( .a ({new_AGEMA_signal_8514, new_AGEMA_signal_8513, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58}), .b ({new_AGEMA_signal_8522, new_AGEMA_signal_8521, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8}), .c ({new_AGEMA_signal_8996, new_AGEMA_signal_8995, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L19_U1 ( .a ({new_AGEMA_signal_8518, new_AGEMA_signal_8517, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63}), .b ({new_AGEMA_signal_8986, new_AGEMA_signal_8985, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_9388, new_AGEMA_signal_9387, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L20_U1 ( .a ({new_AGEMA_signal_9376, new_AGEMA_signal_9375, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}), .b ({new_AGEMA_signal_8520, new_AGEMA_signal_8519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_9744, new_AGEMA_signal_9743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L21_U1 ( .a ({new_AGEMA_signal_8520, new_AGEMA_signal_8519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .b ({new_AGEMA_signal_9380, new_AGEMA_signal_9379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7}), .c ({new_AGEMA_signal_9746, new_AGEMA_signal_9745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L22_U1 ( .a ({new_AGEMA_signal_8984, new_AGEMA_signal_8983, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3}), .b ({new_AGEMA_signal_8524, new_AGEMA_signal_8523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12}), .c ({new_AGEMA_signal_9390, new_AGEMA_signal_9389, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L23_U1 ( .a ({new_AGEMA_signal_8996, new_AGEMA_signal_8995, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18}), .b ({new_AGEMA_signal_8982, new_AGEMA_signal_8981, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_9392, new_AGEMA_signal_9391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L24_U1 ( .a ({new_AGEMA_signal_8992, new_AGEMA_signal_8991, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15}), .b ({new_AGEMA_signal_9382, new_AGEMA_signal_9381, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_9748, new_AGEMA_signal_9747, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L25_U1 ( .a ({new_AGEMA_signal_9378, new_AGEMA_signal_9377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_9384, new_AGEMA_signal_9383, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_9750, new_AGEMA_signal_9749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L26_U1 ( .a ({new_AGEMA_signal_9380, new_AGEMA_signal_9379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7}), .b ({new_AGEMA_signal_9382, new_AGEMA_signal_9381, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_9752, new_AGEMA_signal_9751, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L27_U1 ( .a ({new_AGEMA_signal_8522, new_AGEMA_signal_8521, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8}), .b ({new_AGEMA_signal_9384, new_AGEMA_signal_9383, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_9754, new_AGEMA_signal_9753, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L28_U1 ( .a ({new_AGEMA_signal_9386, new_AGEMA_signal_9385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_8990, new_AGEMA_signal_8989, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14}), .c ({new_AGEMA_signal_9756, new_AGEMA_signal_9755, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L29_U1 ( .a ({new_AGEMA_signal_9386, new_AGEMA_signal_9385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_8994, new_AGEMA_signal_8993, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17}), .c ({new_AGEMA_signal_9758, new_AGEMA_signal_9757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S0_U1 ( .a ({new_AGEMA_signal_9378, new_AGEMA_signal_9377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_9748, new_AGEMA_signal_9747, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24}), .c ({new_AGEMA_signal_10180, new_AGEMA_signal_10179, KeyExpansionIns_tmp[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S1_U1 ( .a ({new_AGEMA_signal_9742, new_AGEMA_signal_9741, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16}), .b ({new_AGEMA_signal_9752, new_AGEMA_signal_9751, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26}), .c ({new_AGEMA_signal_10182, new_AGEMA_signal_10181, KeyExpansionIns_tmp[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S2_U1 ( .a ({new_AGEMA_signal_9388, new_AGEMA_signal_9387, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19}), .b ({new_AGEMA_signal_9756, new_AGEMA_signal_9755, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28}), .c ({new_AGEMA_signal_10184, new_AGEMA_signal_10183, KeyExpansionIns_tmp[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S3_U1 ( .a ({new_AGEMA_signal_9378, new_AGEMA_signal_9377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_9746, new_AGEMA_signal_9745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21}), .c ({new_AGEMA_signal_10186, new_AGEMA_signal_10185, KeyExpansionIns_tmp[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S4_U1 ( .a ({new_AGEMA_signal_9744, new_AGEMA_signal_9743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20}), .b ({new_AGEMA_signal_9390, new_AGEMA_signal_9389, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22}), .c ({new_AGEMA_signal_10188, new_AGEMA_signal_10187, KeyExpansionIns_tmp[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S5_U1 ( .a ({new_AGEMA_signal_9750, new_AGEMA_signal_9749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25}), .b ({new_AGEMA_signal_9758, new_AGEMA_signal_9757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29}), .c ({new_AGEMA_signal_10190, new_AGEMA_signal_10189, KeyExpansionIns_tmp[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S6_U1 ( .a ({new_AGEMA_signal_9740, new_AGEMA_signal_9739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13}), .b ({new_AGEMA_signal_9754, new_AGEMA_signal_9753, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27}), .c ({new_AGEMA_signal_10192, new_AGEMA_signal_10191, KeyExpansionIns_tmp[17]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S7_U1 ( .a ({new_AGEMA_signal_9378, new_AGEMA_signal_9377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_9392, new_AGEMA_signal_9391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23}), .c ({new_AGEMA_signal_9760, new_AGEMA_signal_9759, KeyExpansionIns_tmp[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M46_U1 ( .a ({new_AGEMA_signal_8052, new_AGEMA_signal_8051, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_5750, new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .clk (clk), .r ({Fresh[1934], Fresh[1933], Fresh[1932]}), .c ({new_AGEMA_signal_8528, new_AGEMA_signal_8527, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M47_U1 ( .a ({new_AGEMA_signal_7860, new_AGEMA_signal_7859, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_6090, new_AGEMA_signal_6089, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8}), .clk (clk), .r ({Fresh[1937], Fresh[1936], Fresh[1935]}), .c ({new_AGEMA_signal_8054, new_AGEMA_signal_8053, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M48_U1 ( .a ({new_AGEMA_signal_7858, new_AGEMA_signal_7857, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, RoundKey[0]}), .clk (clk), .r ({Fresh[1940], Fresh[1939], Fresh[1938]}), .c ({new_AGEMA_signal_8056, new_AGEMA_signal_8055, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M49_U1 ( .a ({new_AGEMA_signal_8050, new_AGEMA_signal_8049, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_5758, new_AGEMA_signal_5757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .clk (clk), .r ({Fresh[1943], Fresh[1942], Fresh[1941]}), .c ({new_AGEMA_signal_8530, new_AGEMA_signal_8529, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M50_U1 ( .a ({new_AGEMA_signal_7856, new_AGEMA_signal_7855, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_5752, new_AGEMA_signal_5751, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}), .clk (clk), .r ({Fresh[1946], Fresh[1945], Fresh[1944]}), .c ({new_AGEMA_signal_8058, new_AGEMA_signal_8057, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M51_U1 ( .a ({new_AGEMA_signal_7854, new_AGEMA_signal_7853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_6096, new_AGEMA_signal_6095, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}), .clk (clk), .r ({Fresh[1949], Fresh[1948], Fresh[1947]}), .c ({new_AGEMA_signal_8060, new_AGEMA_signal_8059, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M52_U1 ( .a ({new_AGEMA_signal_8048, new_AGEMA_signal_8047, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_5756, new_AGEMA_signal_5755, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15}), .clk (clk), .r ({Fresh[1952], Fresh[1951], Fresh[1950]}), .c ({new_AGEMA_signal_8532, new_AGEMA_signal_8531, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M53_U1 ( .a ({new_AGEMA_signal_8526, new_AGEMA_signal_8525, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_5764, new_AGEMA_signal_5763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27}), .clk (clk), .r ({Fresh[1955], Fresh[1954], Fresh[1953]}), .c ({new_AGEMA_signal_8998, new_AGEMA_signal_8997, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M54_U1 ( .a ({new_AGEMA_signal_8046, new_AGEMA_signal_8045, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_6092, new_AGEMA_signal_6091, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}), .clk (clk), .r ({Fresh[1958], Fresh[1957], Fresh[1956]}), .c ({new_AGEMA_signal_8534, new_AGEMA_signal_8533, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M55_U1 ( .a ({new_AGEMA_signal_8052, new_AGEMA_signal_8051, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_5754, new_AGEMA_signal_5753, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13}), .clk (clk), .r ({Fresh[1961], Fresh[1960], Fresh[1959]}), .c ({new_AGEMA_signal_8536, new_AGEMA_signal_8535, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M56_U1 ( .a ({new_AGEMA_signal_7860, new_AGEMA_signal_7859, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_6100, new_AGEMA_signal_6099, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23}), .clk (clk), .r ({Fresh[1964], Fresh[1963], Fresh[1962]}), .c ({new_AGEMA_signal_8062, new_AGEMA_signal_8061, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M57_U1 ( .a ({new_AGEMA_signal_7858, new_AGEMA_signal_7857, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_5760, new_AGEMA_signal_5759, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}), .clk (clk), .r ({Fresh[1967], Fresh[1966], Fresh[1965]}), .c ({new_AGEMA_signal_8064, new_AGEMA_signal_8063, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M58_U1 ( .a ({new_AGEMA_signal_8050, new_AGEMA_signal_8049, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_5362, new_AGEMA_signal_5361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .clk (clk), .r ({Fresh[1970], Fresh[1969], Fresh[1968]}), .c ({new_AGEMA_signal_8538, new_AGEMA_signal_8537, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M59_U1 ( .a ({new_AGEMA_signal_7856, new_AGEMA_signal_7855, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_5762, new_AGEMA_signal_5761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}), .clk (clk), .r ({Fresh[1973], Fresh[1972], Fresh[1971]}), .c ({new_AGEMA_signal_8066, new_AGEMA_signal_8065, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M60_U1 ( .a ({new_AGEMA_signal_7854, new_AGEMA_signal_7853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_6098, new_AGEMA_signal_6097, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}), .clk (clk), .r ({Fresh[1976], Fresh[1975], Fresh[1974]}), .c ({new_AGEMA_signal_8068, new_AGEMA_signal_8067, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M61_U1 ( .a ({new_AGEMA_signal_8048, new_AGEMA_signal_8047, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_5358, new_AGEMA_signal_5357, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .clk (clk), .r ({Fresh[1979], Fresh[1978], Fresh[1977]}), .c ({new_AGEMA_signal_8540, new_AGEMA_signal_8539, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M62_U1 ( .a ({new_AGEMA_signal_8526, new_AGEMA_signal_8525, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_5364, new_AGEMA_signal_5363, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}), .clk (clk), .r ({Fresh[1982], Fresh[1981], Fresh[1980]}), .c ({new_AGEMA_signal_9000, new_AGEMA_signal_8999, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M63_U1 ( .a ({new_AGEMA_signal_8046, new_AGEMA_signal_8045, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_5360, new_AGEMA_signal_5359, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .clk (clk), .r ({Fresh[1985], Fresh[1984], Fresh[1983]}), .c ({new_AGEMA_signal_8542, new_AGEMA_signal_8541, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L0_U1 ( .a ({new_AGEMA_signal_8540, new_AGEMA_signal_8539, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}), .b ({new_AGEMA_signal_9000, new_AGEMA_signal_8999, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62}), .c ({new_AGEMA_signal_9394, new_AGEMA_signal_9393, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L1_U1 ( .a ({new_AGEMA_signal_8058, new_AGEMA_signal_8057, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_8062, new_AGEMA_signal_8061, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56}), .c ({new_AGEMA_signal_8544, new_AGEMA_signal_8543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L2_U1 ( .a ({new_AGEMA_signal_8528, new_AGEMA_signal_8527, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_8056, new_AGEMA_signal_8055, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48}), .c ({new_AGEMA_signal_9002, new_AGEMA_signal_9001, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L3_U1 ( .a ({new_AGEMA_signal_8054, new_AGEMA_signal_8053, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47}), .b ({new_AGEMA_signal_8536, new_AGEMA_signal_8535, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55}), .c ({new_AGEMA_signal_9004, new_AGEMA_signal_9003, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L4_U1 ( .a ({new_AGEMA_signal_8534, new_AGEMA_signal_8533, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54}), .b ({new_AGEMA_signal_8538, new_AGEMA_signal_8537, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58}), .c ({new_AGEMA_signal_9006, new_AGEMA_signal_9005, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L5_U1 ( .a ({new_AGEMA_signal_8530, new_AGEMA_signal_8529, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49}), .b ({new_AGEMA_signal_8540, new_AGEMA_signal_8539, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_9008, new_AGEMA_signal_9007, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L6_U1 ( .a ({new_AGEMA_signal_9000, new_AGEMA_signal_8999, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62}), .b ({new_AGEMA_signal_9008, new_AGEMA_signal_9007, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5}), .c ({new_AGEMA_signal_9396, new_AGEMA_signal_9395, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L7_U1 ( .a ({new_AGEMA_signal_8528, new_AGEMA_signal_8527, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_9004, new_AGEMA_signal_9003, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3}), .c ({new_AGEMA_signal_9398, new_AGEMA_signal_9397, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L8_U1 ( .a ({new_AGEMA_signal_8060, new_AGEMA_signal_8059, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51}), .b ({new_AGEMA_signal_8066, new_AGEMA_signal_8065, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59}), .c ({new_AGEMA_signal_8546, new_AGEMA_signal_8545, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L9_U1 ( .a ({new_AGEMA_signal_8532, new_AGEMA_signal_8531, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_8998, new_AGEMA_signal_8997, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53}), .c ({new_AGEMA_signal_9400, new_AGEMA_signal_9399, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L10_U1 ( .a ({new_AGEMA_signal_8998, new_AGEMA_signal_8997, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53}), .b ({new_AGEMA_signal_9006, new_AGEMA_signal_9005, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_9402, new_AGEMA_signal_9401, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L11_U1 ( .a ({new_AGEMA_signal_8068, new_AGEMA_signal_8067, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60}), .b ({new_AGEMA_signal_9002, new_AGEMA_signal_9001, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_9404, new_AGEMA_signal_9403, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L12_U1 ( .a ({new_AGEMA_signal_8056, new_AGEMA_signal_8055, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48}), .b ({new_AGEMA_signal_8060, new_AGEMA_signal_8059, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51}), .c ({new_AGEMA_signal_8548, new_AGEMA_signal_8547, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L13_U1 ( .a ({new_AGEMA_signal_8058, new_AGEMA_signal_8057, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_9394, new_AGEMA_signal_9393, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_9762, new_AGEMA_signal_9761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L14_U1 ( .a ({new_AGEMA_signal_8532, new_AGEMA_signal_8531, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_8540, new_AGEMA_signal_8539, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_9010, new_AGEMA_signal_9009, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L15_U1 ( .a ({new_AGEMA_signal_8536, new_AGEMA_signal_8535, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55}), .b ({new_AGEMA_signal_8544, new_AGEMA_signal_8543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_9012, new_AGEMA_signal_9011, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L16_U1 ( .a ({new_AGEMA_signal_8062, new_AGEMA_signal_8061, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56}), .b ({new_AGEMA_signal_9394, new_AGEMA_signal_9393, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_9764, new_AGEMA_signal_9763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L17_U1 ( .a ({new_AGEMA_signal_8064, new_AGEMA_signal_8063, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57}), .b ({new_AGEMA_signal_8544, new_AGEMA_signal_8543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_9014, new_AGEMA_signal_9013, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L18_U1 ( .a ({new_AGEMA_signal_8538, new_AGEMA_signal_8537, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58}), .b ({new_AGEMA_signal_8546, new_AGEMA_signal_8545, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8}), .c ({new_AGEMA_signal_9016, new_AGEMA_signal_9015, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L19_U1 ( .a ({new_AGEMA_signal_8542, new_AGEMA_signal_8541, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63}), .b ({new_AGEMA_signal_9006, new_AGEMA_signal_9005, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_9406, new_AGEMA_signal_9405, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L20_U1 ( .a ({new_AGEMA_signal_9394, new_AGEMA_signal_9393, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}), .b ({new_AGEMA_signal_8544, new_AGEMA_signal_8543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_9766, new_AGEMA_signal_9765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L21_U1 ( .a ({new_AGEMA_signal_8544, new_AGEMA_signal_8543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .b ({new_AGEMA_signal_9398, new_AGEMA_signal_9397, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7}), .c ({new_AGEMA_signal_9768, new_AGEMA_signal_9767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L22_U1 ( .a ({new_AGEMA_signal_9004, new_AGEMA_signal_9003, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3}), .b ({new_AGEMA_signal_8548, new_AGEMA_signal_8547, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12}), .c ({new_AGEMA_signal_9408, new_AGEMA_signal_9407, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L23_U1 ( .a ({new_AGEMA_signal_9016, new_AGEMA_signal_9015, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18}), .b ({new_AGEMA_signal_9002, new_AGEMA_signal_9001, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_9410, new_AGEMA_signal_9409, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L24_U1 ( .a ({new_AGEMA_signal_9012, new_AGEMA_signal_9011, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15}), .b ({new_AGEMA_signal_9400, new_AGEMA_signal_9399, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_9770, new_AGEMA_signal_9769, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L25_U1 ( .a ({new_AGEMA_signal_9396, new_AGEMA_signal_9395, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_9402, new_AGEMA_signal_9401, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_9772, new_AGEMA_signal_9771, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L26_U1 ( .a ({new_AGEMA_signal_9398, new_AGEMA_signal_9397, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7}), .b ({new_AGEMA_signal_9400, new_AGEMA_signal_9399, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_9774, new_AGEMA_signal_9773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L27_U1 ( .a ({new_AGEMA_signal_8546, new_AGEMA_signal_8545, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8}), .b ({new_AGEMA_signal_9402, new_AGEMA_signal_9401, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_9776, new_AGEMA_signal_9775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L28_U1 ( .a ({new_AGEMA_signal_9404, new_AGEMA_signal_9403, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_9010, new_AGEMA_signal_9009, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14}), .c ({new_AGEMA_signal_9778, new_AGEMA_signal_9777, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L29_U1 ( .a ({new_AGEMA_signal_9404, new_AGEMA_signal_9403, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_9014, new_AGEMA_signal_9013, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17}), .c ({new_AGEMA_signal_9780, new_AGEMA_signal_9779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S0_U1 ( .a ({new_AGEMA_signal_9396, new_AGEMA_signal_9395, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_9770, new_AGEMA_signal_9769, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24}), .c ({new_AGEMA_signal_10194, new_AGEMA_signal_10193, KeyExpansionIns_tmp[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S1_U1 ( .a ({new_AGEMA_signal_9764, new_AGEMA_signal_9763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16}), .b ({new_AGEMA_signal_9774, new_AGEMA_signal_9773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26}), .c ({new_AGEMA_signal_10196, new_AGEMA_signal_10195, KeyExpansionIns_tmp[14]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S2_U1 ( .a ({new_AGEMA_signal_9406, new_AGEMA_signal_9405, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19}), .b ({new_AGEMA_signal_9778, new_AGEMA_signal_9777, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28}), .c ({new_AGEMA_signal_10198, new_AGEMA_signal_10197, KeyExpansionIns_tmp[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S3_U1 ( .a ({new_AGEMA_signal_9396, new_AGEMA_signal_9395, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_9768, new_AGEMA_signal_9767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21}), .c ({new_AGEMA_signal_10200, new_AGEMA_signal_10199, KeyExpansionIns_tmp[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S4_U1 ( .a ({new_AGEMA_signal_9766, new_AGEMA_signal_9765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20}), .b ({new_AGEMA_signal_9408, new_AGEMA_signal_9407, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22}), .c ({new_AGEMA_signal_10202, new_AGEMA_signal_10201, KeyExpansionIns_tmp[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S5_U1 ( .a ({new_AGEMA_signal_9772, new_AGEMA_signal_9771, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25}), .b ({new_AGEMA_signal_9780, new_AGEMA_signal_9779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29}), .c ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, KeyExpansionIns_tmp[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S6_U1 ( .a ({new_AGEMA_signal_9762, new_AGEMA_signal_9761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13}), .b ({new_AGEMA_signal_9776, new_AGEMA_signal_9775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27}), .c ({new_AGEMA_signal_10206, new_AGEMA_signal_10205, KeyExpansionIns_tmp[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S7_U1 ( .a ({new_AGEMA_signal_9396, new_AGEMA_signal_9395, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_9410, new_AGEMA_signal_9409, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23}), .c ({new_AGEMA_signal_9782, new_AGEMA_signal_9781, KeyExpansionIns_tmp[8]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M46_U1 ( .a ({new_AGEMA_signal_8076, new_AGEMA_signal_8075, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .clk (clk), .r ({Fresh[1988], Fresh[1987], Fresh[1986]}), .c ({new_AGEMA_signal_8552, new_AGEMA_signal_8551, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M47_U1 ( .a ({new_AGEMA_signal_7868, new_AGEMA_signal_7867, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_6116, new_AGEMA_signal_6115, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8}), .clk (clk), .r ({Fresh[1991], Fresh[1990], Fresh[1989]}), .c ({new_AGEMA_signal_8078, new_AGEMA_signal_8077, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M48_U1 ( .a ({new_AGEMA_signal_7866, new_AGEMA_signal_7865, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, RoundKey[24]}), .clk (clk), .r ({Fresh[1994], Fresh[1993], Fresh[1992]}), .c ({new_AGEMA_signal_8080, new_AGEMA_signal_8079, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M49_U1 ( .a ({new_AGEMA_signal_8074, new_AGEMA_signal_8073, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_5774, new_AGEMA_signal_5773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .clk (clk), .r ({Fresh[1997], Fresh[1996], Fresh[1995]}), .c ({new_AGEMA_signal_8554, new_AGEMA_signal_8553, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M50_U1 ( .a ({new_AGEMA_signal_7864, new_AGEMA_signal_7863, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_5768, new_AGEMA_signal_5767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}), .clk (clk), .r ({Fresh[2000], Fresh[1999], Fresh[1998]}), .c ({new_AGEMA_signal_8082, new_AGEMA_signal_8081, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M51_U1 ( .a ({new_AGEMA_signal_7862, new_AGEMA_signal_7861, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_6122, new_AGEMA_signal_6121, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}), .clk (clk), .r ({Fresh[2003], Fresh[2002], Fresh[2001]}), .c ({new_AGEMA_signal_8084, new_AGEMA_signal_8083, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M52_U1 ( .a ({new_AGEMA_signal_8072, new_AGEMA_signal_8071, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_5772, new_AGEMA_signal_5771, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15}), .clk (clk), .r ({Fresh[2006], Fresh[2005], Fresh[2004]}), .c ({new_AGEMA_signal_8556, new_AGEMA_signal_8555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M53_U1 ( .a ({new_AGEMA_signal_8550, new_AGEMA_signal_8549, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_5780, new_AGEMA_signal_5779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27}), .clk (clk), .r ({Fresh[2009], Fresh[2008], Fresh[2007]}), .c ({new_AGEMA_signal_9018, new_AGEMA_signal_9017, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M54_U1 ( .a ({new_AGEMA_signal_8070, new_AGEMA_signal_8069, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_6118, new_AGEMA_signal_6117, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}), .clk (clk), .r ({Fresh[2012], Fresh[2011], Fresh[2010]}), .c ({new_AGEMA_signal_8558, new_AGEMA_signal_8557, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M55_U1 ( .a ({new_AGEMA_signal_8076, new_AGEMA_signal_8075, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_5770, new_AGEMA_signal_5769, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13}), .clk (clk), .r ({Fresh[2015], Fresh[2014], Fresh[2013]}), .c ({new_AGEMA_signal_8560, new_AGEMA_signal_8559, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M56_U1 ( .a ({new_AGEMA_signal_7868, new_AGEMA_signal_7867, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_6126, new_AGEMA_signal_6125, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23}), .clk (clk), .r ({Fresh[2018], Fresh[2017], Fresh[2016]}), .c ({new_AGEMA_signal_8086, new_AGEMA_signal_8085, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M57_U1 ( .a ({new_AGEMA_signal_7866, new_AGEMA_signal_7865, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_5776, new_AGEMA_signal_5775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}), .clk (clk), .r ({Fresh[2021], Fresh[2020], Fresh[2019]}), .c ({new_AGEMA_signal_8088, new_AGEMA_signal_8087, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M58_U1 ( .a ({new_AGEMA_signal_8074, new_AGEMA_signal_8073, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_5382, new_AGEMA_signal_5381, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .clk (clk), .r ({Fresh[2024], Fresh[2023], Fresh[2022]}), .c ({new_AGEMA_signal_8562, new_AGEMA_signal_8561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M59_U1 ( .a ({new_AGEMA_signal_7864, new_AGEMA_signal_7863, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_5778, new_AGEMA_signal_5777, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}), .clk (clk), .r ({Fresh[2027], Fresh[2026], Fresh[2025]}), .c ({new_AGEMA_signal_8090, new_AGEMA_signal_8089, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M60_U1 ( .a ({new_AGEMA_signal_7862, new_AGEMA_signal_7861, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_6124, new_AGEMA_signal_6123, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}), .clk (clk), .r ({Fresh[2030], Fresh[2029], Fresh[2028]}), .c ({new_AGEMA_signal_8092, new_AGEMA_signal_8091, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M61_U1 ( .a ({new_AGEMA_signal_8072, new_AGEMA_signal_8071, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_5378, new_AGEMA_signal_5377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .clk (clk), .r ({Fresh[2033], Fresh[2032], Fresh[2031]}), .c ({new_AGEMA_signal_8564, new_AGEMA_signal_8563, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M62_U1 ( .a ({new_AGEMA_signal_8550, new_AGEMA_signal_8549, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_5384, new_AGEMA_signal_5383, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}), .clk (clk), .r ({Fresh[2036], Fresh[2035], Fresh[2034]}), .c ({new_AGEMA_signal_9020, new_AGEMA_signal_9019, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M63_U1 ( .a ({new_AGEMA_signal_8070, new_AGEMA_signal_8069, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_5380, new_AGEMA_signal_5379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .clk (clk), .r ({Fresh[2039], Fresh[2038], Fresh[2037]}), .c ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L0_U1 ( .a ({new_AGEMA_signal_8564, new_AGEMA_signal_8563, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}), .b ({new_AGEMA_signal_9020, new_AGEMA_signal_9019, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62}), .c ({new_AGEMA_signal_9412, new_AGEMA_signal_9411, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L1_U1 ( .a ({new_AGEMA_signal_8082, new_AGEMA_signal_8081, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_8086, new_AGEMA_signal_8085, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56}), .c ({new_AGEMA_signal_8568, new_AGEMA_signal_8567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L2_U1 ( .a ({new_AGEMA_signal_8552, new_AGEMA_signal_8551, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_8080, new_AGEMA_signal_8079, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48}), .c ({new_AGEMA_signal_9022, new_AGEMA_signal_9021, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L3_U1 ( .a ({new_AGEMA_signal_8078, new_AGEMA_signal_8077, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47}), .b ({new_AGEMA_signal_8560, new_AGEMA_signal_8559, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55}), .c ({new_AGEMA_signal_9024, new_AGEMA_signal_9023, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L4_U1 ( .a ({new_AGEMA_signal_8558, new_AGEMA_signal_8557, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54}), .b ({new_AGEMA_signal_8562, new_AGEMA_signal_8561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58}), .c ({new_AGEMA_signal_9026, new_AGEMA_signal_9025, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L5_U1 ( .a ({new_AGEMA_signal_8554, new_AGEMA_signal_8553, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49}), .b ({new_AGEMA_signal_8564, new_AGEMA_signal_8563, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_9028, new_AGEMA_signal_9027, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L6_U1 ( .a ({new_AGEMA_signal_9020, new_AGEMA_signal_9019, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62}), .b ({new_AGEMA_signal_9028, new_AGEMA_signal_9027, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5}), .c ({new_AGEMA_signal_9414, new_AGEMA_signal_9413, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L7_U1 ( .a ({new_AGEMA_signal_8552, new_AGEMA_signal_8551, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_9024, new_AGEMA_signal_9023, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3}), .c ({new_AGEMA_signal_9416, new_AGEMA_signal_9415, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L8_U1 ( .a ({new_AGEMA_signal_8084, new_AGEMA_signal_8083, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51}), .b ({new_AGEMA_signal_8090, new_AGEMA_signal_8089, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59}), .c ({new_AGEMA_signal_8570, new_AGEMA_signal_8569, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L9_U1 ( .a ({new_AGEMA_signal_8556, new_AGEMA_signal_8555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_9018, new_AGEMA_signal_9017, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53}), .c ({new_AGEMA_signal_9418, new_AGEMA_signal_9417, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L10_U1 ( .a ({new_AGEMA_signal_9018, new_AGEMA_signal_9017, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53}), .b ({new_AGEMA_signal_9026, new_AGEMA_signal_9025, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_9420, new_AGEMA_signal_9419, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L11_U1 ( .a ({new_AGEMA_signal_8092, new_AGEMA_signal_8091, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60}), .b ({new_AGEMA_signal_9022, new_AGEMA_signal_9021, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_9422, new_AGEMA_signal_9421, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L12_U1 ( .a ({new_AGEMA_signal_8080, new_AGEMA_signal_8079, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48}), .b ({new_AGEMA_signal_8084, new_AGEMA_signal_8083, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51}), .c ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L13_U1 ( .a ({new_AGEMA_signal_8082, new_AGEMA_signal_8081, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_9412, new_AGEMA_signal_9411, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_9784, new_AGEMA_signal_9783, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L14_U1 ( .a ({new_AGEMA_signal_8556, new_AGEMA_signal_8555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_8564, new_AGEMA_signal_8563, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_9030, new_AGEMA_signal_9029, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L15_U1 ( .a ({new_AGEMA_signal_8560, new_AGEMA_signal_8559, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55}), .b ({new_AGEMA_signal_8568, new_AGEMA_signal_8567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_9032, new_AGEMA_signal_9031, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L16_U1 ( .a ({new_AGEMA_signal_8086, new_AGEMA_signal_8085, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56}), .b ({new_AGEMA_signal_9412, new_AGEMA_signal_9411, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_9786, new_AGEMA_signal_9785, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L17_U1 ( .a ({new_AGEMA_signal_8088, new_AGEMA_signal_8087, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57}), .b ({new_AGEMA_signal_8568, new_AGEMA_signal_8567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_9034, new_AGEMA_signal_9033, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L18_U1 ( .a ({new_AGEMA_signal_8562, new_AGEMA_signal_8561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58}), .b ({new_AGEMA_signal_8570, new_AGEMA_signal_8569, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8}), .c ({new_AGEMA_signal_9036, new_AGEMA_signal_9035, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L19_U1 ( .a ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63}), .b ({new_AGEMA_signal_9026, new_AGEMA_signal_9025, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_9424, new_AGEMA_signal_9423, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L20_U1 ( .a ({new_AGEMA_signal_9412, new_AGEMA_signal_9411, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}), .b ({new_AGEMA_signal_8568, new_AGEMA_signal_8567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_9788, new_AGEMA_signal_9787, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L21_U1 ( .a ({new_AGEMA_signal_8568, new_AGEMA_signal_8567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .b ({new_AGEMA_signal_9416, new_AGEMA_signal_9415, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7}), .c ({new_AGEMA_signal_9790, new_AGEMA_signal_9789, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L22_U1 ( .a ({new_AGEMA_signal_9024, new_AGEMA_signal_9023, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3}), .b ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12}), .c ({new_AGEMA_signal_9426, new_AGEMA_signal_9425, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L23_U1 ( .a ({new_AGEMA_signal_9036, new_AGEMA_signal_9035, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18}), .b ({new_AGEMA_signal_9022, new_AGEMA_signal_9021, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_9428, new_AGEMA_signal_9427, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L24_U1 ( .a ({new_AGEMA_signal_9032, new_AGEMA_signal_9031, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15}), .b ({new_AGEMA_signal_9418, new_AGEMA_signal_9417, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_9792, new_AGEMA_signal_9791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L25_U1 ( .a ({new_AGEMA_signal_9414, new_AGEMA_signal_9413, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_9420, new_AGEMA_signal_9419, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_9794, new_AGEMA_signal_9793, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L26_U1 ( .a ({new_AGEMA_signal_9416, new_AGEMA_signal_9415, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7}), .b ({new_AGEMA_signal_9418, new_AGEMA_signal_9417, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_9796, new_AGEMA_signal_9795, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L27_U1 ( .a ({new_AGEMA_signal_8570, new_AGEMA_signal_8569, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8}), .b ({new_AGEMA_signal_9420, new_AGEMA_signal_9419, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_9798, new_AGEMA_signal_9797, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L28_U1 ( .a ({new_AGEMA_signal_9422, new_AGEMA_signal_9421, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_9030, new_AGEMA_signal_9029, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14}), .c ({new_AGEMA_signal_9800, new_AGEMA_signal_9799, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L29_U1 ( .a ({new_AGEMA_signal_9422, new_AGEMA_signal_9421, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_9034, new_AGEMA_signal_9033, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17}), .c ({new_AGEMA_signal_9802, new_AGEMA_signal_9801, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S0_U1 ( .a ({new_AGEMA_signal_9414, new_AGEMA_signal_9413, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_9792, new_AGEMA_signal_9791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24}), .c ({new_AGEMA_signal_10208, new_AGEMA_signal_10207, KeyExpansionIns_tmp[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S1_U1 ( .a ({new_AGEMA_signal_9786, new_AGEMA_signal_9785, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16}), .b ({new_AGEMA_signal_9796, new_AGEMA_signal_9795, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26}), .c ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, KeyExpansionIns_tmp[6]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S2_U1 ( .a ({new_AGEMA_signal_9424, new_AGEMA_signal_9423, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19}), .b ({new_AGEMA_signal_9800, new_AGEMA_signal_9799, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28}), .c ({new_AGEMA_signal_10212, new_AGEMA_signal_10211, KeyExpansionIns_tmp[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S3_U1 ( .a ({new_AGEMA_signal_9414, new_AGEMA_signal_9413, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_9790, new_AGEMA_signal_9789, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21}), .c ({new_AGEMA_signal_10214, new_AGEMA_signal_10213, KeyExpansionIns_tmp[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S4_U1 ( .a ({new_AGEMA_signal_9788, new_AGEMA_signal_9787, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20}), .b ({new_AGEMA_signal_9426, new_AGEMA_signal_9425, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22}), .c ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, KeyExpansionIns_tmp[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S5_U1 ( .a ({new_AGEMA_signal_9794, new_AGEMA_signal_9793, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25}), .b ({new_AGEMA_signal_9802, new_AGEMA_signal_9801, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29}), .c ({new_AGEMA_signal_10218, new_AGEMA_signal_10217, KeyExpansionIns_tmp[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S6_U1 ( .a ({new_AGEMA_signal_9784, new_AGEMA_signal_9783, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13}), .b ({new_AGEMA_signal_9798, new_AGEMA_signal_9797, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27}), .c ({new_AGEMA_signal_10220, new_AGEMA_signal_10219, KeyExpansionIns_tmp[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S7_U1 ( .a ({new_AGEMA_signal_9414, new_AGEMA_signal_9413, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_9428, new_AGEMA_signal_9427, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23}), .c ({new_AGEMA_signal_9804, new_AGEMA_signal_9803, KeyExpansionIns_tmp[0]}) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12316, new_AGEMA_signal_12315, RoundReg_Inst_ff_SDE_0_next_state}), .Q ({new_AGEMA_signal_4550, new_AGEMA_signal_4549, RoundInput[0]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12664, new_AGEMA_signal_12663, RoundReg_Inst_ff_SDE_1_next_state}), .Q ({new_AGEMA_signal_4784, new_AGEMA_signal_4783, RoundInput[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12320, new_AGEMA_signal_12319, RoundReg_Inst_ff_SDE_2_next_state}), .Q ({new_AGEMA_signal_4850, new_AGEMA_signal_4849, RoundInput[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12668, new_AGEMA_signal_12667, RoundReg_Inst_ff_SDE_3_next_state}), .Q ({new_AGEMA_signal_4916, new_AGEMA_signal_4915, RoundInput[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12672, new_AGEMA_signal_12671, RoundReg_Inst_ff_SDE_4_next_state}), .Q ({new_AGEMA_signal_4982, new_AGEMA_signal_4981, RoundInput[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12324, new_AGEMA_signal_12323, RoundReg_Inst_ff_SDE_5_next_state}), .Q ({new_AGEMA_signal_5048, new_AGEMA_signal_5047, RoundInput[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12328, new_AGEMA_signal_12327, RoundReg_Inst_ff_SDE_6_next_state}), .Q ({new_AGEMA_signal_5114, new_AGEMA_signal_5113, RoundInput[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12332, new_AGEMA_signal_12331, RoundReg_Inst_ff_SDE_7_next_state}), .Q ({new_AGEMA_signal_5180, new_AGEMA_signal_5179, RoundInput[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12336, new_AGEMA_signal_12335, RoundReg_Inst_ff_SDE_8_next_state}), .Q ({new_AGEMA_signal_5246, new_AGEMA_signal_5245, RoundInput[8]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12676, new_AGEMA_signal_12675, RoundReg_Inst_ff_SDE_9_next_state}), .Q ({new_AGEMA_signal_5312, new_AGEMA_signal_5311, RoundInput[9]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12340, new_AGEMA_signal_12339, RoundReg_Inst_ff_SDE_10_next_state}), .Q ({new_AGEMA_signal_4616, new_AGEMA_signal_4615, RoundInput[10]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12680, new_AGEMA_signal_12679, RoundReg_Inst_ff_SDE_11_next_state}), .Q ({new_AGEMA_signal_4682, new_AGEMA_signal_4681, RoundInput[11]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12684, new_AGEMA_signal_12683, RoundReg_Inst_ff_SDE_12_next_state}), .Q ({new_AGEMA_signal_4736, new_AGEMA_signal_4735, RoundInput[12]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12344, new_AGEMA_signal_12343, RoundReg_Inst_ff_SDE_13_next_state}), .Q ({new_AGEMA_signal_4742, new_AGEMA_signal_4741, RoundInput[13]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12348, new_AGEMA_signal_12347, RoundReg_Inst_ff_SDE_14_next_state}), .Q ({new_AGEMA_signal_4748, new_AGEMA_signal_4747, RoundInput[14]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12352, new_AGEMA_signal_12351, RoundReg_Inst_ff_SDE_15_next_state}), .Q ({new_AGEMA_signal_4754, new_AGEMA_signal_4753, RoundInput[15]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12356, new_AGEMA_signal_12355, RoundReg_Inst_ff_SDE_16_next_state}), .Q ({new_AGEMA_signal_4760, new_AGEMA_signal_4759, RoundInput[16]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12688, new_AGEMA_signal_12687, RoundReg_Inst_ff_SDE_17_next_state}), .Q ({new_AGEMA_signal_4766, new_AGEMA_signal_4765, RoundInput[17]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12360, new_AGEMA_signal_12359, RoundReg_Inst_ff_SDE_18_next_state}), .Q ({new_AGEMA_signal_4772, new_AGEMA_signal_4771, RoundInput[18]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12692, new_AGEMA_signal_12691, RoundReg_Inst_ff_SDE_19_next_state}), .Q ({new_AGEMA_signal_4778, new_AGEMA_signal_4777, RoundInput[19]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12696, new_AGEMA_signal_12695, RoundReg_Inst_ff_SDE_20_next_state}), .Q ({new_AGEMA_signal_4790, new_AGEMA_signal_4789, RoundInput[20]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12364, new_AGEMA_signal_12363, RoundReg_Inst_ff_SDE_21_next_state}), .Q ({new_AGEMA_signal_4796, new_AGEMA_signal_4795, RoundInput[21]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12368, new_AGEMA_signal_12367, RoundReg_Inst_ff_SDE_22_next_state}), .Q ({new_AGEMA_signal_4802, new_AGEMA_signal_4801, RoundInput[22]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12372, new_AGEMA_signal_12371, RoundReg_Inst_ff_SDE_23_next_state}), .Q ({new_AGEMA_signal_4808, new_AGEMA_signal_4807, RoundInput[23]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12376, new_AGEMA_signal_12375, RoundReg_Inst_ff_SDE_24_next_state}), .Q ({new_AGEMA_signal_4814, new_AGEMA_signal_4813, RoundInput[24]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12700, new_AGEMA_signal_12699, RoundReg_Inst_ff_SDE_25_next_state}), .Q ({new_AGEMA_signal_4820, new_AGEMA_signal_4819, RoundInput[25]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12380, new_AGEMA_signal_12379, RoundReg_Inst_ff_SDE_26_next_state}), .Q ({new_AGEMA_signal_4826, new_AGEMA_signal_4825, RoundInput[26]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12704, new_AGEMA_signal_12703, RoundReg_Inst_ff_SDE_27_next_state}), .Q ({new_AGEMA_signal_4832, new_AGEMA_signal_4831, RoundInput[27]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12708, new_AGEMA_signal_12707, RoundReg_Inst_ff_SDE_28_next_state}), .Q ({new_AGEMA_signal_4838, new_AGEMA_signal_4837, RoundInput[28]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12384, new_AGEMA_signal_12383, RoundReg_Inst_ff_SDE_29_next_state}), .Q ({new_AGEMA_signal_4844, new_AGEMA_signal_4843, RoundInput[29]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12388, new_AGEMA_signal_12387, RoundReg_Inst_ff_SDE_30_next_state}), .Q ({new_AGEMA_signal_4856, new_AGEMA_signal_4855, RoundInput[30]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12392, new_AGEMA_signal_12391, RoundReg_Inst_ff_SDE_31_next_state}), .Q ({new_AGEMA_signal_4862, new_AGEMA_signal_4861, RoundInput[31]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12396, new_AGEMA_signal_12395, RoundReg_Inst_ff_SDE_32_next_state}), .Q ({new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundInput[32]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12712, new_AGEMA_signal_12711, RoundReg_Inst_ff_SDE_33_next_state}), .Q ({new_AGEMA_signal_4874, new_AGEMA_signal_4873, RoundInput[33]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12400, new_AGEMA_signal_12399, RoundReg_Inst_ff_SDE_34_next_state}), .Q ({new_AGEMA_signal_4880, new_AGEMA_signal_4879, RoundInput[34]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12716, new_AGEMA_signal_12715, RoundReg_Inst_ff_SDE_35_next_state}), .Q ({new_AGEMA_signal_4886, new_AGEMA_signal_4885, RoundInput[35]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12720, new_AGEMA_signal_12719, RoundReg_Inst_ff_SDE_36_next_state}), .Q ({new_AGEMA_signal_4892, new_AGEMA_signal_4891, RoundInput[36]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12404, new_AGEMA_signal_12403, RoundReg_Inst_ff_SDE_37_next_state}), .Q ({new_AGEMA_signal_4898, new_AGEMA_signal_4897, RoundInput[37]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12408, new_AGEMA_signal_12407, RoundReg_Inst_ff_SDE_38_next_state}), .Q ({new_AGEMA_signal_4904, new_AGEMA_signal_4903, RoundInput[38]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12412, new_AGEMA_signal_12411, RoundReg_Inst_ff_SDE_39_next_state}), .Q ({new_AGEMA_signal_4910, new_AGEMA_signal_4909, RoundInput[39]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12416, new_AGEMA_signal_12415, RoundReg_Inst_ff_SDE_40_next_state}), .Q ({new_AGEMA_signal_4922, new_AGEMA_signal_4921, RoundInput[40]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12724, new_AGEMA_signal_12723, RoundReg_Inst_ff_SDE_41_next_state}), .Q ({new_AGEMA_signal_4928, new_AGEMA_signal_4927, RoundInput[41]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12420, new_AGEMA_signal_12419, RoundReg_Inst_ff_SDE_42_next_state}), .Q ({new_AGEMA_signal_4934, new_AGEMA_signal_4933, RoundInput[42]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12728, new_AGEMA_signal_12727, RoundReg_Inst_ff_SDE_43_next_state}), .Q ({new_AGEMA_signal_4940, new_AGEMA_signal_4939, RoundInput[43]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12732, new_AGEMA_signal_12731, RoundReg_Inst_ff_SDE_44_next_state}), .Q ({new_AGEMA_signal_4946, new_AGEMA_signal_4945, RoundInput[44]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12424, new_AGEMA_signal_12423, RoundReg_Inst_ff_SDE_45_next_state}), .Q ({new_AGEMA_signal_4952, new_AGEMA_signal_4951, RoundInput[45]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12428, new_AGEMA_signal_12427, RoundReg_Inst_ff_SDE_46_next_state}), .Q ({new_AGEMA_signal_4958, new_AGEMA_signal_4957, RoundInput[46]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12432, new_AGEMA_signal_12431, RoundReg_Inst_ff_SDE_47_next_state}), .Q ({new_AGEMA_signal_4964, new_AGEMA_signal_4963, RoundInput[47]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12436, new_AGEMA_signal_12435, RoundReg_Inst_ff_SDE_48_next_state}), .Q ({new_AGEMA_signal_4970, new_AGEMA_signal_4969, RoundInput[48]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12736, new_AGEMA_signal_12735, RoundReg_Inst_ff_SDE_49_next_state}), .Q ({new_AGEMA_signal_4976, new_AGEMA_signal_4975, RoundInput[49]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12440, new_AGEMA_signal_12439, RoundReg_Inst_ff_SDE_50_next_state}), .Q ({new_AGEMA_signal_4988, new_AGEMA_signal_4987, RoundInput[50]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12740, new_AGEMA_signal_12739, RoundReg_Inst_ff_SDE_51_next_state}), .Q ({new_AGEMA_signal_4994, new_AGEMA_signal_4993, RoundInput[51]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12744, new_AGEMA_signal_12743, RoundReg_Inst_ff_SDE_52_next_state}), .Q ({new_AGEMA_signal_5000, new_AGEMA_signal_4999, RoundInput[52]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12444, new_AGEMA_signal_12443, RoundReg_Inst_ff_SDE_53_next_state}), .Q ({new_AGEMA_signal_5006, new_AGEMA_signal_5005, RoundInput[53]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12448, new_AGEMA_signal_12447, RoundReg_Inst_ff_SDE_54_next_state}), .Q ({new_AGEMA_signal_5012, new_AGEMA_signal_5011, RoundInput[54]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12452, new_AGEMA_signal_12451, RoundReg_Inst_ff_SDE_55_next_state}), .Q ({new_AGEMA_signal_5018, new_AGEMA_signal_5017, RoundInput[55]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12456, new_AGEMA_signal_12455, RoundReg_Inst_ff_SDE_56_next_state}), .Q ({new_AGEMA_signal_5024, new_AGEMA_signal_5023, RoundInput[56]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12748, new_AGEMA_signal_12747, RoundReg_Inst_ff_SDE_57_next_state}), .Q ({new_AGEMA_signal_5030, new_AGEMA_signal_5029, RoundInput[57]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12460, new_AGEMA_signal_12459, RoundReg_Inst_ff_SDE_58_next_state}), .Q ({new_AGEMA_signal_5036, new_AGEMA_signal_5035, RoundInput[58]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12752, new_AGEMA_signal_12751, RoundReg_Inst_ff_SDE_59_next_state}), .Q ({new_AGEMA_signal_5042, new_AGEMA_signal_5041, RoundInput[59]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12756, new_AGEMA_signal_12755, RoundReg_Inst_ff_SDE_60_next_state}), .Q ({new_AGEMA_signal_5054, new_AGEMA_signal_5053, RoundInput[60]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12464, new_AGEMA_signal_12463, RoundReg_Inst_ff_SDE_61_next_state}), .Q ({new_AGEMA_signal_5060, new_AGEMA_signal_5059, RoundInput[61]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12468, new_AGEMA_signal_12467, RoundReg_Inst_ff_SDE_62_next_state}), .Q ({new_AGEMA_signal_5066, new_AGEMA_signal_5065, RoundInput[62]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12472, new_AGEMA_signal_12471, RoundReg_Inst_ff_SDE_63_next_state}), .Q ({new_AGEMA_signal_5072, new_AGEMA_signal_5071, RoundInput[63]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12476, new_AGEMA_signal_12475, RoundReg_Inst_ff_SDE_64_next_state}), .Q ({new_AGEMA_signal_5078, new_AGEMA_signal_5077, RoundInput[64]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12760, new_AGEMA_signal_12759, RoundReg_Inst_ff_SDE_65_next_state}), .Q ({new_AGEMA_signal_5084, new_AGEMA_signal_5083, RoundInput[65]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12480, new_AGEMA_signal_12479, RoundReg_Inst_ff_SDE_66_next_state}), .Q ({new_AGEMA_signal_5090, new_AGEMA_signal_5089, RoundInput[66]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12764, new_AGEMA_signal_12763, RoundReg_Inst_ff_SDE_67_next_state}), .Q ({new_AGEMA_signal_5096, new_AGEMA_signal_5095, RoundInput[67]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12768, new_AGEMA_signal_12767, RoundReg_Inst_ff_SDE_68_next_state}), .Q ({new_AGEMA_signal_5102, new_AGEMA_signal_5101, RoundInput[68]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12484, new_AGEMA_signal_12483, RoundReg_Inst_ff_SDE_69_next_state}), .Q ({new_AGEMA_signal_5108, new_AGEMA_signal_5107, RoundInput[69]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12488, new_AGEMA_signal_12487, RoundReg_Inst_ff_SDE_70_next_state}), .Q ({new_AGEMA_signal_5120, new_AGEMA_signal_5119, RoundInput[70]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12492, new_AGEMA_signal_12491, RoundReg_Inst_ff_SDE_71_next_state}), .Q ({new_AGEMA_signal_5126, new_AGEMA_signal_5125, RoundInput[71]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12496, new_AGEMA_signal_12495, RoundReg_Inst_ff_SDE_72_next_state}), .Q ({new_AGEMA_signal_5132, new_AGEMA_signal_5131, RoundInput[72]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12772, new_AGEMA_signal_12771, RoundReg_Inst_ff_SDE_73_next_state}), .Q ({new_AGEMA_signal_5138, new_AGEMA_signal_5137, RoundInput[73]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12500, new_AGEMA_signal_12499, RoundReg_Inst_ff_SDE_74_next_state}), .Q ({new_AGEMA_signal_5144, new_AGEMA_signal_5143, RoundInput[74]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12776, new_AGEMA_signal_12775, RoundReg_Inst_ff_SDE_75_next_state}), .Q ({new_AGEMA_signal_5150, new_AGEMA_signal_5149, RoundInput[75]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12780, new_AGEMA_signal_12779, RoundReg_Inst_ff_SDE_76_next_state}), .Q ({new_AGEMA_signal_5156, new_AGEMA_signal_5155, RoundInput[76]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12504, new_AGEMA_signal_12503, RoundReg_Inst_ff_SDE_77_next_state}), .Q ({new_AGEMA_signal_5162, new_AGEMA_signal_5161, RoundInput[77]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12508, new_AGEMA_signal_12507, RoundReg_Inst_ff_SDE_78_next_state}), .Q ({new_AGEMA_signal_5168, new_AGEMA_signal_5167, RoundInput[78]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12512, new_AGEMA_signal_12511, RoundReg_Inst_ff_SDE_79_next_state}), .Q ({new_AGEMA_signal_5174, new_AGEMA_signal_5173, RoundInput[79]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12516, new_AGEMA_signal_12515, RoundReg_Inst_ff_SDE_80_next_state}), .Q ({new_AGEMA_signal_5186, new_AGEMA_signal_5185, RoundInput[80]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12784, new_AGEMA_signal_12783, RoundReg_Inst_ff_SDE_81_next_state}), .Q ({new_AGEMA_signal_5192, new_AGEMA_signal_5191, RoundInput[81]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12520, new_AGEMA_signal_12519, RoundReg_Inst_ff_SDE_82_next_state}), .Q ({new_AGEMA_signal_5198, new_AGEMA_signal_5197, RoundInput[82]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12788, new_AGEMA_signal_12787, RoundReg_Inst_ff_SDE_83_next_state}), .Q ({new_AGEMA_signal_5204, new_AGEMA_signal_5203, RoundInput[83]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12792, new_AGEMA_signal_12791, RoundReg_Inst_ff_SDE_84_next_state}), .Q ({new_AGEMA_signal_5210, new_AGEMA_signal_5209, RoundInput[84]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12524, new_AGEMA_signal_12523, RoundReg_Inst_ff_SDE_85_next_state}), .Q ({new_AGEMA_signal_5216, new_AGEMA_signal_5215, RoundInput[85]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12528, new_AGEMA_signal_12527, RoundReg_Inst_ff_SDE_86_next_state}), .Q ({new_AGEMA_signal_5222, new_AGEMA_signal_5221, RoundInput[86]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12532, new_AGEMA_signal_12531, RoundReg_Inst_ff_SDE_87_next_state}), .Q ({new_AGEMA_signal_5228, new_AGEMA_signal_5227, RoundInput[87]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12536, new_AGEMA_signal_12535, RoundReg_Inst_ff_SDE_88_next_state}), .Q ({new_AGEMA_signal_5234, new_AGEMA_signal_5233, RoundInput[88]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12796, new_AGEMA_signal_12795, RoundReg_Inst_ff_SDE_89_next_state}), .Q ({new_AGEMA_signal_5240, new_AGEMA_signal_5239, RoundInput[89]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12540, new_AGEMA_signal_12539, RoundReg_Inst_ff_SDE_90_next_state}), .Q ({new_AGEMA_signal_5252, new_AGEMA_signal_5251, RoundInput[90]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12800, new_AGEMA_signal_12799, RoundReg_Inst_ff_SDE_91_next_state}), .Q ({new_AGEMA_signal_5258, new_AGEMA_signal_5257, RoundInput[91]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12804, new_AGEMA_signal_12803, RoundReg_Inst_ff_SDE_92_next_state}), .Q ({new_AGEMA_signal_5264, new_AGEMA_signal_5263, RoundInput[92]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12544, new_AGEMA_signal_12543, RoundReg_Inst_ff_SDE_93_next_state}), .Q ({new_AGEMA_signal_5270, new_AGEMA_signal_5269, RoundInput[93]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12548, new_AGEMA_signal_12547, RoundReg_Inst_ff_SDE_94_next_state}), .Q ({new_AGEMA_signal_5276, new_AGEMA_signal_5275, RoundInput[94]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12552, new_AGEMA_signal_12551, RoundReg_Inst_ff_SDE_95_next_state}), .Q ({new_AGEMA_signal_5282, new_AGEMA_signal_5281, RoundInput[95]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12556, new_AGEMA_signal_12555, RoundReg_Inst_ff_SDE_96_next_state}), .Q ({new_AGEMA_signal_5288, new_AGEMA_signal_5287, RoundInput[96]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12808, new_AGEMA_signal_12807, RoundReg_Inst_ff_SDE_97_next_state}), .Q ({new_AGEMA_signal_5294, new_AGEMA_signal_5293, RoundInput[97]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12560, new_AGEMA_signal_12559, RoundReg_Inst_ff_SDE_98_next_state}), .Q ({new_AGEMA_signal_5300, new_AGEMA_signal_5299, RoundInput[98]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12812, new_AGEMA_signal_12811, RoundReg_Inst_ff_SDE_99_next_state}), .Q ({new_AGEMA_signal_5306, new_AGEMA_signal_5305, RoundInput[99]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12816, new_AGEMA_signal_12815, RoundReg_Inst_ff_SDE_100_next_state}), .Q ({new_AGEMA_signal_4556, new_AGEMA_signal_4555, RoundInput[100]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12564, new_AGEMA_signal_12563, RoundReg_Inst_ff_SDE_101_next_state}), .Q ({new_AGEMA_signal_4562, new_AGEMA_signal_4561, RoundInput[101]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12568, new_AGEMA_signal_12567, RoundReg_Inst_ff_SDE_102_next_state}), .Q ({new_AGEMA_signal_4568, new_AGEMA_signal_4567, RoundInput[102]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12572, new_AGEMA_signal_12571, RoundReg_Inst_ff_SDE_103_next_state}), .Q ({new_AGEMA_signal_4574, new_AGEMA_signal_4573, RoundInput[103]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12576, new_AGEMA_signal_12575, RoundReg_Inst_ff_SDE_104_next_state}), .Q ({new_AGEMA_signal_4580, new_AGEMA_signal_4579, RoundInput[104]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, RoundReg_Inst_ff_SDE_105_next_state}), .Q ({new_AGEMA_signal_4586, new_AGEMA_signal_4585, RoundInput[105]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12580, new_AGEMA_signal_12579, RoundReg_Inst_ff_SDE_106_next_state}), .Q ({new_AGEMA_signal_4592, new_AGEMA_signal_4591, RoundInput[106]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12824, new_AGEMA_signal_12823, RoundReg_Inst_ff_SDE_107_next_state}), .Q ({new_AGEMA_signal_4598, new_AGEMA_signal_4597, RoundInput[107]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12828, new_AGEMA_signal_12827, RoundReg_Inst_ff_SDE_108_next_state}), .Q ({new_AGEMA_signal_4604, new_AGEMA_signal_4603, RoundInput[108]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12584, new_AGEMA_signal_12583, RoundReg_Inst_ff_SDE_109_next_state}), .Q ({new_AGEMA_signal_4610, new_AGEMA_signal_4609, RoundInput[109]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12588, new_AGEMA_signal_12587, RoundReg_Inst_ff_SDE_110_next_state}), .Q ({new_AGEMA_signal_4622, new_AGEMA_signal_4621, RoundInput[110]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12592, new_AGEMA_signal_12591, RoundReg_Inst_ff_SDE_111_next_state}), .Q ({new_AGEMA_signal_4628, new_AGEMA_signal_4627, RoundInput[111]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12596, new_AGEMA_signal_12595, RoundReg_Inst_ff_SDE_112_next_state}), .Q ({new_AGEMA_signal_4634, new_AGEMA_signal_4633, RoundInput[112]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, RoundReg_Inst_ff_SDE_113_next_state}), .Q ({new_AGEMA_signal_4640, new_AGEMA_signal_4639, RoundInput[113]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12600, new_AGEMA_signal_12599, RoundReg_Inst_ff_SDE_114_next_state}), .Q ({new_AGEMA_signal_4646, new_AGEMA_signal_4645, RoundInput[114]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12836, new_AGEMA_signal_12835, RoundReg_Inst_ff_SDE_115_next_state}), .Q ({new_AGEMA_signal_4652, new_AGEMA_signal_4651, RoundInput[115]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12840, new_AGEMA_signal_12839, RoundReg_Inst_ff_SDE_116_next_state}), .Q ({new_AGEMA_signal_4658, new_AGEMA_signal_4657, RoundInput[116]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12604, new_AGEMA_signal_12603, RoundReg_Inst_ff_SDE_117_next_state}), .Q ({new_AGEMA_signal_4664, new_AGEMA_signal_4663, RoundInput[117]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12608, new_AGEMA_signal_12607, RoundReg_Inst_ff_SDE_118_next_state}), .Q ({new_AGEMA_signal_4670, new_AGEMA_signal_4669, RoundInput[118]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12612, new_AGEMA_signal_12611, RoundReg_Inst_ff_SDE_119_next_state}), .Q ({new_AGEMA_signal_4676, new_AGEMA_signal_4675, RoundInput[119]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12616, new_AGEMA_signal_12615, RoundReg_Inst_ff_SDE_120_next_state}), .Q ({new_AGEMA_signal_4688, new_AGEMA_signal_4687, RoundInput[120]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12844, new_AGEMA_signal_12843, RoundReg_Inst_ff_SDE_121_next_state}), .Q ({new_AGEMA_signal_4694, new_AGEMA_signal_4693, RoundInput[121]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12620, new_AGEMA_signal_12619, RoundReg_Inst_ff_SDE_122_next_state}), .Q ({new_AGEMA_signal_4700, new_AGEMA_signal_4699, RoundInput[122]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12848, new_AGEMA_signal_12847, RoundReg_Inst_ff_SDE_123_next_state}), .Q ({new_AGEMA_signal_4706, new_AGEMA_signal_4705, RoundInput[123]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12852, new_AGEMA_signal_12851, RoundReg_Inst_ff_SDE_124_next_state}), .Q ({new_AGEMA_signal_4712, new_AGEMA_signal_4711, RoundInput[124]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12624, new_AGEMA_signal_12623, RoundReg_Inst_ff_SDE_125_next_state}), .Q ({new_AGEMA_signal_4718, new_AGEMA_signal_4717, RoundInput[125]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12628, new_AGEMA_signal_12627, RoundReg_Inst_ff_SDE_126_next_state}), .Q ({new_AGEMA_signal_4724, new_AGEMA_signal_4723, RoundInput[126]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12632, new_AGEMA_signal_12631, RoundReg_Inst_ff_SDE_127_next_state}), .Q ({new_AGEMA_signal_4730, new_AGEMA_signal_4729, RoundInput[127]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11648, new_AGEMA_signal_11647, KeyReg_Inst_ff_SDE_0_next_state}), .Q ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, RoundKey[0]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12090, new_AGEMA_signal_12089, KeyReg_Inst_ff_SDE_1_next_state}), .Q ({new_AGEMA_signal_4786, new_AGEMA_signal_4785, RoundKey[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12094, new_AGEMA_signal_12093, KeyReg_Inst_ff_SDE_2_next_state}), .Q ({new_AGEMA_signal_4852, new_AGEMA_signal_4851, RoundKey[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12098, new_AGEMA_signal_12097, KeyReg_Inst_ff_SDE_3_next_state}), .Q ({new_AGEMA_signal_4918, new_AGEMA_signal_4917, RoundKey[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12102, new_AGEMA_signal_12101, KeyReg_Inst_ff_SDE_4_next_state}), .Q ({new_AGEMA_signal_4984, new_AGEMA_signal_4983, RoundKey[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12106, new_AGEMA_signal_12105, KeyReg_Inst_ff_SDE_5_next_state}), .Q ({new_AGEMA_signal_5050, new_AGEMA_signal_5049, RoundKey[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12110, new_AGEMA_signal_12109, KeyReg_Inst_ff_SDE_6_next_state}), .Q ({new_AGEMA_signal_5116, new_AGEMA_signal_5115, RoundKey[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12114, new_AGEMA_signal_12113, KeyReg_Inst_ff_SDE_7_next_state}), .Q ({new_AGEMA_signal_5182, new_AGEMA_signal_5181, RoundKey[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11652, new_AGEMA_signal_11651, KeyReg_Inst_ff_SDE_8_next_state}), .Q ({new_AGEMA_signal_5248, new_AGEMA_signal_5247, RoundKey[8]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12118, new_AGEMA_signal_12117, KeyReg_Inst_ff_SDE_9_next_state}), .Q ({new_AGEMA_signal_5314, new_AGEMA_signal_5313, RoundKey[9]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12122, new_AGEMA_signal_12121, KeyReg_Inst_ff_SDE_10_next_state}), .Q ({new_AGEMA_signal_4618, new_AGEMA_signal_4617, RoundKey[10]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12126, new_AGEMA_signal_12125, KeyReg_Inst_ff_SDE_11_next_state}), .Q ({new_AGEMA_signal_4684, new_AGEMA_signal_4683, RoundKey[11]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12130, new_AGEMA_signal_12129, KeyReg_Inst_ff_SDE_12_next_state}), .Q ({new_AGEMA_signal_4738, new_AGEMA_signal_4737, RoundKey[12]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12134, new_AGEMA_signal_12133, KeyReg_Inst_ff_SDE_13_next_state}), .Q ({new_AGEMA_signal_4744, new_AGEMA_signal_4743, RoundKey[13]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12138, new_AGEMA_signal_12137, KeyReg_Inst_ff_SDE_14_next_state}), .Q ({new_AGEMA_signal_4750, new_AGEMA_signal_4749, RoundKey[14]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12142, new_AGEMA_signal_12141, KeyReg_Inst_ff_SDE_15_next_state}), .Q ({new_AGEMA_signal_4756, new_AGEMA_signal_4755, RoundKey[15]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11656, new_AGEMA_signal_11655, KeyReg_Inst_ff_SDE_16_next_state}), .Q ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, RoundKey[16]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12146, new_AGEMA_signal_12145, KeyReg_Inst_ff_SDE_17_next_state}), .Q ({new_AGEMA_signal_4768, new_AGEMA_signal_4767, RoundKey[17]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12150, new_AGEMA_signal_12149, KeyReg_Inst_ff_SDE_18_next_state}), .Q ({new_AGEMA_signal_4774, new_AGEMA_signal_4773, RoundKey[18]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12154, new_AGEMA_signal_12153, KeyReg_Inst_ff_SDE_19_next_state}), .Q ({new_AGEMA_signal_4780, new_AGEMA_signal_4779, RoundKey[19]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12158, new_AGEMA_signal_12157, KeyReg_Inst_ff_SDE_20_next_state}), .Q ({new_AGEMA_signal_4792, new_AGEMA_signal_4791, RoundKey[20]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12162, new_AGEMA_signal_12161, KeyReg_Inst_ff_SDE_21_next_state}), .Q ({new_AGEMA_signal_4798, new_AGEMA_signal_4797, RoundKey[21]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12166, new_AGEMA_signal_12165, KeyReg_Inst_ff_SDE_22_next_state}), .Q ({new_AGEMA_signal_4804, new_AGEMA_signal_4803, RoundKey[22]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12170, new_AGEMA_signal_12169, KeyReg_Inst_ff_SDE_23_next_state}), .Q ({new_AGEMA_signal_4810, new_AGEMA_signal_4809, RoundKey[23]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12174, new_AGEMA_signal_12173, KeyReg_Inst_ff_SDE_24_next_state}), .Q ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, RoundKey[24]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12636, new_AGEMA_signal_12635, KeyReg_Inst_ff_SDE_25_next_state}), .Q ({new_AGEMA_signal_4822, new_AGEMA_signal_4821, RoundKey[25]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12640, new_AGEMA_signal_12639, KeyReg_Inst_ff_SDE_26_next_state}), .Q ({new_AGEMA_signal_4828, new_AGEMA_signal_4827, RoundKey[26]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12644, new_AGEMA_signal_12643, KeyReg_Inst_ff_SDE_27_next_state}), .Q ({new_AGEMA_signal_4834, new_AGEMA_signal_4833, RoundKey[27]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12648, new_AGEMA_signal_12647, KeyReg_Inst_ff_SDE_28_next_state}), .Q ({new_AGEMA_signal_4840, new_AGEMA_signal_4839, RoundKey[28]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12652, new_AGEMA_signal_12651, KeyReg_Inst_ff_SDE_29_next_state}), .Q ({new_AGEMA_signal_4846, new_AGEMA_signal_4845, RoundKey[29]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12656, new_AGEMA_signal_12655, KeyReg_Inst_ff_SDE_30_next_state}), .Q ({new_AGEMA_signal_4858, new_AGEMA_signal_4857, RoundKey[30]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12660, new_AGEMA_signal_12659, KeyReg_Inst_ff_SDE_31_next_state}), .Q ({new_AGEMA_signal_4864, new_AGEMA_signal_4863, RoundKey[31]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11200, new_AGEMA_signal_11199, KeyReg_Inst_ff_SDE_32_next_state}), .Q ({new_AGEMA_signal_4870, new_AGEMA_signal_4869, RoundKey[32]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11660, new_AGEMA_signal_11659, KeyReg_Inst_ff_SDE_33_next_state}), .Q ({new_AGEMA_signal_4876, new_AGEMA_signal_4875, RoundKey[33]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11664, new_AGEMA_signal_11663, KeyReg_Inst_ff_SDE_34_next_state}), .Q ({new_AGEMA_signal_4882, new_AGEMA_signal_4881, RoundKey[34]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11668, new_AGEMA_signal_11667, KeyReg_Inst_ff_SDE_35_next_state}), .Q ({new_AGEMA_signal_4888, new_AGEMA_signal_4887, RoundKey[35]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11672, new_AGEMA_signal_11671, KeyReg_Inst_ff_SDE_36_next_state}), .Q ({new_AGEMA_signal_4894, new_AGEMA_signal_4893, RoundKey[36]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11676, new_AGEMA_signal_11675, KeyReg_Inst_ff_SDE_37_next_state}), .Q ({new_AGEMA_signal_4900, new_AGEMA_signal_4899, RoundKey[37]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11680, new_AGEMA_signal_11679, KeyReg_Inst_ff_SDE_38_next_state}), .Q ({new_AGEMA_signal_4906, new_AGEMA_signal_4905, RoundKey[38]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11684, new_AGEMA_signal_11683, KeyReg_Inst_ff_SDE_39_next_state}), .Q ({new_AGEMA_signal_4912, new_AGEMA_signal_4911, RoundKey[39]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11204, new_AGEMA_signal_11203, KeyReg_Inst_ff_SDE_40_next_state}), .Q ({new_AGEMA_signal_4924, new_AGEMA_signal_4923, RoundKey[40]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11688, new_AGEMA_signal_11687, KeyReg_Inst_ff_SDE_41_next_state}), .Q ({new_AGEMA_signal_4930, new_AGEMA_signal_4929, RoundKey[41]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11692, new_AGEMA_signal_11691, KeyReg_Inst_ff_SDE_42_next_state}), .Q ({new_AGEMA_signal_4936, new_AGEMA_signal_4935, RoundKey[42]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11696, new_AGEMA_signal_11695, KeyReg_Inst_ff_SDE_43_next_state}), .Q ({new_AGEMA_signal_4942, new_AGEMA_signal_4941, RoundKey[43]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11700, new_AGEMA_signal_11699, KeyReg_Inst_ff_SDE_44_next_state}), .Q ({new_AGEMA_signal_4948, new_AGEMA_signal_4947, RoundKey[44]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11704, new_AGEMA_signal_11703, KeyReg_Inst_ff_SDE_45_next_state}), .Q ({new_AGEMA_signal_4954, new_AGEMA_signal_4953, RoundKey[45]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11708, new_AGEMA_signal_11707, KeyReg_Inst_ff_SDE_46_next_state}), .Q ({new_AGEMA_signal_4960, new_AGEMA_signal_4959, RoundKey[46]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11712, new_AGEMA_signal_11711, KeyReg_Inst_ff_SDE_47_next_state}), .Q ({new_AGEMA_signal_4966, new_AGEMA_signal_4965, RoundKey[47]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11208, new_AGEMA_signal_11207, KeyReg_Inst_ff_SDE_48_next_state}), .Q ({new_AGEMA_signal_4972, new_AGEMA_signal_4971, RoundKey[48]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11716, new_AGEMA_signal_11715, KeyReg_Inst_ff_SDE_49_next_state}), .Q ({new_AGEMA_signal_4978, new_AGEMA_signal_4977, RoundKey[49]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11720, new_AGEMA_signal_11719, KeyReg_Inst_ff_SDE_50_next_state}), .Q ({new_AGEMA_signal_4990, new_AGEMA_signal_4989, RoundKey[50]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11724, new_AGEMA_signal_11723, KeyReg_Inst_ff_SDE_51_next_state}), .Q ({new_AGEMA_signal_4996, new_AGEMA_signal_4995, RoundKey[51]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11728, new_AGEMA_signal_11727, KeyReg_Inst_ff_SDE_52_next_state}), .Q ({new_AGEMA_signal_5002, new_AGEMA_signal_5001, RoundKey[52]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11732, new_AGEMA_signal_11731, KeyReg_Inst_ff_SDE_53_next_state}), .Q ({new_AGEMA_signal_5008, new_AGEMA_signal_5007, RoundKey[53]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11736, new_AGEMA_signal_11735, KeyReg_Inst_ff_SDE_54_next_state}), .Q ({new_AGEMA_signal_5014, new_AGEMA_signal_5013, RoundKey[54]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11740, new_AGEMA_signal_11739, KeyReg_Inst_ff_SDE_55_next_state}), .Q ({new_AGEMA_signal_5020, new_AGEMA_signal_5019, RoundKey[55]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11744, new_AGEMA_signal_11743, KeyReg_Inst_ff_SDE_56_next_state}), .Q ({new_AGEMA_signal_5026, new_AGEMA_signal_5025, RoundKey[56]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12178, new_AGEMA_signal_12177, KeyReg_Inst_ff_SDE_57_next_state}), .Q ({new_AGEMA_signal_5032, new_AGEMA_signal_5031, RoundKey[57]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12182, new_AGEMA_signal_12181, KeyReg_Inst_ff_SDE_58_next_state}), .Q ({new_AGEMA_signal_5038, new_AGEMA_signal_5037, RoundKey[58]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12186, new_AGEMA_signal_12185, KeyReg_Inst_ff_SDE_59_next_state}), .Q ({new_AGEMA_signal_5044, new_AGEMA_signal_5043, RoundKey[59]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12190, new_AGEMA_signal_12189, KeyReg_Inst_ff_SDE_60_next_state}), .Q ({new_AGEMA_signal_5056, new_AGEMA_signal_5055, RoundKey[60]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12194, new_AGEMA_signal_12193, KeyReg_Inst_ff_SDE_61_next_state}), .Q ({new_AGEMA_signal_5062, new_AGEMA_signal_5061, RoundKey[61]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12198, new_AGEMA_signal_12197, KeyReg_Inst_ff_SDE_62_next_state}), .Q ({new_AGEMA_signal_5068, new_AGEMA_signal_5067, RoundKey[62]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_12202, new_AGEMA_signal_12201, KeyReg_Inst_ff_SDE_63_next_state}), .Q ({new_AGEMA_signal_5074, new_AGEMA_signal_5073, RoundKey[63]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10780, new_AGEMA_signal_10779, KeyReg_Inst_ff_SDE_64_next_state}), .Q ({new_AGEMA_signal_5080, new_AGEMA_signal_5079, RoundKey[64]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11212, new_AGEMA_signal_11211, KeyReg_Inst_ff_SDE_65_next_state}), .Q ({new_AGEMA_signal_5086, new_AGEMA_signal_5085, RoundKey[65]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11216, new_AGEMA_signal_11215, KeyReg_Inst_ff_SDE_66_next_state}), .Q ({new_AGEMA_signal_5092, new_AGEMA_signal_5091, RoundKey[66]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11220, new_AGEMA_signal_11219, KeyReg_Inst_ff_SDE_67_next_state}), .Q ({new_AGEMA_signal_5098, new_AGEMA_signal_5097, RoundKey[67]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11224, new_AGEMA_signal_11223, KeyReg_Inst_ff_SDE_68_next_state}), .Q ({new_AGEMA_signal_5104, new_AGEMA_signal_5103, RoundKey[68]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11228, new_AGEMA_signal_11227, KeyReg_Inst_ff_SDE_69_next_state}), .Q ({new_AGEMA_signal_5110, new_AGEMA_signal_5109, RoundKey[69]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11232, new_AGEMA_signal_11231, KeyReg_Inst_ff_SDE_70_next_state}), .Q ({new_AGEMA_signal_5122, new_AGEMA_signal_5121, RoundKey[70]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11236, new_AGEMA_signal_11235, KeyReg_Inst_ff_SDE_71_next_state}), .Q ({new_AGEMA_signal_5128, new_AGEMA_signal_5127, RoundKey[71]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10784, new_AGEMA_signal_10783, KeyReg_Inst_ff_SDE_72_next_state}), .Q ({new_AGEMA_signal_5134, new_AGEMA_signal_5133, RoundKey[72]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11240, new_AGEMA_signal_11239, KeyReg_Inst_ff_SDE_73_next_state}), .Q ({new_AGEMA_signal_5140, new_AGEMA_signal_5139, RoundKey[73]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11244, new_AGEMA_signal_11243, KeyReg_Inst_ff_SDE_74_next_state}), .Q ({new_AGEMA_signal_5146, new_AGEMA_signal_5145, RoundKey[74]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11248, new_AGEMA_signal_11247, KeyReg_Inst_ff_SDE_75_next_state}), .Q ({new_AGEMA_signal_5152, new_AGEMA_signal_5151, RoundKey[75]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11252, new_AGEMA_signal_11251, KeyReg_Inst_ff_SDE_76_next_state}), .Q ({new_AGEMA_signal_5158, new_AGEMA_signal_5157, RoundKey[76]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11256, new_AGEMA_signal_11255, KeyReg_Inst_ff_SDE_77_next_state}), .Q ({new_AGEMA_signal_5164, new_AGEMA_signal_5163, RoundKey[77]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11260, new_AGEMA_signal_11259, KeyReg_Inst_ff_SDE_78_next_state}), .Q ({new_AGEMA_signal_5170, new_AGEMA_signal_5169, RoundKey[78]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11264, new_AGEMA_signal_11263, KeyReg_Inst_ff_SDE_79_next_state}), .Q ({new_AGEMA_signal_5176, new_AGEMA_signal_5175, RoundKey[79]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10788, new_AGEMA_signal_10787, KeyReg_Inst_ff_SDE_80_next_state}), .Q ({new_AGEMA_signal_5188, new_AGEMA_signal_5187, RoundKey[80]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11268, new_AGEMA_signal_11267, KeyReg_Inst_ff_SDE_81_next_state}), .Q ({new_AGEMA_signal_5194, new_AGEMA_signal_5193, RoundKey[81]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11272, new_AGEMA_signal_11271, KeyReg_Inst_ff_SDE_82_next_state}), .Q ({new_AGEMA_signal_5200, new_AGEMA_signal_5199, RoundKey[82]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11276, new_AGEMA_signal_11275, KeyReg_Inst_ff_SDE_83_next_state}), .Q ({new_AGEMA_signal_5206, new_AGEMA_signal_5205, RoundKey[83]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11280, new_AGEMA_signal_11279, KeyReg_Inst_ff_SDE_84_next_state}), .Q ({new_AGEMA_signal_5212, new_AGEMA_signal_5211, RoundKey[84]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11284, new_AGEMA_signal_11283, KeyReg_Inst_ff_SDE_85_next_state}), .Q ({new_AGEMA_signal_5218, new_AGEMA_signal_5217, RoundKey[85]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11288, new_AGEMA_signal_11287, KeyReg_Inst_ff_SDE_86_next_state}), .Q ({new_AGEMA_signal_5224, new_AGEMA_signal_5223, RoundKey[86]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11292, new_AGEMA_signal_11291, KeyReg_Inst_ff_SDE_87_next_state}), .Q ({new_AGEMA_signal_5230, new_AGEMA_signal_5229, RoundKey[87]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11296, new_AGEMA_signal_11295, KeyReg_Inst_ff_SDE_88_next_state}), .Q ({new_AGEMA_signal_5236, new_AGEMA_signal_5235, RoundKey[88]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11748, new_AGEMA_signal_11747, KeyReg_Inst_ff_SDE_89_next_state}), .Q ({new_AGEMA_signal_5242, new_AGEMA_signal_5241, RoundKey[89]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11752, new_AGEMA_signal_11751, KeyReg_Inst_ff_SDE_90_next_state}), .Q ({new_AGEMA_signal_5254, new_AGEMA_signal_5253, RoundKey[90]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11756, new_AGEMA_signal_11755, KeyReg_Inst_ff_SDE_91_next_state}), .Q ({new_AGEMA_signal_5260, new_AGEMA_signal_5259, RoundKey[91]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11760, new_AGEMA_signal_11759, KeyReg_Inst_ff_SDE_92_next_state}), .Q ({new_AGEMA_signal_5266, new_AGEMA_signal_5265, RoundKey[92]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11764, new_AGEMA_signal_11763, KeyReg_Inst_ff_SDE_93_next_state}), .Q ({new_AGEMA_signal_5272, new_AGEMA_signal_5271, RoundKey[93]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11768, new_AGEMA_signal_11767, KeyReg_Inst_ff_SDE_94_next_state}), .Q ({new_AGEMA_signal_5278, new_AGEMA_signal_5277, RoundKey[94]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11772, new_AGEMA_signal_11771, KeyReg_Inst_ff_SDE_95_next_state}), .Q ({new_AGEMA_signal_5284, new_AGEMA_signal_5283, RoundKey[95]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10448, new_AGEMA_signal_10447, KeyReg_Inst_ff_SDE_96_next_state}), .Q ({new_AGEMA_signal_5290, new_AGEMA_signal_5289, RoundKey[96]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10792, new_AGEMA_signal_10791, KeyReg_Inst_ff_SDE_97_next_state}), .Q ({new_AGEMA_signal_5296, new_AGEMA_signal_5295, RoundKey[97]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10796, new_AGEMA_signal_10795, KeyReg_Inst_ff_SDE_98_next_state}), .Q ({new_AGEMA_signal_5302, new_AGEMA_signal_5301, RoundKey[98]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10800, new_AGEMA_signal_10799, KeyReg_Inst_ff_SDE_99_next_state}), .Q ({new_AGEMA_signal_5308, new_AGEMA_signal_5307, RoundKey[99]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10804, new_AGEMA_signal_10803, KeyReg_Inst_ff_SDE_100_next_state}), .Q ({new_AGEMA_signal_4558, new_AGEMA_signal_4557, RoundKey[100]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10808, new_AGEMA_signal_10807, KeyReg_Inst_ff_SDE_101_next_state}), .Q ({new_AGEMA_signal_4564, new_AGEMA_signal_4563, RoundKey[101]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10812, new_AGEMA_signal_10811, KeyReg_Inst_ff_SDE_102_next_state}), .Q ({new_AGEMA_signal_4570, new_AGEMA_signal_4569, RoundKey[102]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10816, new_AGEMA_signal_10815, KeyReg_Inst_ff_SDE_103_next_state}), .Q ({new_AGEMA_signal_4576, new_AGEMA_signal_4575, RoundKey[103]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10452, new_AGEMA_signal_10451, KeyReg_Inst_ff_SDE_104_next_state}), .Q ({new_AGEMA_signal_4582, new_AGEMA_signal_4581, RoundKey[104]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10820, new_AGEMA_signal_10819, KeyReg_Inst_ff_SDE_105_next_state}), .Q ({new_AGEMA_signal_4588, new_AGEMA_signal_4587, RoundKey[105]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10824, new_AGEMA_signal_10823, KeyReg_Inst_ff_SDE_106_next_state}), .Q ({new_AGEMA_signal_4594, new_AGEMA_signal_4593, RoundKey[106]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10828, new_AGEMA_signal_10827, KeyReg_Inst_ff_SDE_107_next_state}), .Q ({new_AGEMA_signal_4600, new_AGEMA_signal_4599, RoundKey[107]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10832, new_AGEMA_signal_10831, KeyReg_Inst_ff_SDE_108_next_state}), .Q ({new_AGEMA_signal_4606, new_AGEMA_signal_4605, RoundKey[108]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10836, new_AGEMA_signal_10835, KeyReg_Inst_ff_SDE_109_next_state}), .Q ({new_AGEMA_signal_4612, new_AGEMA_signal_4611, RoundKey[109]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10840, new_AGEMA_signal_10839, KeyReg_Inst_ff_SDE_110_next_state}), .Q ({new_AGEMA_signal_4624, new_AGEMA_signal_4623, RoundKey[110]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10844, new_AGEMA_signal_10843, KeyReg_Inst_ff_SDE_111_next_state}), .Q ({new_AGEMA_signal_4630, new_AGEMA_signal_4629, RoundKey[111]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, KeyReg_Inst_ff_SDE_112_next_state}), .Q ({new_AGEMA_signal_4636, new_AGEMA_signal_4635, RoundKey[112]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10848, new_AGEMA_signal_10847, KeyReg_Inst_ff_SDE_113_next_state}), .Q ({new_AGEMA_signal_4642, new_AGEMA_signal_4641, RoundKey[113]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10852, new_AGEMA_signal_10851, KeyReg_Inst_ff_SDE_114_next_state}), .Q ({new_AGEMA_signal_4648, new_AGEMA_signal_4647, RoundKey[114]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10856, new_AGEMA_signal_10855, KeyReg_Inst_ff_SDE_115_next_state}), .Q ({new_AGEMA_signal_4654, new_AGEMA_signal_4653, RoundKey[115]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10860, new_AGEMA_signal_10859, KeyReg_Inst_ff_SDE_116_next_state}), .Q ({new_AGEMA_signal_4660, new_AGEMA_signal_4659, RoundKey[116]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10864, new_AGEMA_signal_10863, KeyReg_Inst_ff_SDE_117_next_state}), .Q ({new_AGEMA_signal_4666, new_AGEMA_signal_4665, RoundKey[117]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10868, new_AGEMA_signal_10867, KeyReg_Inst_ff_SDE_118_next_state}), .Q ({new_AGEMA_signal_4672, new_AGEMA_signal_4671, RoundKey[118]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10872, new_AGEMA_signal_10871, KeyReg_Inst_ff_SDE_119_next_state}), .Q ({new_AGEMA_signal_4678, new_AGEMA_signal_4677, RoundKey[119]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_10876, new_AGEMA_signal_10875, KeyReg_Inst_ff_SDE_120_next_state}), .Q ({new_AGEMA_signal_4690, new_AGEMA_signal_4689, RoundKey[120]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11300, new_AGEMA_signal_11299, KeyReg_Inst_ff_SDE_121_next_state}), .Q ({new_AGEMA_signal_4696, new_AGEMA_signal_4695, RoundKey[121]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11304, new_AGEMA_signal_11303, KeyReg_Inst_ff_SDE_122_next_state}), .Q ({new_AGEMA_signal_4702, new_AGEMA_signal_4701, RoundKey[122]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11308, new_AGEMA_signal_11307, KeyReg_Inst_ff_SDE_123_next_state}), .Q ({new_AGEMA_signal_4708, new_AGEMA_signal_4707, RoundKey[123]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11312, new_AGEMA_signal_11311, KeyReg_Inst_ff_SDE_124_next_state}), .Q ({new_AGEMA_signal_4714, new_AGEMA_signal_4713, RoundKey[124]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11316, new_AGEMA_signal_11315, KeyReg_Inst_ff_SDE_125_next_state}), .Q ({new_AGEMA_signal_4720, new_AGEMA_signal_4719, RoundKey[125]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11320, new_AGEMA_signal_11319, KeyReg_Inst_ff_SDE_126_next_state}), .Q ({new_AGEMA_signal_4726, new_AGEMA_signal_4725, RoundKey[126]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_11324, new_AGEMA_signal_11323, KeyReg_Inst_ff_SDE_127_next_state}), .Q ({new_AGEMA_signal_4732, new_AGEMA_signal_4731, RoundKey[127]}) ) ;
    DFF_X1 RoundCounterIns_count_reg_0__FF_FF ( .CK (clk_gated), .D (RoundCounterIns_N7), .Q (RoundCounter[0]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_1__FF_FF ( .CK (clk_gated), .D (RoundCounterIns_N8), .Q (RoundCounter[1]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_2__FF_FF ( .CK (clk_gated), .D (RoundCounterIns_n1), .Q (RoundCounter[2]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_3__FF_FF ( .CK (clk_gated), .D (RoundCounterIns_N10), .Q (RoundCounter[3]), .QN () ) ;
endmodule
