////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module AES in file /AGEMA/Designs/AES_serial/AGEMA/sbox_opt3/AES.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module AES_HPC2_ClockGating_d3 (plaintext_s0, key_s0, clk, start, plaintext_s1, plaintext_s2, plaintext_s3, key_s1, key_s2, key_s3, Fresh, ciphertext_s0, done, ciphertext_s1, ciphertext_s2, ciphertext_s3, Synch);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input start ;
    input [127:0] plaintext_s1 ;
    input [127:0] plaintext_s2 ;
    input [127:0] plaintext_s3 ;
    input [127:0] key_s1 ;
    input [127:0] key_s2 ;
    input [127:0] key_s3 ;
    input [203:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    output [127:0] ciphertext_s2 ;
    output [127:0] ciphertext_s3 ;
    output Synch ;
    wire nReset ;
    wire selMC ;
    wire selSR ;
    wire selXOR ;
    wire enRCon ;
    wire finalStep ;
    wire intFinal ;
    wire intselXOR ;
    wire notFirst ;
    wire n10 ;
    wire n9 ;
    wire n12 ;
    wire n13 ;
    wire ctrl_n16 ;
    wire ctrl_n15 ;
    wire ctrl_n14 ;
    wire ctrl_n11 ;
    wire ctrl_n10 ;
    wire ctrl_n9 ;
    wire ctrl_n8 ;
    wire ctrl_n7 ;
    wire ctrl_n5 ;
    wire ctrl_n4 ;
    wire ctrl_n2 ;
    wire ctrl_n12 ;
    wire ctrl_n6 ;
    wire ctrl_N14 ;
    wire ctrl_seq4Out_1_ ;
    wire ctrl_seq4In_1_ ;
    wire ctrl_nRstSeq4 ;
    wire ctrl_n13 ;
    wire ctrl_seq6Out_4_ ;
    wire ctrl_seq6In_1_ ;
    wire ctrl_seq6In_2_ ;
    wire ctrl_seq6In_3_ ;
    wire ctrl_seq6In_4_ ;
    wire ctrl_seq6_SFF_0_QD ;
    wire ctrl_seq6_SFF_1_QD ;
    wire ctrl_seq6_SFF_2_QD ;
    wire ctrl_seq6_SFF_3_QD ;
    wire ctrl_seq6_SFF_4_QD ;
    wire ctrl_seq4_SFF_0_QD ;
    wire ctrl_seq4_SFF_1_QD ;
    wire stateArray_n33 ;
    wire stateArray_n32 ;
    wire stateArray_n31 ;
    wire stateArray_n30 ;
    wire stateArray_n29 ;
    wire stateArray_n28 ;
    wire stateArray_n27 ;
    wire stateArray_n26 ;
    wire stateArray_n25 ;
    wire stateArray_n24 ;
    wire stateArray_n23 ;
    wire stateArray_n22 ;
    wire stateArray_n21 ;
    wire stateArray_n20 ;
    wire stateArray_n19 ;
    wire stateArray_n18 ;
    wire stateArray_n17 ;
    wire stateArray_n16 ;
    wire stateArray_n15 ;
    wire stateArray_n14 ;
    wire stateArray_n13 ;
    wire stateArray_S00reg_gff_1_SFF_0_QD ;
    wire stateArray_S00reg_gff_1_SFF_1_QD ;
    wire stateArray_S00reg_gff_1_SFF_2_QD ;
    wire stateArray_S00reg_gff_1_SFF_3_QD ;
    wire stateArray_S00reg_gff_1_SFF_4_QD ;
    wire stateArray_S00reg_gff_1_SFF_5_QD ;
    wire stateArray_S00reg_gff_1_SFF_6_QD ;
    wire stateArray_S00reg_gff_1_SFF_7_QD ;
    wire stateArray_S01reg_gff_1_SFF_0_QD ;
    wire stateArray_S01reg_gff_1_SFF_1_QD ;
    wire stateArray_S01reg_gff_1_SFF_2_QD ;
    wire stateArray_S01reg_gff_1_SFF_3_QD ;
    wire stateArray_S01reg_gff_1_SFF_4_QD ;
    wire stateArray_S01reg_gff_1_SFF_5_QD ;
    wire stateArray_S01reg_gff_1_SFF_6_QD ;
    wire stateArray_S01reg_gff_1_SFF_7_QD ;
    wire stateArray_S02reg_gff_1_SFF_0_QD ;
    wire stateArray_S02reg_gff_1_SFF_1_QD ;
    wire stateArray_S02reg_gff_1_SFF_2_QD ;
    wire stateArray_S02reg_gff_1_SFF_3_QD ;
    wire stateArray_S02reg_gff_1_SFF_4_QD ;
    wire stateArray_S02reg_gff_1_SFF_5_QD ;
    wire stateArray_S02reg_gff_1_SFF_6_QD ;
    wire stateArray_S02reg_gff_1_SFF_7_QD ;
    wire stateArray_S03reg_gff_1_SFF_0_QD ;
    wire stateArray_S03reg_gff_1_SFF_1_QD ;
    wire stateArray_S03reg_gff_1_SFF_2_QD ;
    wire stateArray_S03reg_gff_1_SFF_3_QD ;
    wire stateArray_S03reg_gff_1_SFF_4_QD ;
    wire stateArray_S03reg_gff_1_SFF_5_QD ;
    wire stateArray_S03reg_gff_1_SFF_6_QD ;
    wire stateArray_S03reg_gff_1_SFF_7_QD ;
    wire stateArray_S10reg_gff_1_SFF_0_QD ;
    wire stateArray_S10reg_gff_1_SFF_1_QD ;
    wire stateArray_S10reg_gff_1_SFF_2_QD ;
    wire stateArray_S10reg_gff_1_SFF_3_QD ;
    wire stateArray_S10reg_gff_1_SFF_4_QD ;
    wire stateArray_S10reg_gff_1_SFF_5_QD ;
    wire stateArray_S10reg_gff_1_SFF_6_QD ;
    wire stateArray_S10reg_gff_1_SFF_7_QD ;
    wire stateArray_S11reg_gff_1_SFF_0_QD ;
    wire stateArray_S11reg_gff_1_SFF_1_QD ;
    wire stateArray_S11reg_gff_1_SFF_2_QD ;
    wire stateArray_S11reg_gff_1_SFF_3_QD ;
    wire stateArray_S11reg_gff_1_SFF_4_QD ;
    wire stateArray_S11reg_gff_1_SFF_5_QD ;
    wire stateArray_S11reg_gff_1_SFF_6_QD ;
    wire stateArray_S11reg_gff_1_SFF_7_QD ;
    wire stateArray_S12reg_gff_1_SFF_0_QD ;
    wire stateArray_S12reg_gff_1_SFF_1_QD ;
    wire stateArray_S12reg_gff_1_SFF_2_QD ;
    wire stateArray_S12reg_gff_1_SFF_3_QD ;
    wire stateArray_S12reg_gff_1_SFF_4_QD ;
    wire stateArray_S12reg_gff_1_SFF_5_QD ;
    wire stateArray_S12reg_gff_1_SFF_6_QD ;
    wire stateArray_S12reg_gff_1_SFF_7_QD ;
    wire stateArray_S13reg_gff_1_SFF_0_QD ;
    wire stateArray_S13reg_gff_1_SFF_1_QD ;
    wire stateArray_S13reg_gff_1_SFF_2_QD ;
    wire stateArray_S13reg_gff_1_SFF_3_QD ;
    wire stateArray_S13reg_gff_1_SFF_4_QD ;
    wire stateArray_S13reg_gff_1_SFF_5_QD ;
    wire stateArray_S13reg_gff_1_SFF_6_QD ;
    wire stateArray_S13reg_gff_1_SFF_7_QD ;
    wire stateArray_S20reg_gff_1_SFF_0_QD ;
    wire stateArray_S20reg_gff_1_SFF_1_QD ;
    wire stateArray_S20reg_gff_1_SFF_2_QD ;
    wire stateArray_S20reg_gff_1_SFF_3_QD ;
    wire stateArray_S20reg_gff_1_SFF_4_QD ;
    wire stateArray_S20reg_gff_1_SFF_5_QD ;
    wire stateArray_S20reg_gff_1_SFF_6_QD ;
    wire stateArray_S20reg_gff_1_SFF_7_QD ;
    wire stateArray_S21reg_gff_1_SFF_0_QD ;
    wire stateArray_S21reg_gff_1_SFF_1_QD ;
    wire stateArray_S21reg_gff_1_SFF_2_QD ;
    wire stateArray_S21reg_gff_1_SFF_3_QD ;
    wire stateArray_S21reg_gff_1_SFF_4_QD ;
    wire stateArray_S21reg_gff_1_SFF_5_QD ;
    wire stateArray_S21reg_gff_1_SFF_6_QD ;
    wire stateArray_S21reg_gff_1_SFF_7_QD ;
    wire stateArray_S22reg_gff_1_SFF_0_QD ;
    wire stateArray_S22reg_gff_1_SFF_1_QD ;
    wire stateArray_S22reg_gff_1_SFF_2_QD ;
    wire stateArray_S22reg_gff_1_SFF_3_QD ;
    wire stateArray_S22reg_gff_1_SFF_4_QD ;
    wire stateArray_S22reg_gff_1_SFF_5_QD ;
    wire stateArray_S22reg_gff_1_SFF_6_QD ;
    wire stateArray_S22reg_gff_1_SFF_7_QD ;
    wire stateArray_S23reg_gff_1_SFF_0_QD ;
    wire stateArray_S23reg_gff_1_SFF_1_QD ;
    wire stateArray_S23reg_gff_1_SFF_2_QD ;
    wire stateArray_S23reg_gff_1_SFF_3_QD ;
    wire stateArray_S23reg_gff_1_SFF_4_QD ;
    wire stateArray_S23reg_gff_1_SFF_5_QD ;
    wire stateArray_S23reg_gff_1_SFF_6_QD ;
    wire stateArray_S23reg_gff_1_SFF_7_QD ;
    wire stateArray_S30reg_gff_1_SFF_0_QD ;
    wire stateArray_S30reg_gff_1_SFF_1_QD ;
    wire stateArray_S30reg_gff_1_SFF_2_QD ;
    wire stateArray_S30reg_gff_1_SFF_3_QD ;
    wire stateArray_S30reg_gff_1_SFF_4_QD ;
    wire stateArray_S30reg_gff_1_SFF_5_QD ;
    wire stateArray_S30reg_gff_1_SFF_6_QD ;
    wire stateArray_S30reg_gff_1_SFF_7_QD ;
    wire stateArray_S31reg_gff_1_SFF_0_QD ;
    wire stateArray_S31reg_gff_1_SFF_1_QD ;
    wire stateArray_S31reg_gff_1_SFF_2_QD ;
    wire stateArray_S31reg_gff_1_SFF_3_QD ;
    wire stateArray_S31reg_gff_1_SFF_4_QD ;
    wire stateArray_S31reg_gff_1_SFF_5_QD ;
    wire stateArray_S31reg_gff_1_SFF_6_QD ;
    wire stateArray_S31reg_gff_1_SFF_7_QD ;
    wire stateArray_S32reg_gff_1_SFF_0_QD ;
    wire stateArray_S32reg_gff_1_SFF_1_QD ;
    wire stateArray_S32reg_gff_1_SFF_2_QD ;
    wire stateArray_S32reg_gff_1_SFF_3_QD ;
    wire stateArray_S32reg_gff_1_SFF_4_QD ;
    wire stateArray_S32reg_gff_1_SFF_5_QD ;
    wire stateArray_S32reg_gff_1_SFF_6_QD ;
    wire stateArray_S32reg_gff_1_SFF_7_QD ;
    wire stateArray_S33reg_gff_1_SFF_0_QD ;
    wire stateArray_S33reg_gff_1_SFF_1_QD ;
    wire stateArray_S33reg_gff_1_SFF_2_QD ;
    wire stateArray_S33reg_gff_1_SFF_3_QD ;
    wire stateArray_S33reg_gff_1_SFF_4_QD ;
    wire stateArray_S33reg_gff_1_SFF_5_QD ;
    wire stateArray_S33reg_gff_1_SFF_6_QD ;
    wire stateArray_S33reg_gff_1_SFF_7_QD ;
    wire MUX_StateInMC_n7 ;
    wire MUX_StateInMC_n6 ;
    wire MUX_StateInMC_n5 ;
    wire KeyArray_n55 ;
    wire KeyArray_n54 ;
    wire KeyArray_n53 ;
    wire KeyArray_n52 ;
    wire KeyArray_n51 ;
    wire KeyArray_n50 ;
    wire KeyArray_n49 ;
    wire KeyArray_n48 ;
    wire KeyArray_n47 ;
    wire KeyArray_n46 ;
    wire KeyArray_n45 ;
    wire KeyArray_n44 ;
    wire KeyArray_n43 ;
    wire KeyArray_n42 ;
    wire KeyArray_n41 ;
    wire KeyArray_n40 ;
    wire KeyArray_n39 ;
    wire KeyArray_n38 ;
    wire KeyArray_n37 ;
    wire KeyArray_n36 ;
    wire KeyArray_n35 ;
    wire KeyArray_n34 ;
    wire KeyArray_n33 ;
    wire KeyArray_n32 ;
    wire KeyArray_n31 ;
    wire KeyArray_n30 ;
    wire KeyArray_n29 ;
    wire KeyArray_n28 ;
    wire KeyArray_n27 ;
    wire KeyArray_n26 ;
    wire KeyArray_n25 ;
    wire KeyArray_n24 ;
    wire KeyArray_n23 ;
    wire KeyArray_n22 ;
    wire KeyArray_outS01ser_0_ ;
    wire KeyArray_outS01ser_1_ ;
    wire KeyArray_outS01ser_2_ ;
    wire KeyArray_outS01ser_3_ ;
    wire KeyArray_outS01ser_4_ ;
    wire KeyArray_outS01ser_5_ ;
    wire KeyArray_outS01ser_6_ ;
    wire KeyArray_outS01ser_7_ ;
    wire KeyArray_S00reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S00reg_gff_1_SFF_0_QD ;
    wire KeyArray_S00reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_1_QD ;
    wire KeyArray_S00reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_2_QD ;
    wire KeyArray_S00reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_3_QD ;
    wire KeyArray_S00reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_4_QD ;
    wire KeyArray_S00reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_5_QD ;
    wire KeyArray_S00reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_6_QD ;
    wire KeyArray_S00reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_7_QD ;
    wire KeyArray_S01reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_0_QD ;
    wire KeyArray_S01reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_1_QD ;
    wire KeyArray_S01reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_2_QD ;
    wire KeyArray_S01reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_3_QD ;
    wire KeyArray_S01reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_4_QD ;
    wire KeyArray_S01reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_5_QD ;
    wire KeyArray_S01reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_6_QD ;
    wire KeyArray_S01reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_7_QD ;
    wire KeyArray_S02reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_0_QD ;
    wire KeyArray_S02reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_1_QD ;
    wire KeyArray_S02reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_2_QD ;
    wire KeyArray_S02reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_3_QD ;
    wire KeyArray_S02reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_4_QD ;
    wire KeyArray_S02reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_5_QD ;
    wire KeyArray_S02reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_6_QD ;
    wire KeyArray_S02reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_7_QD ;
    wire KeyArray_S03reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_0_QD ;
    wire KeyArray_S03reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_1_QD ;
    wire KeyArray_S03reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_2_QD ;
    wire KeyArray_S03reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_3_QD ;
    wire KeyArray_S03reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_4_QD ;
    wire KeyArray_S03reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S03reg_gff_1_SFF_5_QD ;
    wire KeyArray_S03reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S03reg_gff_1_SFF_6_QD ;
    wire KeyArray_S03reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S03reg_gff_1_SFF_7_QD ;
    wire KeyArray_S10reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_0_QD ;
    wire KeyArray_S10reg_gff_1_SFF_1_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_1_QD ;
    wire KeyArray_S10reg_gff_1_SFF_2_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_2_QD ;
    wire KeyArray_S10reg_gff_1_SFF_3_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_3_QD ;
    wire KeyArray_S10reg_gff_1_SFF_4_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_4_QD ;
    wire KeyArray_S10reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_5_QD ;
    wire KeyArray_S10reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_6_QD ;
    wire KeyArray_S10reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_7_QD ;
    wire KeyArray_S11reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_0_QD ;
    wire KeyArray_S11reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_1_QD ;
    wire KeyArray_S11reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_2_QD ;
    wire KeyArray_S11reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_3_QD ;
    wire KeyArray_S11reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_4_QD ;
    wire KeyArray_S11reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_5_QD ;
    wire KeyArray_S11reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_6_QD ;
    wire KeyArray_S11reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_7_QD ;
    wire KeyArray_S12reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_0_QD ;
    wire KeyArray_S12reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_1_QD ;
    wire KeyArray_S12reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_2_QD ;
    wire KeyArray_S12reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_3_QD ;
    wire KeyArray_S12reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_4_QD ;
    wire KeyArray_S12reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_5_QD ;
    wire KeyArray_S12reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_6_QD ;
    wire KeyArray_S12reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_7_QD ;
    wire KeyArray_S13reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_0_QD ;
    wire KeyArray_S13reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_1_QD ;
    wire KeyArray_S13reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_2_QD ;
    wire KeyArray_S13reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_3_QD ;
    wire KeyArray_S13reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_4_QD ;
    wire KeyArray_S13reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S13reg_gff_1_SFF_5_QD ;
    wire KeyArray_S13reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S13reg_gff_1_SFF_6_QD ;
    wire KeyArray_S13reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S13reg_gff_1_SFF_7_QD ;
    wire KeyArray_S20reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_0_QD ;
    wire KeyArray_S20reg_gff_1_SFF_1_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_1_QD ;
    wire KeyArray_S20reg_gff_1_SFF_2_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_2_QD ;
    wire KeyArray_S20reg_gff_1_SFF_3_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_3_QD ;
    wire KeyArray_S20reg_gff_1_SFF_4_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_4_QD ;
    wire KeyArray_S20reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_5_QD ;
    wire KeyArray_S20reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_6_QD ;
    wire KeyArray_S20reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_7_QD ;
    wire KeyArray_S21reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_0_QD ;
    wire KeyArray_S21reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_1_QD ;
    wire KeyArray_S21reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_2_QD ;
    wire KeyArray_S21reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_3_QD ;
    wire KeyArray_S21reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_4_QD ;
    wire KeyArray_S21reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_5_QD ;
    wire KeyArray_S21reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_6_QD ;
    wire KeyArray_S21reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_7_QD ;
    wire KeyArray_S22reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_0_QD ;
    wire KeyArray_S22reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_1_QD ;
    wire KeyArray_S22reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_2_QD ;
    wire KeyArray_S22reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_3_QD ;
    wire KeyArray_S22reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_4_QD ;
    wire KeyArray_S22reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_5_QD ;
    wire KeyArray_S22reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_6_QD ;
    wire KeyArray_S22reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_7_QD ;
    wire KeyArray_S23reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_0_QD ;
    wire KeyArray_S23reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_1_QD ;
    wire KeyArray_S23reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_2_QD ;
    wire KeyArray_S23reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_3_QD ;
    wire KeyArray_S23reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_4_QD ;
    wire KeyArray_S23reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S23reg_gff_1_SFF_5_QD ;
    wire KeyArray_S23reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S23reg_gff_1_SFF_6_QD ;
    wire KeyArray_S23reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S23reg_gff_1_SFF_7_QD ;
    wire KeyArray_S30reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_0_QD ;
    wire KeyArray_S30reg_gff_1_SFF_1_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_1_QD ;
    wire KeyArray_S30reg_gff_1_SFF_2_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_2_QD ;
    wire KeyArray_S30reg_gff_1_SFF_3_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_3_QD ;
    wire KeyArray_S30reg_gff_1_SFF_4_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_4_QD ;
    wire KeyArray_S30reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_5_QD ;
    wire KeyArray_S30reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_6_QD ;
    wire KeyArray_S30reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_7_QD ;
    wire KeyArray_S31reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_0_QD ;
    wire KeyArray_S31reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_1_QD ;
    wire KeyArray_S31reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_2_QD ;
    wire KeyArray_S31reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_3_QD ;
    wire KeyArray_S31reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_4_QD ;
    wire KeyArray_S31reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_5_QD ;
    wire KeyArray_S31reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_6_QD ;
    wire KeyArray_S31reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_7_QD ;
    wire KeyArray_S32reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_0_QD ;
    wire KeyArray_S32reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_1_QD ;
    wire KeyArray_S32reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_2_QD ;
    wire KeyArray_S32reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_3_QD ;
    wire KeyArray_S32reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_4_QD ;
    wire KeyArray_S32reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_5_QD ;
    wire KeyArray_S32reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S32reg_gff_1_SFF_6_QD ;
    wire KeyArray_S32reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S32reg_gff_1_SFF_7_QD ;
    wire KeyArray_S33reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_0_QD ;
    wire KeyArray_S33reg_gff_1_SFF_1_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_1_QD ;
    wire KeyArray_S33reg_gff_1_SFF_2_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_2_QD ;
    wire KeyArray_S33reg_gff_1_SFF_3_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_3_QD ;
    wire KeyArray_S33reg_gff_1_SFF_4_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_4_QD ;
    wire KeyArray_S33reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_5_QD ;
    wire KeyArray_S33reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_6_QD ;
    wire KeyArray_S33reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_7_QD ;
    wire MixColumns_line0_n16 ;
    wire MixColumns_line0_n15 ;
    wire MixColumns_line0_n14 ;
    wire MixColumns_line0_n13 ;
    wire MixColumns_line0_n12 ;
    wire MixColumns_line0_n11 ;
    wire MixColumns_line0_n10 ;
    wire MixColumns_line0_n9 ;
    wire MixColumns_line0_n8 ;
    wire MixColumns_line0_n7 ;
    wire MixColumns_line0_n6 ;
    wire MixColumns_line0_n5 ;
    wire MixColumns_line0_n4 ;
    wire MixColumns_line0_n3 ;
    wire MixColumns_line0_n2 ;
    wire MixColumns_line0_n1 ;
    wire MixColumns_line1_n16 ;
    wire MixColumns_line1_n15 ;
    wire MixColumns_line1_n14 ;
    wire MixColumns_line1_n13 ;
    wire MixColumns_line1_n12 ;
    wire MixColumns_line1_n11 ;
    wire MixColumns_line1_n10 ;
    wire MixColumns_line1_n9 ;
    wire MixColumns_line1_n8 ;
    wire MixColumns_line1_n7 ;
    wire MixColumns_line1_n6 ;
    wire MixColumns_line1_n5 ;
    wire MixColumns_line1_n4 ;
    wire MixColumns_line1_n3 ;
    wire MixColumns_line1_n2 ;
    wire MixColumns_line1_n1 ;
    wire MixColumns_line1_S02_1_ ;
    wire MixColumns_line1_S02_3_ ;
    wire MixColumns_line1_S02_4_ ;
    wire MixColumns_line2_n16 ;
    wire MixColumns_line2_n15 ;
    wire MixColumns_line2_n14 ;
    wire MixColumns_line2_n13 ;
    wire MixColumns_line2_n12 ;
    wire MixColumns_line2_n11 ;
    wire MixColumns_line2_n10 ;
    wire MixColumns_line2_n9 ;
    wire MixColumns_line2_n8 ;
    wire MixColumns_line2_n7 ;
    wire MixColumns_line2_n6 ;
    wire MixColumns_line2_n5 ;
    wire MixColumns_line2_n4 ;
    wire MixColumns_line2_n3 ;
    wire MixColumns_line2_n2 ;
    wire MixColumns_line2_n1 ;
    wire MixColumns_line2_S02_1_ ;
    wire MixColumns_line2_S02_3_ ;
    wire MixColumns_line2_S02_4_ ;
    wire MixColumns_line3_n16 ;
    wire MixColumns_line3_n15 ;
    wire MixColumns_line3_n14 ;
    wire MixColumns_line3_n13 ;
    wire MixColumns_line3_n12 ;
    wire MixColumns_line3_n11 ;
    wire MixColumns_line3_n10 ;
    wire MixColumns_line3_n9 ;
    wire MixColumns_line3_n8 ;
    wire MixColumns_line3_n7 ;
    wire MixColumns_line3_n6 ;
    wire MixColumns_line3_n5 ;
    wire MixColumns_line3_n4 ;
    wire MixColumns_line3_n3 ;
    wire MixColumns_line3_n2 ;
    wire MixColumns_line3_n1 ;
    wire MixColumns_line3_S02_1_ ;
    wire MixColumns_line3_S02_3_ ;
    wire MixColumns_line3_S02_4_ ;
    wire MixColumns_line3_timesTHREE_input2_1_ ;
    wire MixColumns_line3_timesTHREE_input2_3_ ;
    wire MixColumns_line3_timesTHREE_input2_4_ ;
    wire calcRCon_n38 ;
    wire calcRCon_n37 ;
    wire calcRCon_n36 ;
    wire calcRCon_n35 ;
    wire calcRCon_n34 ;
    wire calcRCon_n33 ;
    wire calcRCon_n32 ;
    wire calcRCon_n31 ;
    wire calcRCon_n30 ;
    wire calcRCon_n29 ;
    wire calcRCon_n28 ;
    wire calcRCon_n27 ;
    wire calcRCon_n26 ;
    wire calcRCon_n25 ;
    wire calcRCon_n24 ;
    wire calcRCon_n23 ;
    wire calcRCon_n22 ;
    wire calcRCon_n21 ;
    wire calcRCon_n20 ;
    wire calcRCon_n19 ;
    wire calcRCon_n18 ;
    wire calcRCon_n17 ;
    wire calcRCon_n10 ;
    wire calcRCon_n9 ;
    wire calcRCon_n8 ;
    wire calcRCon_n7 ;
    wire calcRCon_n6 ;
    wire calcRCon_n5 ;
    wire calcRCon_n3 ;
    wire calcRCon_n11 ;
    wire calcRCon_n44 ;
    wire calcRCon_n16 ;
    wire calcRCon_n45 ;
    wire calcRCon_n46 ;
    wire calcRCon_n47 ;
    wire calcRCon_n15 ;
    wire calcRCon_n48 ;
    wire calcRCon_n12 ;
    wire calcRCon_n49 ;
    wire calcRCon_n14 ;
    wire calcRCon_n50 ;
    wire calcRCon_n13 ;
    wire calcRCon_s_current_state_0_ ;
    wire calcRCon_s_current_state_1_ ;
    wire calcRCon_s_current_state_2_ ;
    wire calcRCon_s_current_state_3_ ;
    wire calcRCon_s_current_state_4_ ;
    wire calcRCon_s_current_state_5_ ;
    wire calcRCon_s_current_state_6_ ;
    wire calcRCon_n51 ;
    wire Inst_bSbox_L29 ;
    wire Inst_bSbox_L28 ;
    wire Inst_bSbox_L27 ;
    wire Inst_bSbox_L26 ;
    wire Inst_bSbox_L25 ;
    wire Inst_bSbox_L24 ;
    wire Inst_bSbox_L23 ;
    wire Inst_bSbox_L22 ;
    wire Inst_bSbox_L21 ;
    wire Inst_bSbox_L20 ;
    wire Inst_bSbox_L19 ;
    wire Inst_bSbox_L18 ;
    wire Inst_bSbox_L17 ;
    wire Inst_bSbox_L16 ;
    wire Inst_bSbox_L15 ;
    wire Inst_bSbox_L14 ;
    wire Inst_bSbox_L13 ;
    wire Inst_bSbox_L12 ;
    wire Inst_bSbox_L11 ;
    wire Inst_bSbox_L10 ;
    wire Inst_bSbox_L9 ;
    wire Inst_bSbox_L8 ;
    wire Inst_bSbox_L7 ;
    wire Inst_bSbox_L6 ;
    wire Inst_bSbox_L5 ;
    wire Inst_bSbox_L4 ;
    wire Inst_bSbox_L3 ;
    wire Inst_bSbox_L2 ;
    wire Inst_bSbox_L1 ;
    wire Inst_bSbox_L0 ;
    wire Inst_bSbox_M63 ;
    wire Inst_bSbox_M62 ;
    wire Inst_bSbox_M61 ;
    wire Inst_bSbox_M60 ;
    wire Inst_bSbox_M59 ;
    wire Inst_bSbox_M58 ;
    wire Inst_bSbox_M57 ;
    wire Inst_bSbox_M56 ;
    wire Inst_bSbox_M55 ;
    wire Inst_bSbox_M54 ;
    wire Inst_bSbox_M53 ;
    wire Inst_bSbox_M52 ;
    wire Inst_bSbox_M51 ;
    wire Inst_bSbox_M50 ;
    wire Inst_bSbox_M49 ;
    wire Inst_bSbox_M48 ;
    wire Inst_bSbox_M47 ;
    wire Inst_bSbox_M46 ;
    wire Inst_bSbox_M45 ;
    wire Inst_bSbox_M44 ;
    wire Inst_bSbox_M43 ;
    wire Inst_bSbox_M42 ;
    wire Inst_bSbox_M41 ;
    wire Inst_bSbox_M40 ;
    wire Inst_bSbox_M39 ;
    wire Inst_bSbox_M38 ;
    wire Inst_bSbox_M37 ;
    wire Inst_bSbox_M36 ;
    wire Inst_bSbox_M35 ;
    wire Inst_bSbox_M34 ;
    wire Inst_bSbox_M33 ;
    wire Inst_bSbox_M32 ;
    wire Inst_bSbox_M31 ;
    wire Inst_bSbox_M30 ;
    wire Inst_bSbox_M29 ;
    wire Inst_bSbox_M28 ;
    wire Inst_bSbox_M27 ;
    wire Inst_bSbox_M26 ;
    wire Inst_bSbox_M25 ;
    wire Inst_bSbox_M24 ;
    wire Inst_bSbox_M23 ;
    wire Inst_bSbox_M22 ;
    wire Inst_bSbox_M21 ;
    wire Inst_bSbox_M20 ;
    wire Inst_bSbox_M19 ;
    wire Inst_bSbox_M18 ;
    wire Inst_bSbox_M17 ;
    wire Inst_bSbox_M16 ;
    wire Inst_bSbox_M15 ;
    wire Inst_bSbox_M14 ;
    wire Inst_bSbox_M13 ;
    wire Inst_bSbox_M12 ;
    wire Inst_bSbox_M11 ;
    wire Inst_bSbox_M10 ;
    wire Inst_bSbox_M9 ;
    wire Inst_bSbox_M8 ;
    wire Inst_bSbox_M7 ;
    wire Inst_bSbox_M6 ;
    wire Inst_bSbox_M5 ;
    wire Inst_bSbox_M4 ;
    wire Inst_bSbox_M3 ;
    wire Inst_bSbox_M2 ;
    wire Inst_bSbox_M1 ;
    wire Inst_bSbox_T27 ;
    wire Inst_bSbox_T26 ;
    wire Inst_bSbox_T25 ;
    wire Inst_bSbox_T24 ;
    wire Inst_bSbox_T23 ;
    wire Inst_bSbox_T22 ;
    wire Inst_bSbox_T21 ;
    wire Inst_bSbox_T20 ;
    wire Inst_bSbox_T19 ;
    wire Inst_bSbox_T18 ;
    wire Inst_bSbox_T17 ;
    wire Inst_bSbox_T16 ;
    wire Inst_bSbox_T15 ;
    wire Inst_bSbox_T14 ;
    wire Inst_bSbox_T13 ;
    wire Inst_bSbox_T12 ;
    wire Inst_bSbox_T11 ;
    wire Inst_bSbox_T10 ;
    wire Inst_bSbox_T9 ;
    wire Inst_bSbox_T8 ;
    wire Inst_bSbox_T7 ;
    wire Inst_bSbox_T6 ;
    wire Inst_bSbox_T5 ;
    wire Inst_bSbox_T4 ;
    wire Inst_bSbox_T3 ;
    wire Inst_bSbox_T2 ;
    wire Inst_bSbox_T1 ;
    wire [7:0] SboxOut ;
    wire [7:0] StateOutXORroundKey ;
    wire [7:0] StateIn ;
    wire [31:0] StateInMC ;
    wire [31:0] MCout ;
    wire [7:0] keyStateIn ;
    wire [7:0] roundConstant ;
    wire [7:0] keySBIn ;
    wire [7:0] SboxIn ;
    wire [7:0] stateArray_input_MC ;
    wire [7:0] stateArray_outS30ser_MC ;
    wire [7:0] stateArray_outS20ser_MC ;
    wire [7:0] stateArray_outS10ser_MC ;
    wire [7:0] stateArray_inS33ser ;
    wire [7:0] stateArray_inS32ser ;
    wire [7:0] stateArray_inS31ser ;
    wire [7:0] stateArray_inS30ser ;
    wire [7:0] stateArray_inS23ser ;
    wire [7:0] stateArray_inS22ser ;
    wire [7:0] stateArray_inS21ser ;
    wire [7:0] stateArray_inS20ser ;
    wire [7:0] stateArray_inS13ser ;
    wire [7:0] stateArray_inS12ser ;
    wire [7:0] stateArray_inS11ser ;
    wire [7:0] stateArray_inS10ser ;
    wire [7:0] stateArray_inS03ser ;
    wire [7:0] stateArray_inS02ser ;
    wire [7:0] stateArray_inS01ser ;
    wire [7:0] stateArray_inS00ser ;
    wire [7:0] KeyArray_outS01ser_p ;
    wire [7:0] KeyArray_outS01ser_XOR_00 ;
    wire [7:0] KeyArray_outS33ser ;
    wire [7:0] KeyArray_inS33ser ;
    wire [7:0] KeyArray_outS32ser ;
    wire [7:0] KeyArray_inS32ser ;
    wire [7:0] KeyArray_outS31ser ;
    wire [7:0] KeyArray_inS31ser ;
    wire [7:0] KeyArray_outS30ser ;
    wire [7:0] KeyArray_inS30par ;
    wire [7:0] KeyArray_inS30ser ;
    wire [7:0] KeyArray_outS23ser ;
    wire [7:0] KeyArray_inS23ser ;
    wire [7:0] KeyArray_outS22ser ;
    wire [7:0] KeyArray_inS22ser ;
    wire [7:0] KeyArray_outS21ser ;
    wire [7:0] KeyArray_inS21ser ;
    wire [7:0] KeyArray_outS20ser ;
    wire [7:0] KeyArray_inS20ser ;
    wire [7:0] KeyArray_inS13ser ;
    wire [7:0] KeyArray_outS12ser ;
    wire [7:0] KeyArray_inS12ser ;
    wire [7:0] KeyArray_outS11ser ;
    wire [7:0] KeyArray_inS11ser ;
    wire [7:0] KeyArray_outS10ser ;
    wire [7:0] KeyArray_inS10ser ;
    wire [7:0] KeyArray_outS03ser ;
    wire [7:0] KeyArray_inS03ser ;
    wire [7:0] KeyArray_outS02ser ;
    wire [7:0] KeyArray_inS02ser ;
    wire [7:0] KeyArray_inS01ser ;
    wire [7:0] KeyArray_inS00ser ;
    wire [7:0] MixColumns_line0_S13 ;
    wire [4:1] MixColumns_line0_S02 ;
    wire [4:1] MixColumns_line0_timesTHREE_input2 ;
    wire [7:0] MixColumns_line1_S13 ;
    wire [4:1] MixColumns_line1_timesTHREE_input2 ;
    wire [7:0] MixColumns_line2_S13 ;
    wire [4:1] MixColumns_line2_timesTHREE_input2 ;
    wire [7:0] MixColumns_line3_S13 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4373 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4379 ;
    wire new_AGEMA_signal_4380 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4497 ;
    wire new_AGEMA_signal_4498 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire clk_gated ;

    /* cells in depth 0 */
    INV_X1 U28 ( .A (selSR), .ZN (n12) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U29 ( .a ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, new_AGEMA_signal_1985, keyStateIn[0]}), .c ({new_AGEMA_signal_1990, new_AGEMA_signal_1989, new_AGEMA_signal_1988, StateOutXORroundKey[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U30 ( .a ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .b ({new_AGEMA_signal_1996, new_AGEMA_signal_1995, new_AGEMA_signal_1994, keyStateIn[1]}), .c ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, new_AGEMA_signal_1997, StateOutXORroundKey[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U31 ( .a ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .b ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, new_AGEMA_signal_2003, keyStateIn[2]}), .c ({new_AGEMA_signal_2008, new_AGEMA_signal_2007, new_AGEMA_signal_2006, StateOutXORroundKey[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U32 ( .a ({ciphertext_s3[123], ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}), .b ({new_AGEMA_signal_2014, new_AGEMA_signal_2013, new_AGEMA_signal_2012, keyStateIn[3]}), .c ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, new_AGEMA_signal_2015, StateOutXORroundKey[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U33 ( .a ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, new_AGEMA_signal_2021, keyStateIn[4]}), .c ({new_AGEMA_signal_2026, new_AGEMA_signal_2025, new_AGEMA_signal_2024, StateOutXORroundKey[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U34 ( .a ({ciphertext_s3[125], ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .b ({new_AGEMA_signal_2032, new_AGEMA_signal_2031, new_AGEMA_signal_2030, keyStateIn[5]}), .c ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, new_AGEMA_signal_2033, StateOutXORroundKey[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U35 ( .a ({ciphertext_s3[126], ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .b ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, new_AGEMA_signal_2039, keyStateIn[6]}), .c ({new_AGEMA_signal_2044, new_AGEMA_signal_2043, new_AGEMA_signal_2042, StateOutXORroundKey[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U36 ( .a ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_2050, new_AGEMA_signal_2049, new_AGEMA_signal_2048, keyStateIn[7]}), .c ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, new_AGEMA_signal_2051, StateOutXORroundKey[7]}) ) ;
    NAND2_X1 U37 ( .A1 (intFinal), .A2 (finalStep), .ZN (n13) ) ;
    NOR2_X1 U38 ( .A1 (n10), .A2 (n13), .ZN (done) ) ;
    AND2_X1 U39 ( .A1 (notFirst), .A2 (selXOR), .ZN (intselXOR) ) ;
    INV_X1 U40 ( .A (start), .ZN (n9) ) ;
    NOR2_X1 ctrl_U20 ( .A1 (ctrl_n16), .A2 (ctrl_n4), .ZN (ctrl_nRstSeq4) ) ;
    XNOR2_X1 ctrl_U19 ( .A (ctrl_seq6Out_4_), .B (ctrl_seq6In_1_), .ZN (ctrl_n13) ) ;
    NOR2_X1 ctrl_U18 ( .A1 (ctrl_n15), .A2 (ctrl_n14), .ZN (finalStep) ) ;
    NAND2_X1 ctrl_U17 ( .A1 (ctrl_seq4In_1_), .A2 (ctrl_n2), .ZN (ctrl_n14) ) ;
    INV_X1 ctrl_U16 ( .A (ctrl_n16), .ZN (ctrl_n15) ) ;
    INV_X1 ctrl_U15 ( .A (ctrl_seq4Out_1_), .ZN (ctrl_n2) ) ;
    NAND2_X1 ctrl_U14 ( .A1 (ctrl_n11), .A2 (ctrl_n10), .ZN (ctrl_N14) ) ;
    NAND2_X1 ctrl_U13 ( .A1 (selXOR), .A2 (ctrl_n6), .ZN (ctrl_n11) ) ;
    NOR2_X1 ctrl_U12 ( .A1 (ctrl_seq6In_3_), .A2 (ctrl_seq6Out_4_), .ZN (ctrl_n7) ) ;
    NOR2_X1 ctrl_U11 ( .A1 (ctrl_seq6In_1_), .A2 (ctrl_seq6In_4_), .ZN (ctrl_n8) ) ;
    NOR2_X1 ctrl_U10 ( .A1 (ctrl_n4), .A2 (ctrl_n5), .ZN (selXOR) ) ;
    NOR2_X1 ctrl_U9 ( .A1 (ctrl_seq4Out_1_), .A2 (ctrl_seq4In_1_), .ZN (ctrl_n5) ) ;
    INV_X1 ctrl_U8 ( .A (nReset), .ZN (ctrl_n4) ) ;
    NAND2_X1 ctrl_U7 ( .A1 (ctrl_n8), .A2 (ctrl_n7), .ZN (ctrl_n9) ) ;
    NOR2_X1 ctrl_U6 ( .A1 (ctrl_seq6In_2_), .A2 (ctrl_n9), .ZN (ctrl_n16) ) ;
    NAND2_X1 ctrl_U5 ( .A1 (nReset), .A2 (ctrl_n16), .ZN (ctrl_n10) ) ;
    INV_X1 ctrl_U4 ( .A (ctrl_n10), .ZN (selSR) ) ;
    NOR2_X1 ctrl_U3 ( .A1 (ctrl_n12), .A2 (ctrl_n4), .ZN (selMC) ) ;
    MUX2_X1 ctrl_seq6_SFF_0_MUXInst_U1 ( .S (nReset), .A (1'b1), .B (ctrl_n13), .Z (ctrl_seq6_SFF_0_QD) ) ;
    MUX2_X1 ctrl_seq6_SFF_1_MUXInst_U1 ( .S (nReset), .A (1'b0), .B (ctrl_seq6In_1_), .Z (ctrl_seq6_SFF_1_QD) ) ;
    MUX2_X1 ctrl_seq6_SFF_2_MUXInst_U1 ( .S (nReset), .A (1'b1), .B (ctrl_seq6In_2_), .Z (ctrl_seq6_SFF_2_QD) ) ;
    MUX2_X1 ctrl_seq6_SFF_3_MUXInst_U1 ( .S (nReset), .A (1'b0), .B (ctrl_seq6In_3_), .Z (ctrl_seq6_SFF_3_QD) ) ;
    MUX2_X1 ctrl_seq6_SFF_4_MUXInst_U1 ( .S (nReset), .A (1'b1), .B (ctrl_seq6In_4_), .Z (ctrl_seq6_SFF_4_QD) ) ;
    MUX2_X1 ctrl_seq4_SFF_0_MUXInst_U1 ( .S (ctrl_nRstSeq4), .A (1'b1), .B (ctrl_n2), .Z (ctrl_seq4_SFF_0_QD) ) ;
    MUX2_X1 ctrl_seq4_SFF_1_MUXInst_U1 ( .S (ctrl_nRstSeq4), .A (1'b0), .B (ctrl_seq4In_1_), .Z (ctrl_seq4_SFF_1_QD) ) ;
    INV_X1 ctrl_CSselMC_reg_U1 ( .A (ctrl_n6), .ZN (ctrl_n12) ) ;
    INV_X1 stateArray_U21 ( .A (selMC), .ZN (stateArray_n24) ) ;
    INV_X1 stateArray_U20 ( .A (stateArray_n24), .ZN (stateArray_n22) ) ;
    INV_X1 stateArray_U19 ( .A (nReset), .ZN (stateArray_n33) ) ;
    INV_X1 stateArray_U18 ( .A (stateArray_n33), .ZN (stateArray_n25) ) ;
    INV_X1 stateArray_U17 ( .A (stateArray_n21), .ZN (stateArray_n13) ) ;
    INV_X1 stateArray_U16 ( .A (stateArray_n24), .ZN (stateArray_n23) ) ;
    INV_X1 stateArray_U15 ( .A (stateArray_n33), .ZN (stateArray_n29) ) ;
    INV_X1 stateArray_U14 ( .A (stateArray_n21), .ZN (stateArray_n17) ) ;
    INV_X1 stateArray_U13 ( .A (stateArray_n33), .ZN (stateArray_n31) ) ;
    INV_X1 stateArray_U12 ( .A (stateArray_n21), .ZN (stateArray_n19) ) ;
    INV_X1 stateArray_U11 ( .A (stateArray_n33), .ZN (stateArray_n27) ) ;
    INV_X1 stateArray_U10 ( .A (stateArray_n21), .ZN (stateArray_n15) ) ;
    INV_X1 stateArray_U9 ( .A (stateArray_n33), .ZN (stateArray_n32) ) ;
    INV_X1 stateArray_U8 ( .A (stateArray_n21), .ZN (stateArray_n20) ) ;
    INV_X1 stateArray_U7 ( .A (stateArray_n33), .ZN (stateArray_n30) ) ;
    INV_X1 stateArray_U6 ( .A (stateArray_n21), .ZN (stateArray_n18) ) ;
    INV_X1 stateArray_U5 ( .A (stateArray_n33), .ZN (stateArray_n28) ) ;
    INV_X1 stateArray_U4 ( .A (stateArray_n21), .ZN (stateArray_n16) ) ;
    INV_X1 stateArray_U3 ( .A (stateArray_n33), .ZN (stateArray_n26) ) ;
    INV_X1 stateArray_U2 ( .A (stateArray_n21), .ZN (stateArray_n14) ) ;
    INV_X1 stateArray_U1 ( .A (selSR), .ZN (stateArray_n21) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S00reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2506, new_AGEMA_signal_2505, new_AGEMA_signal_2504, stateArray_inS00ser[0]}), .a ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_5416, new_AGEMA_signal_5415, new_AGEMA_signal_5414, stateArray_S00reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S00reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, new_AGEMA_signal_2513, stateArray_inS00ser[1]}), .a ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_5419, new_AGEMA_signal_5418, new_AGEMA_signal_5417, stateArray_S00reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S00reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2524, new_AGEMA_signal_2523, new_AGEMA_signal_2522, stateArray_inS00ser[2]}), .a ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_5422, new_AGEMA_signal_5421, new_AGEMA_signal_5420, stateArray_S00reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S00reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, new_AGEMA_signal_2531, stateArray_inS00ser[3]}), .a ({ciphertext_s3[123], ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_5425, new_AGEMA_signal_5424, new_AGEMA_signal_5423, stateArray_S00reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S00reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2542, new_AGEMA_signal_2541, new_AGEMA_signal_2540, stateArray_inS00ser[4]}), .a ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_5428, new_AGEMA_signal_5427, new_AGEMA_signal_5426, stateArray_S00reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S00reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, new_AGEMA_signal_2549, stateArray_inS00ser[5]}), .a ({ciphertext_s3[125], ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_5431, new_AGEMA_signal_5430, new_AGEMA_signal_5429, stateArray_S00reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S00reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2560, new_AGEMA_signal_2559, new_AGEMA_signal_2558, stateArray_inS00ser[6]}), .a ({ciphertext_s3[126], ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .c ({new_AGEMA_signal_5434, new_AGEMA_signal_5433, new_AGEMA_signal_5432, stateArray_S00reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S00reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, new_AGEMA_signal_2567, stateArray_inS00ser[7]}), .a ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .c ({new_AGEMA_signal_5437, new_AGEMA_signal_5436, new_AGEMA_signal_5435, stateArray_S00reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S01reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2578, new_AGEMA_signal_2577, new_AGEMA_signal_2576, stateArray_inS01ser[0]}), .a ({ciphertext_s3[112], ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_5440, new_AGEMA_signal_5439, new_AGEMA_signal_5438, stateArray_S01reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S01reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, new_AGEMA_signal_2585, stateArray_inS01ser[1]}), .a ({ciphertext_s3[113], ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_5443, new_AGEMA_signal_5442, new_AGEMA_signal_5441, stateArray_S01reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S01reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2596, new_AGEMA_signal_2595, new_AGEMA_signal_2594, stateArray_inS01ser[2]}), .a ({ciphertext_s3[114], ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_5446, new_AGEMA_signal_5445, new_AGEMA_signal_5444, stateArray_S01reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S01reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, new_AGEMA_signal_2603, stateArray_inS01ser[3]}), .a ({ciphertext_s3[115], ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}), .c ({new_AGEMA_signal_5449, new_AGEMA_signal_5448, new_AGEMA_signal_5447, stateArray_S01reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S01reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2614, new_AGEMA_signal_2613, new_AGEMA_signal_2612, stateArray_inS01ser[4]}), .a ({ciphertext_s3[116], ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .c ({new_AGEMA_signal_5452, new_AGEMA_signal_5451, new_AGEMA_signal_5450, stateArray_S01reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S01reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, new_AGEMA_signal_2621, stateArray_inS01ser[5]}), .a ({ciphertext_s3[117], ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}), .c ({new_AGEMA_signal_5455, new_AGEMA_signal_5454, new_AGEMA_signal_5453, stateArray_S01reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S01reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2632, new_AGEMA_signal_2631, new_AGEMA_signal_2630, stateArray_inS01ser[6]}), .a ({ciphertext_s3[118], ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}), .c ({new_AGEMA_signal_5458, new_AGEMA_signal_5457, new_AGEMA_signal_5456, stateArray_S01reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S01reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, new_AGEMA_signal_2639, stateArray_inS01ser[7]}), .a ({ciphertext_s3[119], ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .c ({new_AGEMA_signal_5461, new_AGEMA_signal_5460, new_AGEMA_signal_5459, stateArray_S01reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S02reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2650, new_AGEMA_signal_2649, new_AGEMA_signal_2648, stateArray_inS02ser[0]}), .a ({ciphertext_s3[104], ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_5464, new_AGEMA_signal_5463, new_AGEMA_signal_5462, stateArray_S02reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S02reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, new_AGEMA_signal_2657, stateArray_inS02ser[1]}), .a ({ciphertext_s3[105], ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_5467, new_AGEMA_signal_5466, new_AGEMA_signal_5465, stateArray_S02reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S02reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2668, new_AGEMA_signal_2667, new_AGEMA_signal_2666, stateArray_inS02ser[2]}), .a ({ciphertext_s3[106], ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_5470, new_AGEMA_signal_5469, new_AGEMA_signal_5468, stateArray_S02reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S02reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, new_AGEMA_signal_2675, stateArray_inS02ser[3]}), .a ({ciphertext_s3[107], ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}), .c ({new_AGEMA_signal_5473, new_AGEMA_signal_5472, new_AGEMA_signal_5471, stateArray_S02reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S02reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2686, new_AGEMA_signal_2685, new_AGEMA_signal_2684, stateArray_inS02ser[4]}), .a ({ciphertext_s3[108], ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .c ({new_AGEMA_signal_5476, new_AGEMA_signal_5475, new_AGEMA_signal_5474, stateArray_S02reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S02reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, new_AGEMA_signal_2693, stateArray_inS02ser[5]}), .a ({ciphertext_s3[109], ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}), .c ({new_AGEMA_signal_5479, new_AGEMA_signal_5478, new_AGEMA_signal_5477, stateArray_S02reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S02reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, new_AGEMA_signal_2702, stateArray_inS02ser[6]}), .a ({ciphertext_s3[110], ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}), .c ({new_AGEMA_signal_5482, new_AGEMA_signal_5481, new_AGEMA_signal_5480, stateArray_S02reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S02reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, new_AGEMA_signal_2711, stateArray_inS02ser[7]}), .a ({ciphertext_s3[111], ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .c ({new_AGEMA_signal_5485, new_AGEMA_signal_5484, new_AGEMA_signal_5483, stateArray_S02reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S03reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_5176, new_AGEMA_signal_5175, new_AGEMA_signal_5174, stateArray_inS03ser[0]}), .a ({ciphertext_s3[96], ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_5488, new_AGEMA_signal_5487, new_AGEMA_signal_5486, stateArray_S03reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S03reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_5182, new_AGEMA_signal_5181, new_AGEMA_signal_5180, stateArray_inS03ser[1]}), .a ({ciphertext_s3[97], ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_5491, new_AGEMA_signal_5490, new_AGEMA_signal_5489, stateArray_S03reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S03reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_5188, new_AGEMA_signal_5187, new_AGEMA_signal_5186, stateArray_inS03ser[2]}), .a ({ciphertext_s3[98], ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_5494, new_AGEMA_signal_5493, new_AGEMA_signal_5492, stateArray_S03reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S03reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_5194, new_AGEMA_signal_5193, new_AGEMA_signal_5192, stateArray_inS03ser[3]}), .a ({ciphertext_s3[99], ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}), .c ({new_AGEMA_signal_5497, new_AGEMA_signal_5496, new_AGEMA_signal_5495, stateArray_S03reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S03reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_5200, new_AGEMA_signal_5199, new_AGEMA_signal_5198, stateArray_inS03ser[4]}), .a ({ciphertext_s3[100], ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .c ({new_AGEMA_signal_5500, new_AGEMA_signal_5499, new_AGEMA_signal_5498, stateArray_S03reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S03reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_5206, new_AGEMA_signal_5205, new_AGEMA_signal_5204, stateArray_inS03ser[5]}), .a ({ciphertext_s3[101], ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}), .c ({new_AGEMA_signal_5503, new_AGEMA_signal_5502, new_AGEMA_signal_5501, stateArray_S03reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S03reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_5212, new_AGEMA_signal_5211, new_AGEMA_signal_5210, stateArray_inS03ser[6]}), .a ({ciphertext_s3[102], ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}), .c ({new_AGEMA_signal_5506, new_AGEMA_signal_5505, new_AGEMA_signal_5504, stateArray_S03reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S03reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_5218, new_AGEMA_signal_5217, new_AGEMA_signal_5216, stateArray_inS03ser[7]}), .a ({ciphertext_s3[103], ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .c ({new_AGEMA_signal_5509, new_AGEMA_signal_5508, new_AGEMA_signal_5507, stateArray_S03reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S10reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2722, new_AGEMA_signal_2721, new_AGEMA_signal_2720, stateArray_inS10ser[0]}), .a ({ciphertext_s3[80], ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_5512, new_AGEMA_signal_5511, new_AGEMA_signal_5510, stateArray_S10reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S10reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, new_AGEMA_signal_2729, stateArray_inS10ser[1]}), .a ({ciphertext_s3[81], ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_5515, new_AGEMA_signal_5514, new_AGEMA_signal_5513, stateArray_S10reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S10reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2740, new_AGEMA_signal_2739, new_AGEMA_signal_2738, stateArray_inS10ser[2]}), .a ({ciphertext_s3[82], ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_5518, new_AGEMA_signal_5517, new_AGEMA_signal_5516, stateArray_S10reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S10reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, new_AGEMA_signal_2747, stateArray_inS10ser[3]}), .a ({ciphertext_s3[83], ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}), .c ({new_AGEMA_signal_5521, new_AGEMA_signal_5520, new_AGEMA_signal_5519, stateArray_S10reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S10reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2758, new_AGEMA_signal_2757, new_AGEMA_signal_2756, stateArray_inS10ser[4]}), .a ({ciphertext_s3[84], ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .c ({new_AGEMA_signal_5524, new_AGEMA_signal_5523, new_AGEMA_signal_5522, stateArray_S10reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S10reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, new_AGEMA_signal_2765, stateArray_inS10ser[5]}), .a ({ciphertext_s3[85], ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}), .c ({new_AGEMA_signal_5527, new_AGEMA_signal_5526, new_AGEMA_signal_5525, stateArray_S10reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S10reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2776, new_AGEMA_signal_2775, new_AGEMA_signal_2774, stateArray_inS10ser[6]}), .a ({ciphertext_s3[86], ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}), .c ({new_AGEMA_signal_5530, new_AGEMA_signal_5529, new_AGEMA_signal_5528, stateArray_S10reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S10reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, new_AGEMA_signal_2783, stateArray_inS10ser[7]}), .a ({ciphertext_s3[87], ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .c ({new_AGEMA_signal_5533, new_AGEMA_signal_5532, new_AGEMA_signal_5531, stateArray_S10reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S11reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2794, new_AGEMA_signal_2793, new_AGEMA_signal_2792, stateArray_inS11ser[0]}), .a ({ciphertext_s3[72], ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_5536, new_AGEMA_signal_5535, new_AGEMA_signal_5534, stateArray_S11reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S11reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, new_AGEMA_signal_2801, stateArray_inS11ser[1]}), .a ({ciphertext_s3[73], ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_5539, new_AGEMA_signal_5538, new_AGEMA_signal_5537, stateArray_S11reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S11reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2812, new_AGEMA_signal_2811, new_AGEMA_signal_2810, stateArray_inS11ser[2]}), .a ({ciphertext_s3[74], ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_5542, new_AGEMA_signal_5541, new_AGEMA_signal_5540, stateArray_S11reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S11reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, new_AGEMA_signal_2819, stateArray_inS11ser[3]}), .a ({ciphertext_s3[75], ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}), .c ({new_AGEMA_signal_5545, new_AGEMA_signal_5544, new_AGEMA_signal_5543, stateArray_S11reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S11reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2830, new_AGEMA_signal_2829, new_AGEMA_signal_2828, stateArray_inS11ser[4]}), .a ({ciphertext_s3[76], ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .c ({new_AGEMA_signal_5548, new_AGEMA_signal_5547, new_AGEMA_signal_5546, stateArray_S11reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S11reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, new_AGEMA_signal_2837, stateArray_inS11ser[5]}), .a ({ciphertext_s3[77], ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}), .c ({new_AGEMA_signal_5551, new_AGEMA_signal_5550, new_AGEMA_signal_5549, stateArray_S11reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S11reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2848, new_AGEMA_signal_2847, new_AGEMA_signal_2846, stateArray_inS11ser[6]}), .a ({ciphertext_s3[78], ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}), .c ({new_AGEMA_signal_5554, new_AGEMA_signal_5553, new_AGEMA_signal_5552, stateArray_S11reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S11reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, new_AGEMA_signal_2855, stateArray_inS11ser[7]}), .a ({ciphertext_s3[79], ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .c ({new_AGEMA_signal_5557, new_AGEMA_signal_5556, new_AGEMA_signal_5555, stateArray_S11reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S12reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2866, new_AGEMA_signal_2865, new_AGEMA_signal_2864, stateArray_inS12ser[0]}), .a ({ciphertext_s3[64], ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_5560, new_AGEMA_signal_5559, new_AGEMA_signal_5558, stateArray_S12reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S12reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, new_AGEMA_signal_2873, stateArray_inS12ser[1]}), .a ({ciphertext_s3[65], ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_5563, new_AGEMA_signal_5562, new_AGEMA_signal_5561, stateArray_S12reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S12reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2884, new_AGEMA_signal_2883, new_AGEMA_signal_2882, stateArray_inS12ser[2]}), .a ({ciphertext_s3[66], ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_5566, new_AGEMA_signal_5565, new_AGEMA_signal_5564, stateArray_S12reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S12reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, new_AGEMA_signal_2891, stateArray_inS12ser[3]}), .a ({ciphertext_s3[67], ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}), .c ({new_AGEMA_signal_5569, new_AGEMA_signal_5568, new_AGEMA_signal_5567, stateArray_S12reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S12reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2902, new_AGEMA_signal_2901, new_AGEMA_signal_2900, stateArray_inS12ser[4]}), .a ({ciphertext_s3[68], ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .c ({new_AGEMA_signal_5572, new_AGEMA_signal_5571, new_AGEMA_signal_5570, stateArray_S12reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S12reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, new_AGEMA_signal_2909, stateArray_inS12ser[5]}), .a ({ciphertext_s3[69], ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}), .c ({new_AGEMA_signal_5575, new_AGEMA_signal_5574, new_AGEMA_signal_5573, stateArray_S12reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S12reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2920, new_AGEMA_signal_2919, new_AGEMA_signal_2918, stateArray_inS12ser[6]}), .a ({ciphertext_s3[70], ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}), .c ({new_AGEMA_signal_5578, new_AGEMA_signal_5577, new_AGEMA_signal_5576, stateArray_S12reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S12reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, new_AGEMA_signal_2927, stateArray_inS12ser[7]}), .a ({ciphertext_s3[71], ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .c ({new_AGEMA_signal_5581, new_AGEMA_signal_5580, new_AGEMA_signal_5579, stateArray_S12reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S13reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_5224, new_AGEMA_signal_5223, new_AGEMA_signal_5222, stateArray_inS13ser[0]}), .a ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_5584, new_AGEMA_signal_5583, new_AGEMA_signal_5582, stateArray_S13reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S13reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_5230, new_AGEMA_signal_5229, new_AGEMA_signal_5228, stateArray_inS13ser[1]}), .a ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_5587, new_AGEMA_signal_5586, new_AGEMA_signal_5585, stateArray_S13reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S13reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_5236, new_AGEMA_signal_5235, new_AGEMA_signal_5234, stateArray_inS13ser[2]}), .a ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_5590, new_AGEMA_signal_5589, new_AGEMA_signal_5588, stateArray_S13reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S13reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_5242, new_AGEMA_signal_5241, new_AGEMA_signal_5240, stateArray_inS13ser[3]}), .a ({ciphertext_s3[91], ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_5593, new_AGEMA_signal_5592, new_AGEMA_signal_5591, stateArray_S13reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S13reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_5248, new_AGEMA_signal_5247, new_AGEMA_signal_5246, stateArray_inS13ser[4]}), .a ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_5596, new_AGEMA_signal_5595, new_AGEMA_signal_5594, stateArray_S13reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S13reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_5254, new_AGEMA_signal_5253, new_AGEMA_signal_5252, stateArray_inS13ser[5]}), .a ({ciphertext_s3[93], ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_5599, new_AGEMA_signal_5598, new_AGEMA_signal_5597, stateArray_S13reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S13reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_5260, new_AGEMA_signal_5259, new_AGEMA_signal_5258, stateArray_inS13ser[6]}), .a ({ciphertext_s3[94], ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .c ({new_AGEMA_signal_5602, new_AGEMA_signal_5601, new_AGEMA_signal_5600, stateArray_S13reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S13reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_5266, new_AGEMA_signal_5265, new_AGEMA_signal_5264, stateArray_inS13ser[7]}), .a ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .c ({new_AGEMA_signal_5605, new_AGEMA_signal_5604, new_AGEMA_signal_5603, stateArray_S13reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S20reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2938, new_AGEMA_signal_2937, new_AGEMA_signal_2936, stateArray_inS20ser[0]}), .a ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_5608, new_AGEMA_signal_5607, new_AGEMA_signal_5606, stateArray_S20reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S20reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, new_AGEMA_signal_2945, stateArray_inS20ser[1]}), .a ({ciphertext_s3[41], ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_5611, new_AGEMA_signal_5610, new_AGEMA_signal_5609, stateArray_S20reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S20reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2956, new_AGEMA_signal_2955, new_AGEMA_signal_2954, stateArray_inS20ser[2]}), .a ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5614, new_AGEMA_signal_5613, new_AGEMA_signal_5612, stateArray_S20reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S20reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, new_AGEMA_signal_2963, stateArray_inS20ser[3]}), .a ({ciphertext_s3[43], ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .c ({new_AGEMA_signal_5617, new_AGEMA_signal_5616, new_AGEMA_signal_5615, stateArray_S20reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S20reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2974, new_AGEMA_signal_2973, new_AGEMA_signal_2972, stateArray_inS20ser[4]}), .a ({ciphertext_s3[44], ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .c ({new_AGEMA_signal_5620, new_AGEMA_signal_5619, new_AGEMA_signal_5618, stateArray_S20reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S20reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, new_AGEMA_signal_2981, stateArray_inS20ser[5]}), .a ({ciphertext_s3[45], ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .c ({new_AGEMA_signal_5623, new_AGEMA_signal_5622, new_AGEMA_signal_5621, stateArray_S20reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S20reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2992, new_AGEMA_signal_2991, new_AGEMA_signal_2990, stateArray_inS20ser[6]}), .a ({ciphertext_s3[46], ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .c ({new_AGEMA_signal_5626, new_AGEMA_signal_5625, new_AGEMA_signal_5624, stateArray_S20reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S20reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, new_AGEMA_signal_2999, stateArray_inS20ser[7]}), .a ({ciphertext_s3[47], ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .c ({new_AGEMA_signal_5629, new_AGEMA_signal_5628, new_AGEMA_signal_5627, stateArray_S20reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S21reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_3010, new_AGEMA_signal_3009, new_AGEMA_signal_3008, stateArray_inS21ser[0]}), .a ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_5632, new_AGEMA_signal_5631, new_AGEMA_signal_5630, stateArray_S21reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S21reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, new_AGEMA_signal_3017, stateArray_inS21ser[1]}), .a ({ciphertext_s3[33], ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_5635, new_AGEMA_signal_5634, new_AGEMA_signal_5633, stateArray_S21reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S21reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_3028, new_AGEMA_signal_3027, new_AGEMA_signal_3026, stateArray_inS21ser[2]}), .a ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5638, new_AGEMA_signal_5637, new_AGEMA_signal_5636, stateArray_S21reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S21reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, new_AGEMA_signal_3035, stateArray_inS21ser[3]}), .a ({ciphertext_s3[35], ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .c ({new_AGEMA_signal_5641, new_AGEMA_signal_5640, new_AGEMA_signal_5639, stateArray_S21reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S21reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_3046, new_AGEMA_signal_3045, new_AGEMA_signal_3044, stateArray_inS21ser[4]}), .a ({ciphertext_s3[36], ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .c ({new_AGEMA_signal_5644, new_AGEMA_signal_5643, new_AGEMA_signal_5642, stateArray_S21reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S21reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, new_AGEMA_signal_3053, stateArray_inS21ser[5]}), .a ({ciphertext_s3[37], ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .c ({new_AGEMA_signal_5647, new_AGEMA_signal_5646, new_AGEMA_signal_5645, stateArray_S21reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S21reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_3064, new_AGEMA_signal_3063, new_AGEMA_signal_3062, stateArray_inS21ser[6]}), .a ({ciphertext_s3[38], ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .c ({new_AGEMA_signal_5650, new_AGEMA_signal_5649, new_AGEMA_signal_5648, stateArray_S21reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S21reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_3073, new_AGEMA_signal_3072, new_AGEMA_signal_3071, stateArray_inS21ser[7]}), .a ({ciphertext_s3[39], ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .c ({new_AGEMA_signal_5653, new_AGEMA_signal_5652, new_AGEMA_signal_5651, stateArray_S21reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S22reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3082, new_AGEMA_signal_3081, new_AGEMA_signal_3080, stateArray_inS22ser[0]}), .a ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_5656, new_AGEMA_signal_5655, new_AGEMA_signal_5654, stateArray_S22reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S22reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, new_AGEMA_signal_3089, stateArray_inS22ser[1]}), .a ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_5659, new_AGEMA_signal_5658, new_AGEMA_signal_5657, stateArray_S22reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S22reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3100, new_AGEMA_signal_3099, new_AGEMA_signal_3098, stateArray_inS22ser[2]}), .a ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_5662, new_AGEMA_signal_5661, new_AGEMA_signal_5660, stateArray_S22reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S22reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, new_AGEMA_signal_3107, stateArray_inS22ser[3]}), .a ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_5665, new_AGEMA_signal_5664, new_AGEMA_signal_5663, stateArray_S22reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S22reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3118, new_AGEMA_signal_3117, new_AGEMA_signal_3116, stateArray_inS22ser[4]}), .a ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_5668, new_AGEMA_signal_5667, new_AGEMA_signal_5666, stateArray_S22reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S22reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, new_AGEMA_signal_3125, stateArray_inS22ser[5]}), .a ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_5671, new_AGEMA_signal_5670, new_AGEMA_signal_5669, stateArray_S22reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S22reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3136, new_AGEMA_signal_3135, new_AGEMA_signal_3134, stateArray_inS22ser[6]}), .a ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .c ({new_AGEMA_signal_5674, new_AGEMA_signal_5673, new_AGEMA_signal_5672, stateArray_S22reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S22reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, new_AGEMA_signal_3143, stateArray_inS22ser[7]}), .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .c ({new_AGEMA_signal_5677, new_AGEMA_signal_5676, new_AGEMA_signal_5675, stateArray_S22reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S23reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_5272, new_AGEMA_signal_5271, new_AGEMA_signal_5270, stateArray_inS23ser[0]}), .a ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_5680, new_AGEMA_signal_5679, new_AGEMA_signal_5678, stateArray_S23reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S23reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_5278, new_AGEMA_signal_5277, new_AGEMA_signal_5276, stateArray_inS23ser[1]}), .a ({ciphertext_s3[49], ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_5683, new_AGEMA_signal_5682, new_AGEMA_signal_5681, stateArray_S23reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S23reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_5284, new_AGEMA_signal_5283, new_AGEMA_signal_5282, stateArray_inS23ser[2]}), .a ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_5686, new_AGEMA_signal_5685, new_AGEMA_signal_5684, stateArray_S23reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S23reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_5290, new_AGEMA_signal_5289, new_AGEMA_signal_5288, stateArray_inS23ser[3]}), .a ({ciphertext_s3[51], ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .c ({new_AGEMA_signal_5689, new_AGEMA_signal_5688, new_AGEMA_signal_5687, stateArray_S23reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S23reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_5296, new_AGEMA_signal_5295, new_AGEMA_signal_5294, stateArray_inS23ser[4]}), .a ({ciphertext_s3[52], ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .c ({new_AGEMA_signal_5692, new_AGEMA_signal_5691, new_AGEMA_signal_5690, stateArray_S23reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S23reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_5302, new_AGEMA_signal_5301, new_AGEMA_signal_5300, stateArray_inS23ser[5]}), .a ({ciphertext_s3[53], ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .c ({new_AGEMA_signal_5695, new_AGEMA_signal_5694, new_AGEMA_signal_5693, stateArray_S23reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S23reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_5308, new_AGEMA_signal_5307, new_AGEMA_signal_5306, stateArray_inS23ser[6]}), .a ({ciphertext_s3[54], ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .c ({new_AGEMA_signal_5698, new_AGEMA_signal_5697, new_AGEMA_signal_5696, stateArray_S23reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S23reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_5314, new_AGEMA_signal_5313, new_AGEMA_signal_5312, stateArray_inS23ser[7]}), .a ({ciphertext_s3[55], ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .c ({new_AGEMA_signal_5701, new_AGEMA_signal_5700, new_AGEMA_signal_5699, stateArray_S23reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S30reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_3154, new_AGEMA_signal_3153, new_AGEMA_signal_3152, stateArray_inS30ser[0]}), .a ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_5704, new_AGEMA_signal_5703, new_AGEMA_signal_5702, stateArray_S30reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S30reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, new_AGEMA_signal_3161, stateArray_inS30ser[1]}), .a ({ciphertext_s3[1], ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_5707, new_AGEMA_signal_5706, new_AGEMA_signal_5705, stateArray_S30reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S30reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_3172, new_AGEMA_signal_3171, new_AGEMA_signal_3170, stateArray_inS30ser[2]}), .a ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_5710, new_AGEMA_signal_5709, new_AGEMA_signal_5708, stateArray_S30reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S30reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, new_AGEMA_signal_3179, stateArray_inS30ser[3]}), .a ({ciphertext_s3[3], ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .c ({new_AGEMA_signal_5713, new_AGEMA_signal_5712, new_AGEMA_signal_5711, stateArray_S30reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S30reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_3190, new_AGEMA_signal_3189, new_AGEMA_signal_3188, stateArray_inS30ser[4]}), .a ({ciphertext_s3[4], ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .c ({new_AGEMA_signal_5716, new_AGEMA_signal_5715, new_AGEMA_signal_5714, stateArray_S30reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S30reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, new_AGEMA_signal_3197, stateArray_inS30ser[5]}), .a ({ciphertext_s3[5], ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .c ({new_AGEMA_signal_5719, new_AGEMA_signal_5718, new_AGEMA_signal_5717, stateArray_S30reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S30reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_3208, new_AGEMA_signal_3207, new_AGEMA_signal_3206, stateArray_inS30ser[6]}), .a ({ciphertext_s3[6], ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .c ({new_AGEMA_signal_5722, new_AGEMA_signal_5721, new_AGEMA_signal_5720, stateArray_S30reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S30reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, new_AGEMA_signal_3215, stateArray_inS30ser[7]}), .a ({ciphertext_s3[7], ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .c ({new_AGEMA_signal_5725, new_AGEMA_signal_5724, new_AGEMA_signal_5723, stateArray_S30reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S31reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_3226, new_AGEMA_signal_3225, new_AGEMA_signal_3224, stateArray_inS31ser[0]}), .a ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_5728, new_AGEMA_signal_5727, new_AGEMA_signal_5726, stateArray_S31reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S31reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, new_AGEMA_signal_3233, stateArray_inS31ser[1]}), .a ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_5731, new_AGEMA_signal_5730, new_AGEMA_signal_5729, stateArray_S31reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S31reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_3244, new_AGEMA_signal_3243, new_AGEMA_signal_3242, stateArray_inS31ser[2]}), .a ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5734, new_AGEMA_signal_5733, new_AGEMA_signal_5732, stateArray_S31reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S31reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, new_AGEMA_signal_3251, stateArray_inS31ser[3]}), .a ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_5737, new_AGEMA_signal_5736, new_AGEMA_signal_5735, stateArray_S31reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S31reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_3262, new_AGEMA_signal_3261, new_AGEMA_signal_3260, stateArray_inS31ser[4]}), .a ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_5740, new_AGEMA_signal_5739, new_AGEMA_signal_5738, stateArray_S31reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S31reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, new_AGEMA_signal_3269, stateArray_inS31ser[5]}), .a ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_5743, new_AGEMA_signal_5742, new_AGEMA_signal_5741, stateArray_S31reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S31reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_3280, new_AGEMA_signal_3279, new_AGEMA_signal_3278, stateArray_inS31ser[6]}), .a ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .c ({new_AGEMA_signal_5746, new_AGEMA_signal_5745, new_AGEMA_signal_5744, stateArray_S31reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S31reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, new_AGEMA_signal_3287, stateArray_inS31ser[7]}), .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .c ({new_AGEMA_signal_5749, new_AGEMA_signal_5748, new_AGEMA_signal_5747, stateArray_S31reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S32reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_3298, new_AGEMA_signal_3297, new_AGEMA_signal_3296, stateArray_inS32ser[0]}), .a ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_5752, new_AGEMA_signal_5751, new_AGEMA_signal_5750, stateArray_S32reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S32reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, new_AGEMA_signal_3305, stateArray_inS32ser[1]}), .a ({ciphertext_s3[17], ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_5755, new_AGEMA_signal_5754, new_AGEMA_signal_5753, stateArray_S32reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S32reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_3316, new_AGEMA_signal_3315, new_AGEMA_signal_3314, stateArray_inS32ser[2]}), .a ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_5758, new_AGEMA_signal_5757, new_AGEMA_signal_5756, stateArray_S32reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S32reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, new_AGEMA_signal_3323, stateArray_inS32ser[3]}), .a ({ciphertext_s3[19], ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .c ({new_AGEMA_signal_5761, new_AGEMA_signal_5760, new_AGEMA_signal_5759, stateArray_S32reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S32reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_3334, new_AGEMA_signal_3333, new_AGEMA_signal_3332, stateArray_inS32ser[4]}), .a ({ciphertext_s3[20], ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .c ({new_AGEMA_signal_5764, new_AGEMA_signal_5763, new_AGEMA_signal_5762, stateArray_S32reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S32reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, new_AGEMA_signal_3341, stateArray_inS32ser[5]}), .a ({ciphertext_s3[21], ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .c ({new_AGEMA_signal_5767, new_AGEMA_signal_5766, new_AGEMA_signal_5765, stateArray_S32reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S32reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_3352, new_AGEMA_signal_3351, new_AGEMA_signal_3350, stateArray_inS32ser[6]}), .a ({ciphertext_s3[22], ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .c ({new_AGEMA_signal_5770, new_AGEMA_signal_5769, new_AGEMA_signal_5768, stateArray_S32reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S32reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, new_AGEMA_signal_3359, stateArray_inS32ser[7]}), .a ({ciphertext_s3[23], ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .c ({new_AGEMA_signal_5773, new_AGEMA_signal_5772, new_AGEMA_signal_5771, stateArray_S32reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS00ser_mux_inst_0_U1 ( .s (stateArray_n32), .b ({plaintext_s3[120], plaintext_s2[120], plaintext_s1[120], plaintext_s0[120]}), .a ({ciphertext_s3[112], ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_2506, new_AGEMA_signal_2505, new_AGEMA_signal_2504, stateArray_inS00ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS00ser_mux_inst_1_U1 ( .s (stateArray_n32), .b ({plaintext_s3[121], plaintext_s2[121], plaintext_s1[121], plaintext_s0[121]}), .a ({ciphertext_s3[113], ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, new_AGEMA_signal_2513, stateArray_inS00ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS00ser_mux_inst_2_U1 ( .s (stateArray_n32), .b ({plaintext_s3[122], plaintext_s2[122], plaintext_s1[122], plaintext_s0[122]}), .a ({ciphertext_s3[114], ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_2524, new_AGEMA_signal_2523, new_AGEMA_signal_2522, stateArray_inS00ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS00ser_mux_inst_3_U1 ( .s (stateArray_n32), .b ({plaintext_s3[123], plaintext_s2[123], plaintext_s1[123], plaintext_s0[123]}), .a ({ciphertext_s3[115], ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}), .c ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, new_AGEMA_signal_2531, stateArray_inS00ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS00ser_mux_inst_4_U1 ( .s (stateArray_n32), .b ({plaintext_s3[124], plaintext_s2[124], plaintext_s1[124], plaintext_s0[124]}), .a ({ciphertext_s3[116], ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .c ({new_AGEMA_signal_2542, new_AGEMA_signal_2541, new_AGEMA_signal_2540, stateArray_inS00ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS00ser_mux_inst_5_U1 ( .s (stateArray_n32), .b ({plaintext_s3[125], plaintext_s2[125], plaintext_s1[125], plaintext_s0[125]}), .a ({ciphertext_s3[117], ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}), .c ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, new_AGEMA_signal_2549, stateArray_inS00ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS00ser_mux_inst_6_U1 ( .s (stateArray_n32), .b ({plaintext_s3[126], plaintext_s2[126], plaintext_s1[126], plaintext_s0[126]}), .a ({ciphertext_s3[118], ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}), .c ({new_AGEMA_signal_2560, new_AGEMA_signal_2559, new_AGEMA_signal_2558, stateArray_inS00ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS00ser_mux_inst_7_U1 ( .s (stateArray_n32), .b ({plaintext_s3[127], plaintext_s2[127], plaintext_s1[127], plaintext_s0[127]}), .a ({ciphertext_s3[119], ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .c ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, new_AGEMA_signal_2567, stateArray_inS00ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS01ser_mux_inst_0_U1 ( .s (stateArray_n32), .b ({plaintext_s3[112], plaintext_s2[112], plaintext_s1[112], plaintext_s0[112]}), .a ({ciphertext_s3[104], ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_2578, new_AGEMA_signal_2577, new_AGEMA_signal_2576, stateArray_inS01ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS01ser_mux_inst_1_U1 ( .s (stateArray_n32), .b ({plaintext_s3[113], plaintext_s2[113], plaintext_s1[113], plaintext_s0[113]}), .a ({ciphertext_s3[105], ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, new_AGEMA_signal_2585, stateArray_inS01ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS01ser_mux_inst_2_U1 ( .s (stateArray_n32), .b ({plaintext_s3[114], plaintext_s2[114], plaintext_s1[114], plaintext_s0[114]}), .a ({ciphertext_s3[106], ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_2596, new_AGEMA_signal_2595, new_AGEMA_signal_2594, stateArray_inS01ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS01ser_mux_inst_3_U1 ( .s (stateArray_n32), .b ({plaintext_s3[115], plaintext_s2[115], plaintext_s1[115], plaintext_s0[115]}), .a ({ciphertext_s3[107], ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}), .c ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, new_AGEMA_signal_2603, stateArray_inS01ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS01ser_mux_inst_4_U1 ( .s (stateArray_n32), .b ({plaintext_s3[116], plaintext_s2[116], plaintext_s1[116], plaintext_s0[116]}), .a ({ciphertext_s3[108], ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .c ({new_AGEMA_signal_2614, new_AGEMA_signal_2613, new_AGEMA_signal_2612, stateArray_inS01ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS01ser_mux_inst_5_U1 ( .s (stateArray_n32), .b ({plaintext_s3[117], plaintext_s2[117], plaintext_s1[117], plaintext_s0[117]}), .a ({ciphertext_s3[109], ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}), .c ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, new_AGEMA_signal_2621, stateArray_inS01ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS01ser_mux_inst_6_U1 ( .s (stateArray_n32), .b ({plaintext_s3[118], plaintext_s2[118], plaintext_s1[118], plaintext_s0[118]}), .a ({ciphertext_s3[110], ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}), .c ({new_AGEMA_signal_2632, new_AGEMA_signal_2631, new_AGEMA_signal_2630, stateArray_inS01ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS01ser_mux_inst_7_U1 ( .s (stateArray_n32), .b ({plaintext_s3[119], plaintext_s2[119], plaintext_s1[119], plaintext_s0[119]}), .a ({ciphertext_s3[111], ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .c ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, new_AGEMA_signal_2639, stateArray_inS01ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS02ser_mux_inst_0_U1 ( .s (stateArray_n31), .b ({plaintext_s3[104], plaintext_s2[104], plaintext_s1[104], plaintext_s0[104]}), .a ({ciphertext_s3[96], ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_2650, new_AGEMA_signal_2649, new_AGEMA_signal_2648, stateArray_inS02ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS02ser_mux_inst_1_U1 ( .s (stateArray_n31), .b ({plaintext_s3[105], plaintext_s2[105], plaintext_s1[105], plaintext_s0[105]}), .a ({ciphertext_s3[97], ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, new_AGEMA_signal_2657, stateArray_inS02ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS02ser_mux_inst_2_U1 ( .s (stateArray_n31), .b ({plaintext_s3[106], plaintext_s2[106], plaintext_s1[106], plaintext_s0[106]}), .a ({ciphertext_s3[98], ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_2668, new_AGEMA_signal_2667, new_AGEMA_signal_2666, stateArray_inS02ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS02ser_mux_inst_3_U1 ( .s (stateArray_n31), .b ({plaintext_s3[107], plaintext_s2[107], plaintext_s1[107], plaintext_s0[107]}), .a ({ciphertext_s3[99], ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}), .c ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, new_AGEMA_signal_2675, stateArray_inS02ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS02ser_mux_inst_4_U1 ( .s (stateArray_n31), .b ({plaintext_s3[108], plaintext_s2[108], plaintext_s1[108], plaintext_s0[108]}), .a ({ciphertext_s3[100], ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .c ({new_AGEMA_signal_2686, new_AGEMA_signal_2685, new_AGEMA_signal_2684, stateArray_inS02ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS02ser_mux_inst_5_U1 ( .s (stateArray_n31), .b ({plaintext_s3[109], plaintext_s2[109], plaintext_s1[109], plaintext_s0[109]}), .a ({ciphertext_s3[101], ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}), .c ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, new_AGEMA_signal_2693, stateArray_inS02ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS02ser_mux_inst_6_U1 ( .s (stateArray_n31), .b ({plaintext_s3[110], plaintext_s2[110], plaintext_s1[110], plaintext_s0[110]}), .a ({ciphertext_s3[102], ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}), .c ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, new_AGEMA_signal_2702, stateArray_inS02ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS02ser_mux_inst_7_U1 ( .s (stateArray_n31), .b ({plaintext_s3[111], plaintext_s2[111], plaintext_s1[111], plaintext_s0[111]}), .a ({ciphertext_s3[103], ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .c ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, new_AGEMA_signal_2711, stateArray_inS02ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS10_MC_mux_inst_0_U1 ( .s (stateArray_n23), .b ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .a ({new_AGEMA_signal_4678, new_AGEMA_signal_4677, new_AGEMA_signal_4676, StateInMC[24]}), .c ({new_AGEMA_signal_5062, new_AGEMA_signal_5061, new_AGEMA_signal_5060, stateArray_outS10ser_MC[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS10_MC_mux_inst_1_U1 ( .s (stateArray_n23), .b ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .a ({new_AGEMA_signal_4681, new_AGEMA_signal_4680, new_AGEMA_signal_4679, StateInMC[25]}), .c ({new_AGEMA_signal_5065, new_AGEMA_signal_5064, new_AGEMA_signal_5063, stateArray_outS10ser_MC[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS10_MC_mux_inst_2_U1 ( .s (stateArray_n23), .b ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .a ({new_AGEMA_signal_4684, new_AGEMA_signal_4683, new_AGEMA_signal_4682, StateInMC[26]}), .c ({new_AGEMA_signal_5068, new_AGEMA_signal_5067, new_AGEMA_signal_5066, stateArray_outS10ser_MC[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS10_MC_mux_inst_3_U1 ( .s (stateArray_n23), .b ({ciphertext_s3[91], ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}), .a ({new_AGEMA_signal_4687, new_AGEMA_signal_4686, new_AGEMA_signal_4685, StateInMC[27]}), .c ({new_AGEMA_signal_5071, new_AGEMA_signal_5070, new_AGEMA_signal_5069, stateArray_outS10ser_MC[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS10_MC_mux_inst_4_U1 ( .s (stateArray_n23), .b ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .a ({new_AGEMA_signal_4690, new_AGEMA_signal_4689, new_AGEMA_signal_4688, StateInMC[28]}), .c ({new_AGEMA_signal_5074, new_AGEMA_signal_5073, new_AGEMA_signal_5072, stateArray_outS10ser_MC[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS10_MC_mux_inst_5_U1 ( .s (stateArray_n23), .b ({ciphertext_s3[93], ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .a ({new_AGEMA_signal_4693, new_AGEMA_signal_4692, new_AGEMA_signal_4691, StateInMC[29]}), .c ({new_AGEMA_signal_5077, new_AGEMA_signal_5076, new_AGEMA_signal_5075, stateArray_outS10ser_MC[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS10_MC_mux_inst_6_U1 ( .s (stateArray_n23), .b ({ciphertext_s3[94], ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .a ({new_AGEMA_signal_4696, new_AGEMA_signal_4695, new_AGEMA_signal_4694, StateInMC[30]}), .c ({new_AGEMA_signal_5080, new_AGEMA_signal_5079, new_AGEMA_signal_5078, stateArray_outS10ser_MC[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS10_MC_mux_inst_7_U1 ( .s (stateArray_n23), .b ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .a ({new_AGEMA_signal_4699, new_AGEMA_signal_4698, new_AGEMA_signal_4697, StateInMC[31]}), .c ({new_AGEMA_signal_5083, new_AGEMA_signal_5082, new_AGEMA_signal_5081, stateArray_outS10ser_MC[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS03ser_mux_inst_0_U1 ( .s (stateArray_n31), .b ({plaintext_s3[96], plaintext_s2[96], plaintext_s1[96], plaintext_s0[96]}), .a ({new_AGEMA_signal_5062, new_AGEMA_signal_5061, new_AGEMA_signal_5060, stateArray_outS10ser_MC[0]}), .c ({new_AGEMA_signal_5176, new_AGEMA_signal_5175, new_AGEMA_signal_5174, stateArray_inS03ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS03ser_mux_inst_1_U1 ( .s (stateArray_n31), .b ({plaintext_s3[97], plaintext_s2[97], plaintext_s1[97], plaintext_s0[97]}), .a ({new_AGEMA_signal_5065, new_AGEMA_signal_5064, new_AGEMA_signal_5063, stateArray_outS10ser_MC[1]}), .c ({new_AGEMA_signal_5182, new_AGEMA_signal_5181, new_AGEMA_signal_5180, stateArray_inS03ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS03ser_mux_inst_2_U1 ( .s (stateArray_n31), .b ({plaintext_s3[98], plaintext_s2[98], plaintext_s1[98], plaintext_s0[98]}), .a ({new_AGEMA_signal_5068, new_AGEMA_signal_5067, new_AGEMA_signal_5066, stateArray_outS10ser_MC[2]}), .c ({new_AGEMA_signal_5188, new_AGEMA_signal_5187, new_AGEMA_signal_5186, stateArray_inS03ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS03ser_mux_inst_3_U1 ( .s (stateArray_n31), .b ({plaintext_s3[99], plaintext_s2[99], plaintext_s1[99], plaintext_s0[99]}), .a ({new_AGEMA_signal_5071, new_AGEMA_signal_5070, new_AGEMA_signal_5069, stateArray_outS10ser_MC[3]}), .c ({new_AGEMA_signal_5194, new_AGEMA_signal_5193, new_AGEMA_signal_5192, stateArray_inS03ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS03ser_mux_inst_4_U1 ( .s (stateArray_n31), .b ({plaintext_s3[100], plaintext_s2[100], plaintext_s1[100], plaintext_s0[100]}), .a ({new_AGEMA_signal_5074, new_AGEMA_signal_5073, new_AGEMA_signal_5072, stateArray_outS10ser_MC[4]}), .c ({new_AGEMA_signal_5200, new_AGEMA_signal_5199, new_AGEMA_signal_5198, stateArray_inS03ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS03ser_mux_inst_5_U1 ( .s (stateArray_n31), .b ({plaintext_s3[101], plaintext_s2[101], plaintext_s1[101], plaintext_s0[101]}), .a ({new_AGEMA_signal_5077, new_AGEMA_signal_5076, new_AGEMA_signal_5075, stateArray_outS10ser_MC[5]}), .c ({new_AGEMA_signal_5206, new_AGEMA_signal_5205, new_AGEMA_signal_5204, stateArray_inS03ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS03ser_mux_inst_6_U1 ( .s (stateArray_n31), .b ({plaintext_s3[102], plaintext_s2[102], plaintext_s1[102], plaintext_s0[102]}), .a ({new_AGEMA_signal_5080, new_AGEMA_signal_5079, new_AGEMA_signal_5078, stateArray_outS10ser_MC[6]}), .c ({new_AGEMA_signal_5212, new_AGEMA_signal_5211, new_AGEMA_signal_5210, stateArray_inS03ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS03ser_mux_inst_7_U1 ( .s (stateArray_n31), .b ({plaintext_s3[103], plaintext_s2[103], plaintext_s1[103], plaintext_s0[103]}), .a ({new_AGEMA_signal_5083, new_AGEMA_signal_5082, new_AGEMA_signal_5081, stateArray_outS10ser_MC[7]}), .c ({new_AGEMA_signal_5218, new_AGEMA_signal_5217, new_AGEMA_signal_5216, stateArray_inS03ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS10ser_mux_inst_0_U1 ( .s (stateArray_n30), .b ({plaintext_s3[88], plaintext_s2[88], plaintext_s1[88], plaintext_s0[88]}), .a ({ciphertext_s3[80], ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_2722, new_AGEMA_signal_2721, new_AGEMA_signal_2720, stateArray_inS10ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS10ser_mux_inst_1_U1 ( .s (stateArray_n30), .b ({plaintext_s3[89], plaintext_s2[89], plaintext_s1[89], plaintext_s0[89]}), .a ({ciphertext_s3[81], ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, new_AGEMA_signal_2729, stateArray_inS10ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS10ser_mux_inst_2_U1 ( .s (stateArray_n30), .b ({plaintext_s3[90], plaintext_s2[90], plaintext_s1[90], plaintext_s0[90]}), .a ({ciphertext_s3[82], ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_2740, new_AGEMA_signal_2739, new_AGEMA_signal_2738, stateArray_inS10ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS10ser_mux_inst_3_U1 ( .s (stateArray_n30), .b ({plaintext_s3[91], plaintext_s2[91], plaintext_s1[91], plaintext_s0[91]}), .a ({ciphertext_s3[83], ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}), .c ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, new_AGEMA_signal_2747, stateArray_inS10ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS10ser_mux_inst_4_U1 ( .s (stateArray_n30), .b ({plaintext_s3[92], plaintext_s2[92], plaintext_s1[92], plaintext_s0[92]}), .a ({ciphertext_s3[84], ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .c ({new_AGEMA_signal_2758, new_AGEMA_signal_2757, new_AGEMA_signal_2756, stateArray_inS10ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS10ser_mux_inst_5_U1 ( .s (stateArray_n30), .b ({plaintext_s3[93], plaintext_s2[93], plaintext_s1[93], plaintext_s0[93]}), .a ({ciphertext_s3[85], ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}), .c ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, new_AGEMA_signal_2765, stateArray_inS10ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS10ser_mux_inst_6_U1 ( .s (stateArray_n30), .b ({plaintext_s3[94], plaintext_s2[94], plaintext_s1[94], plaintext_s0[94]}), .a ({ciphertext_s3[86], ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}), .c ({new_AGEMA_signal_2776, new_AGEMA_signal_2775, new_AGEMA_signal_2774, stateArray_inS10ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS10ser_mux_inst_7_U1 ( .s (stateArray_n30), .b ({plaintext_s3[95], plaintext_s2[95], plaintext_s1[95], plaintext_s0[95]}), .a ({ciphertext_s3[87], ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .c ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, new_AGEMA_signal_2783, stateArray_inS10ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS11ser_mux_inst_0_U1 ( .s (stateArray_n30), .b ({plaintext_s3[80], plaintext_s2[80], plaintext_s1[80], plaintext_s0[80]}), .a ({ciphertext_s3[72], ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_2794, new_AGEMA_signal_2793, new_AGEMA_signal_2792, stateArray_inS11ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS11ser_mux_inst_1_U1 ( .s (stateArray_n30), .b ({plaintext_s3[81], plaintext_s2[81], plaintext_s1[81], plaintext_s0[81]}), .a ({ciphertext_s3[73], ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, new_AGEMA_signal_2801, stateArray_inS11ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS11ser_mux_inst_2_U1 ( .s (stateArray_n30), .b ({plaintext_s3[82], plaintext_s2[82], plaintext_s1[82], plaintext_s0[82]}), .a ({ciphertext_s3[74], ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_2812, new_AGEMA_signal_2811, new_AGEMA_signal_2810, stateArray_inS11ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS11ser_mux_inst_3_U1 ( .s (stateArray_n30), .b ({plaintext_s3[83], plaintext_s2[83], plaintext_s1[83], plaintext_s0[83]}), .a ({ciphertext_s3[75], ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}), .c ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, new_AGEMA_signal_2819, stateArray_inS11ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS11ser_mux_inst_4_U1 ( .s (stateArray_n30), .b ({plaintext_s3[84], plaintext_s2[84], plaintext_s1[84], plaintext_s0[84]}), .a ({ciphertext_s3[76], ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .c ({new_AGEMA_signal_2830, new_AGEMA_signal_2829, new_AGEMA_signal_2828, stateArray_inS11ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS11ser_mux_inst_5_U1 ( .s (stateArray_n30), .b ({plaintext_s3[85], plaintext_s2[85], plaintext_s1[85], plaintext_s0[85]}), .a ({ciphertext_s3[77], ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}), .c ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, new_AGEMA_signal_2837, stateArray_inS11ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS11ser_mux_inst_6_U1 ( .s (stateArray_n30), .b ({plaintext_s3[86], plaintext_s2[86], plaintext_s1[86], plaintext_s0[86]}), .a ({ciphertext_s3[78], ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}), .c ({new_AGEMA_signal_2848, new_AGEMA_signal_2847, new_AGEMA_signal_2846, stateArray_inS11ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS11ser_mux_inst_7_U1 ( .s (stateArray_n30), .b ({plaintext_s3[87], plaintext_s2[87], plaintext_s1[87], plaintext_s0[87]}), .a ({ciphertext_s3[79], ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .c ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, new_AGEMA_signal_2855, stateArray_inS11ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS12ser_mux_inst_0_U1 ( .s (stateArray_n29), .b ({plaintext_s3[72], plaintext_s2[72], plaintext_s1[72], plaintext_s0[72]}), .a ({ciphertext_s3[64], ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_2866, new_AGEMA_signal_2865, new_AGEMA_signal_2864, stateArray_inS12ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS12ser_mux_inst_1_U1 ( .s (stateArray_n29), .b ({plaintext_s3[73], plaintext_s2[73], plaintext_s1[73], plaintext_s0[73]}), .a ({ciphertext_s3[65], ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, new_AGEMA_signal_2873, stateArray_inS12ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS12ser_mux_inst_2_U1 ( .s (stateArray_n29), .b ({plaintext_s3[74], plaintext_s2[74], plaintext_s1[74], plaintext_s0[74]}), .a ({ciphertext_s3[66], ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_2884, new_AGEMA_signal_2883, new_AGEMA_signal_2882, stateArray_inS12ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS12ser_mux_inst_3_U1 ( .s (stateArray_n29), .b ({plaintext_s3[75], plaintext_s2[75], plaintext_s1[75], plaintext_s0[75]}), .a ({ciphertext_s3[67], ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}), .c ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, new_AGEMA_signal_2891, stateArray_inS12ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS12ser_mux_inst_4_U1 ( .s (stateArray_n29), .b ({plaintext_s3[76], plaintext_s2[76], plaintext_s1[76], plaintext_s0[76]}), .a ({ciphertext_s3[68], ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .c ({new_AGEMA_signal_2902, new_AGEMA_signal_2901, new_AGEMA_signal_2900, stateArray_inS12ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS12ser_mux_inst_5_U1 ( .s (stateArray_n29), .b ({plaintext_s3[77], plaintext_s2[77], plaintext_s1[77], plaintext_s0[77]}), .a ({ciphertext_s3[69], ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}), .c ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, new_AGEMA_signal_2909, stateArray_inS12ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS12ser_mux_inst_6_U1 ( .s (stateArray_n29), .b ({plaintext_s3[78], plaintext_s2[78], plaintext_s1[78], plaintext_s0[78]}), .a ({ciphertext_s3[70], ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}), .c ({new_AGEMA_signal_2920, new_AGEMA_signal_2919, new_AGEMA_signal_2918, stateArray_inS12ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS12ser_mux_inst_7_U1 ( .s (stateArray_n29), .b ({plaintext_s3[79], plaintext_s2[79], plaintext_s1[79], plaintext_s0[79]}), .a ({ciphertext_s3[71], ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .c ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, new_AGEMA_signal_2927, stateArray_inS12ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS20_MC_mux_inst_0_U1 ( .s (stateArray_n23), .b ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .a ({new_AGEMA_signal_4654, new_AGEMA_signal_4653, new_AGEMA_signal_4652, StateInMC[16]}), .c ({new_AGEMA_signal_5086, new_AGEMA_signal_5085, new_AGEMA_signal_5084, stateArray_outS20ser_MC[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS20_MC_mux_inst_1_U1 ( .s (stateArray_n23), .b ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .a ({new_AGEMA_signal_4657, new_AGEMA_signal_4656, new_AGEMA_signal_4655, StateInMC[17]}), .c ({new_AGEMA_signal_5089, new_AGEMA_signal_5088, new_AGEMA_signal_5087, stateArray_outS20ser_MC[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS20_MC_mux_inst_2_U1 ( .s (stateArray_n23), .b ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .a ({new_AGEMA_signal_4660, new_AGEMA_signal_4659, new_AGEMA_signal_4658, StateInMC[18]}), .c ({new_AGEMA_signal_5092, new_AGEMA_signal_5091, new_AGEMA_signal_5090, stateArray_outS20ser_MC[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS20_MC_mux_inst_3_U1 ( .s (stateArray_n23), .b ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .a ({new_AGEMA_signal_4663, new_AGEMA_signal_4662, new_AGEMA_signal_4661, StateInMC[19]}), .c ({new_AGEMA_signal_5095, new_AGEMA_signal_5094, new_AGEMA_signal_5093, stateArray_outS20ser_MC[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS20_MC_mux_inst_4_U1 ( .s (stateArray_n23), .b ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .a ({new_AGEMA_signal_4666, new_AGEMA_signal_4665, new_AGEMA_signal_4664, StateInMC[20]}), .c ({new_AGEMA_signal_5098, new_AGEMA_signal_5097, new_AGEMA_signal_5096, stateArray_outS20ser_MC[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS20_MC_mux_inst_5_U1 ( .s (stateArray_n23), .b ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .a ({new_AGEMA_signal_4669, new_AGEMA_signal_4668, new_AGEMA_signal_4667, StateInMC[21]}), .c ({new_AGEMA_signal_5101, new_AGEMA_signal_5100, new_AGEMA_signal_5099, stateArray_outS20ser_MC[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS20_MC_mux_inst_6_U1 ( .s (stateArray_n23), .b ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .a ({new_AGEMA_signal_4672, new_AGEMA_signal_4671, new_AGEMA_signal_4670, StateInMC[22]}), .c ({new_AGEMA_signal_5104, new_AGEMA_signal_5103, new_AGEMA_signal_5102, stateArray_outS20ser_MC[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS20_MC_mux_inst_7_U1 ( .s (stateArray_n23), .b ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .a ({new_AGEMA_signal_4675, new_AGEMA_signal_4674, new_AGEMA_signal_4673, StateInMC[23]}), .c ({new_AGEMA_signal_5107, new_AGEMA_signal_5106, new_AGEMA_signal_5105, stateArray_outS20ser_MC[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS13ser_mux_inst_0_U1 ( .s (stateArray_n29), .b ({plaintext_s3[64], plaintext_s2[64], plaintext_s1[64], plaintext_s0[64]}), .a ({new_AGEMA_signal_5086, new_AGEMA_signal_5085, new_AGEMA_signal_5084, stateArray_outS20ser_MC[0]}), .c ({new_AGEMA_signal_5224, new_AGEMA_signal_5223, new_AGEMA_signal_5222, stateArray_inS13ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS13ser_mux_inst_1_U1 ( .s (stateArray_n29), .b ({plaintext_s3[65], plaintext_s2[65], plaintext_s1[65], plaintext_s0[65]}), .a ({new_AGEMA_signal_5089, new_AGEMA_signal_5088, new_AGEMA_signal_5087, stateArray_outS20ser_MC[1]}), .c ({new_AGEMA_signal_5230, new_AGEMA_signal_5229, new_AGEMA_signal_5228, stateArray_inS13ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS13ser_mux_inst_2_U1 ( .s (stateArray_n29), .b ({plaintext_s3[66], plaintext_s2[66], plaintext_s1[66], plaintext_s0[66]}), .a ({new_AGEMA_signal_5092, new_AGEMA_signal_5091, new_AGEMA_signal_5090, stateArray_outS20ser_MC[2]}), .c ({new_AGEMA_signal_5236, new_AGEMA_signal_5235, new_AGEMA_signal_5234, stateArray_inS13ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS13ser_mux_inst_3_U1 ( .s (stateArray_n29), .b ({plaintext_s3[67], plaintext_s2[67], plaintext_s1[67], plaintext_s0[67]}), .a ({new_AGEMA_signal_5095, new_AGEMA_signal_5094, new_AGEMA_signal_5093, stateArray_outS20ser_MC[3]}), .c ({new_AGEMA_signal_5242, new_AGEMA_signal_5241, new_AGEMA_signal_5240, stateArray_inS13ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS13ser_mux_inst_4_U1 ( .s (stateArray_n29), .b ({plaintext_s3[68], plaintext_s2[68], plaintext_s1[68], plaintext_s0[68]}), .a ({new_AGEMA_signal_5098, new_AGEMA_signal_5097, new_AGEMA_signal_5096, stateArray_outS20ser_MC[4]}), .c ({new_AGEMA_signal_5248, new_AGEMA_signal_5247, new_AGEMA_signal_5246, stateArray_inS13ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS13ser_mux_inst_5_U1 ( .s (stateArray_n29), .b ({plaintext_s3[69], plaintext_s2[69], plaintext_s1[69], plaintext_s0[69]}), .a ({new_AGEMA_signal_5101, new_AGEMA_signal_5100, new_AGEMA_signal_5099, stateArray_outS20ser_MC[5]}), .c ({new_AGEMA_signal_5254, new_AGEMA_signal_5253, new_AGEMA_signal_5252, stateArray_inS13ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS13ser_mux_inst_6_U1 ( .s (stateArray_n29), .b ({plaintext_s3[70], plaintext_s2[70], plaintext_s1[70], plaintext_s0[70]}), .a ({new_AGEMA_signal_5104, new_AGEMA_signal_5103, new_AGEMA_signal_5102, stateArray_outS20ser_MC[6]}), .c ({new_AGEMA_signal_5260, new_AGEMA_signal_5259, new_AGEMA_signal_5258, stateArray_inS13ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS13ser_mux_inst_7_U1 ( .s (stateArray_n29), .b ({plaintext_s3[71], plaintext_s2[71], plaintext_s1[71], plaintext_s0[71]}), .a ({new_AGEMA_signal_5107, new_AGEMA_signal_5106, new_AGEMA_signal_5105, stateArray_outS20ser_MC[7]}), .c ({new_AGEMA_signal_5266, new_AGEMA_signal_5265, new_AGEMA_signal_5264, stateArray_inS13ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS20ser_mux_inst_0_U1 ( .s (stateArray_n28), .b ({plaintext_s3[56], plaintext_s2[56], plaintext_s1[56], plaintext_s0[56]}), .a ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_2938, new_AGEMA_signal_2937, new_AGEMA_signal_2936, stateArray_inS20ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS20ser_mux_inst_1_U1 ( .s (stateArray_n28), .b ({plaintext_s3[57], plaintext_s2[57], plaintext_s1[57], plaintext_s0[57]}), .a ({ciphertext_s3[49], ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, new_AGEMA_signal_2945, stateArray_inS20ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS20ser_mux_inst_2_U1 ( .s (stateArray_n28), .b ({plaintext_s3[58], plaintext_s2[58], plaintext_s1[58], plaintext_s0[58]}), .a ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_2956, new_AGEMA_signal_2955, new_AGEMA_signal_2954, stateArray_inS20ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS20ser_mux_inst_3_U1 ( .s (stateArray_n28), .b ({plaintext_s3[59], plaintext_s2[59], plaintext_s1[59], plaintext_s0[59]}), .a ({ciphertext_s3[51], ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .c ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, new_AGEMA_signal_2963, stateArray_inS20ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS20ser_mux_inst_4_U1 ( .s (stateArray_n28), .b ({plaintext_s3[60], plaintext_s2[60], plaintext_s1[60], plaintext_s0[60]}), .a ({ciphertext_s3[52], ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .c ({new_AGEMA_signal_2974, new_AGEMA_signal_2973, new_AGEMA_signal_2972, stateArray_inS20ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS20ser_mux_inst_5_U1 ( .s (stateArray_n28), .b ({plaintext_s3[61], plaintext_s2[61], plaintext_s1[61], plaintext_s0[61]}), .a ({ciphertext_s3[53], ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .c ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, new_AGEMA_signal_2981, stateArray_inS20ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS20ser_mux_inst_6_U1 ( .s (stateArray_n28), .b ({plaintext_s3[62], plaintext_s2[62], plaintext_s1[62], plaintext_s0[62]}), .a ({ciphertext_s3[54], ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .c ({new_AGEMA_signal_2992, new_AGEMA_signal_2991, new_AGEMA_signal_2990, stateArray_inS20ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS20ser_mux_inst_7_U1 ( .s (stateArray_n28), .b ({plaintext_s3[63], plaintext_s2[63], plaintext_s1[63], plaintext_s0[63]}), .a ({ciphertext_s3[55], ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .c ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, new_AGEMA_signal_2999, stateArray_inS20ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS21ser_mux_inst_0_U1 ( .s (stateArray_n28), .b ({plaintext_s3[48], plaintext_s2[48], plaintext_s1[48], plaintext_s0[48]}), .a ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_3010, new_AGEMA_signal_3009, new_AGEMA_signal_3008, stateArray_inS21ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS21ser_mux_inst_1_U1 ( .s (stateArray_n28), .b ({plaintext_s3[49], plaintext_s2[49], plaintext_s1[49], plaintext_s0[49]}), .a ({ciphertext_s3[41], ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, new_AGEMA_signal_3017, stateArray_inS21ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS21ser_mux_inst_2_U1 ( .s (stateArray_n28), .b ({plaintext_s3[50], plaintext_s2[50], plaintext_s1[50], plaintext_s0[50]}), .a ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_3028, new_AGEMA_signal_3027, new_AGEMA_signal_3026, stateArray_inS21ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS21ser_mux_inst_3_U1 ( .s (stateArray_n28), .b ({plaintext_s3[51], plaintext_s2[51], plaintext_s1[51], plaintext_s0[51]}), .a ({ciphertext_s3[43], ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .c ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, new_AGEMA_signal_3035, stateArray_inS21ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS21ser_mux_inst_4_U1 ( .s (stateArray_n28), .b ({plaintext_s3[52], plaintext_s2[52], plaintext_s1[52], plaintext_s0[52]}), .a ({ciphertext_s3[44], ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .c ({new_AGEMA_signal_3046, new_AGEMA_signal_3045, new_AGEMA_signal_3044, stateArray_inS21ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS21ser_mux_inst_5_U1 ( .s (stateArray_n28), .b ({plaintext_s3[53], plaintext_s2[53], plaintext_s1[53], plaintext_s0[53]}), .a ({ciphertext_s3[45], ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .c ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, new_AGEMA_signal_3053, stateArray_inS21ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS21ser_mux_inst_6_U1 ( .s (stateArray_n28), .b ({plaintext_s3[54], plaintext_s2[54], plaintext_s1[54], plaintext_s0[54]}), .a ({ciphertext_s3[46], ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .c ({new_AGEMA_signal_3064, new_AGEMA_signal_3063, new_AGEMA_signal_3062, stateArray_inS21ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS21ser_mux_inst_7_U1 ( .s (stateArray_n28), .b ({plaintext_s3[55], plaintext_s2[55], plaintext_s1[55], plaintext_s0[55]}), .a ({ciphertext_s3[47], ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .c ({new_AGEMA_signal_3073, new_AGEMA_signal_3072, new_AGEMA_signal_3071, stateArray_inS21ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS22ser_mux_inst_0_U1 ( .s (stateArray_n27), .b ({plaintext_s3[40], plaintext_s2[40], plaintext_s1[40], plaintext_s0[40]}), .a ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_3082, new_AGEMA_signal_3081, new_AGEMA_signal_3080, stateArray_inS22ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS22ser_mux_inst_1_U1 ( .s (stateArray_n27), .b ({plaintext_s3[41], plaintext_s2[41], plaintext_s1[41], plaintext_s0[41]}), .a ({ciphertext_s3[33], ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, new_AGEMA_signal_3089, stateArray_inS22ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS22ser_mux_inst_2_U1 ( .s (stateArray_n27), .b ({plaintext_s3[42], plaintext_s2[42], plaintext_s1[42], plaintext_s0[42]}), .a ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_3100, new_AGEMA_signal_3099, new_AGEMA_signal_3098, stateArray_inS22ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS22ser_mux_inst_3_U1 ( .s (stateArray_n27), .b ({plaintext_s3[43], plaintext_s2[43], plaintext_s1[43], plaintext_s0[43]}), .a ({ciphertext_s3[35], ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .c ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, new_AGEMA_signal_3107, stateArray_inS22ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS22ser_mux_inst_4_U1 ( .s (stateArray_n27), .b ({plaintext_s3[44], plaintext_s2[44], plaintext_s1[44], plaintext_s0[44]}), .a ({ciphertext_s3[36], ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .c ({new_AGEMA_signal_3118, new_AGEMA_signal_3117, new_AGEMA_signal_3116, stateArray_inS22ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS22ser_mux_inst_5_U1 ( .s (stateArray_n27), .b ({plaintext_s3[45], plaintext_s2[45], plaintext_s1[45], plaintext_s0[45]}), .a ({ciphertext_s3[37], ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .c ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, new_AGEMA_signal_3125, stateArray_inS22ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS22ser_mux_inst_6_U1 ( .s (stateArray_n27), .b ({plaintext_s3[46], plaintext_s2[46], plaintext_s1[46], plaintext_s0[46]}), .a ({ciphertext_s3[38], ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .c ({new_AGEMA_signal_3136, new_AGEMA_signal_3135, new_AGEMA_signal_3134, stateArray_inS22ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS22ser_mux_inst_7_U1 ( .s (stateArray_n27), .b ({plaintext_s3[47], plaintext_s2[47], plaintext_s1[47], plaintext_s0[47]}), .a ({ciphertext_s3[39], ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .c ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, new_AGEMA_signal_3143, stateArray_inS22ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS30_MC_mux_inst_0_U1 ( .s (stateArray_n22), .b ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .a ({new_AGEMA_signal_4630, new_AGEMA_signal_4629, new_AGEMA_signal_4628, StateInMC[8]}), .c ({new_AGEMA_signal_5110, new_AGEMA_signal_5109, new_AGEMA_signal_5108, stateArray_outS30ser_MC[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS30_MC_mux_inst_1_U1 ( .s (stateArray_n22), .b ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .a ({new_AGEMA_signal_4633, new_AGEMA_signal_4632, new_AGEMA_signal_4631, StateInMC[9]}), .c ({new_AGEMA_signal_5113, new_AGEMA_signal_5112, new_AGEMA_signal_5111, stateArray_outS30ser_MC[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS30_MC_mux_inst_2_U1 ( .s (stateArray_n22), .b ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .a ({new_AGEMA_signal_4636, new_AGEMA_signal_4635, new_AGEMA_signal_4634, StateInMC[10]}), .c ({new_AGEMA_signal_5116, new_AGEMA_signal_5115, new_AGEMA_signal_5114, stateArray_outS30ser_MC[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS30_MC_mux_inst_3_U1 ( .s (stateArray_n22), .b ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .a ({new_AGEMA_signal_4639, new_AGEMA_signal_4638, new_AGEMA_signal_4637, StateInMC[11]}), .c ({new_AGEMA_signal_5119, new_AGEMA_signal_5118, new_AGEMA_signal_5117, stateArray_outS30ser_MC[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS30_MC_mux_inst_4_U1 ( .s (stateArray_n22), .b ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .a ({new_AGEMA_signal_4642, new_AGEMA_signal_4641, new_AGEMA_signal_4640, StateInMC[12]}), .c ({new_AGEMA_signal_5122, new_AGEMA_signal_5121, new_AGEMA_signal_5120, stateArray_outS30ser_MC[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS30_MC_mux_inst_5_U1 ( .s (stateArray_n22), .b ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .a ({new_AGEMA_signal_4645, new_AGEMA_signal_4644, new_AGEMA_signal_4643, StateInMC[13]}), .c ({new_AGEMA_signal_5125, new_AGEMA_signal_5124, new_AGEMA_signal_5123, stateArray_outS30ser_MC[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS30_MC_mux_inst_6_U1 ( .s (stateArray_n22), .b ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .a ({new_AGEMA_signal_4648, new_AGEMA_signal_4647, new_AGEMA_signal_4646, StateInMC[14]}), .c ({new_AGEMA_signal_5128, new_AGEMA_signal_5127, new_AGEMA_signal_5126, stateArray_outS30ser_MC[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_outS30_MC_mux_inst_7_U1 ( .s (stateArray_n22), .b ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .a ({new_AGEMA_signal_4651, new_AGEMA_signal_4650, new_AGEMA_signal_4649, StateInMC[15]}), .c ({new_AGEMA_signal_5131, new_AGEMA_signal_5130, new_AGEMA_signal_5129, stateArray_outS30ser_MC[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS23ser_mux_inst_0_U1 ( .s (stateArray_n27), .b ({plaintext_s3[32], plaintext_s2[32], plaintext_s1[32], plaintext_s0[32]}), .a ({new_AGEMA_signal_5110, new_AGEMA_signal_5109, new_AGEMA_signal_5108, stateArray_outS30ser_MC[0]}), .c ({new_AGEMA_signal_5272, new_AGEMA_signal_5271, new_AGEMA_signal_5270, stateArray_inS23ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS23ser_mux_inst_1_U1 ( .s (stateArray_n27), .b ({plaintext_s3[33], plaintext_s2[33], plaintext_s1[33], plaintext_s0[33]}), .a ({new_AGEMA_signal_5113, new_AGEMA_signal_5112, new_AGEMA_signal_5111, stateArray_outS30ser_MC[1]}), .c ({new_AGEMA_signal_5278, new_AGEMA_signal_5277, new_AGEMA_signal_5276, stateArray_inS23ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS23ser_mux_inst_2_U1 ( .s (stateArray_n27), .b ({plaintext_s3[34], plaintext_s2[34], plaintext_s1[34], plaintext_s0[34]}), .a ({new_AGEMA_signal_5116, new_AGEMA_signal_5115, new_AGEMA_signal_5114, stateArray_outS30ser_MC[2]}), .c ({new_AGEMA_signal_5284, new_AGEMA_signal_5283, new_AGEMA_signal_5282, stateArray_inS23ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS23ser_mux_inst_3_U1 ( .s (stateArray_n27), .b ({plaintext_s3[35], plaintext_s2[35], plaintext_s1[35], plaintext_s0[35]}), .a ({new_AGEMA_signal_5119, new_AGEMA_signal_5118, new_AGEMA_signal_5117, stateArray_outS30ser_MC[3]}), .c ({new_AGEMA_signal_5290, new_AGEMA_signal_5289, new_AGEMA_signal_5288, stateArray_inS23ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS23ser_mux_inst_4_U1 ( .s (stateArray_n27), .b ({plaintext_s3[36], plaintext_s2[36], plaintext_s1[36], plaintext_s0[36]}), .a ({new_AGEMA_signal_5122, new_AGEMA_signal_5121, new_AGEMA_signal_5120, stateArray_outS30ser_MC[4]}), .c ({new_AGEMA_signal_5296, new_AGEMA_signal_5295, new_AGEMA_signal_5294, stateArray_inS23ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS23ser_mux_inst_5_U1 ( .s (stateArray_n27), .b ({plaintext_s3[37], plaintext_s2[37], plaintext_s1[37], plaintext_s0[37]}), .a ({new_AGEMA_signal_5125, new_AGEMA_signal_5124, new_AGEMA_signal_5123, stateArray_outS30ser_MC[5]}), .c ({new_AGEMA_signal_5302, new_AGEMA_signal_5301, new_AGEMA_signal_5300, stateArray_inS23ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS23ser_mux_inst_6_U1 ( .s (stateArray_n27), .b ({plaintext_s3[38], plaintext_s2[38], plaintext_s1[38], plaintext_s0[38]}), .a ({new_AGEMA_signal_5128, new_AGEMA_signal_5127, new_AGEMA_signal_5126, stateArray_outS30ser_MC[6]}), .c ({new_AGEMA_signal_5308, new_AGEMA_signal_5307, new_AGEMA_signal_5306, stateArray_inS23ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS23ser_mux_inst_7_U1 ( .s (stateArray_n27), .b ({plaintext_s3[39], plaintext_s2[39], plaintext_s1[39], plaintext_s0[39]}), .a ({new_AGEMA_signal_5131, new_AGEMA_signal_5130, new_AGEMA_signal_5129, stateArray_outS30ser_MC[7]}), .c ({new_AGEMA_signal_5314, new_AGEMA_signal_5313, new_AGEMA_signal_5312, stateArray_inS23ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS30ser_mux_inst_0_U1 ( .s (stateArray_n26), .b ({plaintext_s3[24], plaintext_s2[24], plaintext_s1[24], plaintext_s0[24]}), .a ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_3154, new_AGEMA_signal_3153, new_AGEMA_signal_3152, stateArray_inS30ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS30ser_mux_inst_1_U1 ( .s (stateArray_n26), .b ({plaintext_s3[25], plaintext_s2[25], plaintext_s1[25], plaintext_s0[25]}), .a ({ciphertext_s3[17], ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, new_AGEMA_signal_3161, stateArray_inS30ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS30ser_mux_inst_2_U1 ( .s (stateArray_n26), .b ({plaintext_s3[26], plaintext_s2[26], plaintext_s1[26], plaintext_s0[26]}), .a ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_3172, new_AGEMA_signal_3171, new_AGEMA_signal_3170, stateArray_inS30ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS30ser_mux_inst_3_U1 ( .s (stateArray_n26), .b ({plaintext_s3[27], plaintext_s2[27], plaintext_s1[27], plaintext_s0[27]}), .a ({ciphertext_s3[19], ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .c ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, new_AGEMA_signal_3179, stateArray_inS30ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS30ser_mux_inst_4_U1 ( .s (stateArray_n26), .b ({plaintext_s3[28], plaintext_s2[28], plaintext_s1[28], plaintext_s0[28]}), .a ({ciphertext_s3[20], ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .c ({new_AGEMA_signal_3190, new_AGEMA_signal_3189, new_AGEMA_signal_3188, stateArray_inS30ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS30ser_mux_inst_5_U1 ( .s (stateArray_n26), .b ({plaintext_s3[29], plaintext_s2[29], plaintext_s1[29], plaintext_s0[29]}), .a ({ciphertext_s3[21], ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .c ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, new_AGEMA_signal_3197, stateArray_inS30ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS30ser_mux_inst_6_U1 ( .s (stateArray_n26), .b ({plaintext_s3[30], plaintext_s2[30], plaintext_s1[30], plaintext_s0[30]}), .a ({ciphertext_s3[22], ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .c ({new_AGEMA_signal_3208, new_AGEMA_signal_3207, new_AGEMA_signal_3206, stateArray_inS30ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS30ser_mux_inst_7_U1 ( .s (stateArray_n26), .b ({plaintext_s3[31], plaintext_s2[31], plaintext_s1[31], plaintext_s0[31]}), .a ({ciphertext_s3[23], ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .c ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, new_AGEMA_signal_3215, stateArray_inS30ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS31ser_mux_inst_0_U1 ( .s (stateArray_n26), .b ({plaintext_s3[16], plaintext_s2[16], plaintext_s1[16], plaintext_s0[16]}), .a ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .c ({new_AGEMA_signal_3226, new_AGEMA_signal_3225, new_AGEMA_signal_3224, stateArray_inS31ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS31ser_mux_inst_1_U1 ( .s (stateArray_n26), .b ({plaintext_s3[17], plaintext_s2[17], plaintext_s1[17], plaintext_s0[17]}), .a ({ciphertext_s3[9], ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .c ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, new_AGEMA_signal_3233, stateArray_inS31ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS31ser_mux_inst_2_U1 ( .s (stateArray_n26), .b ({plaintext_s3[18], plaintext_s2[18], plaintext_s1[18], plaintext_s0[18]}), .a ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_3244, new_AGEMA_signal_3243, new_AGEMA_signal_3242, stateArray_inS31ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS31ser_mux_inst_3_U1 ( .s (stateArray_n26), .b ({plaintext_s3[19], plaintext_s2[19], plaintext_s1[19], plaintext_s0[19]}), .a ({ciphertext_s3[11], ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .c ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, new_AGEMA_signal_3251, stateArray_inS31ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS31ser_mux_inst_4_U1 ( .s (stateArray_n26), .b ({plaintext_s3[20], plaintext_s2[20], plaintext_s1[20], plaintext_s0[20]}), .a ({ciphertext_s3[12], ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .c ({new_AGEMA_signal_3262, new_AGEMA_signal_3261, new_AGEMA_signal_3260, stateArray_inS31ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS31ser_mux_inst_5_U1 ( .s (stateArray_n26), .b ({plaintext_s3[21], plaintext_s2[21], plaintext_s1[21], plaintext_s0[21]}), .a ({ciphertext_s3[13], ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .c ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, new_AGEMA_signal_3269, stateArray_inS31ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS31ser_mux_inst_6_U1 ( .s (stateArray_n26), .b ({plaintext_s3[22], plaintext_s2[22], plaintext_s1[22], plaintext_s0[22]}), .a ({ciphertext_s3[14], ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .c ({new_AGEMA_signal_3280, new_AGEMA_signal_3279, new_AGEMA_signal_3278, stateArray_inS31ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS31ser_mux_inst_7_U1 ( .s (stateArray_n26), .b ({plaintext_s3[23], plaintext_s2[23], plaintext_s1[23], plaintext_s0[23]}), .a ({ciphertext_s3[15], ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .c ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, new_AGEMA_signal_3287, stateArray_inS31ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS32ser_mux_inst_0_U1 ( .s (stateArray_n25), .b ({plaintext_s3[8], plaintext_s2[8], plaintext_s1[8], plaintext_s0[8]}), .a ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_3298, new_AGEMA_signal_3297, new_AGEMA_signal_3296, stateArray_inS32ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS32ser_mux_inst_1_U1 ( .s (stateArray_n25), .b ({plaintext_s3[9], plaintext_s2[9], plaintext_s1[9], plaintext_s0[9]}), .a ({ciphertext_s3[1], ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, new_AGEMA_signal_3305, stateArray_inS32ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS32ser_mux_inst_2_U1 ( .s (stateArray_n25), .b ({plaintext_s3[10], plaintext_s2[10], plaintext_s1[10], plaintext_s0[10]}), .a ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_3316, new_AGEMA_signal_3315, new_AGEMA_signal_3314, stateArray_inS32ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS32ser_mux_inst_3_U1 ( .s (stateArray_n25), .b ({plaintext_s3[11], plaintext_s2[11], plaintext_s1[11], plaintext_s0[11]}), .a ({ciphertext_s3[3], ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .c ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, new_AGEMA_signal_3323, stateArray_inS32ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS32ser_mux_inst_4_U1 ( .s (stateArray_n25), .b ({plaintext_s3[12], plaintext_s2[12], plaintext_s1[12], plaintext_s0[12]}), .a ({ciphertext_s3[4], ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .c ({new_AGEMA_signal_3334, new_AGEMA_signal_3333, new_AGEMA_signal_3332, stateArray_inS32ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS32ser_mux_inst_5_U1 ( .s (stateArray_n25), .b ({plaintext_s3[13], plaintext_s2[13], plaintext_s1[13], plaintext_s0[13]}), .a ({ciphertext_s3[5], ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .c ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, new_AGEMA_signal_3341, stateArray_inS32ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS32ser_mux_inst_6_U1 ( .s (stateArray_n25), .b ({plaintext_s3[14], plaintext_s2[14], plaintext_s1[14], plaintext_s0[14]}), .a ({ciphertext_s3[6], ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .c ({new_AGEMA_signal_3352, new_AGEMA_signal_3351, new_AGEMA_signal_3350, stateArray_inS32ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS32ser_mux_inst_7_U1 ( .s (stateArray_n25), .b ({plaintext_s3[15], plaintext_s2[15], plaintext_s1[15], plaintext_s0[15]}), .a ({ciphertext_s3[7], ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .c ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, new_AGEMA_signal_3359, stateArray_inS32ser[7]}) ) ;
    INV_X1 MUX_StateInMC_U3 ( .A (intFinal), .ZN (MUX_StateInMC_n7) ) ;
    INV_X1 MUX_StateInMC_U2 ( .A (MUX_StateInMC_n7), .ZN (MUX_StateInMC_n6) ) ;
    INV_X1 MUX_StateInMC_U1 ( .A (MUX_StateInMC_n7), .ZN (MUX_StateInMC_n5) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_0_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_4513, new_AGEMA_signal_4512, new_AGEMA_signal_4511, MCout[0]}), .a ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_4618, new_AGEMA_signal_4617, new_AGEMA_signal_4616, StateInMC[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_1_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_4585, new_AGEMA_signal_4584, new_AGEMA_signal_4583, MCout[1]}), .a ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_4621, new_AGEMA_signal_4620, new_AGEMA_signal_4619, StateInMC[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_2_U1 ( .s (intFinal), .b ({new_AGEMA_signal_4507, new_AGEMA_signal_4506, new_AGEMA_signal_4505, MCout[2]}), .a ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_4540, new_AGEMA_signal_4539, new_AGEMA_signal_4538, StateInMC[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_3_U1 ( .s (intFinal), .b ({new_AGEMA_signal_4582, new_AGEMA_signal_4581, new_AGEMA_signal_4580, MCout[3]}), .a ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_4624, new_AGEMA_signal_4623, new_AGEMA_signal_4622, StateInMC[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_4_U1 ( .s (intFinal), .b ({new_AGEMA_signal_4579, new_AGEMA_signal_4578, new_AGEMA_signal_4577, MCout[4]}), .a ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_4627, new_AGEMA_signal_4626, new_AGEMA_signal_4625, StateInMC[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_5_U1 ( .s (intFinal), .b ({new_AGEMA_signal_4498, new_AGEMA_signal_4497, new_AGEMA_signal_4496, MCout[5]}), .a ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, new_AGEMA_signal_4541, StateInMC[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_6_U1 ( .s (intFinal), .b ({new_AGEMA_signal_4495, new_AGEMA_signal_4494, new_AGEMA_signal_4493, MCout[6]}), .a ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .c ({new_AGEMA_signal_4546, new_AGEMA_signal_4545, new_AGEMA_signal_4544, StateInMC[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_7_U1 ( .s (intFinal), .b ({new_AGEMA_signal_4492, new_AGEMA_signal_4491, new_AGEMA_signal_4490, MCout[7]}), .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .c ({new_AGEMA_signal_4549, new_AGEMA_signal_4548, new_AGEMA_signal_4547, StateInMC[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_8_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_4489, new_AGEMA_signal_4488, new_AGEMA_signal_4487, MCout[8]}), .a ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_4630, new_AGEMA_signal_4629, new_AGEMA_signal_4628, StateInMC[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_9_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_4576, new_AGEMA_signal_4575, new_AGEMA_signal_4574, MCout[9]}), .a ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_4633, new_AGEMA_signal_4632, new_AGEMA_signal_4631, StateInMC[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_10_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_4483, new_AGEMA_signal_4482, new_AGEMA_signal_4481, MCout[10]}), .a ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_4636, new_AGEMA_signal_4635, new_AGEMA_signal_4634, StateInMC[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_11_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_4573, new_AGEMA_signal_4572, new_AGEMA_signal_4571, MCout[11]}), .a ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_4639, new_AGEMA_signal_4638, new_AGEMA_signal_4637, StateInMC[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_12_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_4570, new_AGEMA_signal_4569, new_AGEMA_signal_4568, MCout[12]}), .a ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_4642, new_AGEMA_signal_4641, new_AGEMA_signal_4640, StateInMC[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_13_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_4474, new_AGEMA_signal_4473, new_AGEMA_signal_4472, MCout[13]}), .a ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_4645, new_AGEMA_signal_4644, new_AGEMA_signal_4643, StateInMC[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_14_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_4471, new_AGEMA_signal_4470, new_AGEMA_signal_4469, MCout[14]}), .a ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .c ({new_AGEMA_signal_4648, new_AGEMA_signal_4647, new_AGEMA_signal_4646, StateInMC[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_15_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_4468, new_AGEMA_signal_4467, new_AGEMA_signal_4466, MCout[15]}), .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .c ({new_AGEMA_signal_4651, new_AGEMA_signal_4650, new_AGEMA_signal_4649, StateInMC[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_16_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_4465, new_AGEMA_signal_4464, new_AGEMA_signal_4463, MCout[16]}), .a ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_4654, new_AGEMA_signal_4653, new_AGEMA_signal_4652, StateInMC[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_17_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_4567, new_AGEMA_signal_4566, new_AGEMA_signal_4565, MCout[17]}), .a ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_4657, new_AGEMA_signal_4656, new_AGEMA_signal_4655, StateInMC[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_18_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_4459, new_AGEMA_signal_4458, new_AGEMA_signal_4457, MCout[18]}), .a ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_4660, new_AGEMA_signal_4659, new_AGEMA_signal_4658, StateInMC[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_19_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_4564, new_AGEMA_signal_4563, new_AGEMA_signal_4562, MCout[19]}), .a ({ciphertext_s3[91], ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_4663, new_AGEMA_signal_4662, new_AGEMA_signal_4661, StateInMC[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_20_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_4561, new_AGEMA_signal_4560, new_AGEMA_signal_4559, MCout[20]}), .a ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_4666, new_AGEMA_signal_4665, new_AGEMA_signal_4664, StateInMC[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_21_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_4450, new_AGEMA_signal_4449, new_AGEMA_signal_4448, MCout[21]}), .a ({ciphertext_s3[93], ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_4669, new_AGEMA_signal_4668, new_AGEMA_signal_4667, StateInMC[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_22_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_4447, new_AGEMA_signal_4446, new_AGEMA_signal_4445, MCout[22]}), .a ({ciphertext_s3[94], ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .c ({new_AGEMA_signal_4672, new_AGEMA_signal_4671, new_AGEMA_signal_4670, StateInMC[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_23_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_4444, new_AGEMA_signal_4443, new_AGEMA_signal_4442, MCout[23]}), .a ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .c ({new_AGEMA_signal_4675, new_AGEMA_signal_4674, new_AGEMA_signal_4673, StateInMC[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_24_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, new_AGEMA_signal_4439, MCout[24]}), .a ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_4678, new_AGEMA_signal_4677, new_AGEMA_signal_4676, StateInMC[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_25_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_4558, new_AGEMA_signal_4557, new_AGEMA_signal_4556, MCout[25]}), .a ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_4681, new_AGEMA_signal_4680, new_AGEMA_signal_4679, StateInMC[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_26_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_4435, new_AGEMA_signal_4434, new_AGEMA_signal_4433, MCout[26]}), .a ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_4684, new_AGEMA_signal_4683, new_AGEMA_signal_4682, StateInMC[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_27_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_4555, new_AGEMA_signal_4554, new_AGEMA_signal_4553, MCout[27]}), .a ({ciphertext_s3[123], ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_4687, new_AGEMA_signal_4686, new_AGEMA_signal_4685, StateInMC[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_28_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, new_AGEMA_signal_4550, MCout[28]}), .a ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_4690, new_AGEMA_signal_4689, new_AGEMA_signal_4688, StateInMC[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_29_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_4426, new_AGEMA_signal_4425, new_AGEMA_signal_4424, MCout[29]}), .a ({ciphertext_s3[125], ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_4693, new_AGEMA_signal_4692, new_AGEMA_signal_4691, StateInMC[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_30_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_4423, new_AGEMA_signal_4422, new_AGEMA_signal_4421, MCout[30]}), .a ({ciphertext_s3[126], ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .c ({new_AGEMA_signal_4696, new_AGEMA_signal_4695, new_AGEMA_signal_4694, StateInMC[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateInMC_mux_inst_31_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_4420, new_AGEMA_signal_4419, new_AGEMA_signal_4418, MCout[31]}), .a ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .c ({new_AGEMA_signal_4699, new_AGEMA_signal_4698, new_AGEMA_signal_4697, StateInMC[31]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U50 ( .a ({new_AGEMA_signal_2056, new_AGEMA_signal_2055, new_AGEMA_signal_2054, KeyArray_outS01ser_7_}), .b ({new_AGEMA_signal_2050, new_AGEMA_signal_2049, new_AGEMA_signal_2048, keyStateIn[7]}), .c ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, new_AGEMA_signal_2057, KeyArray_outS01ser_XOR_00[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U49 ( .a ({new_AGEMA_signal_2062, new_AGEMA_signal_2061, new_AGEMA_signal_2060, KeyArray_outS01ser_6_}), .b ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, new_AGEMA_signal_2039, keyStateIn[6]}), .c ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, new_AGEMA_signal_2063, KeyArray_outS01ser_XOR_00[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U48 ( .a ({new_AGEMA_signal_2068, new_AGEMA_signal_2067, new_AGEMA_signal_2066, KeyArray_outS01ser_5_}), .b ({new_AGEMA_signal_2032, new_AGEMA_signal_2031, new_AGEMA_signal_2030, keyStateIn[5]}), .c ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, new_AGEMA_signal_2069, KeyArray_outS01ser_XOR_00[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U47 ( .a ({new_AGEMA_signal_2074, new_AGEMA_signal_2073, new_AGEMA_signal_2072, KeyArray_outS01ser_4_}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, new_AGEMA_signal_2021, keyStateIn[4]}), .c ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, new_AGEMA_signal_2075, KeyArray_outS01ser_XOR_00[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U46 ( .a ({new_AGEMA_signal_2080, new_AGEMA_signal_2079, new_AGEMA_signal_2078, KeyArray_outS01ser_3_}), .b ({new_AGEMA_signal_2014, new_AGEMA_signal_2013, new_AGEMA_signal_2012, keyStateIn[3]}), .c ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, new_AGEMA_signal_2081, KeyArray_outS01ser_XOR_00[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U45 ( .a ({new_AGEMA_signal_2086, new_AGEMA_signal_2085, new_AGEMA_signal_2084, KeyArray_outS01ser_2_}), .b ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, new_AGEMA_signal_2003, keyStateIn[2]}), .c ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, new_AGEMA_signal_2087, KeyArray_outS01ser_XOR_00[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U44 ( .a ({new_AGEMA_signal_2092, new_AGEMA_signal_2091, new_AGEMA_signal_2090, KeyArray_outS01ser_1_}), .b ({new_AGEMA_signal_1996, new_AGEMA_signal_1995, new_AGEMA_signal_1994, keyStateIn[1]}), .c ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, new_AGEMA_signal_2093, KeyArray_outS01ser_XOR_00[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U43 ( .a ({new_AGEMA_signal_2098, new_AGEMA_signal_2097, new_AGEMA_signal_2096, KeyArray_outS01ser_0_}), .b ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, new_AGEMA_signal_1985, keyStateIn[0]}), .c ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, new_AGEMA_signal_2099, KeyArray_outS01ser_XOR_00[0]}) ) ;
    INV_X1 KeyArray_U26 ( .A (KeyArray_n47), .ZN (KeyArray_n46) ) ;
    INV_X1 KeyArray_U25 ( .A (KeyArray_n47), .ZN (KeyArray_n45) ) ;
    INV_X1 KeyArray_U24 ( .A (KeyArray_n47), .ZN (KeyArray_n44) ) ;
    INV_X1 KeyArray_U23 ( .A (KeyArray_n47), .ZN (KeyArray_n43) ) ;
    INV_X1 KeyArray_U22 ( .A (KeyArray_n47), .ZN (KeyArray_n42) ) ;
    INV_X1 KeyArray_U21 ( .A (KeyArray_n47), .ZN (KeyArray_n41) ) ;
    INV_X1 KeyArray_U20 ( .A (KeyArray_n47), .ZN (KeyArray_n40) ) ;
    INV_X1 KeyArray_U19 ( .A (KeyArray_n47), .ZN (KeyArray_n39) ) ;
    INV_X1 KeyArray_U18 ( .A (nReset), .ZN (KeyArray_n47) ) ;
    INV_X1 KeyArray_U17 ( .A (KeyArray_n38), .ZN (KeyArray_n31) ) ;
    INV_X1 KeyArray_U16 ( .A (KeyArray_n29), .ZN (KeyArray_n23) ) ;
    INV_X1 KeyArray_U15 ( .A (KeyArray_n38), .ZN (KeyArray_n37) ) ;
    INV_X1 KeyArray_U14 ( .A (KeyArray_n29), .ZN (KeyArray_n28) ) ;
    INV_X1 KeyArray_U13 ( .A (KeyArray_n38), .ZN (KeyArray_n36) ) ;
    INV_X1 KeyArray_U12 ( .A (KeyArray_n29), .ZN (KeyArray_n27) ) ;
    INV_X1 KeyArray_U11 ( .A (KeyArray_n38), .ZN (KeyArray_n35) ) ;
    INV_X1 KeyArray_U10 ( .A (KeyArray_n29), .ZN (KeyArray_n26) ) ;
    INV_X1 KeyArray_U9 ( .A (KeyArray_n38), .ZN (KeyArray_n32) ) ;
    INV_X1 KeyArray_U8 ( .A (KeyArray_n29), .ZN (KeyArray_n24) ) ;
    INV_X1 KeyArray_U7 ( .A (KeyArray_n38), .ZN (KeyArray_n33) ) ;
    INV_X1 KeyArray_U6 ( .A (KeyArray_n29), .ZN (KeyArray_n25) ) ;
    INV_X1 KeyArray_U5 ( .A (KeyArray_n38), .ZN (KeyArray_n30) ) ;
    INV_X1 KeyArray_U4 ( .A (KeyArray_n29), .ZN (KeyArray_n22) ) ;
    INV_X1 KeyArray_U3 ( .A (KeyArray_n38), .ZN (KeyArray_n34) ) ;
    INV_X1 KeyArray_U2 ( .A (selMC), .ZN (KeyArray_n38) ) ;
    INV_X1 KeyArray_U1 ( .A (n12), .ZN (KeyArray_n29) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_0_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, new_AGEMA_signal_1985, keyStateIn[0]}), .a ({new_AGEMA_signal_5839, new_AGEMA_signal_5838, new_AGEMA_signal_5837, KeyArray_S00reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_6163, new_AGEMA_signal_6162, new_AGEMA_signal_6161, KeyArray_S00reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_5779, new_AGEMA_signal_5778, new_AGEMA_signal_5777, KeyArray_inS00ser[0]}), .a ({new_AGEMA_signal_3511, new_AGEMA_signal_3510, new_AGEMA_signal_3509, KeyArray_outS10ser[0]}), .c ({new_AGEMA_signal_5839, new_AGEMA_signal_5838, new_AGEMA_signal_5837, KeyArray_S00reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_1_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_1996, new_AGEMA_signal_1995, new_AGEMA_signal_1994, keyStateIn[1]}), .a ({new_AGEMA_signal_5842, new_AGEMA_signal_5841, new_AGEMA_signal_5840, KeyArray_S00reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_6166, new_AGEMA_signal_6165, new_AGEMA_signal_6164, KeyArray_S00reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_5785, new_AGEMA_signal_5784, new_AGEMA_signal_5783, KeyArray_inS00ser[1]}), .a ({new_AGEMA_signal_3520, new_AGEMA_signal_3519, new_AGEMA_signal_3518, KeyArray_outS10ser[1]}), .c ({new_AGEMA_signal_5842, new_AGEMA_signal_5841, new_AGEMA_signal_5840, KeyArray_S00reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_2_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, new_AGEMA_signal_2003, keyStateIn[2]}), .a ({new_AGEMA_signal_5845, new_AGEMA_signal_5844, new_AGEMA_signal_5843, KeyArray_S00reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_6169, new_AGEMA_signal_6168, new_AGEMA_signal_6167, KeyArray_S00reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_5791, new_AGEMA_signal_5790, new_AGEMA_signal_5789, KeyArray_inS00ser[2]}), .a ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, new_AGEMA_signal_3527, KeyArray_outS10ser[2]}), .c ({new_AGEMA_signal_5845, new_AGEMA_signal_5844, new_AGEMA_signal_5843, KeyArray_S00reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_3_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2014, new_AGEMA_signal_2013, new_AGEMA_signal_2012, keyStateIn[3]}), .a ({new_AGEMA_signal_5848, new_AGEMA_signal_5847, new_AGEMA_signal_5846, KeyArray_S00reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_6172, new_AGEMA_signal_6171, new_AGEMA_signal_6170, KeyArray_S00reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_5797, new_AGEMA_signal_5796, new_AGEMA_signal_5795, KeyArray_inS00ser[3]}), .a ({new_AGEMA_signal_3538, new_AGEMA_signal_3537, new_AGEMA_signal_3536, KeyArray_outS10ser[3]}), .c ({new_AGEMA_signal_5848, new_AGEMA_signal_5847, new_AGEMA_signal_5846, KeyArray_S00reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_4_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, new_AGEMA_signal_2021, keyStateIn[4]}), .a ({new_AGEMA_signal_5851, new_AGEMA_signal_5850, new_AGEMA_signal_5849, KeyArray_S00reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_6175, new_AGEMA_signal_6174, new_AGEMA_signal_6173, KeyArray_S00reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_5803, new_AGEMA_signal_5802, new_AGEMA_signal_5801, KeyArray_inS00ser[4]}), .a ({new_AGEMA_signal_3547, new_AGEMA_signal_3546, new_AGEMA_signal_3545, KeyArray_outS10ser[4]}), .c ({new_AGEMA_signal_5851, new_AGEMA_signal_5850, new_AGEMA_signal_5849, KeyArray_S00reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_5_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2032, new_AGEMA_signal_2031, new_AGEMA_signal_2030, keyStateIn[5]}), .a ({new_AGEMA_signal_5854, new_AGEMA_signal_5853, new_AGEMA_signal_5852, KeyArray_S00reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_6178, new_AGEMA_signal_6177, new_AGEMA_signal_6176, KeyArray_S00reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_5809, new_AGEMA_signal_5808, new_AGEMA_signal_5807, KeyArray_inS00ser[5]}), .a ({new_AGEMA_signal_3556, new_AGEMA_signal_3555, new_AGEMA_signal_3554, KeyArray_outS10ser[5]}), .c ({new_AGEMA_signal_5854, new_AGEMA_signal_5853, new_AGEMA_signal_5852, KeyArray_S00reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_6_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, new_AGEMA_signal_2039, keyStateIn[6]}), .a ({new_AGEMA_signal_5857, new_AGEMA_signal_5856, new_AGEMA_signal_5855, KeyArray_S00reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_6181, new_AGEMA_signal_6180, new_AGEMA_signal_6179, KeyArray_S00reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_5815, new_AGEMA_signal_5814, new_AGEMA_signal_5813, KeyArray_inS00ser[6]}), .a ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, new_AGEMA_signal_3563, KeyArray_outS10ser[6]}), .c ({new_AGEMA_signal_5857, new_AGEMA_signal_5856, new_AGEMA_signal_5855, KeyArray_S00reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_7_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2050, new_AGEMA_signal_2049, new_AGEMA_signal_2048, keyStateIn[7]}), .a ({new_AGEMA_signal_5860, new_AGEMA_signal_5859, new_AGEMA_signal_5858, KeyArray_S00reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_6184, new_AGEMA_signal_6183, new_AGEMA_signal_6182, KeyArray_S00reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_5821, new_AGEMA_signal_5820, new_AGEMA_signal_5819, KeyArray_inS00ser[7]}), .a ({new_AGEMA_signal_3574, new_AGEMA_signal_3573, new_AGEMA_signal_3572, KeyArray_outS10ser[7]}), .c ({new_AGEMA_signal_5860, new_AGEMA_signal_5859, new_AGEMA_signal_5858, KeyArray_S00reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_0_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2098, new_AGEMA_signal_2097, new_AGEMA_signal_2096, KeyArray_outS01ser_0_}), .a ({new_AGEMA_signal_4702, new_AGEMA_signal_4701, new_AGEMA_signal_4700, KeyArray_S01reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_5863, new_AGEMA_signal_5862, new_AGEMA_signal_5861, KeyArray_S01reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3370, new_AGEMA_signal_3369, new_AGEMA_signal_3368, KeyArray_inS01ser[0]}), .a ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, new_AGEMA_signal_3581, KeyArray_outS11ser[0]}), .c ({new_AGEMA_signal_4702, new_AGEMA_signal_4701, new_AGEMA_signal_4700, KeyArray_S01reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_1_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2092, new_AGEMA_signal_2091, new_AGEMA_signal_2090, KeyArray_outS01ser_1_}), .a ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, new_AGEMA_signal_4703, KeyArray_S01reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_5866, new_AGEMA_signal_5865, new_AGEMA_signal_5864, KeyArray_S01reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3379, new_AGEMA_signal_3378, new_AGEMA_signal_3377, KeyArray_inS01ser[1]}), .a ({new_AGEMA_signal_3592, new_AGEMA_signal_3591, new_AGEMA_signal_3590, KeyArray_outS11ser[1]}), .c ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, new_AGEMA_signal_4703, KeyArray_S01reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_2_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2086, new_AGEMA_signal_2085, new_AGEMA_signal_2084, KeyArray_outS01ser_2_}), .a ({new_AGEMA_signal_4708, new_AGEMA_signal_4707, new_AGEMA_signal_4706, KeyArray_S01reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_5869, new_AGEMA_signal_5868, new_AGEMA_signal_5867, KeyArray_S01reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3388, new_AGEMA_signal_3387, new_AGEMA_signal_3386, KeyArray_inS01ser[2]}), .a ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, new_AGEMA_signal_3599, KeyArray_outS11ser[2]}), .c ({new_AGEMA_signal_4708, new_AGEMA_signal_4707, new_AGEMA_signal_4706, KeyArray_S01reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_3_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2080, new_AGEMA_signal_2079, new_AGEMA_signal_2078, KeyArray_outS01ser_3_}), .a ({new_AGEMA_signal_4711, new_AGEMA_signal_4710, new_AGEMA_signal_4709, KeyArray_S01reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_5872, new_AGEMA_signal_5871, new_AGEMA_signal_5870, KeyArray_S01reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, new_AGEMA_signal_3395, KeyArray_inS01ser[3]}), .a ({new_AGEMA_signal_3610, new_AGEMA_signal_3609, new_AGEMA_signal_3608, KeyArray_outS11ser[3]}), .c ({new_AGEMA_signal_4711, new_AGEMA_signal_4710, new_AGEMA_signal_4709, KeyArray_S01reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_4_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2074, new_AGEMA_signal_2073, new_AGEMA_signal_2072, KeyArray_outS01ser_4_}), .a ({new_AGEMA_signal_4714, new_AGEMA_signal_4713, new_AGEMA_signal_4712, KeyArray_S01reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_5875, new_AGEMA_signal_5874, new_AGEMA_signal_5873, KeyArray_S01reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3406, new_AGEMA_signal_3405, new_AGEMA_signal_3404, KeyArray_inS01ser[4]}), .a ({new_AGEMA_signal_3619, new_AGEMA_signal_3618, new_AGEMA_signal_3617, KeyArray_outS11ser[4]}), .c ({new_AGEMA_signal_4714, new_AGEMA_signal_4713, new_AGEMA_signal_4712, KeyArray_S01reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_5_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2068, new_AGEMA_signal_2067, new_AGEMA_signal_2066, KeyArray_outS01ser_5_}), .a ({new_AGEMA_signal_4717, new_AGEMA_signal_4716, new_AGEMA_signal_4715, KeyArray_S01reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_5878, new_AGEMA_signal_5877, new_AGEMA_signal_5876, KeyArray_S01reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3415, new_AGEMA_signal_3414, new_AGEMA_signal_3413, KeyArray_inS01ser[5]}), .a ({new_AGEMA_signal_3628, new_AGEMA_signal_3627, new_AGEMA_signal_3626, KeyArray_outS11ser[5]}), .c ({new_AGEMA_signal_4717, new_AGEMA_signal_4716, new_AGEMA_signal_4715, KeyArray_S01reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_6_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2062, new_AGEMA_signal_2061, new_AGEMA_signal_2060, KeyArray_outS01ser_6_}), .a ({new_AGEMA_signal_4720, new_AGEMA_signal_4719, new_AGEMA_signal_4718, KeyArray_S01reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_5881, new_AGEMA_signal_5880, new_AGEMA_signal_5879, KeyArray_S01reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3424, new_AGEMA_signal_3423, new_AGEMA_signal_3422, KeyArray_inS01ser[6]}), .a ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, new_AGEMA_signal_3635, KeyArray_outS11ser[6]}), .c ({new_AGEMA_signal_4720, new_AGEMA_signal_4719, new_AGEMA_signal_4718, KeyArray_S01reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_7_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2056, new_AGEMA_signal_2055, new_AGEMA_signal_2054, KeyArray_outS01ser_7_}), .a ({new_AGEMA_signal_4723, new_AGEMA_signal_4722, new_AGEMA_signal_4721, KeyArray_S01reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_5884, new_AGEMA_signal_5883, new_AGEMA_signal_5882, KeyArray_S01reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, new_AGEMA_signal_3431, KeyArray_inS01ser[7]}), .a ({new_AGEMA_signal_3646, new_AGEMA_signal_3645, new_AGEMA_signal_3644, KeyArray_outS11ser[7]}), .c ({new_AGEMA_signal_4723, new_AGEMA_signal_4722, new_AGEMA_signal_4721, KeyArray_S01reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_0_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, new_AGEMA_signal_3365, KeyArray_outS02ser[0]}), .a ({new_AGEMA_signal_4726, new_AGEMA_signal_4725, new_AGEMA_signal_4724, KeyArray_S02reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_5887, new_AGEMA_signal_5886, new_AGEMA_signal_5885, KeyArray_S02reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_3442, new_AGEMA_signal_3441, new_AGEMA_signal_3440, KeyArray_inS02ser[0]}), .a ({new_AGEMA_signal_3655, new_AGEMA_signal_3654, new_AGEMA_signal_3653, KeyArray_outS12ser[0]}), .c ({new_AGEMA_signal_4726, new_AGEMA_signal_4725, new_AGEMA_signal_4724, KeyArray_S02reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_1_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_3376, new_AGEMA_signal_3375, new_AGEMA_signal_3374, KeyArray_outS02ser[1]}), .a ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, new_AGEMA_signal_4727, KeyArray_S02reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_5890, new_AGEMA_signal_5889, new_AGEMA_signal_5888, KeyArray_S02reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_3451, new_AGEMA_signal_3450, new_AGEMA_signal_3449, KeyArray_inS02ser[1]}), .a ({new_AGEMA_signal_3664, new_AGEMA_signal_3663, new_AGEMA_signal_3662, KeyArray_outS12ser[1]}), .c ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, new_AGEMA_signal_4727, KeyArray_S02reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_2_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, new_AGEMA_signal_3383, KeyArray_outS02ser[2]}), .a ({new_AGEMA_signal_4732, new_AGEMA_signal_4731, new_AGEMA_signal_4730, KeyArray_S02reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_5893, new_AGEMA_signal_5892, new_AGEMA_signal_5891, KeyArray_S02reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_3460, new_AGEMA_signal_3459, new_AGEMA_signal_3458, KeyArray_inS02ser[2]}), .a ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, new_AGEMA_signal_3671, KeyArray_outS12ser[2]}), .c ({new_AGEMA_signal_4732, new_AGEMA_signal_4731, new_AGEMA_signal_4730, KeyArray_S02reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_3_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_3394, new_AGEMA_signal_3393, new_AGEMA_signal_3392, KeyArray_outS02ser[3]}), .a ({new_AGEMA_signal_4735, new_AGEMA_signal_4734, new_AGEMA_signal_4733, KeyArray_S02reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_5896, new_AGEMA_signal_5895, new_AGEMA_signal_5894, KeyArray_S02reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, new_AGEMA_signal_3467, KeyArray_inS02ser[3]}), .a ({new_AGEMA_signal_3682, new_AGEMA_signal_3681, new_AGEMA_signal_3680, KeyArray_outS12ser[3]}), .c ({new_AGEMA_signal_4735, new_AGEMA_signal_4734, new_AGEMA_signal_4733, KeyArray_S02reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_4_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, new_AGEMA_signal_3401, KeyArray_outS02ser[4]}), .a ({new_AGEMA_signal_4738, new_AGEMA_signal_4737, new_AGEMA_signal_4736, KeyArray_S02reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_5899, new_AGEMA_signal_5898, new_AGEMA_signal_5897, KeyArray_S02reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_3478, new_AGEMA_signal_3477, new_AGEMA_signal_3476, KeyArray_inS02ser[4]}), .a ({new_AGEMA_signal_3691, new_AGEMA_signal_3690, new_AGEMA_signal_3689, KeyArray_outS12ser[4]}), .c ({new_AGEMA_signal_4738, new_AGEMA_signal_4737, new_AGEMA_signal_4736, KeyArray_S02reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_5_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_3412, new_AGEMA_signal_3411, new_AGEMA_signal_3410, KeyArray_outS02ser[5]}), .a ({new_AGEMA_signal_4741, new_AGEMA_signal_4740, new_AGEMA_signal_4739, KeyArray_S02reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_5902, new_AGEMA_signal_5901, new_AGEMA_signal_5900, KeyArray_S02reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_3487, new_AGEMA_signal_3486, new_AGEMA_signal_3485, KeyArray_inS02ser[5]}), .a ({new_AGEMA_signal_3700, new_AGEMA_signal_3699, new_AGEMA_signal_3698, KeyArray_outS12ser[5]}), .c ({new_AGEMA_signal_4741, new_AGEMA_signal_4740, new_AGEMA_signal_4739, KeyArray_S02reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_6_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, new_AGEMA_signal_3419, KeyArray_outS02ser[6]}), .a ({new_AGEMA_signal_4744, new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyArray_S02reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_5905, new_AGEMA_signal_5904, new_AGEMA_signal_5903, KeyArray_S02reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_3496, new_AGEMA_signal_3495, new_AGEMA_signal_3494, KeyArray_inS02ser[6]}), .a ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, new_AGEMA_signal_3707, KeyArray_outS12ser[6]}), .c ({new_AGEMA_signal_4744, new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyArray_S02reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_7_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_3430, new_AGEMA_signal_3429, new_AGEMA_signal_3428, KeyArray_outS02ser[7]}), .a ({new_AGEMA_signal_4747, new_AGEMA_signal_4746, new_AGEMA_signal_4745, KeyArray_S02reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_5908, new_AGEMA_signal_5907, new_AGEMA_signal_5906, KeyArray_S02reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, new_AGEMA_signal_3503, KeyArray_inS02ser[7]}), .a ({new_AGEMA_signal_3718, new_AGEMA_signal_3717, new_AGEMA_signal_3716, KeyArray_outS12ser[7]}), .c ({new_AGEMA_signal_4747, new_AGEMA_signal_4746, new_AGEMA_signal_4745, KeyArray_S02reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_0_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_3439, new_AGEMA_signal_3438, new_AGEMA_signal_3437, KeyArray_outS03ser[0]}), .a ({new_AGEMA_signal_4750, new_AGEMA_signal_4749, new_AGEMA_signal_4748, KeyArray_S03reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_5911, new_AGEMA_signal_5910, new_AGEMA_signal_5909, KeyArray_S03reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_3514, new_AGEMA_signal_3513, new_AGEMA_signal_3512, KeyArray_inS03ser[0]}), .a ({new_AGEMA_signal_3727, new_AGEMA_signal_3726, new_AGEMA_signal_3725, keySBIn[0]}), .c ({new_AGEMA_signal_4750, new_AGEMA_signal_4749, new_AGEMA_signal_4748, KeyArray_S03reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_1_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_3448, new_AGEMA_signal_3447, new_AGEMA_signal_3446, KeyArray_outS03ser[1]}), .a ({new_AGEMA_signal_4753, new_AGEMA_signal_4752, new_AGEMA_signal_4751, KeyArray_S03reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_5914, new_AGEMA_signal_5913, new_AGEMA_signal_5912, KeyArray_S03reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_3523, new_AGEMA_signal_3522, new_AGEMA_signal_3521, KeyArray_inS03ser[1]}), .a ({new_AGEMA_signal_3736, new_AGEMA_signal_3735, new_AGEMA_signal_3734, keySBIn[1]}), .c ({new_AGEMA_signal_4753, new_AGEMA_signal_4752, new_AGEMA_signal_4751, KeyArray_S03reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_2_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, new_AGEMA_signal_3455, KeyArray_outS03ser[2]}), .a ({new_AGEMA_signal_4756, new_AGEMA_signal_4755, new_AGEMA_signal_4754, KeyArray_S03reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_5917, new_AGEMA_signal_5916, new_AGEMA_signal_5915, KeyArray_S03reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_3532, new_AGEMA_signal_3531, new_AGEMA_signal_3530, KeyArray_inS03ser[2]}), .a ({new_AGEMA_signal_3745, new_AGEMA_signal_3744, new_AGEMA_signal_3743, keySBIn[2]}), .c ({new_AGEMA_signal_4756, new_AGEMA_signal_4755, new_AGEMA_signal_4754, KeyArray_S03reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_3_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_3466, new_AGEMA_signal_3465, new_AGEMA_signal_3464, KeyArray_outS03ser[3]}), .a ({new_AGEMA_signal_4759, new_AGEMA_signal_4758, new_AGEMA_signal_4757, KeyArray_S03reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_5920, new_AGEMA_signal_5919, new_AGEMA_signal_5918, KeyArray_S03reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, new_AGEMA_signal_3539, KeyArray_inS03ser[3]}), .a ({new_AGEMA_signal_3754, new_AGEMA_signal_3753, new_AGEMA_signal_3752, keySBIn[3]}), .c ({new_AGEMA_signal_4759, new_AGEMA_signal_4758, new_AGEMA_signal_4757, KeyArray_S03reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_4_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, new_AGEMA_signal_3473, KeyArray_outS03ser[4]}), .a ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, new_AGEMA_signal_4760, KeyArray_S03reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_5923, new_AGEMA_signal_5922, new_AGEMA_signal_5921, KeyArray_S03reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_3550, new_AGEMA_signal_3549, new_AGEMA_signal_3548, KeyArray_inS03ser[4]}), .a ({new_AGEMA_signal_3763, new_AGEMA_signal_3762, new_AGEMA_signal_3761, keySBIn[4]}), .c ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, new_AGEMA_signal_4760, KeyArray_S03reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_5_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_3484, new_AGEMA_signal_3483, new_AGEMA_signal_3482, KeyArray_outS03ser[5]}), .a ({new_AGEMA_signal_4765, new_AGEMA_signal_4764, new_AGEMA_signal_4763, KeyArray_S03reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_5926, new_AGEMA_signal_5925, new_AGEMA_signal_5924, KeyArray_S03reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_3559, new_AGEMA_signal_3558, new_AGEMA_signal_3557, KeyArray_inS03ser[5]}), .a ({new_AGEMA_signal_3772, new_AGEMA_signal_3771, new_AGEMA_signal_3770, keySBIn[5]}), .c ({new_AGEMA_signal_4765, new_AGEMA_signal_4764, new_AGEMA_signal_4763, KeyArray_S03reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_6_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, new_AGEMA_signal_3491, KeyArray_outS03ser[6]}), .a ({new_AGEMA_signal_4768, new_AGEMA_signal_4767, new_AGEMA_signal_4766, KeyArray_S03reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_5929, new_AGEMA_signal_5928, new_AGEMA_signal_5927, KeyArray_S03reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_3568, new_AGEMA_signal_3567, new_AGEMA_signal_3566, KeyArray_inS03ser[6]}), .a ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, new_AGEMA_signal_3779, keySBIn[6]}), .c ({new_AGEMA_signal_4768, new_AGEMA_signal_4767, new_AGEMA_signal_4766, KeyArray_S03reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_7_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_3502, new_AGEMA_signal_3501, new_AGEMA_signal_3500, KeyArray_outS03ser[7]}), .a ({new_AGEMA_signal_4771, new_AGEMA_signal_4770, new_AGEMA_signal_4769, KeyArray_S03reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_5932, new_AGEMA_signal_5931, new_AGEMA_signal_5930, KeyArray_S03reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, new_AGEMA_signal_3575, KeyArray_inS03ser[7]}), .a ({new_AGEMA_signal_3790, new_AGEMA_signal_3789, new_AGEMA_signal_3788, keySBIn[7]}), .c ({new_AGEMA_signal_4771, new_AGEMA_signal_4770, new_AGEMA_signal_4769, KeyArray_S03reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_0_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_3511, new_AGEMA_signal_3510, new_AGEMA_signal_3509, KeyArray_outS10ser[0]}), .a ({new_AGEMA_signal_4774, new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyArray_S10reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_5935, new_AGEMA_signal_5934, new_AGEMA_signal_5933, KeyArray_S10reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_3586, new_AGEMA_signal_3585, new_AGEMA_signal_3584, KeyArray_inS10ser[0]}), .a ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, new_AGEMA_signal_3797, KeyArray_outS20ser[0]}), .c ({new_AGEMA_signal_4774, new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyArray_S10reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_1_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_3520, new_AGEMA_signal_3519, new_AGEMA_signal_3518, KeyArray_outS10ser[1]}), .a ({new_AGEMA_signal_4777, new_AGEMA_signal_4776, new_AGEMA_signal_4775, KeyArray_S10reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_5938, new_AGEMA_signal_5937, new_AGEMA_signal_5936, KeyArray_S10reg_gff_1_SFF_1_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_3595, new_AGEMA_signal_3594, new_AGEMA_signal_3593, KeyArray_inS10ser[1]}), .a ({new_AGEMA_signal_3808, new_AGEMA_signal_3807, new_AGEMA_signal_3806, KeyArray_outS20ser[1]}), .c ({new_AGEMA_signal_4777, new_AGEMA_signal_4776, new_AGEMA_signal_4775, KeyArray_S10reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_2_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, new_AGEMA_signal_3527, KeyArray_outS10ser[2]}), .a ({new_AGEMA_signal_4780, new_AGEMA_signal_4779, new_AGEMA_signal_4778, KeyArray_S10reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_5941, new_AGEMA_signal_5940, new_AGEMA_signal_5939, KeyArray_S10reg_gff_1_SFF_2_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_3604, new_AGEMA_signal_3603, new_AGEMA_signal_3602, KeyArray_inS10ser[2]}), .a ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, new_AGEMA_signal_3815, KeyArray_outS20ser[2]}), .c ({new_AGEMA_signal_4780, new_AGEMA_signal_4779, new_AGEMA_signal_4778, KeyArray_S10reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_3_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_3538, new_AGEMA_signal_3537, new_AGEMA_signal_3536, KeyArray_outS10ser[3]}), .a ({new_AGEMA_signal_4783, new_AGEMA_signal_4782, new_AGEMA_signal_4781, KeyArray_S10reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_5944, new_AGEMA_signal_5943, new_AGEMA_signal_5942, KeyArray_S10reg_gff_1_SFF_3_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, new_AGEMA_signal_3611, KeyArray_inS10ser[3]}), .a ({new_AGEMA_signal_3826, new_AGEMA_signal_3825, new_AGEMA_signal_3824, KeyArray_outS20ser[3]}), .c ({new_AGEMA_signal_4783, new_AGEMA_signal_4782, new_AGEMA_signal_4781, KeyArray_S10reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_4_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_3547, new_AGEMA_signal_3546, new_AGEMA_signal_3545, KeyArray_outS10ser[4]}), .a ({new_AGEMA_signal_4786, new_AGEMA_signal_4785, new_AGEMA_signal_4784, KeyArray_S10reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_5947, new_AGEMA_signal_5946, new_AGEMA_signal_5945, KeyArray_S10reg_gff_1_SFF_4_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_3622, new_AGEMA_signal_3621, new_AGEMA_signal_3620, KeyArray_inS10ser[4]}), .a ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, new_AGEMA_signal_3833, KeyArray_outS20ser[4]}), .c ({new_AGEMA_signal_4786, new_AGEMA_signal_4785, new_AGEMA_signal_4784, KeyArray_S10reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_5_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_3556, new_AGEMA_signal_3555, new_AGEMA_signal_3554, KeyArray_outS10ser[5]}), .a ({new_AGEMA_signal_4789, new_AGEMA_signal_4788, new_AGEMA_signal_4787, KeyArray_S10reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_5950, new_AGEMA_signal_5949, new_AGEMA_signal_5948, KeyArray_S10reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_3631, new_AGEMA_signal_3630, new_AGEMA_signal_3629, KeyArray_inS10ser[5]}), .a ({new_AGEMA_signal_3844, new_AGEMA_signal_3843, new_AGEMA_signal_3842, KeyArray_outS20ser[5]}), .c ({new_AGEMA_signal_4789, new_AGEMA_signal_4788, new_AGEMA_signal_4787, KeyArray_S10reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_6_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, new_AGEMA_signal_3563, KeyArray_outS10ser[6]}), .a ({new_AGEMA_signal_4792, new_AGEMA_signal_4791, new_AGEMA_signal_4790, KeyArray_S10reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_5953, new_AGEMA_signal_5952, new_AGEMA_signal_5951, KeyArray_S10reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_3640, new_AGEMA_signal_3639, new_AGEMA_signal_3638, KeyArray_inS10ser[6]}), .a ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, new_AGEMA_signal_3851, KeyArray_outS20ser[6]}), .c ({new_AGEMA_signal_4792, new_AGEMA_signal_4791, new_AGEMA_signal_4790, KeyArray_S10reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_7_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_3574, new_AGEMA_signal_3573, new_AGEMA_signal_3572, KeyArray_outS10ser[7]}), .a ({new_AGEMA_signal_4795, new_AGEMA_signal_4794, new_AGEMA_signal_4793, KeyArray_S10reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_5956, new_AGEMA_signal_5955, new_AGEMA_signal_5954, KeyArray_S10reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_3649, new_AGEMA_signal_3648, new_AGEMA_signal_3647, KeyArray_inS10ser[7]}), .a ({new_AGEMA_signal_3862, new_AGEMA_signal_3861, new_AGEMA_signal_3860, KeyArray_outS20ser[7]}), .c ({new_AGEMA_signal_4795, new_AGEMA_signal_4794, new_AGEMA_signal_4793, KeyArray_S10reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_0_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, new_AGEMA_signal_3581, KeyArray_outS11ser[0]}), .a ({new_AGEMA_signal_4798, new_AGEMA_signal_4797, new_AGEMA_signal_4796, KeyArray_S11reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_5959, new_AGEMA_signal_5958, new_AGEMA_signal_5957, KeyArray_S11reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_3658, new_AGEMA_signal_3657, new_AGEMA_signal_3656, KeyArray_inS11ser[0]}), .a ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, new_AGEMA_signal_3869, KeyArray_outS21ser[0]}), .c ({new_AGEMA_signal_4798, new_AGEMA_signal_4797, new_AGEMA_signal_4796, KeyArray_S11reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_1_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_3592, new_AGEMA_signal_3591, new_AGEMA_signal_3590, KeyArray_outS11ser[1]}), .a ({new_AGEMA_signal_4801, new_AGEMA_signal_4800, new_AGEMA_signal_4799, KeyArray_S11reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_5962, new_AGEMA_signal_5961, new_AGEMA_signal_5960, KeyArray_S11reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_3667, new_AGEMA_signal_3666, new_AGEMA_signal_3665, KeyArray_inS11ser[1]}), .a ({new_AGEMA_signal_3880, new_AGEMA_signal_3879, new_AGEMA_signal_3878, KeyArray_outS21ser[1]}), .c ({new_AGEMA_signal_4801, new_AGEMA_signal_4800, new_AGEMA_signal_4799, KeyArray_S11reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_2_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, new_AGEMA_signal_3599, KeyArray_outS11ser[2]}), .a ({new_AGEMA_signal_4804, new_AGEMA_signal_4803, new_AGEMA_signal_4802, KeyArray_S11reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_5965, new_AGEMA_signal_5964, new_AGEMA_signal_5963, KeyArray_S11reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_3676, new_AGEMA_signal_3675, new_AGEMA_signal_3674, KeyArray_inS11ser[2]}), .a ({new_AGEMA_signal_3889, new_AGEMA_signal_3888, new_AGEMA_signal_3887, KeyArray_outS21ser[2]}), .c ({new_AGEMA_signal_4804, new_AGEMA_signal_4803, new_AGEMA_signal_4802, KeyArray_S11reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_3_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_3610, new_AGEMA_signal_3609, new_AGEMA_signal_3608, KeyArray_outS11ser[3]}), .a ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, new_AGEMA_signal_4805, KeyArray_S11reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_5968, new_AGEMA_signal_5967, new_AGEMA_signal_5966, KeyArray_S11reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_3685, new_AGEMA_signal_3684, new_AGEMA_signal_3683, KeyArray_inS11ser[3]}), .a ({new_AGEMA_signal_3898, new_AGEMA_signal_3897, new_AGEMA_signal_3896, KeyArray_outS21ser[3]}), .c ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, new_AGEMA_signal_4805, KeyArray_S11reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_4_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_3619, new_AGEMA_signal_3618, new_AGEMA_signal_3617, KeyArray_outS11ser[4]}), .a ({new_AGEMA_signal_4810, new_AGEMA_signal_4809, new_AGEMA_signal_4808, KeyArray_S11reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_5971, new_AGEMA_signal_5970, new_AGEMA_signal_5969, KeyArray_S11reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_3694, new_AGEMA_signal_3693, new_AGEMA_signal_3692, KeyArray_inS11ser[4]}), .a ({new_AGEMA_signal_3907, new_AGEMA_signal_3906, new_AGEMA_signal_3905, KeyArray_outS21ser[4]}), .c ({new_AGEMA_signal_4810, new_AGEMA_signal_4809, new_AGEMA_signal_4808, KeyArray_S11reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_5_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_3628, new_AGEMA_signal_3627, new_AGEMA_signal_3626, KeyArray_outS11ser[5]}), .a ({new_AGEMA_signal_4813, new_AGEMA_signal_4812, new_AGEMA_signal_4811, KeyArray_S11reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_5974, new_AGEMA_signal_5973, new_AGEMA_signal_5972, KeyArray_S11reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_3703, new_AGEMA_signal_3702, new_AGEMA_signal_3701, KeyArray_inS11ser[5]}), .a ({new_AGEMA_signal_3916, new_AGEMA_signal_3915, new_AGEMA_signal_3914, KeyArray_outS21ser[5]}), .c ({new_AGEMA_signal_4813, new_AGEMA_signal_4812, new_AGEMA_signal_4811, KeyArray_S11reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_6_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, new_AGEMA_signal_3635, KeyArray_outS11ser[6]}), .a ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, new_AGEMA_signal_4814, KeyArray_S11reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_5977, new_AGEMA_signal_5976, new_AGEMA_signal_5975, KeyArray_S11reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_3712, new_AGEMA_signal_3711, new_AGEMA_signal_3710, KeyArray_inS11ser[6]}), .a ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, new_AGEMA_signal_3923, KeyArray_outS21ser[6]}), .c ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, new_AGEMA_signal_4814, KeyArray_S11reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_7_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_3646, new_AGEMA_signal_3645, new_AGEMA_signal_3644, KeyArray_outS11ser[7]}), .a ({new_AGEMA_signal_4819, new_AGEMA_signal_4818, new_AGEMA_signal_4817, KeyArray_S11reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_5980, new_AGEMA_signal_5979, new_AGEMA_signal_5978, KeyArray_S11reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_3721, new_AGEMA_signal_3720, new_AGEMA_signal_3719, KeyArray_inS11ser[7]}), .a ({new_AGEMA_signal_3934, new_AGEMA_signal_3933, new_AGEMA_signal_3932, KeyArray_outS21ser[7]}), .c ({new_AGEMA_signal_4819, new_AGEMA_signal_4818, new_AGEMA_signal_4817, KeyArray_S11reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_0_U1 ( .s (n12), .b ({new_AGEMA_signal_3655, new_AGEMA_signal_3654, new_AGEMA_signal_3653, KeyArray_outS12ser[0]}), .a ({new_AGEMA_signal_4822, new_AGEMA_signal_4821, new_AGEMA_signal_4820, KeyArray_S12reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_5317, new_AGEMA_signal_5316, new_AGEMA_signal_5315, KeyArray_S12reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_3730, new_AGEMA_signal_3729, new_AGEMA_signal_3728, KeyArray_inS12ser[0]}), .a ({new_AGEMA_signal_3943, new_AGEMA_signal_3942, new_AGEMA_signal_3941, KeyArray_outS22ser[0]}), .c ({new_AGEMA_signal_4822, new_AGEMA_signal_4821, new_AGEMA_signal_4820, KeyArray_S12reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_1_U1 ( .s (n12), .b ({new_AGEMA_signal_3664, new_AGEMA_signal_3663, new_AGEMA_signal_3662, KeyArray_outS12ser[1]}), .a ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, new_AGEMA_signal_4823, KeyArray_S12reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_5320, new_AGEMA_signal_5319, new_AGEMA_signal_5318, KeyArray_S12reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_3739, new_AGEMA_signal_3738, new_AGEMA_signal_3737, KeyArray_inS12ser[1]}), .a ({new_AGEMA_signal_3952, new_AGEMA_signal_3951, new_AGEMA_signal_3950, KeyArray_outS22ser[1]}), .c ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, new_AGEMA_signal_4823, KeyArray_S12reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_2_U1 ( .s (n12), .b ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, new_AGEMA_signal_3671, KeyArray_outS12ser[2]}), .a ({new_AGEMA_signal_4828, new_AGEMA_signal_4827, new_AGEMA_signal_4826, KeyArray_S12reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_5323, new_AGEMA_signal_5322, new_AGEMA_signal_5321, KeyArray_S12reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_3748, new_AGEMA_signal_3747, new_AGEMA_signal_3746, KeyArray_inS12ser[2]}), .a ({new_AGEMA_signal_3961, new_AGEMA_signal_3960, new_AGEMA_signal_3959, KeyArray_outS22ser[2]}), .c ({new_AGEMA_signal_4828, new_AGEMA_signal_4827, new_AGEMA_signal_4826, KeyArray_S12reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_3_U1 ( .s (n12), .b ({new_AGEMA_signal_3682, new_AGEMA_signal_3681, new_AGEMA_signal_3680, KeyArray_outS12ser[3]}), .a ({new_AGEMA_signal_4831, new_AGEMA_signal_4830, new_AGEMA_signal_4829, KeyArray_S12reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_5326, new_AGEMA_signal_5325, new_AGEMA_signal_5324, KeyArray_S12reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, new_AGEMA_signal_3755, KeyArray_inS12ser[3]}), .a ({new_AGEMA_signal_3970, new_AGEMA_signal_3969, new_AGEMA_signal_3968, KeyArray_outS22ser[3]}), .c ({new_AGEMA_signal_4831, new_AGEMA_signal_4830, new_AGEMA_signal_4829, KeyArray_S12reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_4_U1 ( .s (n12), .b ({new_AGEMA_signal_3691, new_AGEMA_signal_3690, new_AGEMA_signal_3689, KeyArray_outS12ser[4]}), .a ({new_AGEMA_signal_4834, new_AGEMA_signal_4833, new_AGEMA_signal_4832, KeyArray_S12reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_5329, new_AGEMA_signal_5328, new_AGEMA_signal_5327, KeyArray_S12reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_3766, new_AGEMA_signal_3765, new_AGEMA_signal_3764, KeyArray_inS12ser[4]}), .a ({new_AGEMA_signal_3979, new_AGEMA_signal_3978, new_AGEMA_signal_3977, KeyArray_outS22ser[4]}), .c ({new_AGEMA_signal_4834, new_AGEMA_signal_4833, new_AGEMA_signal_4832, KeyArray_S12reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_5_U1 ( .s (n12), .b ({new_AGEMA_signal_3700, new_AGEMA_signal_3699, new_AGEMA_signal_3698, KeyArray_outS12ser[5]}), .a ({new_AGEMA_signal_4837, new_AGEMA_signal_4836, new_AGEMA_signal_4835, KeyArray_S12reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_5332, new_AGEMA_signal_5331, new_AGEMA_signal_5330, KeyArray_S12reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, new_AGEMA_signal_3773, KeyArray_inS12ser[5]}), .a ({new_AGEMA_signal_3988, new_AGEMA_signal_3987, new_AGEMA_signal_3986, KeyArray_outS22ser[5]}), .c ({new_AGEMA_signal_4837, new_AGEMA_signal_4836, new_AGEMA_signal_4835, KeyArray_S12reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_6_U1 ( .s (n12), .b ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, new_AGEMA_signal_3707, KeyArray_outS12ser[6]}), .a ({new_AGEMA_signal_4840, new_AGEMA_signal_4839, new_AGEMA_signal_4838, KeyArray_S12reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_5335, new_AGEMA_signal_5334, new_AGEMA_signal_5333, KeyArray_S12reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_3784, new_AGEMA_signal_3783, new_AGEMA_signal_3782, KeyArray_inS12ser[6]}), .a ({new_AGEMA_signal_3997, new_AGEMA_signal_3996, new_AGEMA_signal_3995, KeyArray_outS22ser[6]}), .c ({new_AGEMA_signal_4840, new_AGEMA_signal_4839, new_AGEMA_signal_4838, KeyArray_S12reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_7_U1 ( .s (n12), .b ({new_AGEMA_signal_3718, new_AGEMA_signal_3717, new_AGEMA_signal_3716, KeyArray_outS12ser[7]}), .a ({new_AGEMA_signal_4843, new_AGEMA_signal_4842, new_AGEMA_signal_4841, KeyArray_S12reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_5338, new_AGEMA_signal_5337, new_AGEMA_signal_5336, KeyArray_S12reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, new_AGEMA_signal_3791, KeyArray_inS12ser[7]}), .a ({new_AGEMA_signal_4006, new_AGEMA_signal_4005, new_AGEMA_signal_4004, KeyArray_outS22ser[7]}), .c ({new_AGEMA_signal_4843, new_AGEMA_signal_4842, new_AGEMA_signal_4841, KeyArray_S12reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_0_U1 ( .s (n12), .b ({new_AGEMA_signal_3727, new_AGEMA_signal_3726, new_AGEMA_signal_3725, keySBIn[0]}), .a ({new_AGEMA_signal_4846, new_AGEMA_signal_4845, new_AGEMA_signal_4844, KeyArray_S13reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_5341, new_AGEMA_signal_5340, new_AGEMA_signal_5339, KeyArray_S13reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_3802, new_AGEMA_signal_3801, new_AGEMA_signal_3800, KeyArray_inS13ser[0]}), .a ({new_AGEMA_signal_4015, new_AGEMA_signal_4014, new_AGEMA_signal_4013, KeyArray_outS23ser[0]}), .c ({new_AGEMA_signal_4846, new_AGEMA_signal_4845, new_AGEMA_signal_4844, KeyArray_S13reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_1_U1 ( .s (n12), .b ({new_AGEMA_signal_3736, new_AGEMA_signal_3735, new_AGEMA_signal_3734, keySBIn[1]}), .a ({new_AGEMA_signal_4849, new_AGEMA_signal_4848, new_AGEMA_signal_4847, KeyArray_S13reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_5344, new_AGEMA_signal_5343, new_AGEMA_signal_5342, KeyArray_S13reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, new_AGEMA_signal_3809, KeyArray_inS13ser[1]}), .a ({new_AGEMA_signal_4024, new_AGEMA_signal_4023, new_AGEMA_signal_4022, KeyArray_outS23ser[1]}), .c ({new_AGEMA_signal_4849, new_AGEMA_signal_4848, new_AGEMA_signal_4847, KeyArray_S13reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_2_U1 ( .s (n12), .b ({new_AGEMA_signal_3745, new_AGEMA_signal_3744, new_AGEMA_signal_3743, keySBIn[2]}), .a ({new_AGEMA_signal_4852, new_AGEMA_signal_4851, new_AGEMA_signal_4850, KeyArray_S13reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_5347, new_AGEMA_signal_5346, new_AGEMA_signal_5345, KeyArray_S13reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_3820, new_AGEMA_signal_3819, new_AGEMA_signal_3818, KeyArray_inS13ser[2]}), .a ({new_AGEMA_signal_4033, new_AGEMA_signal_4032, new_AGEMA_signal_4031, KeyArray_outS23ser[2]}), .c ({new_AGEMA_signal_4852, new_AGEMA_signal_4851, new_AGEMA_signal_4850, KeyArray_S13reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_3_U1 ( .s (n12), .b ({new_AGEMA_signal_3754, new_AGEMA_signal_3753, new_AGEMA_signal_3752, keySBIn[3]}), .a ({new_AGEMA_signal_4855, new_AGEMA_signal_4854, new_AGEMA_signal_4853, KeyArray_S13reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_5350, new_AGEMA_signal_5349, new_AGEMA_signal_5348, KeyArray_S13reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, new_AGEMA_signal_3827, KeyArray_inS13ser[3]}), .a ({new_AGEMA_signal_4042, new_AGEMA_signal_4041, new_AGEMA_signal_4040, KeyArray_outS23ser[3]}), .c ({new_AGEMA_signal_4855, new_AGEMA_signal_4854, new_AGEMA_signal_4853, KeyArray_S13reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_4_U1 ( .s (n12), .b ({new_AGEMA_signal_3763, new_AGEMA_signal_3762, new_AGEMA_signal_3761, keySBIn[4]}), .a ({new_AGEMA_signal_4858, new_AGEMA_signal_4857, new_AGEMA_signal_4856, KeyArray_S13reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_5353, new_AGEMA_signal_5352, new_AGEMA_signal_5351, KeyArray_S13reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_3838, new_AGEMA_signal_3837, new_AGEMA_signal_3836, KeyArray_inS13ser[4]}), .a ({new_AGEMA_signal_4051, new_AGEMA_signal_4050, new_AGEMA_signal_4049, KeyArray_outS23ser[4]}), .c ({new_AGEMA_signal_4858, new_AGEMA_signal_4857, new_AGEMA_signal_4856, KeyArray_S13reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_5_U1 ( .s (n12), .b ({new_AGEMA_signal_3772, new_AGEMA_signal_3771, new_AGEMA_signal_3770, keySBIn[5]}), .a ({new_AGEMA_signal_4861, new_AGEMA_signal_4860, new_AGEMA_signal_4859, KeyArray_S13reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_5356, new_AGEMA_signal_5355, new_AGEMA_signal_5354, KeyArray_S13reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_3847, new_AGEMA_signal_3846, new_AGEMA_signal_3845, KeyArray_inS13ser[5]}), .a ({new_AGEMA_signal_4060, new_AGEMA_signal_4059, new_AGEMA_signal_4058, KeyArray_outS23ser[5]}), .c ({new_AGEMA_signal_4861, new_AGEMA_signal_4860, new_AGEMA_signal_4859, KeyArray_S13reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_6_U1 ( .s (n12), .b ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, new_AGEMA_signal_3779, keySBIn[6]}), .a ({new_AGEMA_signal_4864, new_AGEMA_signal_4863, new_AGEMA_signal_4862, KeyArray_S13reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_5359, new_AGEMA_signal_5358, new_AGEMA_signal_5357, KeyArray_S13reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_3856, new_AGEMA_signal_3855, new_AGEMA_signal_3854, KeyArray_inS13ser[6]}), .a ({new_AGEMA_signal_4069, new_AGEMA_signal_4068, new_AGEMA_signal_4067, KeyArray_outS23ser[6]}), .c ({new_AGEMA_signal_4864, new_AGEMA_signal_4863, new_AGEMA_signal_4862, KeyArray_S13reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_7_U1 ( .s (n12), .b ({new_AGEMA_signal_3790, new_AGEMA_signal_3789, new_AGEMA_signal_3788, keySBIn[7]}), .a ({new_AGEMA_signal_4867, new_AGEMA_signal_4866, new_AGEMA_signal_4865, KeyArray_S13reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_5362, new_AGEMA_signal_5361, new_AGEMA_signal_5360, KeyArray_S13reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_3865, new_AGEMA_signal_3864, new_AGEMA_signal_3863, KeyArray_inS13ser[7]}), .a ({new_AGEMA_signal_4078, new_AGEMA_signal_4077, new_AGEMA_signal_4076, KeyArray_outS23ser[7]}), .c ({new_AGEMA_signal_4867, new_AGEMA_signal_4866, new_AGEMA_signal_4865, KeyArray_S13reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_0_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, new_AGEMA_signal_3797, KeyArray_outS20ser[0]}), .a ({new_AGEMA_signal_4870, new_AGEMA_signal_4869, new_AGEMA_signal_4868, KeyArray_S20reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_5983, new_AGEMA_signal_5982, new_AGEMA_signal_5981, KeyArray_S20reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_3874, new_AGEMA_signal_3873, new_AGEMA_signal_3872, KeyArray_inS20ser[0]}), .a ({new_AGEMA_signal_4087, new_AGEMA_signal_4086, new_AGEMA_signal_4085, KeyArray_outS30ser[0]}), .c ({new_AGEMA_signal_4870, new_AGEMA_signal_4869, new_AGEMA_signal_4868, KeyArray_S20reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_1_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_3808, new_AGEMA_signal_3807, new_AGEMA_signal_3806, KeyArray_outS20ser[1]}), .a ({new_AGEMA_signal_4873, new_AGEMA_signal_4872, new_AGEMA_signal_4871, KeyArray_S20reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_5986, new_AGEMA_signal_5985, new_AGEMA_signal_5984, KeyArray_S20reg_gff_1_SFF_1_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, new_AGEMA_signal_3881, KeyArray_inS20ser[1]}), .a ({new_AGEMA_signal_4096, new_AGEMA_signal_4095, new_AGEMA_signal_4094, KeyArray_outS30ser[1]}), .c ({new_AGEMA_signal_4873, new_AGEMA_signal_4872, new_AGEMA_signal_4871, KeyArray_S20reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_2_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, new_AGEMA_signal_3815, KeyArray_outS20ser[2]}), .a ({new_AGEMA_signal_4876, new_AGEMA_signal_4875, new_AGEMA_signal_4874, KeyArray_S20reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_5989, new_AGEMA_signal_5988, new_AGEMA_signal_5987, KeyArray_S20reg_gff_1_SFF_2_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_3892, new_AGEMA_signal_3891, new_AGEMA_signal_3890, KeyArray_inS20ser[2]}), .a ({new_AGEMA_signal_4105, new_AGEMA_signal_4104, new_AGEMA_signal_4103, KeyArray_outS30ser[2]}), .c ({new_AGEMA_signal_4876, new_AGEMA_signal_4875, new_AGEMA_signal_4874, KeyArray_S20reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_3_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_3826, new_AGEMA_signal_3825, new_AGEMA_signal_3824, KeyArray_outS20ser[3]}), .a ({new_AGEMA_signal_4879, new_AGEMA_signal_4878, new_AGEMA_signal_4877, KeyArray_S20reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_5992, new_AGEMA_signal_5991, new_AGEMA_signal_5990, KeyArray_S20reg_gff_1_SFF_3_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_3901, new_AGEMA_signal_3900, new_AGEMA_signal_3899, KeyArray_inS20ser[3]}), .a ({new_AGEMA_signal_4114, new_AGEMA_signal_4113, new_AGEMA_signal_4112, KeyArray_outS30ser[3]}), .c ({new_AGEMA_signal_4879, new_AGEMA_signal_4878, new_AGEMA_signal_4877, KeyArray_S20reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_4_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, new_AGEMA_signal_3833, KeyArray_outS20ser[4]}), .a ({new_AGEMA_signal_4882, new_AGEMA_signal_4881, new_AGEMA_signal_4880, KeyArray_S20reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_5995, new_AGEMA_signal_5994, new_AGEMA_signal_5993, KeyArray_S20reg_gff_1_SFF_4_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_3910, new_AGEMA_signal_3909, new_AGEMA_signal_3908, KeyArray_inS20ser[4]}), .a ({new_AGEMA_signal_4123, new_AGEMA_signal_4122, new_AGEMA_signal_4121, KeyArray_outS30ser[4]}), .c ({new_AGEMA_signal_4882, new_AGEMA_signal_4881, new_AGEMA_signal_4880, KeyArray_S20reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_5_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_3844, new_AGEMA_signal_3843, new_AGEMA_signal_3842, KeyArray_outS20ser[5]}), .a ({new_AGEMA_signal_4885, new_AGEMA_signal_4884, new_AGEMA_signal_4883, KeyArray_S20reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_5998, new_AGEMA_signal_5997, new_AGEMA_signal_5996, KeyArray_S20reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_3919, new_AGEMA_signal_3918, new_AGEMA_signal_3917, KeyArray_inS20ser[5]}), .a ({new_AGEMA_signal_4132, new_AGEMA_signal_4131, new_AGEMA_signal_4130, KeyArray_outS30ser[5]}), .c ({new_AGEMA_signal_4885, new_AGEMA_signal_4884, new_AGEMA_signal_4883, KeyArray_S20reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_6_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, new_AGEMA_signal_3851, KeyArray_outS20ser[6]}), .a ({new_AGEMA_signal_4888, new_AGEMA_signal_4887, new_AGEMA_signal_4886, KeyArray_S20reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_6001, new_AGEMA_signal_6000, new_AGEMA_signal_5999, KeyArray_S20reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_3928, new_AGEMA_signal_3927, new_AGEMA_signal_3926, KeyArray_inS20ser[6]}), .a ({new_AGEMA_signal_4141, new_AGEMA_signal_4140, new_AGEMA_signal_4139, KeyArray_outS30ser[6]}), .c ({new_AGEMA_signal_4888, new_AGEMA_signal_4887, new_AGEMA_signal_4886, KeyArray_S20reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_7_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_3862, new_AGEMA_signal_3861, new_AGEMA_signal_3860, KeyArray_outS20ser[7]}), .a ({new_AGEMA_signal_4891, new_AGEMA_signal_4890, new_AGEMA_signal_4889, KeyArray_S20reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_6004, new_AGEMA_signal_6003, new_AGEMA_signal_6002, KeyArray_S20reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_3937, new_AGEMA_signal_3936, new_AGEMA_signal_3935, KeyArray_inS20ser[7]}), .a ({new_AGEMA_signal_4150, new_AGEMA_signal_4149, new_AGEMA_signal_4148, KeyArray_outS30ser[7]}), .c ({new_AGEMA_signal_4891, new_AGEMA_signal_4890, new_AGEMA_signal_4889, KeyArray_S20reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_0_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, new_AGEMA_signal_3869, KeyArray_outS21ser[0]}), .a ({new_AGEMA_signal_4894, new_AGEMA_signal_4893, new_AGEMA_signal_4892, KeyArray_S21reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_6007, new_AGEMA_signal_6006, new_AGEMA_signal_6005, KeyArray_S21reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_3946, new_AGEMA_signal_3945, new_AGEMA_signal_3944, KeyArray_inS21ser[0]}), .a ({new_AGEMA_signal_4159, new_AGEMA_signal_4158, new_AGEMA_signal_4157, KeyArray_outS31ser[0]}), .c ({new_AGEMA_signal_4894, new_AGEMA_signal_4893, new_AGEMA_signal_4892, KeyArray_S21reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_1_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_3880, new_AGEMA_signal_3879, new_AGEMA_signal_3878, KeyArray_outS21ser[1]}), .a ({new_AGEMA_signal_4897, new_AGEMA_signal_4896, new_AGEMA_signal_4895, KeyArray_S21reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_6010, new_AGEMA_signal_6009, new_AGEMA_signal_6008, KeyArray_S21reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_3955, new_AGEMA_signal_3954, new_AGEMA_signal_3953, KeyArray_inS21ser[1]}), .a ({new_AGEMA_signal_4168, new_AGEMA_signal_4167, new_AGEMA_signal_4166, KeyArray_outS31ser[1]}), .c ({new_AGEMA_signal_4897, new_AGEMA_signal_4896, new_AGEMA_signal_4895, KeyArray_S21reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_2_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_3889, new_AGEMA_signal_3888, new_AGEMA_signal_3887, KeyArray_outS21ser[2]}), .a ({new_AGEMA_signal_4900, new_AGEMA_signal_4899, new_AGEMA_signal_4898, KeyArray_S21reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_6013, new_AGEMA_signal_6012, new_AGEMA_signal_6011, KeyArray_S21reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_3964, new_AGEMA_signal_3963, new_AGEMA_signal_3962, KeyArray_inS21ser[2]}), .a ({new_AGEMA_signal_4177, new_AGEMA_signal_4176, new_AGEMA_signal_4175, KeyArray_outS31ser[2]}), .c ({new_AGEMA_signal_4900, new_AGEMA_signal_4899, new_AGEMA_signal_4898, KeyArray_S21reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_3_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_3898, new_AGEMA_signal_3897, new_AGEMA_signal_3896, KeyArray_outS21ser[3]}), .a ({new_AGEMA_signal_4903, new_AGEMA_signal_4902, new_AGEMA_signal_4901, KeyArray_S21reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_6016, new_AGEMA_signal_6015, new_AGEMA_signal_6014, KeyArray_S21reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_3973, new_AGEMA_signal_3972, new_AGEMA_signal_3971, KeyArray_inS21ser[3]}), .a ({new_AGEMA_signal_4186, new_AGEMA_signal_4185, new_AGEMA_signal_4184, KeyArray_outS31ser[3]}), .c ({new_AGEMA_signal_4903, new_AGEMA_signal_4902, new_AGEMA_signal_4901, KeyArray_S21reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_4_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_3907, new_AGEMA_signal_3906, new_AGEMA_signal_3905, KeyArray_outS21ser[4]}), .a ({new_AGEMA_signal_4906, new_AGEMA_signal_4905, new_AGEMA_signal_4904, KeyArray_S21reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_6019, new_AGEMA_signal_6018, new_AGEMA_signal_6017, KeyArray_S21reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_3982, new_AGEMA_signal_3981, new_AGEMA_signal_3980, KeyArray_inS21ser[4]}), .a ({new_AGEMA_signal_4195, new_AGEMA_signal_4194, new_AGEMA_signal_4193, KeyArray_outS31ser[4]}), .c ({new_AGEMA_signal_4906, new_AGEMA_signal_4905, new_AGEMA_signal_4904, KeyArray_S21reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_5_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_3916, new_AGEMA_signal_3915, new_AGEMA_signal_3914, KeyArray_outS21ser[5]}), .a ({new_AGEMA_signal_4909, new_AGEMA_signal_4908, new_AGEMA_signal_4907, KeyArray_S21reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_6022, new_AGEMA_signal_6021, new_AGEMA_signal_6020, KeyArray_S21reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_3991, new_AGEMA_signal_3990, new_AGEMA_signal_3989, KeyArray_inS21ser[5]}), .a ({new_AGEMA_signal_4204, new_AGEMA_signal_4203, new_AGEMA_signal_4202, KeyArray_outS31ser[5]}), .c ({new_AGEMA_signal_4909, new_AGEMA_signal_4908, new_AGEMA_signal_4907, KeyArray_S21reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_6_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, new_AGEMA_signal_3923, KeyArray_outS21ser[6]}), .a ({new_AGEMA_signal_4912, new_AGEMA_signal_4911, new_AGEMA_signal_4910, KeyArray_S21reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_6025, new_AGEMA_signal_6024, new_AGEMA_signal_6023, KeyArray_S21reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_4000, new_AGEMA_signal_3999, new_AGEMA_signal_3998, KeyArray_inS21ser[6]}), .a ({new_AGEMA_signal_4213, new_AGEMA_signal_4212, new_AGEMA_signal_4211, KeyArray_outS31ser[6]}), .c ({new_AGEMA_signal_4912, new_AGEMA_signal_4911, new_AGEMA_signal_4910, KeyArray_S21reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_7_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_3934, new_AGEMA_signal_3933, new_AGEMA_signal_3932, KeyArray_outS21ser[7]}), .a ({new_AGEMA_signal_4915, new_AGEMA_signal_4914, new_AGEMA_signal_4913, KeyArray_S21reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_6028, new_AGEMA_signal_6027, new_AGEMA_signal_6026, KeyArray_S21reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_4009, new_AGEMA_signal_4008, new_AGEMA_signal_4007, KeyArray_inS21ser[7]}), .a ({new_AGEMA_signal_4222, new_AGEMA_signal_4221, new_AGEMA_signal_4220, KeyArray_outS31ser[7]}), .c ({new_AGEMA_signal_4915, new_AGEMA_signal_4914, new_AGEMA_signal_4913, KeyArray_S21reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_0_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_3943, new_AGEMA_signal_3942, new_AGEMA_signal_3941, KeyArray_outS22ser[0]}), .a ({new_AGEMA_signal_4918, new_AGEMA_signal_4917, new_AGEMA_signal_4916, KeyArray_S22reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_6031, new_AGEMA_signal_6030, new_AGEMA_signal_6029, KeyArray_S22reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_4018, new_AGEMA_signal_4017, new_AGEMA_signal_4016, KeyArray_inS22ser[0]}), .a ({new_AGEMA_signal_4231, new_AGEMA_signal_4230, new_AGEMA_signal_4229, KeyArray_outS32ser[0]}), .c ({new_AGEMA_signal_4918, new_AGEMA_signal_4917, new_AGEMA_signal_4916, KeyArray_S22reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_1_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_3952, new_AGEMA_signal_3951, new_AGEMA_signal_3950, KeyArray_outS22ser[1]}), .a ({new_AGEMA_signal_4921, new_AGEMA_signal_4920, new_AGEMA_signal_4919, KeyArray_S22reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_6034, new_AGEMA_signal_6033, new_AGEMA_signal_6032, KeyArray_S22reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, new_AGEMA_signal_4025, KeyArray_inS22ser[1]}), .a ({new_AGEMA_signal_4240, new_AGEMA_signal_4239, new_AGEMA_signal_4238, KeyArray_outS32ser[1]}), .c ({new_AGEMA_signal_4921, new_AGEMA_signal_4920, new_AGEMA_signal_4919, KeyArray_S22reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_2_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_3961, new_AGEMA_signal_3960, new_AGEMA_signal_3959, KeyArray_outS22ser[2]}), .a ({new_AGEMA_signal_4924, new_AGEMA_signal_4923, new_AGEMA_signal_4922, KeyArray_S22reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_6037, new_AGEMA_signal_6036, new_AGEMA_signal_6035, KeyArray_S22reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_4036, new_AGEMA_signal_4035, new_AGEMA_signal_4034, KeyArray_inS22ser[2]}), .a ({new_AGEMA_signal_4249, new_AGEMA_signal_4248, new_AGEMA_signal_4247, KeyArray_outS32ser[2]}), .c ({new_AGEMA_signal_4924, new_AGEMA_signal_4923, new_AGEMA_signal_4922, KeyArray_S22reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_3_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_3970, new_AGEMA_signal_3969, new_AGEMA_signal_3968, KeyArray_outS22ser[3]}), .a ({new_AGEMA_signal_4927, new_AGEMA_signal_4926, new_AGEMA_signal_4925, KeyArray_S22reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_6040, new_AGEMA_signal_6039, new_AGEMA_signal_6038, KeyArray_S22reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, new_AGEMA_signal_4043, KeyArray_inS22ser[3]}), .a ({new_AGEMA_signal_4258, new_AGEMA_signal_4257, new_AGEMA_signal_4256, KeyArray_outS32ser[3]}), .c ({new_AGEMA_signal_4927, new_AGEMA_signal_4926, new_AGEMA_signal_4925, KeyArray_S22reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_4_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_3979, new_AGEMA_signal_3978, new_AGEMA_signal_3977, KeyArray_outS22ser[4]}), .a ({new_AGEMA_signal_4930, new_AGEMA_signal_4929, new_AGEMA_signal_4928, KeyArray_S22reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_6043, new_AGEMA_signal_6042, new_AGEMA_signal_6041, KeyArray_S22reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_4054, new_AGEMA_signal_4053, new_AGEMA_signal_4052, KeyArray_inS22ser[4]}), .a ({new_AGEMA_signal_4267, new_AGEMA_signal_4266, new_AGEMA_signal_4265, KeyArray_outS32ser[4]}), .c ({new_AGEMA_signal_4930, new_AGEMA_signal_4929, new_AGEMA_signal_4928, KeyArray_S22reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_5_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_3988, new_AGEMA_signal_3987, new_AGEMA_signal_3986, KeyArray_outS22ser[5]}), .a ({new_AGEMA_signal_4933, new_AGEMA_signal_4932, new_AGEMA_signal_4931, KeyArray_S22reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_6046, new_AGEMA_signal_6045, new_AGEMA_signal_6044, KeyArray_S22reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_4063, new_AGEMA_signal_4062, new_AGEMA_signal_4061, KeyArray_inS22ser[5]}), .a ({new_AGEMA_signal_4276, new_AGEMA_signal_4275, new_AGEMA_signal_4274, KeyArray_outS32ser[5]}), .c ({new_AGEMA_signal_4933, new_AGEMA_signal_4932, new_AGEMA_signal_4931, KeyArray_S22reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_6_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_3997, new_AGEMA_signal_3996, new_AGEMA_signal_3995, KeyArray_outS22ser[6]}), .a ({new_AGEMA_signal_4936, new_AGEMA_signal_4935, new_AGEMA_signal_4934, KeyArray_S22reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_6049, new_AGEMA_signal_6048, new_AGEMA_signal_6047, KeyArray_S22reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_4072, new_AGEMA_signal_4071, new_AGEMA_signal_4070, KeyArray_inS22ser[6]}), .a ({new_AGEMA_signal_4285, new_AGEMA_signal_4284, new_AGEMA_signal_4283, KeyArray_outS32ser[6]}), .c ({new_AGEMA_signal_4936, new_AGEMA_signal_4935, new_AGEMA_signal_4934, KeyArray_S22reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_7_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_4006, new_AGEMA_signal_4005, new_AGEMA_signal_4004, KeyArray_outS22ser[7]}), .a ({new_AGEMA_signal_4939, new_AGEMA_signal_4938, new_AGEMA_signal_4937, KeyArray_S22reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_6052, new_AGEMA_signal_6051, new_AGEMA_signal_6050, KeyArray_S22reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_4081, new_AGEMA_signal_4080, new_AGEMA_signal_4079, KeyArray_inS22ser[7]}), .a ({new_AGEMA_signal_4294, new_AGEMA_signal_4293, new_AGEMA_signal_4292, KeyArray_outS32ser[7]}), .c ({new_AGEMA_signal_4939, new_AGEMA_signal_4938, new_AGEMA_signal_4937, KeyArray_S22reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_0_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_4015, new_AGEMA_signal_4014, new_AGEMA_signal_4013, KeyArray_outS23ser[0]}), .a ({new_AGEMA_signal_4942, new_AGEMA_signal_4941, new_AGEMA_signal_4940, KeyArray_S23reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_6055, new_AGEMA_signal_6054, new_AGEMA_signal_6053, KeyArray_S23reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_4090, new_AGEMA_signal_4089, new_AGEMA_signal_4088, KeyArray_inS23ser[0]}), .a ({new_AGEMA_signal_4303, new_AGEMA_signal_4302, new_AGEMA_signal_4301, KeyArray_outS33ser[0]}), .c ({new_AGEMA_signal_4942, new_AGEMA_signal_4941, new_AGEMA_signal_4940, KeyArray_S23reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_1_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_4024, new_AGEMA_signal_4023, new_AGEMA_signal_4022, KeyArray_outS23ser[1]}), .a ({new_AGEMA_signal_4945, new_AGEMA_signal_4944, new_AGEMA_signal_4943, KeyArray_S23reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_6058, new_AGEMA_signal_6057, new_AGEMA_signal_6056, KeyArray_S23reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_4099, new_AGEMA_signal_4098, new_AGEMA_signal_4097, KeyArray_inS23ser[1]}), .a ({new_AGEMA_signal_4312, new_AGEMA_signal_4311, new_AGEMA_signal_4310, KeyArray_outS33ser[1]}), .c ({new_AGEMA_signal_4945, new_AGEMA_signal_4944, new_AGEMA_signal_4943, KeyArray_S23reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_2_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_4033, new_AGEMA_signal_4032, new_AGEMA_signal_4031, KeyArray_outS23ser[2]}), .a ({new_AGEMA_signal_4948, new_AGEMA_signal_4947, new_AGEMA_signal_4946, KeyArray_S23reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_6061, new_AGEMA_signal_6060, new_AGEMA_signal_6059, KeyArray_S23reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_4108, new_AGEMA_signal_4107, new_AGEMA_signal_4106, KeyArray_inS23ser[2]}), .a ({new_AGEMA_signal_4321, new_AGEMA_signal_4320, new_AGEMA_signal_4319, KeyArray_outS33ser[2]}), .c ({new_AGEMA_signal_4948, new_AGEMA_signal_4947, new_AGEMA_signal_4946, KeyArray_S23reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_3_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_4042, new_AGEMA_signal_4041, new_AGEMA_signal_4040, KeyArray_outS23ser[3]}), .a ({new_AGEMA_signal_4951, new_AGEMA_signal_4950, new_AGEMA_signal_4949, KeyArray_S23reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_6064, new_AGEMA_signal_6063, new_AGEMA_signal_6062, KeyArray_S23reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_4117, new_AGEMA_signal_4116, new_AGEMA_signal_4115, KeyArray_inS23ser[3]}), .a ({new_AGEMA_signal_4330, new_AGEMA_signal_4329, new_AGEMA_signal_4328, KeyArray_outS33ser[3]}), .c ({new_AGEMA_signal_4951, new_AGEMA_signal_4950, new_AGEMA_signal_4949, KeyArray_S23reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_4_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_4051, new_AGEMA_signal_4050, new_AGEMA_signal_4049, KeyArray_outS23ser[4]}), .a ({new_AGEMA_signal_4954, new_AGEMA_signal_4953, new_AGEMA_signal_4952, KeyArray_S23reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_6067, new_AGEMA_signal_6066, new_AGEMA_signal_6065, KeyArray_S23reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_4126, new_AGEMA_signal_4125, new_AGEMA_signal_4124, KeyArray_inS23ser[4]}), .a ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, new_AGEMA_signal_4337, KeyArray_outS33ser[4]}), .c ({new_AGEMA_signal_4954, new_AGEMA_signal_4953, new_AGEMA_signal_4952, KeyArray_S23reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_5_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_4060, new_AGEMA_signal_4059, new_AGEMA_signal_4058, KeyArray_outS23ser[5]}), .a ({new_AGEMA_signal_4957, new_AGEMA_signal_4956, new_AGEMA_signal_4955, KeyArray_S23reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_6070, new_AGEMA_signal_6069, new_AGEMA_signal_6068, KeyArray_S23reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_4135, new_AGEMA_signal_4134, new_AGEMA_signal_4133, KeyArray_inS23ser[5]}), .a ({new_AGEMA_signal_4348, new_AGEMA_signal_4347, new_AGEMA_signal_4346, KeyArray_outS33ser[5]}), .c ({new_AGEMA_signal_4957, new_AGEMA_signal_4956, new_AGEMA_signal_4955, KeyArray_S23reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_6_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_4069, new_AGEMA_signal_4068, new_AGEMA_signal_4067, KeyArray_outS23ser[6]}), .a ({new_AGEMA_signal_4960, new_AGEMA_signal_4959, new_AGEMA_signal_4958, KeyArray_S23reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_6073, new_AGEMA_signal_6072, new_AGEMA_signal_6071, KeyArray_S23reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_4144, new_AGEMA_signal_4143, new_AGEMA_signal_4142, KeyArray_inS23ser[6]}), .a ({new_AGEMA_signal_4357, new_AGEMA_signal_4356, new_AGEMA_signal_4355, KeyArray_outS33ser[6]}), .c ({new_AGEMA_signal_4960, new_AGEMA_signal_4959, new_AGEMA_signal_4958, KeyArray_S23reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_7_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_4078, new_AGEMA_signal_4077, new_AGEMA_signal_4076, KeyArray_outS23ser[7]}), .a ({new_AGEMA_signal_4963, new_AGEMA_signal_4962, new_AGEMA_signal_4961, KeyArray_S23reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_6076, new_AGEMA_signal_6075, new_AGEMA_signal_6074, KeyArray_S23reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_4153, new_AGEMA_signal_4152, new_AGEMA_signal_4151, KeyArray_inS23ser[7]}), .a ({new_AGEMA_signal_4366, new_AGEMA_signal_4365, new_AGEMA_signal_4364, KeyArray_outS33ser[7]}), .c ({new_AGEMA_signal_4963, new_AGEMA_signal_4962, new_AGEMA_signal_4961, KeyArray_S23reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_0_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_4159, new_AGEMA_signal_4158, new_AGEMA_signal_4157, KeyArray_outS31ser[0]}), .a ({new_AGEMA_signal_4966, new_AGEMA_signal_4965, new_AGEMA_signal_4964, KeyArray_S31reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_6079, new_AGEMA_signal_6078, new_AGEMA_signal_6077, KeyArray_S31reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_4234, new_AGEMA_signal_4233, new_AGEMA_signal_4232, KeyArray_inS31ser[0]}), .a ({new_AGEMA_signal_2098, new_AGEMA_signal_2097, new_AGEMA_signal_2096, KeyArray_outS01ser_0_}), .c ({new_AGEMA_signal_4966, new_AGEMA_signal_4965, new_AGEMA_signal_4964, KeyArray_S31reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_1_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_4168, new_AGEMA_signal_4167, new_AGEMA_signal_4166, KeyArray_outS31ser[1]}), .a ({new_AGEMA_signal_4969, new_AGEMA_signal_4968, new_AGEMA_signal_4967, KeyArray_S31reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_6082, new_AGEMA_signal_6081, new_AGEMA_signal_6080, KeyArray_S31reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_4243, new_AGEMA_signal_4242, new_AGEMA_signal_4241, KeyArray_inS31ser[1]}), .a ({new_AGEMA_signal_2092, new_AGEMA_signal_2091, new_AGEMA_signal_2090, KeyArray_outS01ser_1_}), .c ({new_AGEMA_signal_4969, new_AGEMA_signal_4968, new_AGEMA_signal_4967, KeyArray_S31reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_2_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_4177, new_AGEMA_signal_4176, new_AGEMA_signal_4175, KeyArray_outS31ser[2]}), .a ({new_AGEMA_signal_4972, new_AGEMA_signal_4971, new_AGEMA_signal_4970, KeyArray_S31reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_6085, new_AGEMA_signal_6084, new_AGEMA_signal_6083, KeyArray_S31reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_4252, new_AGEMA_signal_4251, new_AGEMA_signal_4250, KeyArray_inS31ser[2]}), .a ({new_AGEMA_signal_2086, new_AGEMA_signal_2085, new_AGEMA_signal_2084, KeyArray_outS01ser_2_}), .c ({new_AGEMA_signal_4972, new_AGEMA_signal_4971, new_AGEMA_signal_4970, KeyArray_S31reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_3_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_4186, new_AGEMA_signal_4185, new_AGEMA_signal_4184, KeyArray_outS31ser[3]}), .a ({new_AGEMA_signal_4975, new_AGEMA_signal_4974, new_AGEMA_signal_4973, KeyArray_S31reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_6088, new_AGEMA_signal_6087, new_AGEMA_signal_6086, KeyArray_S31reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_4261, new_AGEMA_signal_4260, new_AGEMA_signal_4259, KeyArray_inS31ser[3]}), .a ({new_AGEMA_signal_2080, new_AGEMA_signal_2079, new_AGEMA_signal_2078, KeyArray_outS01ser_3_}), .c ({new_AGEMA_signal_4975, new_AGEMA_signal_4974, new_AGEMA_signal_4973, KeyArray_S31reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_4_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_4195, new_AGEMA_signal_4194, new_AGEMA_signal_4193, KeyArray_outS31ser[4]}), .a ({new_AGEMA_signal_4978, new_AGEMA_signal_4977, new_AGEMA_signal_4976, KeyArray_S31reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_6091, new_AGEMA_signal_6090, new_AGEMA_signal_6089, KeyArray_S31reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_4270, new_AGEMA_signal_4269, new_AGEMA_signal_4268, KeyArray_inS31ser[4]}), .a ({new_AGEMA_signal_2074, new_AGEMA_signal_2073, new_AGEMA_signal_2072, KeyArray_outS01ser_4_}), .c ({new_AGEMA_signal_4978, new_AGEMA_signal_4977, new_AGEMA_signal_4976, KeyArray_S31reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_5_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_4204, new_AGEMA_signal_4203, new_AGEMA_signal_4202, KeyArray_outS31ser[5]}), .a ({new_AGEMA_signal_4981, new_AGEMA_signal_4980, new_AGEMA_signal_4979, KeyArray_S31reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_6094, new_AGEMA_signal_6093, new_AGEMA_signal_6092, KeyArray_S31reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_4279, new_AGEMA_signal_4278, new_AGEMA_signal_4277, KeyArray_inS31ser[5]}), .a ({new_AGEMA_signal_2068, new_AGEMA_signal_2067, new_AGEMA_signal_2066, KeyArray_outS01ser_5_}), .c ({new_AGEMA_signal_4981, new_AGEMA_signal_4980, new_AGEMA_signal_4979, KeyArray_S31reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_6_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_4213, new_AGEMA_signal_4212, new_AGEMA_signal_4211, KeyArray_outS31ser[6]}), .a ({new_AGEMA_signal_4984, new_AGEMA_signal_4983, new_AGEMA_signal_4982, KeyArray_S31reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_6097, new_AGEMA_signal_6096, new_AGEMA_signal_6095, KeyArray_S31reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_4288, new_AGEMA_signal_4287, new_AGEMA_signal_4286, KeyArray_inS31ser[6]}), .a ({new_AGEMA_signal_2062, new_AGEMA_signal_2061, new_AGEMA_signal_2060, KeyArray_outS01ser_6_}), .c ({new_AGEMA_signal_4984, new_AGEMA_signal_4983, new_AGEMA_signal_4982, KeyArray_S31reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_7_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_4222, new_AGEMA_signal_4221, new_AGEMA_signal_4220, KeyArray_outS31ser[7]}), .a ({new_AGEMA_signal_4987, new_AGEMA_signal_4986, new_AGEMA_signal_4985, KeyArray_S31reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_6100, new_AGEMA_signal_6099, new_AGEMA_signal_6098, KeyArray_S31reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_4297, new_AGEMA_signal_4296, new_AGEMA_signal_4295, KeyArray_inS31ser[7]}), .a ({new_AGEMA_signal_2056, new_AGEMA_signal_2055, new_AGEMA_signal_2054, KeyArray_outS01ser_7_}), .c ({new_AGEMA_signal_4987, new_AGEMA_signal_4986, new_AGEMA_signal_4985, KeyArray_S31reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_0_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_4231, new_AGEMA_signal_4230, new_AGEMA_signal_4229, KeyArray_outS32ser[0]}), .a ({new_AGEMA_signal_4990, new_AGEMA_signal_4989, new_AGEMA_signal_4988, KeyArray_S32reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_6103, new_AGEMA_signal_6102, new_AGEMA_signal_6101, KeyArray_S32reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_4306, new_AGEMA_signal_4305, new_AGEMA_signal_4304, KeyArray_inS32ser[0]}), .a ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, new_AGEMA_signal_3365, KeyArray_outS02ser[0]}), .c ({new_AGEMA_signal_4990, new_AGEMA_signal_4989, new_AGEMA_signal_4988, KeyArray_S32reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_1_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_4240, new_AGEMA_signal_4239, new_AGEMA_signal_4238, KeyArray_outS32ser[1]}), .a ({new_AGEMA_signal_4993, new_AGEMA_signal_4992, new_AGEMA_signal_4991, KeyArray_S32reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_6106, new_AGEMA_signal_6105, new_AGEMA_signal_6104, KeyArray_S32reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_4315, new_AGEMA_signal_4314, new_AGEMA_signal_4313, KeyArray_inS32ser[1]}), .a ({new_AGEMA_signal_3376, new_AGEMA_signal_3375, new_AGEMA_signal_3374, KeyArray_outS02ser[1]}), .c ({new_AGEMA_signal_4993, new_AGEMA_signal_4992, new_AGEMA_signal_4991, KeyArray_S32reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_2_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_4249, new_AGEMA_signal_4248, new_AGEMA_signal_4247, KeyArray_outS32ser[2]}), .a ({new_AGEMA_signal_4996, new_AGEMA_signal_4995, new_AGEMA_signal_4994, KeyArray_S32reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_6109, new_AGEMA_signal_6108, new_AGEMA_signal_6107, KeyArray_S32reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_4324, new_AGEMA_signal_4323, new_AGEMA_signal_4322, KeyArray_inS32ser[2]}), .a ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, new_AGEMA_signal_3383, KeyArray_outS02ser[2]}), .c ({new_AGEMA_signal_4996, new_AGEMA_signal_4995, new_AGEMA_signal_4994, KeyArray_S32reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_3_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_4258, new_AGEMA_signal_4257, new_AGEMA_signal_4256, KeyArray_outS32ser[3]}), .a ({new_AGEMA_signal_4999, new_AGEMA_signal_4998, new_AGEMA_signal_4997, KeyArray_S32reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_6112, new_AGEMA_signal_6111, new_AGEMA_signal_6110, KeyArray_S32reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_4333, new_AGEMA_signal_4332, new_AGEMA_signal_4331, KeyArray_inS32ser[3]}), .a ({new_AGEMA_signal_3394, new_AGEMA_signal_3393, new_AGEMA_signal_3392, KeyArray_outS02ser[3]}), .c ({new_AGEMA_signal_4999, new_AGEMA_signal_4998, new_AGEMA_signal_4997, KeyArray_S32reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_4_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_4267, new_AGEMA_signal_4266, new_AGEMA_signal_4265, KeyArray_outS32ser[4]}), .a ({new_AGEMA_signal_5002, new_AGEMA_signal_5001, new_AGEMA_signal_5000, KeyArray_S32reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_6115, new_AGEMA_signal_6114, new_AGEMA_signal_6113, KeyArray_S32reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_4342, new_AGEMA_signal_4341, new_AGEMA_signal_4340, KeyArray_inS32ser[4]}), .a ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, new_AGEMA_signal_3401, KeyArray_outS02ser[4]}), .c ({new_AGEMA_signal_5002, new_AGEMA_signal_5001, new_AGEMA_signal_5000, KeyArray_S32reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_5_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_4276, new_AGEMA_signal_4275, new_AGEMA_signal_4274, KeyArray_outS32ser[5]}), .a ({new_AGEMA_signal_5005, new_AGEMA_signal_5004, new_AGEMA_signal_5003, KeyArray_S32reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_6118, new_AGEMA_signal_6117, new_AGEMA_signal_6116, KeyArray_S32reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_4351, new_AGEMA_signal_4350, new_AGEMA_signal_4349, KeyArray_inS32ser[5]}), .a ({new_AGEMA_signal_3412, new_AGEMA_signal_3411, new_AGEMA_signal_3410, KeyArray_outS02ser[5]}), .c ({new_AGEMA_signal_5005, new_AGEMA_signal_5004, new_AGEMA_signal_5003, KeyArray_S32reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_6_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_4285, new_AGEMA_signal_4284, new_AGEMA_signal_4283, KeyArray_outS32ser[6]}), .a ({new_AGEMA_signal_5008, new_AGEMA_signal_5007, new_AGEMA_signal_5006, KeyArray_S32reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_6121, new_AGEMA_signal_6120, new_AGEMA_signal_6119, KeyArray_S32reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_4360, new_AGEMA_signal_4359, new_AGEMA_signal_4358, KeyArray_inS32ser[6]}), .a ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, new_AGEMA_signal_3419, KeyArray_outS02ser[6]}), .c ({new_AGEMA_signal_5008, new_AGEMA_signal_5007, new_AGEMA_signal_5006, KeyArray_S32reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_7_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_4294, new_AGEMA_signal_4293, new_AGEMA_signal_4292, KeyArray_outS32ser[7]}), .a ({new_AGEMA_signal_5011, new_AGEMA_signal_5010, new_AGEMA_signal_5009, KeyArray_S32reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_6124, new_AGEMA_signal_6123, new_AGEMA_signal_6122, KeyArray_S32reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_4369, new_AGEMA_signal_4368, new_AGEMA_signal_4367, KeyArray_inS32ser[7]}), .a ({new_AGEMA_signal_3430, new_AGEMA_signal_3429, new_AGEMA_signal_3428, KeyArray_outS02ser[7]}), .c ({new_AGEMA_signal_5011, new_AGEMA_signal_5010, new_AGEMA_signal_5009, KeyArray_S32reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_0_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_4303, new_AGEMA_signal_4302, new_AGEMA_signal_4301, KeyArray_outS33ser[0]}), .a ({new_AGEMA_signal_5014, new_AGEMA_signal_5013, new_AGEMA_signal_5012, KeyArray_S33reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_6127, new_AGEMA_signal_6126, new_AGEMA_signal_6125, KeyArray_S33reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_4375, new_AGEMA_signal_4374, new_AGEMA_signal_4373, KeyArray_inS33ser[0]}), .a ({new_AGEMA_signal_3439, new_AGEMA_signal_3438, new_AGEMA_signal_3437, KeyArray_outS03ser[0]}), .c ({new_AGEMA_signal_5014, new_AGEMA_signal_5013, new_AGEMA_signal_5012, KeyArray_S33reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_1_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_4312, new_AGEMA_signal_4311, new_AGEMA_signal_4310, KeyArray_outS33ser[1]}), .a ({new_AGEMA_signal_5017, new_AGEMA_signal_5016, new_AGEMA_signal_5015, KeyArray_S33reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_6130, new_AGEMA_signal_6129, new_AGEMA_signal_6128, KeyArray_S33reg_gff_1_SFF_1_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_4381, new_AGEMA_signal_4380, new_AGEMA_signal_4379, KeyArray_inS33ser[1]}), .a ({new_AGEMA_signal_3448, new_AGEMA_signal_3447, new_AGEMA_signal_3446, KeyArray_outS03ser[1]}), .c ({new_AGEMA_signal_5017, new_AGEMA_signal_5016, new_AGEMA_signal_5015, KeyArray_S33reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_2_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_4321, new_AGEMA_signal_4320, new_AGEMA_signal_4319, KeyArray_outS33ser[2]}), .a ({new_AGEMA_signal_5020, new_AGEMA_signal_5019, new_AGEMA_signal_5018, KeyArray_S33reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_6133, new_AGEMA_signal_6132, new_AGEMA_signal_6131, KeyArray_S33reg_gff_1_SFF_2_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_4387, new_AGEMA_signal_4386, new_AGEMA_signal_4385, KeyArray_inS33ser[2]}), .a ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, new_AGEMA_signal_3455, KeyArray_outS03ser[2]}), .c ({new_AGEMA_signal_5020, new_AGEMA_signal_5019, new_AGEMA_signal_5018, KeyArray_S33reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_3_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_4330, new_AGEMA_signal_4329, new_AGEMA_signal_4328, KeyArray_outS33ser[3]}), .a ({new_AGEMA_signal_5023, new_AGEMA_signal_5022, new_AGEMA_signal_5021, KeyArray_S33reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_6136, new_AGEMA_signal_6135, new_AGEMA_signal_6134, KeyArray_S33reg_gff_1_SFF_3_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_4393, new_AGEMA_signal_4392, new_AGEMA_signal_4391, KeyArray_inS33ser[3]}), .a ({new_AGEMA_signal_3466, new_AGEMA_signal_3465, new_AGEMA_signal_3464, KeyArray_outS03ser[3]}), .c ({new_AGEMA_signal_5023, new_AGEMA_signal_5022, new_AGEMA_signal_5021, KeyArray_S33reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_4_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, new_AGEMA_signal_4337, KeyArray_outS33ser[4]}), .a ({new_AGEMA_signal_5026, new_AGEMA_signal_5025, new_AGEMA_signal_5024, KeyArray_S33reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_6139, new_AGEMA_signal_6138, new_AGEMA_signal_6137, KeyArray_S33reg_gff_1_SFF_4_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_4399, new_AGEMA_signal_4398, new_AGEMA_signal_4397, KeyArray_inS33ser[4]}), .a ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, new_AGEMA_signal_3473, KeyArray_outS03ser[4]}), .c ({new_AGEMA_signal_5026, new_AGEMA_signal_5025, new_AGEMA_signal_5024, KeyArray_S33reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_5_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_4348, new_AGEMA_signal_4347, new_AGEMA_signal_4346, KeyArray_outS33ser[5]}), .a ({new_AGEMA_signal_5029, new_AGEMA_signal_5028, new_AGEMA_signal_5027, KeyArray_S33reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_6142, new_AGEMA_signal_6141, new_AGEMA_signal_6140, KeyArray_S33reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_4405, new_AGEMA_signal_4404, new_AGEMA_signal_4403, KeyArray_inS33ser[5]}), .a ({new_AGEMA_signal_3484, new_AGEMA_signal_3483, new_AGEMA_signal_3482, KeyArray_outS03ser[5]}), .c ({new_AGEMA_signal_5029, new_AGEMA_signal_5028, new_AGEMA_signal_5027, KeyArray_S33reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_6_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_4357, new_AGEMA_signal_4356, new_AGEMA_signal_4355, KeyArray_outS33ser[6]}), .a ({new_AGEMA_signal_5032, new_AGEMA_signal_5031, new_AGEMA_signal_5030, KeyArray_S33reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_6145, new_AGEMA_signal_6144, new_AGEMA_signal_6143, KeyArray_S33reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_4411, new_AGEMA_signal_4410, new_AGEMA_signal_4409, KeyArray_inS33ser[6]}), .a ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, new_AGEMA_signal_3491, KeyArray_outS03ser[6]}), .c ({new_AGEMA_signal_5032, new_AGEMA_signal_5031, new_AGEMA_signal_5030, KeyArray_S33reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_7_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_4366, new_AGEMA_signal_4365, new_AGEMA_signal_4364, KeyArray_outS33ser[7]}), .a ({new_AGEMA_signal_5035, new_AGEMA_signal_5034, new_AGEMA_signal_5033, KeyArray_S33reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_6148, new_AGEMA_signal_6147, new_AGEMA_signal_6146, KeyArray_S33reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_4417, new_AGEMA_signal_4416, new_AGEMA_signal_4415, KeyArray_inS33ser[7]}), .a ({new_AGEMA_signal_3502, new_AGEMA_signal_3501, new_AGEMA_signal_3500, KeyArray_outS03ser[7]}), .c ({new_AGEMA_signal_5035, new_AGEMA_signal_5034, new_AGEMA_signal_5033, KeyArray_S33reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_selXOR_mux_inst_0_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2098, new_AGEMA_signal_2097, new_AGEMA_signal_2096, KeyArray_outS01ser_0_}), .a ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, new_AGEMA_signal_2099, KeyArray_outS01ser_XOR_00[0]}), .c ({new_AGEMA_signal_5365, new_AGEMA_signal_5364, new_AGEMA_signal_5363, KeyArray_outS01ser_p[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_selXOR_mux_inst_1_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2092, new_AGEMA_signal_2091, new_AGEMA_signal_2090, KeyArray_outS01ser_1_}), .a ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, new_AGEMA_signal_2093, KeyArray_outS01ser_XOR_00[1]}), .c ({new_AGEMA_signal_5368, new_AGEMA_signal_5367, new_AGEMA_signal_5366, KeyArray_outS01ser_p[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_selXOR_mux_inst_2_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2086, new_AGEMA_signal_2085, new_AGEMA_signal_2084, KeyArray_outS01ser_2_}), .a ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, new_AGEMA_signal_2087, KeyArray_outS01ser_XOR_00[2]}), .c ({new_AGEMA_signal_5371, new_AGEMA_signal_5370, new_AGEMA_signal_5369, KeyArray_outS01ser_p[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_selXOR_mux_inst_3_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2080, new_AGEMA_signal_2079, new_AGEMA_signal_2078, KeyArray_outS01ser_3_}), .a ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, new_AGEMA_signal_2081, KeyArray_outS01ser_XOR_00[3]}), .c ({new_AGEMA_signal_5374, new_AGEMA_signal_5373, new_AGEMA_signal_5372, KeyArray_outS01ser_p[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_selXOR_mux_inst_4_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2074, new_AGEMA_signal_2073, new_AGEMA_signal_2072, KeyArray_outS01ser_4_}), .a ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, new_AGEMA_signal_2075, KeyArray_outS01ser_XOR_00[4]}), .c ({new_AGEMA_signal_5377, new_AGEMA_signal_5376, new_AGEMA_signal_5375, KeyArray_outS01ser_p[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_selXOR_mux_inst_5_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2068, new_AGEMA_signal_2067, new_AGEMA_signal_2066, KeyArray_outS01ser_5_}), .a ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, new_AGEMA_signal_2069, KeyArray_outS01ser_XOR_00[5]}), .c ({new_AGEMA_signal_5380, new_AGEMA_signal_5379, new_AGEMA_signal_5378, KeyArray_outS01ser_p[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_selXOR_mux_inst_6_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2062, new_AGEMA_signal_2061, new_AGEMA_signal_2060, KeyArray_outS01ser_6_}), .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, new_AGEMA_signal_2063, KeyArray_outS01ser_XOR_00[6]}), .c ({new_AGEMA_signal_5383, new_AGEMA_signal_5382, new_AGEMA_signal_5381, KeyArray_outS01ser_p[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_selXOR_mux_inst_7_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2056, new_AGEMA_signal_2055, new_AGEMA_signal_2054, KeyArray_outS01ser_7_}), .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, new_AGEMA_signal_2057, KeyArray_outS01ser_XOR_00[7]}), .c ({new_AGEMA_signal_5386, new_AGEMA_signal_5385, new_AGEMA_signal_5384, KeyArray_outS01ser_p[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS00ser_mux_inst_0_U1 ( .s (KeyArray_n46), .b ({key_s3[120], key_s2[120], key_s1[120], key_s0[120]}), .a ({new_AGEMA_signal_5365, new_AGEMA_signal_5364, new_AGEMA_signal_5363, KeyArray_outS01ser_p[0]}), .c ({new_AGEMA_signal_5779, new_AGEMA_signal_5778, new_AGEMA_signal_5777, KeyArray_inS00ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS00ser_mux_inst_1_U1 ( .s (KeyArray_n46), .b ({key_s3[121], key_s2[121], key_s1[121], key_s0[121]}), .a ({new_AGEMA_signal_5368, new_AGEMA_signal_5367, new_AGEMA_signal_5366, KeyArray_outS01ser_p[1]}), .c ({new_AGEMA_signal_5785, new_AGEMA_signal_5784, new_AGEMA_signal_5783, KeyArray_inS00ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS00ser_mux_inst_2_U1 ( .s (KeyArray_n46), .b ({key_s3[122], key_s2[122], key_s1[122], key_s0[122]}), .a ({new_AGEMA_signal_5371, new_AGEMA_signal_5370, new_AGEMA_signal_5369, KeyArray_outS01ser_p[2]}), .c ({new_AGEMA_signal_5791, new_AGEMA_signal_5790, new_AGEMA_signal_5789, KeyArray_inS00ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS00ser_mux_inst_3_U1 ( .s (KeyArray_n46), .b ({key_s3[123], key_s2[123], key_s1[123], key_s0[123]}), .a ({new_AGEMA_signal_5374, new_AGEMA_signal_5373, new_AGEMA_signal_5372, KeyArray_outS01ser_p[3]}), .c ({new_AGEMA_signal_5797, new_AGEMA_signal_5796, new_AGEMA_signal_5795, KeyArray_inS00ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS00ser_mux_inst_4_U1 ( .s (KeyArray_n46), .b ({key_s3[124], key_s2[124], key_s1[124], key_s0[124]}), .a ({new_AGEMA_signal_5377, new_AGEMA_signal_5376, new_AGEMA_signal_5375, KeyArray_outS01ser_p[4]}), .c ({new_AGEMA_signal_5803, new_AGEMA_signal_5802, new_AGEMA_signal_5801, KeyArray_inS00ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS00ser_mux_inst_5_U1 ( .s (KeyArray_n46), .b ({key_s3[125], key_s2[125], key_s1[125], key_s0[125]}), .a ({new_AGEMA_signal_5380, new_AGEMA_signal_5379, new_AGEMA_signal_5378, KeyArray_outS01ser_p[5]}), .c ({new_AGEMA_signal_5809, new_AGEMA_signal_5808, new_AGEMA_signal_5807, KeyArray_inS00ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS00ser_mux_inst_6_U1 ( .s (KeyArray_n46), .b ({key_s3[126], key_s2[126], key_s1[126], key_s0[126]}), .a ({new_AGEMA_signal_5383, new_AGEMA_signal_5382, new_AGEMA_signal_5381, KeyArray_outS01ser_p[6]}), .c ({new_AGEMA_signal_5815, new_AGEMA_signal_5814, new_AGEMA_signal_5813, KeyArray_inS00ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS00ser_mux_inst_7_U1 ( .s (KeyArray_n46), .b ({key_s3[127], key_s2[127], key_s1[127], key_s0[127]}), .a ({new_AGEMA_signal_5386, new_AGEMA_signal_5385, new_AGEMA_signal_5384, KeyArray_outS01ser_p[7]}), .c ({new_AGEMA_signal_5821, new_AGEMA_signal_5820, new_AGEMA_signal_5819, KeyArray_inS00ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS01ser_mux_inst_0_U1 ( .s (KeyArray_n46), .b ({key_s3[112], key_s2[112], key_s1[112], key_s0[112]}), .a ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, new_AGEMA_signal_3365, KeyArray_outS02ser[0]}), .c ({new_AGEMA_signal_3370, new_AGEMA_signal_3369, new_AGEMA_signal_3368, KeyArray_inS01ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS01ser_mux_inst_1_U1 ( .s (KeyArray_n46), .b ({key_s3[113], key_s2[113], key_s1[113], key_s0[113]}), .a ({new_AGEMA_signal_3376, new_AGEMA_signal_3375, new_AGEMA_signal_3374, KeyArray_outS02ser[1]}), .c ({new_AGEMA_signal_3379, new_AGEMA_signal_3378, new_AGEMA_signal_3377, KeyArray_inS01ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS01ser_mux_inst_2_U1 ( .s (KeyArray_n46), .b ({key_s3[114], key_s2[114], key_s1[114], key_s0[114]}), .a ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, new_AGEMA_signal_3383, KeyArray_outS02ser[2]}), .c ({new_AGEMA_signal_3388, new_AGEMA_signal_3387, new_AGEMA_signal_3386, KeyArray_inS01ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS01ser_mux_inst_3_U1 ( .s (KeyArray_n46), .b ({key_s3[115], key_s2[115], key_s1[115], key_s0[115]}), .a ({new_AGEMA_signal_3394, new_AGEMA_signal_3393, new_AGEMA_signal_3392, KeyArray_outS02ser[3]}), .c ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, new_AGEMA_signal_3395, KeyArray_inS01ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS01ser_mux_inst_4_U1 ( .s (KeyArray_n46), .b ({key_s3[116], key_s2[116], key_s1[116], key_s0[116]}), .a ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, new_AGEMA_signal_3401, KeyArray_outS02ser[4]}), .c ({new_AGEMA_signal_3406, new_AGEMA_signal_3405, new_AGEMA_signal_3404, KeyArray_inS01ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS01ser_mux_inst_5_U1 ( .s (KeyArray_n46), .b ({key_s3[117], key_s2[117], key_s1[117], key_s0[117]}), .a ({new_AGEMA_signal_3412, new_AGEMA_signal_3411, new_AGEMA_signal_3410, KeyArray_outS02ser[5]}), .c ({new_AGEMA_signal_3415, new_AGEMA_signal_3414, new_AGEMA_signal_3413, KeyArray_inS01ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS01ser_mux_inst_6_U1 ( .s (KeyArray_n46), .b ({key_s3[118], key_s2[118], key_s1[118], key_s0[118]}), .a ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, new_AGEMA_signal_3419, KeyArray_outS02ser[6]}), .c ({new_AGEMA_signal_3424, new_AGEMA_signal_3423, new_AGEMA_signal_3422, KeyArray_inS01ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS01ser_mux_inst_7_U1 ( .s (KeyArray_n46), .b ({key_s3[119], key_s2[119], key_s1[119], key_s0[119]}), .a ({new_AGEMA_signal_3430, new_AGEMA_signal_3429, new_AGEMA_signal_3428, KeyArray_outS02ser[7]}), .c ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, new_AGEMA_signal_3431, KeyArray_inS01ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS02ser_mux_inst_0_U1 ( .s (KeyArray_n45), .b ({key_s3[104], key_s2[104], key_s1[104], key_s0[104]}), .a ({new_AGEMA_signal_3439, new_AGEMA_signal_3438, new_AGEMA_signal_3437, KeyArray_outS03ser[0]}), .c ({new_AGEMA_signal_3442, new_AGEMA_signal_3441, new_AGEMA_signal_3440, KeyArray_inS02ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS02ser_mux_inst_1_U1 ( .s (KeyArray_n45), .b ({key_s3[105], key_s2[105], key_s1[105], key_s0[105]}), .a ({new_AGEMA_signal_3448, new_AGEMA_signal_3447, new_AGEMA_signal_3446, KeyArray_outS03ser[1]}), .c ({new_AGEMA_signal_3451, new_AGEMA_signal_3450, new_AGEMA_signal_3449, KeyArray_inS02ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS02ser_mux_inst_2_U1 ( .s (KeyArray_n45), .b ({key_s3[106], key_s2[106], key_s1[106], key_s0[106]}), .a ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, new_AGEMA_signal_3455, KeyArray_outS03ser[2]}), .c ({new_AGEMA_signal_3460, new_AGEMA_signal_3459, new_AGEMA_signal_3458, KeyArray_inS02ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS02ser_mux_inst_3_U1 ( .s (KeyArray_n45), .b ({key_s3[107], key_s2[107], key_s1[107], key_s0[107]}), .a ({new_AGEMA_signal_3466, new_AGEMA_signal_3465, new_AGEMA_signal_3464, KeyArray_outS03ser[3]}), .c ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, new_AGEMA_signal_3467, KeyArray_inS02ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS02ser_mux_inst_4_U1 ( .s (KeyArray_n45), .b ({key_s3[108], key_s2[108], key_s1[108], key_s0[108]}), .a ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, new_AGEMA_signal_3473, KeyArray_outS03ser[4]}), .c ({new_AGEMA_signal_3478, new_AGEMA_signal_3477, new_AGEMA_signal_3476, KeyArray_inS02ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS02ser_mux_inst_5_U1 ( .s (KeyArray_n45), .b ({key_s3[109], key_s2[109], key_s1[109], key_s0[109]}), .a ({new_AGEMA_signal_3484, new_AGEMA_signal_3483, new_AGEMA_signal_3482, KeyArray_outS03ser[5]}), .c ({new_AGEMA_signal_3487, new_AGEMA_signal_3486, new_AGEMA_signal_3485, KeyArray_inS02ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS02ser_mux_inst_6_U1 ( .s (KeyArray_n45), .b ({key_s3[110], key_s2[110], key_s1[110], key_s0[110]}), .a ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, new_AGEMA_signal_3491, KeyArray_outS03ser[6]}), .c ({new_AGEMA_signal_3496, new_AGEMA_signal_3495, new_AGEMA_signal_3494, KeyArray_inS02ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS02ser_mux_inst_7_U1 ( .s (KeyArray_n45), .b ({key_s3[111], key_s2[111], key_s1[111], key_s0[111]}), .a ({new_AGEMA_signal_3502, new_AGEMA_signal_3501, new_AGEMA_signal_3500, KeyArray_outS03ser[7]}), .c ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, new_AGEMA_signal_3503, KeyArray_inS02ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS03ser_mux_inst_0_U1 ( .s (KeyArray_n45), .b ({key_s3[96], key_s2[96], key_s1[96], key_s0[96]}), .a ({new_AGEMA_signal_3511, new_AGEMA_signal_3510, new_AGEMA_signal_3509, KeyArray_outS10ser[0]}), .c ({new_AGEMA_signal_3514, new_AGEMA_signal_3513, new_AGEMA_signal_3512, KeyArray_inS03ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS03ser_mux_inst_1_U1 ( .s (KeyArray_n45), .b ({key_s3[97], key_s2[97], key_s1[97], key_s0[97]}), .a ({new_AGEMA_signal_3520, new_AGEMA_signal_3519, new_AGEMA_signal_3518, KeyArray_outS10ser[1]}), .c ({new_AGEMA_signal_3523, new_AGEMA_signal_3522, new_AGEMA_signal_3521, KeyArray_inS03ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS03ser_mux_inst_2_U1 ( .s (KeyArray_n45), .b ({key_s3[98], key_s2[98], key_s1[98], key_s0[98]}), .a ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, new_AGEMA_signal_3527, KeyArray_outS10ser[2]}), .c ({new_AGEMA_signal_3532, new_AGEMA_signal_3531, new_AGEMA_signal_3530, KeyArray_inS03ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS03ser_mux_inst_3_U1 ( .s (KeyArray_n45), .b ({key_s3[99], key_s2[99], key_s1[99], key_s0[99]}), .a ({new_AGEMA_signal_3538, new_AGEMA_signal_3537, new_AGEMA_signal_3536, KeyArray_outS10ser[3]}), .c ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, new_AGEMA_signal_3539, KeyArray_inS03ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS03ser_mux_inst_4_U1 ( .s (KeyArray_n45), .b ({key_s3[100], key_s2[100], key_s1[100], key_s0[100]}), .a ({new_AGEMA_signal_3547, new_AGEMA_signal_3546, new_AGEMA_signal_3545, KeyArray_outS10ser[4]}), .c ({new_AGEMA_signal_3550, new_AGEMA_signal_3549, new_AGEMA_signal_3548, KeyArray_inS03ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS03ser_mux_inst_5_U1 ( .s (KeyArray_n45), .b ({key_s3[101], key_s2[101], key_s1[101], key_s0[101]}), .a ({new_AGEMA_signal_3556, new_AGEMA_signal_3555, new_AGEMA_signal_3554, KeyArray_outS10ser[5]}), .c ({new_AGEMA_signal_3559, new_AGEMA_signal_3558, new_AGEMA_signal_3557, KeyArray_inS03ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS03ser_mux_inst_6_U1 ( .s (KeyArray_n45), .b ({key_s3[102], key_s2[102], key_s1[102], key_s0[102]}), .a ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, new_AGEMA_signal_3563, KeyArray_outS10ser[6]}), .c ({new_AGEMA_signal_3568, new_AGEMA_signal_3567, new_AGEMA_signal_3566, KeyArray_inS03ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS03ser_mux_inst_7_U1 ( .s (KeyArray_n45), .b ({key_s3[103], key_s2[103], key_s1[103], key_s0[103]}), .a ({new_AGEMA_signal_3574, new_AGEMA_signal_3573, new_AGEMA_signal_3572, KeyArray_outS10ser[7]}), .c ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, new_AGEMA_signal_3575, KeyArray_inS03ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS10ser_mux_inst_0_U1 ( .s (KeyArray_n44), .b ({key_s3[88], key_s2[88], key_s1[88], key_s0[88]}), .a ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, new_AGEMA_signal_3581, KeyArray_outS11ser[0]}), .c ({new_AGEMA_signal_3586, new_AGEMA_signal_3585, new_AGEMA_signal_3584, KeyArray_inS10ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS10ser_mux_inst_1_U1 ( .s (KeyArray_n44), .b ({key_s3[89], key_s2[89], key_s1[89], key_s0[89]}), .a ({new_AGEMA_signal_3592, new_AGEMA_signal_3591, new_AGEMA_signal_3590, KeyArray_outS11ser[1]}), .c ({new_AGEMA_signal_3595, new_AGEMA_signal_3594, new_AGEMA_signal_3593, KeyArray_inS10ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS10ser_mux_inst_2_U1 ( .s (KeyArray_n44), .b ({key_s3[90], key_s2[90], key_s1[90], key_s0[90]}), .a ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, new_AGEMA_signal_3599, KeyArray_outS11ser[2]}), .c ({new_AGEMA_signal_3604, new_AGEMA_signal_3603, new_AGEMA_signal_3602, KeyArray_inS10ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS10ser_mux_inst_3_U1 ( .s (KeyArray_n44), .b ({key_s3[91], key_s2[91], key_s1[91], key_s0[91]}), .a ({new_AGEMA_signal_3610, new_AGEMA_signal_3609, new_AGEMA_signal_3608, KeyArray_outS11ser[3]}), .c ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, new_AGEMA_signal_3611, KeyArray_inS10ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS10ser_mux_inst_4_U1 ( .s (KeyArray_n44), .b ({key_s3[92], key_s2[92], key_s1[92], key_s0[92]}), .a ({new_AGEMA_signal_3619, new_AGEMA_signal_3618, new_AGEMA_signal_3617, KeyArray_outS11ser[4]}), .c ({new_AGEMA_signal_3622, new_AGEMA_signal_3621, new_AGEMA_signal_3620, KeyArray_inS10ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS10ser_mux_inst_5_U1 ( .s (KeyArray_n44), .b ({key_s3[93], key_s2[93], key_s1[93], key_s0[93]}), .a ({new_AGEMA_signal_3628, new_AGEMA_signal_3627, new_AGEMA_signal_3626, KeyArray_outS11ser[5]}), .c ({new_AGEMA_signal_3631, new_AGEMA_signal_3630, new_AGEMA_signal_3629, KeyArray_inS10ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS10ser_mux_inst_6_U1 ( .s (KeyArray_n44), .b ({key_s3[94], key_s2[94], key_s1[94], key_s0[94]}), .a ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, new_AGEMA_signal_3635, KeyArray_outS11ser[6]}), .c ({new_AGEMA_signal_3640, new_AGEMA_signal_3639, new_AGEMA_signal_3638, KeyArray_inS10ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS10ser_mux_inst_7_U1 ( .s (KeyArray_n44), .b ({key_s3[95], key_s2[95], key_s1[95], key_s0[95]}), .a ({new_AGEMA_signal_3646, new_AGEMA_signal_3645, new_AGEMA_signal_3644, KeyArray_outS11ser[7]}), .c ({new_AGEMA_signal_3649, new_AGEMA_signal_3648, new_AGEMA_signal_3647, KeyArray_inS10ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS11ser_mux_inst_0_U1 ( .s (KeyArray_n44), .b ({key_s3[80], key_s2[80], key_s1[80], key_s0[80]}), .a ({new_AGEMA_signal_3655, new_AGEMA_signal_3654, new_AGEMA_signal_3653, KeyArray_outS12ser[0]}), .c ({new_AGEMA_signal_3658, new_AGEMA_signal_3657, new_AGEMA_signal_3656, KeyArray_inS11ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS11ser_mux_inst_1_U1 ( .s (KeyArray_n44), .b ({key_s3[81], key_s2[81], key_s1[81], key_s0[81]}), .a ({new_AGEMA_signal_3664, new_AGEMA_signal_3663, new_AGEMA_signal_3662, KeyArray_outS12ser[1]}), .c ({new_AGEMA_signal_3667, new_AGEMA_signal_3666, new_AGEMA_signal_3665, KeyArray_inS11ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS11ser_mux_inst_2_U1 ( .s (KeyArray_n44), .b ({key_s3[82], key_s2[82], key_s1[82], key_s0[82]}), .a ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, new_AGEMA_signal_3671, KeyArray_outS12ser[2]}), .c ({new_AGEMA_signal_3676, new_AGEMA_signal_3675, new_AGEMA_signal_3674, KeyArray_inS11ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS11ser_mux_inst_3_U1 ( .s (KeyArray_n44), .b ({key_s3[83], key_s2[83], key_s1[83], key_s0[83]}), .a ({new_AGEMA_signal_3682, new_AGEMA_signal_3681, new_AGEMA_signal_3680, KeyArray_outS12ser[3]}), .c ({new_AGEMA_signal_3685, new_AGEMA_signal_3684, new_AGEMA_signal_3683, KeyArray_inS11ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS11ser_mux_inst_4_U1 ( .s (KeyArray_n44), .b ({key_s3[84], key_s2[84], key_s1[84], key_s0[84]}), .a ({new_AGEMA_signal_3691, new_AGEMA_signal_3690, new_AGEMA_signal_3689, KeyArray_outS12ser[4]}), .c ({new_AGEMA_signal_3694, new_AGEMA_signal_3693, new_AGEMA_signal_3692, KeyArray_inS11ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS11ser_mux_inst_5_U1 ( .s (KeyArray_n44), .b ({key_s3[85], key_s2[85], key_s1[85], key_s0[85]}), .a ({new_AGEMA_signal_3700, new_AGEMA_signal_3699, new_AGEMA_signal_3698, KeyArray_outS12ser[5]}), .c ({new_AGEMA_signal_3703, new_AGEMA_signal_3702, new_AGEMA_signal_3701, KeyArray_inS11ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS11ser_mux_inst_6_U1 ( .s (KeyArray_n44), .b ({key_s3[86], key_s2[86], key_s1[86], key_s0[86]}), .a ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, new_AGEMA_signal_3707, KeyArray_outS12ser[6]}), .c ({new_AGEMA_signal_3712, new_AGEMA_signal_3711, new_AGEMA_signal_3710, KeyArray_inS11ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS11ser_mux_inst_7_U1 ( .s (KeyArray_n44), .b ({key_s3[87], key_s2[87], key_s1[87], key_s0[87]}), .a ({new_AGEMA_signal_3718, new_AGEMA_signal_3717, new_AGEMA_signal_3716, KeyArray_outS12ser[7]}), .c ({new_AGEMA_signal_3721, new_AGEMA_signal_3720, new_AGEMA_signal_3719, KeyArray_inS11ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS12ser_mux_inst_0_U1 ( .s (KeyArray_n43), .b ({key_s3[72], key_s2[72], key_s1[72], key_s0[72]}), .a ({new_AGEMA_signal_3727, new_AGEMA_signal_3726, new_AGEMA_signal_3725, keySBIn[0]}), .c ({new_AGEMA_signal_3730, new_AGEMA_signal_3729, new_AGEMA_signal_3728, KeyArray_inS12ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS12ser_mux_inst_1_U1 ( .s (KeyArray_n43), .b ({key_s3[73], key_s2[73], key_s1[73], key_s0[73]}), .a ({new_AGEMA_signal_3736, new_AGEMA_signal_3735, new_AGEMA_signal_3734, keySBIn[1]}), .c ({new_AGEMA_signal_3739, new_AGEMA_signal_3738, new_AGEMA_signal_3737, KeyArray_inS12ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS12ser_mux_inst_2_U1 ( .s (KeyArray_n43), .b ({key_s3[74], key_s2[74], key_s1[74], key_s0[74]}), .a ({new_AGEMA_signal_3745, new_AGEMA_signal_3744, new_AGEMA_signal_3743, keySBIn[2]}), .c ({new_AGEMA_signal_3748, new_AGEMA_signal_3747, new_AGEMA_signal_3746, KeyArray_inS12ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS12ser_mux_inst_3_U1 ( .s (KeyArray_n43), .b ({key_s3[75], key_s2[75], key_s1[75], key_s0[75]}), .a ({new_AGEMA_signal_3754, new_AGEMA_signal_3753, new_AGEMA_signal_3752, keySBIn[3]}), .c ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, new_AGEMA_signal_3755, KeyArray_inS12ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS12ser_mux_inst_4_U1 ( .s (KeyArray_n43), .b ({key_s3[76], key_s2[76], key_s1[76], key_s0[76]}), .a ({new_AGEMA_signal_3763, new_AGEMA_signal_3762, new_AGEMA_signal_3761, keySBIn[4]}), .c ({new_AGEMA_signal_3766, new_AGEMA_signal_3765, new_AGEMA_signal_3764, KeyArray_inS12ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS12ser_mux_inst_5_U1 ( .s (KeyArray_n43), .b ({key_s3[77], key_s2[77], key_s1[77], key_s0[77]}), .a ({new_AGEMA_signal_3772, new_AGEMA_signal_3771, new_AGEMA_signal_3770, keySBIn[5]}), .c ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, new_AGEMA_signal_3773, KeyArray_inS12ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS12ser_mux_inst_6_U1 ( .s (KeyArray_n43), .b ({key_s3[78], key_s2[78], key_s1[78], key_s0[78]}), .a ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, new_AGEMA_signal_3779, keySBIn[6]}), .c ({new_AGEMA_signal_3784, new_AGEMA_signal_3783, new_AGEMA_signal_3782, KeyArray_inS12ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS12ser_mux_inst_7_U1 ( .s (KeyArray_n43), .b ({key_s3[79], key_s2[79], key_s1[79], key_s0[79]}), .a ({new_AGEMA_signal_3790, new_AGEMA_signal_3789, new_AGEMA_signal_3788, keySBIn[7]}), .c ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, new_AGEMA_signal_3791, KeyArray_inS12ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS13ser_mux_inst_0_U1 ( .s (KeyArray_n43), .b ({key_s3[64], key_s2[64], key_s1[64], key_s0[64]}), .a ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, new_AGEMA_signal_3797, KeyArray_outS20ser[0]}), .c ({new_AGEMA_signal_3802, new_AGEMA_signal_3801, new_AGEMA_signal_3800, KeyArray_inS13ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS13ser_mux_inst_1_U1 ( .s (KeyArray_n43), .b ({key_s3[65], key_s2[65], key_s1[65], key_s0[65]}), .a ({new_AGEMA_signal_3808, new_AGEMA_signal_3807, new_AGEMA_signal_3806, KeyArray_outS20ser[1]}), .c ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, new_AGEMA_signal_3809, KeyArray_inS13ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS13ser_mux_inst_2_U1 ( .s (KeyArray_n43), .b ({key_s3[66], key_s2[66], key_s1[66], key_s0[66]}), .a ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, new_AGEMA_signal_3815, KeyArray_outS20ser[2]}), .c ({new_AGEMA_signal_3820, new_AGEMA_signal_3819, new_AGEMA_signal_3818, KeyArray_inS13ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS13ser_mux_inst_3_U1 ( .s (KeyArray_n43), .b ({key_s3[67], key_s2[67], key_s1[67], key_s0[67]}), .a ({new_AGEMA_signal_3826, new_AGEMA_signal_3825, new_AGEMA_signal_3824, KeyArray_outS20ser[3]}), .c ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, new_AGEMA_signal_3827, KeyArray_inS13ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS13ser_mux_inst_4_U1 ( .s (KeyArray_n43), .b ({key_s3[68], key_s2[68], key_s1[68], key_s0[68]}), .a ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, new_AGEMA_signal_3833, KeyArray_outS20ser[4]}), .c ({new_AGEMA_signal_3838, new_AGEMA_signal_3837, new_AGEMA_signal_3836, KeyArray_inS13ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS13ser_mux_inst_5_U1 ( .s (KeyArray_n43), .b ({key_s3[69], key_s2[69], key_s1[69], key_s0[69]}), .a ({new_AGEMA_signal_3844, new_AGEMA_signal_3843, new_AGEMA_signal_3842, KeyArray_outS20ser[5]}), .c ({new_AGEMA_signal_3847, new_AGEMA_signal_3846, new_AGEMA_signal_3845, KeyArray_inS13ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS13ser_mux_inst_6_U1 ( .s (KeyArray_n43), .b ({key_s3[70], key_s2[70], key_s1[70], key_s0[70]}), .a ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, new_AGEMA_signal_3851, KeyArray_outS20ser[6]}), .c ({new_AGEMA_signal_3856, new_AGEMA_signal_3855, new_AGEMA_signal_3854, KeyArray_inS13ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS13ser_mux_inst_7_U1 ( .s (KeyArray_n43), .b ({key_s3[71], key_s2[71], key_s1[71], key_s0[71]}), .a ({new_AGEMA_signal_3862, new_AGEMA_signal_3861, new_AGEMA_signal_3860, KeyArray_outS20ser[7]}), .c ({new_AGEMA_signal_3865, new_AGEMA_signal_3864, new_AGEMA_signal_3863, KeyArray_inS13ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS20ser_mux_inst_0_U1 ( .s (KeyArray_n42), .b ({key_s3[56], key_s2[56], key_s1[56], key_s0[56]}), .a ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, new_AGEMA_signal_3869, KeyArray_outS21ser[0]}), .c ({new_AGEMA_signal_3874, new_AGEMA_signal_3873, new_AGEMA_signal_3872, KeyArray_inS20ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS20ser_mux_inst_1_U1 ( .s (KeyArray_n42), .b ({key_s3[57], key_s2[57], key_s1[57], key_s0[57]}), .a ({new_AGEMA_signal_3880, new_AGEMA_signal_3879, new_AGEMA_signal_3878, KeyArray_outS21ser[1]}), .c ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, new_AGEMA_signal_3881, KeyArray_inS20ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS20ser_mux_inst_2_U1 ( .s (KeyArray_n42), .b ({key_s3[58], key_s2[58], key_s1[58], key_s0[58]}), .a ({new_AGEMA_signal_3889, new_AGEMA_signal_3888, new_AGEMA_signal_3887, KeyArray_outS21ser[2]}), .c ({new_AGEMA_signal_3892, new_AGEMA_signal_3891, new_AGEMA_signal_3890, KeyArray_inS20ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS20ser_mux_inst_3_U1 ( .s (KeyArray_n42), .b ({key_s3[59], key_s2[59], key_s1[59], key_s0[59]}), .a ({new_AGEMA_signal_3898, new_AGEMA_signal_3897, new_AGEMA_signal_3896, KeyArray_outS21ser[3]}), .c ({new_AGEMA_signal_3901, new_AGEMA_signal_3900, new_AGEMA_signal_3899, KeyArray_inS20ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS20ser_mux_inst_4_U1 ( .s (KeyArray_n42), .b ({key_s3[60], key_s2[60], key_s1[60], key_s0[60]}), .a ({new_AGEMA_signal_3907, new_AGEMA_signal_3906, new_AGEMA_signal_3905, KeyArray_outS21ser[4]}), .c ({new_AGEMA_signal_3910, new_AGEMA_signal_3909, new_AGEMA_signal_3908, KeyArray_inS20ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS20ser_mux_inst_5_U1 ( .s (KeyArray_n42), .b ({key_s3[61], key_s2[61], key_s1[61], key_s0[61]}), .a ({new_AGEMA_signal_3916, new_AGEMA_signal_3915, new_AGEMA_signal_3914, KeyArray_outS21ser[5]}), .c ({new_AGEMA_signal_3919, new_AGEMA_signal_3918, new_AGEMA_signal_3917, KeyArray_inS20ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS20ser_mux_inst_6_U1 ( .s (KeyArray_n42), .b ({key_s3[62], key_s2[62], key_s1[62], key_s0[62]}), .a ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, new_AGEMA_signal_3923, KeyArray_outS21ser[6]}), .c ({new_AGEMA_signal_3928, new_AGEMA_signal_3927, new_AGEMA_signal_3926, KeyArray_inS20ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS20ser_mux_inst_7_U1 ( .s (KeyArray_n42), .b ({key_s3[63], key_s2[63], key_s1[63], key_s0[63]}), .a ({new_AGEMA_signal_3934, new_AGEMA_signal_3933, new_AGEMA_signal_3932, KeyArray_outS21ser[7]}), .c ({new_AGEMA_signal_3937, new_AGEMA_signal_3936, new_AGEMA_signal_3935, KeyArray_inS20ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS21ser_mux_inst_0_U1 ( .s (KeyArray_n42), .b ({key_s3[48], key_s2[48], key_s1[48], key_s0[48]}), .a ({new_AGEMA_signal_3943, new_AGEMA_signal_3942, new_AGEMA_signal_3941, KeyArray_outS22ser[0]}), .c ({new_AGEMA_signal_3946, new_AGEMA_signal_3945, new_AGEMA_signal_3944, KeyArray_inS21ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS21ser_mux_inst_1_U1 ( .s (KeyArray_n42), .b ({key_s3[49], key_s2[49], key_s1[49], key_s0[49]}), .a ({new_AGEMA_signal_3952, new_AGEMA_signal_3951, new_AGEMA_signal_3950, KeyArray_outS22ser[1]}), .c ({new_AGEMA_signal_3955, new_AGEMA_signal_3954, new_AGEMA_signal_3953, KeyArray_inS21ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS21ser_mux_inst_2_U1 ( .s (KeyArray_n42), .b ({key_s3[50], key_s2[50], key_s1[50], key_s0[50]}), .a ({new_AGEMA_signal_3961, new_AGEMA_signal_3960, new_AGEMA_signal_3959, KeyArray_outS22ser[2]}), .c ({new_AGEMA_signal_3964, new_AGEMA_signal_3963, new_AGEMA_signal_3962, KeyArray_inS21ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS21ser_mux_inst_3_U1 ( .s (KeyArray_n42), .b ({key_s3[51], key_s2[51], key_s1[51], key_s0[51]}), .a ({new_AGEMA_signal_3970, new_AGEMA_signal_3969, new_AGEMA_signal_3968, KeyArray_outS22ser[3]}), .c ({new_AGEMA_signal_3973, new_AGEMA_signal_3972, new_AGEMA_signal_3971, KeyArray_inS21ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS21ser_mux_inst_4_U1 ( .s (KeyArray_n42), .b ({key_s3[52], key_s2[52], key_s1[52], key_s0[52]}), .a ({new_AGEMA_signal_3979, new_AGEMA_signal_3978, new_AGEMA_signal_3977, KeyArray_outS22ser[4]}), .c ({new_AGEMA_signal_3982, new_AGEMA_signal_3981, new_AGEMA_signal_3980, KeyArray_inS21ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS21ser_mux_inst_5_U1 ( .s (KeyArray_n42), .b ({key_s3[53], key_s2[53], key_s1[53], key_s0[53]}), .a ({new_AGEMA_signal_3988, new_AGEMA_signal_3987, new_AGEMA_signal_3986, KeyArray_outS22ser[5]}), .c ({new_AGEMA_signal_3991, new_AGEMA_signal_3990, new_AGEMA_signal_3989, KeyArray_inS21ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS21ser_mux_inst_6_U1 ( .s (KeyArray_n42), .b ({key_s3[54], key_s2[54], key_s1[54], key_s0[54]}), .a ({new_AGEMA_signal_3997, new_AGEMA_signal_3996, new_AGEMA_signal_3995, KeyArray_outS22ser[6]}), .c ({new_AGEMA_signal_4000, new_AGEMA_signal_3999, new_AGEMA_signal_3998, KeyArray_inS21ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS21ser_mux_inst_7_U1 ( .s (KeyArray_n42), .b ({key_s3[55], key_s2[55], key_s1[55], key_s0[55]}), .a ({new_AGEMA_signal_4006, new_AGEMA_signal_4005, new_AGEMA_signal_4004, KeyArray_outS22ser[7]}), .c ({new_AGEMA_signal_4009, new_AGEMA_signal_4008, new_AGEMA_signal_4007, KeyArray_inS21ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS22ser_mux_inst_0_U1 ( .s (KeyArray_n41), .b ({key_s3[40], key_s2[40], key_s1[40], key_s0[40]}), .a ({new_AGEMA_signal_4015, new_AGEMA_signal_4014, new_AGEMA_signal_4013, KeyArray_outS23ser[0]}), .c ({new_AGEMA_signal_4018, new_AGEMA_signal_4017, new_AGEMA_signal_4016, KeyArray_inS22ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS22ser_mux_inst_1_U1 ( .s (KeyArray_n41), .b ({key_s3[41], key_s2[41], key_s1[41], key_s0[41]}), .a ({new_AGEMA_signal_4024, new_AGEMA_signal_4023, new_AGEMA_signal_4022, KeyArray_outS23ser[1]}), .c ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, new_AGEMA_signal_4025, KeyArray_inS22ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS22ser_mux_inst_2_U1 ( .s (KeyArray_n41), .b ({key_s3[42], key_s2[42], key_s1[42], key_s0[42]}), .a ({new_AGEMA_signal_4033, new_AGEMA_signal_4032, new_AGEMA_signal_4031, KeyArray_outS23ser[2]}), .c ({new_AGEMA_signal_4036, new_AGEMA_signal_4035, new_AGEMA_signal_4034, KeyArray_inS22ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS22ser_mux_inst_3_U1 ( .s (KeyArray_n41), .b ({key_s3[43], key_s2[43], key_s1[43], key_s0[43]}), .a ({new_AGEMA_signal_4042, new_AGEMA_signal_4041, new_AGEMA_signal_4040, KeyArray_outS23ser[3]}), .c ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, new_AGEMA_signal_4043, KeyArray_inS22ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS22ser_mux_inst_4_U1 ( .s (KeyArray_n41), .b ({key_s3[44], key_s2[44], key_s1[44], key_s0[44]}), .a ({new_AGEMA_signal_4051, new_AGEMA_signal_4050, new_AGEMA_signal_4049, KeyArray_outS23ser[4]}), .c ({new_AGEMA_signal_4054, new_AGEMA_signal_4053, new_AGEMA_signal_4052, KeyArray_inS22ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS22ser_mux_inst_5_U1 ( .s (KeyArray_n41), .b ({key_s3[45], key_s2[45], key_s1[45], key_s0[45]}), .a ({new_AGEMA_signal_4060, new_AGEMA_signal_4059, new_AGEMA_signal_4058, KeyArray_outS23ser[5]}), .c ({new_AGEMA_signal_4063, new_AGEMA_signal_4062, new_AGEMA_signal_4061, KeyArray_inS22ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS22ser_mux_inst_6_U1 ( .s (KeyArray_n41), .b ({key_s3[46], key_s2[46], key_s1[46], key_s0[46]}), .a ({new_AGEMA_signal_4069, new_AGEMA_signal_4068, new_AGEMA_signal_4067, KeyArray_outS23ser[6]}), .c ({new_AGEMA_signal_4072, new_AGEMA_signal_4071, new_AGEMA_signal_4070, KeyArray_inS22ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS22ser_mux_inst_7_U1 ( .s (KeyArray_n41), .b ({key_s3[47], key_s2[47], key_s1[47], key_s0[47]}), .a ({new_AGEMA_signal_4078, new_AGEMA_signal_4077, new_AGEMA_signal_4076, KeyArray_outS23ser[7]}), .c ({new_AGEMA_signal_4081, new_AGEMA_signal_4080, new_AGEMA_signal_4079, KeyArray_inS22ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS23ser_mux_inst_0_U1 ( .s (KeyArray_n41), .b ({key_s3[32], key_s2[32], key_s1[32], key_s0[32]}), .a ({new_AGEMA_signal_4087, new_AGEMA_signal_4086, new_AGEMA_signal_4085, KeyArray_outS30ser[0]}), .c ({new_AGEMA_signal_4090, new_AGEMA_signal_4089, new_AGEMA_signal_4088, KeyArray_inS23ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS23ser_mux_inst_1_U1 ( .s (KeyArray_n41), .b ({key_s3[33], key_s2[33], key_s1[33], key_s0[33]}), .a ({new_AGEMA_signal_4096, new_AGEMA_signal_4095, new_AGEMA_signal_4094, KeyArray_outS30ser[1]}), .c ({new_AGEMA_signal_4099, new_AGEMA_signal_4098, new_AGEMA_signal_4097, KeyArray_inS23ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS23ser_mux_inst_2_U1 ( .s (KeyArray_n41), .b ({key_s3[34], key_s2[34], key_s1[34], key_s0[34]}), .a ({new_AGEMA_signal_4105, new_AGEMA_signal_4104, new_AGEMA_signal_4103, KeyArray_outS30ser[2]}), .c ({new_AGEMA_signal_4108, new_AGEMA_signal_4107, new_AGEMA_signal_4106, KeyArray_inS23ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS23ser_mux_inst_3_U1 ( .s (KeyArray_n41), .b ({key_s3[35], key_s2[35], key_s1[35], key_s0[35]}), .a ({new_AGEMA_signal_4114, new_AGEMA_signal_4113, new_AGEMA_signal_4112, KeyArray_outS30ser[3]}), .c ({new_AGEMA_signal_4117, new_AGEMA_signal_4116, new_AGEMA_signal_4115, KeyArray_inS23ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS23ser_mux_inst_4_U1 ( .s (KeyArray_n41), .b ({key_s3[36], key_s2[36], key_s1[36], key_s0[36]}), .a ({new_AGEMA_signal_4123, new_AGEMA_signal_4122, new_AGEMA_signal_4121, KeyArray_outS30ser[4]}), .c ({new_AGEMA_signal_4126, new_AGEMA_signal_4125, new_AGEMA_signal_4124, KeyArray_inS23ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS23ser_mux_inst_5_U1 ( .s (KeyArray_n41), .b ({key_s3[37], key_s2[37], key_s1[37], key_s0[37]}), .a ({new_AGEMA_signal_4132, new_AGEMA_signal_4131, new_AGEMA_signal_4130, KeyArray_outS30ser[5]}), .c ({new_AGEMA_signal_4135, new_AGEMA_signal_4134, new_AGEMA_signal_4133, KeyArray_inS23ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS23ser_mux_inst_6_U1 ( .s (KeyArray_n41), .b ({key_s3[38], key_s2[38], key_s1[38], key_s0[38]}), .a ({new_AGEMA_signal_4141, new_AGEMA_signal_4140, new_AGEMA_signal_4139, KeyArray_outS30ser[6]}), .c ({new_AGEMA_signal_4144, new_AGEMA_signal_4143, new_AGEMA_signal_4142, KeyArray_inS23ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS23ser_mux_inst_7_U1 ( .s (KeyArray_n41), .b ({key_s3[39], key_s2[39], key_s1[39], key_s0[39]}), .a ({new_AGEMA_signal_4150, new_AGEMA_signal_4149, new_AGEMA_signal_4148, KeyArray_outS30ser[7]}), .c ({new_AGEMA_signal_4153, new_AGEMA_signal_4152, new_AGEMA_signal_4151, KeyArray_inS23ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS30ser_mux_inst_0_U1 ( .s (KeyArray_n40), .b ({key_s3[24], key_s2[24], key_s1[24], key_s0[24]}), .a ({new_AGEMA_signal_4159, new_AGEMA_signal_4158, new_AGEMA_signal_4157, KeyArray_outS31ser[0]}), .c ({new_AGEMA_signal_4162, new_AGEMA_signal_4161, new_AGEMA_signal_4160, KeyArray_inS30ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS30ser_mux_inst_1_U1 ( .s (KeyArray_n40), .b ({key_s3[25], key_s2[25], key_s1[25], key_s0[25]}), .a ({new_AGEMA_signal_4168, new_AGEMA_signal_4167, new_AGEMA_signal_4166, KeyArray_outS31ser[1]}), .c ({new_AGEMA_signal_4171, new_AGEMA_signal_4170, new_AGEMA_signal_4169, KeyArray_inS30ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS30ser_mux_inst_2_U1 ( .s (KeyArray_n40), .b ({key_s3[26], key_s2[26], key_s1[26], key_s0[26]}), .a ({new_AGEMA_signal_4177, new_AGEMA_signal_4176, new_AGEMA_signal_4175, KeyArray_outS31ser[2]}), .c ({new_AGEMA_signal_4180, new_AGEMA_signal_4179, new_AGEMA_signal_4178, KeyArray_inS30ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS30ser_mux_inst_3_U1 ( .s (KeyArray_n40), .b ({key_s3[27], key_s2[27], key_s1[27], key_s0[27]}), .a ({new_AGEMA_signal_4186, new_AGEMA_signal_4185, new_AGEMA_signal_4184, KeyArray_outS31ser[3]}), .c ({new_AGEMA_signal_4189, new_AGEMA_signal_4188, new_AGEMA_signal_4187, KeyArray_inS30ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS30ser_mux_inst_4_U1 ( .s (KeyArray_n40), .b ({key_s3[28], key_s2[28], key_s1[28], key_s0[28]}), .a ({new_AGEMA_signal_4195, new_AGEMA_signal_4194, new_AGEMA_signal_4193, KeyArray_outS31ser[4]}), .c ({new_AGEMA_signal_4198, new_AGEMA_signal_4197, new_AGEMA_signal_4196, KeyArray_inS30ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS30ser_mux_inst_5_U1 ( .s (KeyArray_n40), .b ({key_s3[29], key_s2[29], key_s1[29], key_s0[29]}), .a ({new_AGEMA_signal_4204, new_AGEMA_signal_4203, new_AGEMA_signal_4202, KeyArray_outS31ser[5]}), .c ({new_AGEMA_signal_4207, new_AGEMA_signal_4206, new_AGEMA_signal_4205, KeyArray_inS30ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS30ser_mux_inst_6_U1 ( .s (KeyArray_n40), .b ({key_s3[30], key_s2[30], key_s1[30], key_s0[30]}), .a ({new_AGEMA_signal_4213, new_AGEMA_signal_4212, new_AGEMA_signal_4211, KeyArray_outS31ser[6]}), .c ({new_AGEMA_signal_4216, new_AGEMA_signal_4215, new_AGEMA_signal_4214, KeyArray_inS30ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS30ser_mux_inst_7_U1 ( .s (KeyArray_n40), .b ({key_s3[31], key_s2[31], key_s1[31], key_s0[31]}), .a ({new_AGEMA_signal_4222, new_AGEMA_signal_4221, new_AGEMA_signal_4220, KeyArray_outS31ser[7]}), .c ({new_AGEMA_signal_4225, new_AGEMA_signal_4224, new_AGEMA_signal_4223, KeyArray_inS30ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS31ser_mux_inst_0_U1 ( .s (KeyArray_n40), .b ({key_s3[16], key_s2[16], key_s1[16], key_s0[16]}), .a ({new_AGEMA_signal_4231, new_AGEMA_signal_4230, new_AGEMA_signal_4229, KeyArray_outS32ser[0]}), .c ({new_AGEMA_signal_4234, new_AGEMA_signal_4233, new_AGEMA_signal_4232, KeyArray_inS31ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS31ser_mux_inst_1_U1 ( .s (KeyArray_n40), .b ({key_s3[17], key_s2[17], key_s1[17], key_s0[17]}), .a ({new_AGEMA_signal_4240, new_AGEMA_signal_4239, new_AGEMA_signal_4238, KeyArray_outS32ser[1]}), .c ({new_AGEMA_signal_4243, new_AGEMA_signal_4242, new_AGEMA_signal_4241, KeyArray_inS31ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS31ser_mux_inst_2_U1 ( .s (KeyArray_n40), .b ({key_s3[18], key_s2[18], key_s1[18], key_s0[18]}), .a ({new_AGEMA_signal_4249, new_AGEMA_signal_4248, new_AGEMA_signal_4247, KeyArray_outS32ser[2]}), .c ({new_AGEMA_signal_4252, new_AGEMA_signal_4251, new_AGEMA_signal_4250, KeyArray_inS31ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS31ser_mux_inst_3_U1 ( .s (KeyArray_n40), .b ({key_s3[19], key_s2[19], key_s1[19], key_s0[19]}), .a ({new_AGEMA_signal_4258, new_AGEMA_signal_4257, new_AGEMA_signal_4256, KeyArray_outS32ser[3]}), .c ({new_AGEMA_signal_4261, new_AGEMA_signal_4260, new_AGEMA_signal_4259, KeyArray_inS31ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS31ser_mux_inst_4_U1 ( .s (KeyArray_n40), .b ({key_s3[20], key_s2[20], key_s1[20], key_s0[20]}), .a ({new_AGEMA_signal_4267, new_AGEMA_signal_4266, new_AGEMA_signal_4265, KeyArray_outS32ser[4]}), .c ({new_AGEMA_signal_4270, new_AGEMA_signal_4269, new_AGEMA_signal_4268, KeyArray_inS31ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS31ser_mux_inst_5_U1 ( .s (KeyArray_n40), .b ({key_s3[21], key_s2[21], key_s1[21], key_s0[21]}), .a ({new_AGEMA_signal_4276, new_AGEMA_signal_4275, new_AGEMA_signal_4274, KeyArray_outS32ser[5]}), .c ({new_AGEMA_signal_4279, new_AGEMA_signal_4278, new_AGEMA_signal_4277, KeyArray_inS31ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS31ser_mux_inst_6_U1 ( .s (KeyArray_n40), .b ({key_s3[22], key_s2[22], key_s1[22], key_s0[22]}), .a ({new_AGEMA_signal_4285, new_AGEMA_signal_4284, new_AGEMA_signal_4283, KeyArray_outS32ser[6]}), .c ({new_AGEMA_signal_4288, new_AGEMA_signal_4287, new_AGEMA_signal_4286, KeyArray_inS31ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS31ser_mux_inst_7_U1 ( .s (KeyArray_n40), .b ({key_s3[23], key_s2[23], key_s1[23], key_s0[23]}), .a ({new_AGEMA_signal_4294, new_AGEMA_signal_4293, new_AGEMA_signal_4292, KeyArray_outS32ser[7]}), .c ({new_AGEMA_signal_4297, new_AGEMA_signal_4296, new_AGEMA_signal_4295, KeyArray_inS31ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS32ser_mux_inst_0_U1 ( .s (KeyArray_n39), .b ({key_s3[8], key_s2[8], key_s1[8], key_s0[8]}), .a ({new_AGEMA_signal_4303, new_AGEMA_signal_4302, new_AGEMA_signal_4301, KeyArray_outS33ser[0]}), .c ({new_AGEMA_signal_4306, new_AGEMA_signal_4305, new_AGEMA_signal_4304, KeyArray_inS32ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS32ser_mux_inst_1_U1 ( .s (KeyArray_n39), .b ({key_s3[9], key_s2[9], key_s1[9], key_s0[9]}), .a ({new_AGEMA_signal_4312, new_AGEMA_signal_4311, new_AGEMA_signal_4310, KeyArray_outS33ser[1]}), .c ({new_AGEMA_signal_4315, new_AGEMA_signal_4314, new_AGEMA_signal_4313, KeyArray_inS32ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS32ser_mux_inst_2_U1 ( .s (KeyArray_n39), .b ({key_s3[10], key_s2[10], key_s1[10], key_s0[10]}), .a ({new_AGEMA_signal_4321, new_AGEMA_signal_4320, new_AGEMA_signal_4319, KeyArray_outS33ser[2]}), .c ({new_AGEMA_signal_4324, new_AGEMA_signal_4323, new_AGEMA_signal_4322, KeyArray_inS32ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS32ser_mux_inst_3_U1 ( .s (KeyArray_n39), .b ({key_s3[11], key_s2[11], key_s1[11], key_s0[11]}), .a ({new_AGEMA_signal_4330, new_AGEMA_signal_4329, new_AGEMA_signal_4328, KeyArray_outS33ser[3]}), .c ({new_AGEMA_signal_4333, new_AGEMA_signal_4332, new_AGEMA_signal_4331, KeyArray_inS32ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS32ser_mux_inst_4_U1 ( .s (KeyArray_n39), .b ({key_s3[12], key_s2[12], key_s1[12], key_s0[12]}), .a ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, new_AGEMA_signal_4337, KeyArray_outS33ser[4]}), .c ({new_AGEMA_signal_4342, new_AGEMA_signal_4341, new_AGEMA_signal_4340, KeyArray_inS32ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS32ser_mux_inst_5_U1 ( .s (KeyArray_n39), .b ({key_s3[13], key_s2[13], key_s1[13], key_s0[13]}), .a ({new_AGEMA_signal_4348, new_AGEMA_signal_4347, new_AGEMA_signal_4346, KeyArray_outS33ser[5]}), .c ({new_AGEMA_signal_4351, new_AGEMA_signal_4350, new_AGEMA_signal_4349, KeyArray_inS32ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS32ser_mux_inst_6_U1 ( .s (KeyArray_n39), .b ({key_s3[14], key_s2[14], key_s1[14], key_s0[14]}), .a ({new_AGEMA_signal_4357, new_AGEMA_signal_4356, new_AGEMA_signal_4355, KeyArray_outS33ser[6]}), .c ({new_AGEMA_signal_4360, new_AGEMA_signal_4359, new_AGEMA_signal_4358, KeyArray_inS32ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS32ser_mux_inst_7_U1 ( .s (KeyArray_n39), .b ({key_s3[15], key_s2[15], key_s1[15], key_s0[15]}), .a ({new_AGEMA_signal_4366, new_AGEMA_signal_4365, new_AGEMA_signal_4364, KeyArray_outS33ser[7]}), .c ({new_AGEMA_signal_4369, new_AGEMA_signal_4368, new_AGEMA_signal_4367, KeyArray_inS32ser[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS33ser_mux_inst_0_U1 ( .s (KeyArray_n39), .b ({key_s3[0], key_s2[0], key_s1[0], key_s0[0]}), .a ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, new_AGEMA_signal_1985, keyStateIn[0]}), .c ({new_AGEMA_signal_4375, new_AGEMA_signal_4374, new_AGEMA_signal_4373, KeyArray_inS33ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS33ser_mux_inst_1_U1 ( .s (KeyArray_n39), .b ({key_s3[1], key_s2[1], key_s1[1], key_s0[1]}), .a ({new_AGEMA_signal_1996, new_AGEMA_signal_1995, new_AGEMA_signal_1994, keyStateIn[1]}), .c ({new_AGEMA_signal_4381, new_AGEMA_signal_4380, new_AGEMA_signal_4379, KeyArray_inS33ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS33ser_mux_inst_2_U1 ( .s (KeyArray_n39), .b ({key_s3[2], key_s2[2], key_s1[2], key_s0[2]}), .a ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, new_AGEMA_signal_2003, keyStateIn[2]}), .c ({new_AGEMA_signal_4387, new_AGEMA_signal_4386, new_AGEMA_signal_4385, KeyArray_inS33ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS33ser_mux_inst_3_U1 ( .s (KeyArray_n39), .b ({key_s3[3], key_s2[3], key_s1[3], key_s0[3]}), .a ({new_AGEMA_signal_2014, new_AGEMA_signal_2013, new_AGEMA_signal_2012, keyStateIn[3]}), .c ({new_AGEMA_signal_4393, new_AGEMA_signal_4392, new_AGEMA_signal_4391, KeyArray_inS33ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS33ser_mux_inst_4_U1 ( .s (KeyArray_n39), .b ({key_s3[4], key_s2[4], key_s1[4], key_s0[4]}), .a ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, new_AGEMA_signal_2021, keyStateIn[4]}), .c ({new_AGEMA_signal_4399, new_AGEMA_signal_4398, new_AGEMA_signal_4397, KeyArray_inS33ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS33ser_mux_inst_5_U1 ( .s (KeyArray_n39), .b ({key_s3[5], key_s2[5], key_s1[5], key_s0[5]}), .a ({new_AGEMA_signal_2032, new_AGEMA_signal_2031, new_AGEMA_signal_2030, keyStateIn[5]}), .c ({new_AGEMA_signal_4405, new_AGEMA_signal_4404, new_AGEMA_signal_4403, KeyArray_inS33ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS33ser_mux_inst_6_U1 ( .s (KeyArray_n39), .b ({key_s3[6], key_s2[6], key_s1[6], key_s0[6]}), .a ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, new_AGEMA_signal_2039, keyStateIn[6]}), .c ({new_AGEMA_signal_4411, new_AGEMA_signal_4410, new_AGEMA_signal_4409, KeyArray_inS33ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_MUX_inS33ser_mux_inst_7_U1 ( .s (KeyArray_n39), .b ({key_s3[7], key_s2[7], key_s1[7], key_s0[7]}), .a ({new_AGEMA_signal_2050, new_AGEMA_signal_2049, new_AGEMA_signal_2048, keyStateIn[7]}), .c ({new_AGEMA_signal_4417, new_AGEMA_signal_4416, new_AGEMA_signal_4415, KeyArray_inS33ser[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U24 ( .a ({new_AGEMA_signal_2404, new_AGEMA_signal_2403, new_AGEMA_signal_2402, MixColumns_line0_n16}), .b ({new_AGEMA_signal_2110, new_AGEMA_signal_2109, new_AGEMA_signal_2108, MixColumns_line0_n15}), .c ({new_AGEMA_signal_4420, new_AGEMA_signal_4419, new_AGEMA_signal_4418, MCout[31]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U23 ( .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .c ({new_AGEMA_signal_2110, new_AGEMA_signal_2109, new_AGEMA_signal_2108, MixColumns_line0_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U22 ( .a ({ciphertext_s3[126], ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .b ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, new_AGEMA_signal_2189, MixColumns_line0_S13[7]}), .c ({new_AGEMA_signal_2404, new_AGEMA_signal_2403, new_AGEMA_signal_2402, MixColumns_line0_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U21 ( .a ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, new_AGEMA_signal_2405, MixColumns_line0_n14}), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, new_AGEMA_signal_2117, MixColumns_line0_n13}), .c ({new_AGEMA_signal_4423, new_AGEMA_signal_4422, new_AGEMA_signal_4421, MCout[30]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U20 ( .a ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .c ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, new_AGEMA_signal_2117, MixColumns_line0_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U19 ( .a ({ciphertext_s3[125], ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .b ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, new_AGEMA_signal_2195, MixColumns_line0_S13[6]}), .c ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, new_AGEMA_signal_2405, MixColumns_line0_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U18 ( .a ({new_AGEMA_signal_2410, new_AGEMA_signal_2409, new_AGEMA_signal_2408, MixColumns_line0_n12}), .b ({new_AGEMA_signal_2128, new_AGEMA_signal_2127, new_AGEMA_signal_2126, MixColumns_line0_n11}), .c ({new_AGEMA_signal_4426, new_AGEMA_signal_4425, new_AGEMA_signal_4424, MCout[29]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U17 ( .a ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_2128, new_AGEMA_signal_2127, new_AGEMA_signal_2126, MixColumns_line0_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U16 ( .a ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .b ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, new_AGEMA_signal_2201, MixColumns_line0_S13[5]}), .c ({new_AGEMA_signal_2410, new_AGEMA_signal_2409, new_AGEMA_signal_2408, MixColumns_line0_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U15 ( .a ({new_AGEMA_signal_4429, new_AGEMA_signal_4428, new_AGEMA_signal_4427, MixColumns_line0_n10}), .b ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, new_AGEMA_signal_2135, MixColumns_line0_n9}), .c ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, new_AGEMA_signal_4550, MCout[28]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U14 ( .a ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, new_AGEMA_signal_2135, MixColumns_line0_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U13 ( .a ({new_AGEMA_signal_2176, new_AGEMA_signal_2175, new_AGEMA_signal_2174, MixColumns_line0_S02[4]}), .b ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, new_AGEMA_signal_2417, MixColumns_line0_S13[4]}), .c ({new_AGEMA_signal_4429, new_AGEMA_signal_4428, new_AGEMA_signal_4427, MixColumns_line0_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U12 ( .a ({new_AGEMA_signal_4432, new_AGEMA_signal_4431, new_AGEMA_signal_4430, MixColumns_line0_n8}), .b ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, new_AGEMA_signal_2144, MixColumns_line0_n7}), .c ({new_AGEMA_signal_4555, new_AGEMA_signal_4554, new_AGEMA_signal_4553, MCout[27]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U11 ( .a ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .b ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, new_AGEMA_signal_2144, MixColumns_line0_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U10 ( .a ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, new_AGEMA_signal_2177, MixColumns_line0_S02[3]}), .b ({new_AGEMA_signal_2422, new_AGEMA_signal_2421, new_AGEMA_signal_2420, MixColumns_line0_S13[3]}), .c ({new_AGEMA_signal_4432, new_AGEMA_signal_4431, new_AGEMA_signal_4430, MixColumns_line0_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U9 ( .a ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, new_AGEMA_signal_2411, MixColumns_line0_n6}), .b ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, new_AGEMA_signal_2153, MixColumns_line0_n5}), .c ({new_AGEMA_signal_4435, new_AGEMA_signal_4434, new_AGEMA_signal_4433, MCout[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U8 ( .a ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, new_AGEMA_signal_2153, MixColumns_line0_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U7 ( .a ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .b ({new_AGEMA_signal_2212, new_AGEMA_signal_2211, new_AGEMA_signal_2210, MixColumns_line0_S13[2]}), .c ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, new_AGEMA_signal_2411, MixColumns_line0_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U6 ( .a ({new_AGEMA_signal_4438, new_AGEMA_signal_4437, new_AGEMA_signal_4436, MixColumns_line0_n4}), .b ({new_AGEMA_signal_2164, new_AGEMA_signal_2163, new_AGEMA_signal_2162, MixColumns_line0_n3}), .c ({new_AGEMA_signal_4558, new_AGEMA_signal_4557, new_AGEMA_signal_4556, MCout[25]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U5 ( .a ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .b ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_2164, new_AGEMA_signal_2163, new_AGEMA_signal_2162, MixColumns_line0_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U4 ( .a ({new_AGEMA_signal_2182, new_AGEMA_signal_2181, new_AGEMA_signal_2180, MixColumns_line0_S02[1]}), .b ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, new_AGEMA_signal_2423, MixColumns_line0_S13[1]}), .c ({new_AGEMA_signal_4438, new_AGEMA_signal_4437, new_AGEMA_signal_4436, MixColumns_line0_n4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U3 ( .a ({new_AGEMA_signal_2416, new_AGEMA_signal_2415, new_AGEMA_signal_2414, MixColumns_line0_n2}), .b ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, new_AGEMA_signal_2171, MixColumns_line0_n1}), .c ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, new_AGEMA_signal_4439, MCout[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U2 ( .a ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, new_AGEMA_signal_2171, MixColumns_line0_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_U1 ( .a ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_2218, new_AGEMA_signal_2217, new_AGEMA_signal_2216, MixColumns_line0_S13[0]}), .c ({new_AGEMA_signal_2416, new_AGEMA_signal_2415, new_AGEMA_signal_2414, MixColumns_line0_n2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_timesTWO_U3 ( .a ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s3[123], ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_2176, new_AGEMA_signal_2175, new_AGEMA_signal_2174, MixColumns_line0_S02[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_timesTWO_U2 ( .a ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, new_AGEMA_signal_2177, MixColumns_line0_S02[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_timesTWO_U1 ( .a ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_2182, new_AGEMA_signal_2181, new_AGEMA_signal_2180, MixColumns_line0_S02[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_timesTHREE_U8 ( .a ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s3[94], ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .c ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, new_AGEMA_signal_2189, MixColumns_line0_S13[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_timesTHREE_U7 ( .a ({ciphertext_s3[94], ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s3[93], ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, new_AGEMA_signal_2195, MixColumns_line0_S13[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_timesTHREE_U6 ( .a ({ciphertext_s3[93], ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, new_AGEMA_signal_2201, MixColumns_line0_S13[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_timesTHREE_U5 ( .a ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .b ({new_AGEMA_signal_2224, new_AGEMA_signal_2223, new_AGEMA_signal_2222, MixColumns_line0_timesTHREE_input2[4]}), .c ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, new_AGEMA_signal_2417, MixColumns_line0_S13[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_timesTHREE_U4 ( .a ({ciphertext_s3[91], ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}), .b ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, new_AGEMA_signal_2225, MixColumns_line0_timesTHREE_input2[3]}), .c ({new_AGEMA_signal_2422, new_AGEMA_signal_2421, new_AGEMA_signal_2420, MixColumns_line0_S13[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_timesTHREE_U3 ( .a ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_2212, new_AGEMA_signal_2211, new_AGEMA_signal_2210, MixColumns_line0_S13[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_timesTHREE_U2 ( .a ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .b ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, new_AGEMA_signal_2228, MixColumns_line0_timesTHREE_input2[1]}), .c ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, new_AGEMA_signal_2423, MixColumns_line0_S13[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_timesTHREE_U1 ( .a ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .b ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .c ({new_AGEMA_signal_2218, new_AGEMA_signal_2217, new_AGEMA_signal_2216, MixColumns_line0_S13[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_timesTHREE_timesTWO_U3 ( .a ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s3[91], ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_2224, new_AGEMA_signal_2223, new_AGEMA_signal_2222, MixColumns_line0_timesTHREE_input2[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_timesTHREE_timesTWO_U2 ( .a ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, new_AGEMA_signal_2225, MixColumns_line0_timesTHREE_input2[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line0_timesTHREE_timesTWO_U1 ( .a ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, new_AGEMA_signal_2228, MixColumns_line0_timesTHREE_input2[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U24 ( .a ({new_AGEMA_signal_2428, new_AGEMA_signal_2427, new_AGEMA_signal_2426, MixColumns_line1_n16}), .b ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, new_AGEMA_signal_2231, MixColumns_line1_n15}), .c ({new_AGEMA_signal_4444, new_AGEMA_signal_4443, new_AGEMA_signal_4442, MCout[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U23 ( .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .c ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, new_AGEMA_signal_2231, MixColumns_line1_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U22 ( .a ({ciphertext_s3[94], ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .b ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, new_AGEMA_signal_2264, MixColumns_line1_S13[7]}), .c ({new_AGEMA_signal_2428, new_AGEMA_signal_2427, new_AGEMA_signal_2426, MixColumns_line1_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U21 ( .a ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, new_AGEMA_signal_2429, MixColumns_line1_n14}), .b ({new_AGEMA_signal_2236, new_AGEMA_signal_2235, new_AGEMA_signal_2234, MixColumns_line1_n13}), .c ({new_AGEMA_signal_4447, new_AGEMA_signal_4446, new_AGEMA_signal_4445, MCout[22]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U20 ( .a ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s3[126], ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .c ({new_AGEMA_signal_2236, new_AGEMA_signal_2235, new_AGEMA_signal_2234, MixColumns_line1_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U19 ( .a ({ciphertext_s3[93], ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .b ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, new_AGEMA_signal_2267, MixColumns_line1_S13[6]}), .c ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, new_AGEMA_signal_2429, MixColumns_line1_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U18 ( .a ({new_AGEMA_signal_2434, new_AGEMA_signal_2433, new_AGEMA_signal_2432, MixColumns_line1_n12}), .b ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, new_AGEMA_signal_2237, MixColumns_line1_n11}), .c ({new_AGEMA_signal_4450, new_AGEMA_signal_4449, new_AGEMA_signal_4448, MCout[21]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U17 ( .a ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s3[125], ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, new_AGEMA_signal_2237, MixColumns_line1_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U16 ( .a ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .b ({new_AGEMA_signal_2272, new_AGEMA_signal_2271, new_AGEMA_signal_2270, MixColumns_line1_S13[5]}), .c ({new_AGEMA_signal_2434, new_AGEMA_signal_2433, new_AGEMA_signal_2432, MixColumns_line1_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U15 ( .a ({new_AGEMA_signal_4453, new_AGEMA_signal_4452, new_AGEMA_signal_4451, MixColumns_line1_n10}), .b ({new_AGEMA_signal_2242, new_AGEMA_signal_2241, new_AGEMA_signal_2240, MixColumns_line1_n9}), .c ({new_AGEMA_signal_4561, new_AGEMA_signal_4560, new_AGEMA_signal_4559, MCout[20]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U14 ( .a ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_2242, new_AGEMA_signal_2241, new_AGEMA_signal_2240, MixColumns_line1_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U13 ( .a ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, new_AGEMA_signal_2255, MixColumns_line1_S02_4_}), .b ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, new_AGEMA_signal_2441, MixColumns_line1_S13[4]}), .c ({new_AGEMA_signal_4453, new_AGEMA_signal_4452, new_AGEMA_signal_4451, MixColumns_line1_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U12 ( .a ({new_AGEMA_signal_4456, new_AGEMA_signal_4455, new_AGEMA_signal_4454, MixColumns_line1_n8}), .b ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, new_AGEMA_signal_2243, MixColumns_line1_n7}), .c ({new_AGEMA_signal_4564, new_AGEMA_signal_4563, new_AGEMA_signal_4562, MCout[19]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U11 ( .a ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .b ({ciphertext_s3[123], ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, new_AGEMA_signal_2243, MixColumns_line1_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U10 ( .a ({new_AGEMA_signal_2260, new_AGEMA_signal_2259, new_AGEMA_signal_2258, MixColumns_line1_S02_3_}), .b ({new_AGEMA_signal_2446, new_AGEMA_signal_2445, new_AGEMA_signal_2444, MixColumns_line1_S13[3]}), .c ({new_AGEMA_signal_4456, new_AGEMA_signal_4455, new_AGEMA_signal_4454, MixColumns_line1_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U9 ( .a ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, new_AGEMA_signal_2435, MixColumns_line1_n6}), .b ({new_AGEMA_signal_2248, new_AGEMA_signal_2247, new_AGEMA_signal_2246, MixColumns_line1_n5}), .c ({new_AGEMA_signal_4459, new_AGEMA_signal_4458, new_AGEMA_signal_4457, MCout[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U8 ( .a ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_2248, new_AGEMA_signal_2247, new_AGEMA_signal_2246, MixColumns_line1_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U7 ( .a ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .b ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, new_AGEMA_signal_2273, MixColumns_line1_S13[2]}), .c ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, new_AGEMA_signal_2435, MixColumns_line1_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U6 ( .a ({new_AGEMA_signal_4462, new_AGEMA_signal_4461, new_AGEMA_signal_4460, MixColumns_line1_n4}), .b ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, new_AGEMA_signal_2249, MixColumns_line1_n3}), .c ({new_AGEMA_signal_4567, new_AGEMA_signal_4566, new_AGEMA_signal_4565, MCout[17]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U5 ( .a ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .b ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, new_AGEMA_signal_2249, MixColumns_line1_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U4 ( .a ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, new_AGEMA_signal_2261, MixColumns_line1_S02_1_}), .b ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, new_AGEMA_signal_2447, MixColumns_line1_S13[1]}), .c ({new_AGEMA_signal_4462, new_AGEMA_signal_4461, new_AGEMA_signal_4460, MixColumns_line1_n4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U3 ( .a ({new_AGEMA_signal_2440, new_AGEMA_signal_2439, new_AGEMA_signal_2438, MixColumns_line1_n2}), .b ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, new_AGEMA_signal_2252, MixColumns_line1_n1}), .c ({new_AGEMA_signal_4465, new_AGEMA_signal_4464, new_AGEMA_signal_4463, MCout[16]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U2 ( .a ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .b ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, new_AGEMA_signal_2252, MixColumns_line1_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_U1 ( .a ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({new_AGEMA_signal_2278, new_AGEMA_signal_2277, new_AGEMA_signal_2276, MixColumns_line1_S13[0]}), .c ({new_AGEMA_signal_2440, new_AGEMA_signal_2439, new_AGEMA_signal_2438, MixColumns_line1_n2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_timesTWO_U3 ( .a ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s3[91], ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, new_AGEMA_signal_2255, MixColumns_line1_S02_4_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_timesTWO_U2 ( .a ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_2260, new_AGEMA_signal_2259, new_AGEMA_signal_2258, MixColumns_line1_S02_3_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_timesTWO_U1 ( .a ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, new_AGEMA_signal_2261, MixColumns_line1_S02_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_timesTHREE_U8 ( .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .c ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, new_AGEMA_signal_2264, MixColumns_line1_S13[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_timesTHREE_U7 ( .a ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, new_AGEMA_signal_2267, MixColumns_line1_S13[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_timesTHREE_U6 ( .a ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_2272, new_AGEMA_signal_2271, new_AGEMA_signal_2270, MixColumns_line1_S13[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_timesTHREE_U5 ( .a ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, new_AGEMA_signal_2279, MixColumns_line1_timesTHREE_input2[4]}), .c ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, new_AGEMA_signal_2441, MixColumns_line1_S13[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_timesTHREE_U4 ( .a ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_2284, new_AGEMA_signal_2283, new_AGEMA_signal_2282, MixColumns_line1_timesTHREE_input2[3]}), .c ({new_AGEMA_signal_2446, new_AGEMA_signal_2445, new_AGEMA_signal_2444, MixColumns_line1_S13[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_timesTHREE_U3 ( .a ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, new_AGEMA_signal_2273, MixColumns_line1_S13[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_timesTHREE_U2 ( .a ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .b ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, new_AGEMA_signal_2285, MixColumns_line1_timesTHREE_input2[1]}), .c ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, new_AGEMA_signal_2447, MixColumns_line1_S13[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_timesTHREE_U1 ( .a ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .c ({new_AGEMA_signal_2278, new_AGEMA_signal_2277, new_AGEMA_signal_2276, MixColumns_line1_S13[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_timesTHREE_timesTWO_U3 ( .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, new_AGEMA_signal_2279, MixColumns_line1_timesTHREE_input2[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_timesTHREE_timesTWO_U2 ( .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_2284, new_AGEMA_signal_2283, new_AGEMA_signal_2282, MixColumns_line1_timesTHREE_input2[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line1_timesTHREE_timesTWO_U1 ( .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, new_AGEMA_signal_2285, MixColumns_line1_timesTHREE_input2[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U24 ( .a ({new_AGEMA_signal_2452, new_AGEMA_signal_2451, new_AGEMA_signal_2450, MixColumns_line2_n16}), .b ({new_AGEMA_signal_2290, new_AGEMA_signal_2289, new_AGEMA_signal_2288, MixColumns_line2_n15}), .c ({new_AGEMA_signal_4468, new_AGEMA_signal_4467, new_AGEMA_signal_4466, MCout[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U23 ( .a ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .c ({new_AGEMA_signal_2290, new_AGEMA_signal_2289, new_AGEMA_signal_2288, MixColumns_line2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U22 ( .a ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, new_AGEMA_signal_2321, MixColumns_line2_S13[7]}), .c ({new_AGEMA_signal_2452, new_AGEMA_signal_2451, new_AGEMA_signal_2450, MixColumns_line2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U21 ( .a ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, new_AGEMA_signal_2453, MixColumns_line2_n14}), .b ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, new_AGEMA_signal_2291, MixColumns_line2_n13}), .c ({new_AGEMA_signal_4471, new_AGEMA_signal_4470, new_AGEMA_signal_4469, MCout[14]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U20 ( .a ({ciphertext_s3[126], ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s3[94], ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .c ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, new_AGEMA_signal_2291, MixColumns_line2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U19 ( .a ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .b ({new_AGEMA_signal_2326, new_AGEMA_signal_2325, new_AGEMA_signal_2324, MixColumns_line2_S13[6]}), .c ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, new_AGEMA_signal_2453, MixColumns_line2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U18 ( .a ({new_AGEMA_signal_2458, new_AGEMA_signal_2457, new_AGEMA_signal_2456, MixColumns_line2_n12}), .b ({new_AGEMA_signal_2296, new_AGEMA_signal_2295, new_AGEMA_signal_2294, MixColumns_line2_n11}), .c ({new_AGEMA_signal_4474, new_AGEMA_signal_4473, new_AGEMA_signal_4472, MCout[13]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U17 ( .a ({ciphertext_s3[125], ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s3[93], ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_2296, new_AGEMA_signal_2295, new_AGEMA_signal_2294, MixColumns_line2_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U16 ( .a ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, new_AGEMA_signal_2327, MixColumns_line2_S13[5]}), .c ({new_AGEMA_signal_2458, new_AGEMA_signal_2457, new_AGEMA_signal_2456, MixColumns_line2_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U15 ( .a ({new_AGEMA_signal_4477, new_AGEMA_signal_4476, new_AGEMA_signal_4475, MixColumns_line2_n10}), .b ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, new_AGEMA_signal_2297, MixColumns_line2_n9}), .c ({new_AGEMA_signal_4570, new_AGEMA_signal_4569, new_AGEMA_signal_4568, MCout[12]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U14 ( .a ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, new_AGEMA_signal_2297, MixColumns_line2_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U13 ( .a ({new_AGEMA_signal_2314, new_AGEMA_signal_2313, new_AGEMA_signal_2312, MixColumns_line2_S02_4_}), .b ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, new_AGEMA_signal_2465, MixColumns_line2_S13[4]}), .c ({new_AGEMA_signal_4477, new_AGEMA_signal_4476, new_AGEMA_signal_4475, MixColumns_line2_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U12 ( .a ({new_AGEMA_signal_4480, new_AGEMA_signal_4479, new_AGEMA_signal_4478, MixColumns_line2_n8}), .b ({new_AGEMA_signal_2302, new_AGEMA_signal_2301, new_AGEMA_signal_2300, MixColumns_line2_n7}), .c ({new_AGEMA_signal_4573, new_AGEMA_signal_4572, new_AGEMA_signal_4571, MCout[11]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U11 ( .a ({ciphertext_s3[123], ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}), .b ({ciphertext_s3[91], ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_2302, new_AGEMA_signal_2301, new_AGEMA_signal_2300, MixColumns_line2_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U10 ( .a ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, new_AGEMA_signal_2315, MixColumns_line2_S02_3_}), .b ({new_AGEMA_signal_2470, new_AGEMA_signal_2469, new_AGEMA_signal_2468, MixColumns_line2_S13[3]}), .c ({new_AGEMA_signal_4480, new_AGEMA_signal_4479, new_AGEMA_signal_4478, MixColumns_line2_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U9 ( .a ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, new_AGEMA_signal_2459, MixColumns_line2_n6}), .b ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, new_AGEMA_signal_2303, MixColumns_line2_n5}), .c ({new_AGEMA_signal_4483, new_AGEMA_signal_4482, new_AGEMA_signal_4481, MCout[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U8 ( .a ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, new_AGEMA_signal_2303, MixColumns_line2_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U7 ( .a ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .b ({new_AGEMA_signal_2332, new_AGEMA_signal_2331, new_AGEMA_signal_2330, MixColumns_line2_S13[2]}), .c ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, new_AGEMA_signal_2459, MixColumns_line2_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U6 ( .a ({new_AGEMA_signal_4486, new_AGEMA_signal_4485, new_AGEMA_signal_4484, MixColumns_line2_n4}), .b ({new_AGEMA_signal_2308, new_AGEMA_signal_2307, new_AGEMA_signal_2306, MixColumns_line2_n3}), .c ({new_AGEMA_signal_4576, new_AGEMA_signal_4575, new_AGEMA_signal_4574, MCout[9]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U5 ( .a ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .b ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_2308, new_AGEMA_signal_2307, new_AGEMA_signal_2306, MixColumns_line2_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U4 ( .a ({new_AGEMA_signal_2320, new_AGEMA_signal_2319, new_AGEMA_signal_2318, MixColumns_line2_S02_1_}), .b ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, new_AGEMA_signal_2471, MixColumns_line2_S13[1]}), .c ({new_AGEMA_signal_4486, new_AGEMA_signal_4485, new_AGEMA_signal_4484, MixColumns_line2_n4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U3 ( .a ({new_AGEMA_signal_2464, new_AGEMA_signal_2463, new_AGEMA_signal_2462, MixColumns_line2_n2}), .b ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, new_AGEMA_signal_2309, MixColumns_line2_n1}), .c ({new_AGEMA_signal_4489, new_AGEMA_signal_4488, new_AGEMA_signal_4487, MCout[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U2 ( .a ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .b ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, new_AGEMA_signal_2309, MixColumns_line2_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_U1 ( .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, new_AGEMA_signal_2333, MixColumns_line2_S13[0]}), .c ({new_AGEMA_signal_2464, new_AGEMA_signal_2463, new_AGEMA_signal_2462, MixColumns_line2_n2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_timesTWO_U3 ( .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_2314, new_AGEMA_signal_2313, new_AGEMA_signal_2312, MixColumns_line2_S02_4_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_timesTWO_U2 ( .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, new_AGEMA_signal_2315, MixColumns_line2_S02_3_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_timesTWO_U1 ( .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_2320, new_AGEMA_signal_2319, new_AGEMA_signal_2318, MixColumns_line2_S02_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_timesTHREE_U8 ( .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .c ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, new_AGEMA_signal_2321, MixColumns_line2_S13[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_timesTHREE_U7 ( .a ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_2326, new_AGEMA_signal_2325, new_AGEMA_signal_2324, MixColumns_line2_S13[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_timesTHREE_U6 ( .a ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, new_AGEMA_signal_2327, MixColumns_line2_S13[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_timesTHREE_U5 ( .a ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_2338, new_AGEMA_signal_2337, new_AGEMA_signal_2336, MixColumns_line2_timesTHREE_input2[4]}), .c ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, new_AGEMA_signal_2465, MixColumns_line2_S13[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_timesTHREE_U4 ( .a ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, new_AGEMA_signal_2339, MixColumns_line2_timesTHREE_input2[3]}), .c ({new_AGEMA_signal_2470, new_AGEMA_signal_2469, new_AGEMA_signal_2468, MixColumns_line2_S13[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_timesTHREE_U3 ( .a ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_2332, new_AGEMA_signal_2331, new_AGEMA_signal_2330, MixColumns_line2_S13[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_timesTHREE_U2 ( .a ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .b ({new_AGEMA_signal_2344, new_AGEMA_signal_2343, new_AGEMA_signal_2342, MixColumns_line2_timesTHREE_input2[1]}), .c ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, new_AGEMA_signal_2471, MixColumns_line2_S13[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_timesTHREE_U1 ( .a ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .c ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, new_AGEMA_signal_2333, MixColumns_line2_S13[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_timesTHREE_timesTWO_U3 ( .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_2338, new_AGEMA_signal_2337, new_AGEMA_signal_2336, MixColumns_line2_timesTHREE_input2[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_timesTHREE_timesTWO_U2 ( .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, new_AGEMA_signal_2339, MixColumns_line2_timesTHREE_input2[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line2_timesTHREE_timesTWO_U1 ( .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_2344, new_AGEMA_signal_2343, new_AGEMA_signal_2342, MixColumns_line2_timesTHREE_input2[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U24 ( .a ({new_AGEMA_signal_2476, new_AGEMA_signal_2475, new_AGEMA_signal_2474, MixColumns_line3_n16}), .b ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, new_AGEMA_signal_2345, MixColumns_line3_n15}), .c ({new_AGEMA_signal_4492, new_AGEMA_signal_4491, new_AGEMA_signal_4490, MCout[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U23 ( .a ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .c ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, new_AGEMA_signal_2345, MixColumns_line3_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U22 ( .a ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_2380, new_AGEMA_signal_2379, new_AGEMA_signal_2378, MixColumns_line3_S13[7]}), .c ({new_AGEMA_signal_2476, new_AGEMA_signal_2475, new_AGEMA_signal_2474, MixColumns_line3_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U21 ( .a ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, new_AGEMA_signal_2477, MixColumns_line3_n14}), .b ({new_AGEMA_signal_2350, new_AGEMA_signal_2349, new_AGEMA_signal_2348, MixColumns_line3_n13}), .c ({new_AGEMA_signal_4495, new_AGEMA_signal_4494, new_AGEMA_signal_4493, MCout[6]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U20 ( .a ({ciphertext_s3[94], ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .c ({new_AGEMA_signal_2350, new_AGEMA_signal_2349, new_AGEMA_signal_2348, MixColumns_line3_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U19 ( .a ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .b ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, new_AGEMA_signal_2381, MixColumns_line3_S13[6]}), .c ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, new_AGEMA_signal_2477, MixColumns_line3_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U18 ( .a ({new_AGEMA_signal_2482, new_AGEMA_signal_2481, new_AGEMA_signal_2480, MixColumns_line3_n12}), .b ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, new_AGEMA_signal_2351, MixColumns_line3_n11}), .c ({new_AGEMA_signal_4498, new_AGEMA_signal_4497, new_AGEMA_signal_4496, MCout[5]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U17 ( .a ({ciphertext_s3[93], ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, new_AGEMA_signal_2351, MixColumns_line3_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U16 ( .a ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_2386, new_AGEMA_signal_2385, new_AGEMA_signal_2384, MixColumns_line3_S13[5]}), .c ({new_AGEMA_signal_2482, new_AGEMA_signal_2481, new_AGEMA_signal_2480, MixColumns_line3_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U15 ( .a ({new_AGEMA_signal_4501, new_AGEMA_signal_4500, new_AGEMA_signal_4499, MixColumns_line3_n10}), .b ({new_AGEMA_signal_2356, new_AGEMA_signal_2355, new_AGEMA_signal_2354, MixColumns_line3_n9}), .c ({new_AGEMA_signal_4579, new_AGEMA_signal_4578, new_AGEMA_signal_4577, MCout[4]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U14 ( .a ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_2356, new_AGEMA_signal_2355, new_AGEMA_signal_2354, MixColumns_line3_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U13 ( .a ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, new_AGEMA_signal_2369, MixColumns_line3_S02_4_}), .b ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, new_AGEMA_signal_2489, MixColumns_line3_S13[4]}), .c ({new_AGEMA_signal_4501, new_AGEMA_signal_4500, new_AGEMA_signal_4499, MixColumns_line3_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U12 ( .a ({new_AGEMA_signal_4504, new_AGEMA_signal_4503, new_AGEMA_signal_4502, MixColumns_line3_n8}), .b ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, new_AGEMA_signal_2357, MixColumns_line3_n7}), .c ({new_AGEMA_signal_4582, new_AGEMA_signal_4581, new_AGEMA_signal_4580, MCout[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U11 ( .a ({ciphertext_s3[91], ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}), .b ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, new_AGEMA_signal_2357, MixColumns_line3_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U10 ( .a ({new_AGEMA_signal_2374, new_AGEMA_signal_2373, new_AGEMA_signal_2372, MixColumns_line3_S02_3_}), .b ({new_AGEMA_signal_2494, new_AGEMA_signal_2493, new_AGEMA_signal_2492, MixColumns_line3_S13[3]}), .c ({new_AGEMA_signal_4504, new_AGEMA_signal_4503, new_AGEMA_signal_4502, MixColumns_line3_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U9 ( .a ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, new_AGEMA_signal_2483, MixColumns_line3_n6}), .b ({new_AGEMA_signal_2362, new_AGEMA_signal_2361, new_AGEMA_signal_2360, MixColumns_line3_n5}), .c ({new_AGEMA_signal_4507, new_AGEMA_signal_4506, new_AGEMA_signal_4505, MCout[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U8 ( .a ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_2362, new_AGEMA_signal_2361, new_AGEMA_signal_2360, MixColumns_line3_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U7 ( .a ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .b ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, new_AGEMA_signal_2387, MixColumns_line3_S13[2]}), .c ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, new_AGEMA_signal_2483, MixColumns_line3_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U6 ( .a ({new_AGEMA_signal_4510, new_AGEMA_signal_4509, new_AGEMA_signal_4508, MixColumns_line3_n4}), .b ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, new_AGEMA_signal_2363, MixColumns_line3_n3}), .c ({new_AGEMA_signal_4585, new_AGEMA_signal_4584, new_AGEMA_signal_4583, MCout[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U5 ( .a ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .b ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, new_AGEMA_signal_2363, MixColumns_line3_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U4 ( .a ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, new_AGEMA_signal_2375, MixColumns_line3_S02_1_}), .b ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, new_AGEMA_signal_2495, MixColumns_line3_S13[1]}), .c ({new_AGEMA_signal_4510, new_AGEMA_signal_4509, new_AGEMA_signal_4508, MixColumns_line3_n4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U3 ( .a ({new_AGEMA_signal_2488, new_AGEMA_signal_2487, new_AGEMA_signal_2486, MixColumns_line3_n2}), .b ({new_AGEMA_signal_2368, new_AGEMA_signal_2367, new_AGEMA_signal_2366, MixColumns_line3_n1}), .c ({new_AGEMA_signal_4513, new_AGEMA_signal_4512, new_AGEMA_signal_4511, MCout[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U2 ( .a ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_2368, new_AGEMA_signal_2367, new_AGEMA_signal_2366, MixColumns_line3_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_U1 ( .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_2392, new_AGEMA_signal_2391, new_AGEMA_signal_2390, MixColumns_line3_S13[0]}), .c ({new_AGEMA_signal_2488, new_AGEMA_signal_2487, new_AGEMA_signal_2486, MixColumns_line3_n2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_timesTWO_U3 ( .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, new_AGEMA_signal_2369, MixColumns_line3_S02_4_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_timesTWO_U2 ( .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_2374, new_AGEMA_signal_2373, new_AGEMA_signal_2372, MixColumns_line3_S02_3_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_timesTWO_U1 ( .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, new_AGEMA_signal_2375, MixColumns_line3_S02_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_timesTHREE_U8 ( .a ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s3[126], ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .c ({new_AGEMA_signal_2380, new_AGEMA_signal_2379, new_AGEMA_signal_2378, MixColumns_line3_S13[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_timesTHREE_U7 ( .a ({ciphertext_s3[126], ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s3[125], ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, new_AGEMA_signal_2381, MixColumns_line3_S13[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_timesTHREE_U6 ( .a ({ciphertext_s3[125], ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_2386, new_AGEMA_signal_2385, new_AGEMA_signal_2384, MixColumns_line3_S13[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_timesTHREE_U5 ( .a ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .b ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, new_AGEMA_signal_2393, MixColumns_line3_timesTHREE_input2_4_}), .c ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, new_AGEMA_signal_2489, MixColumns_line3_S13[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_timesTHREE_U4 ( .a ({ciphertext_s3[123], ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}), .b ({new_AGEMA_signal_2398, new_AGEMA_signal_2397, new_AGEMA_signal_2396, MixColumns_line3_timesTHREE_input2_3_}), .c ({new_AGEMA_signal_2494, new_AGEMA_signal_2493, new_AGEMA_signal_2492, MixColumns_line3_S13[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_timesTHREE_U3 ( .a ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, new_AGEMA_signal_2387, MixColumns_line3_S13[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_timesTHREE_U2 ( .a ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .b ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, new_AGEMA_signal_2399, MixColumns_line3_timesTHREE_input2_1_}), .c ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, new_AGEMA_signal_2495, MixColumns_line3_S13[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_timesTHREE_U1 ( .a ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .b ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .c ({new_AGEMA_signal_2392, new_AGEMA_signal_2391, new_AGEMA_signal_2390, MixColumns_line3_S13[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_timesTHREE_timesTWO_U3 ( .a ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s3[123], ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, new_AGEMA_signal_2393, MixColumns_line3_timesTHREE_input2_4_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_timesTHREE_timesTWO_U2 ( .a ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_2398, new_AGEMA_signal_2397, new_AGEMA_signal_2396, MixColumns_line3_timesTHREE_input2_3_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumns_line3_timesTHREE_timesTWO_U1 ( .a ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, new_AGEMA_signal_2399, MixColumns_line3_timesTHREE_input2_1_}) ) ;
    NOR2_X1 calcRCon_U46 ( .A1 (calcRCon_n11), .A2 (calcRCon_n38), .ZN (roundConstant[7]) ) ;
    NOR2_X1 calcRCon_U45 ( .A1 (calcRCon_n16), .A2 (calcRCon_n38), .ZN (roundConstant[6]) ) ;
    AND2_X1 calcRCon_U44 ( .A1 (calcRCon_s_current_state_5_), .A2 (enRCon), .ZN (roundConstant[5]) ) ;
    AND2_X1 calcRCon_U43 ( .A1 (calcRCon_s_current_state_4_), .A2 (enRCon), .ZN (roundConstant[4]) ) ;
    NOR2_X1 calcRCon_U42 ( .A1 (calcRCon_n15), .A2 (calcRCon_n38), .ZN (roundConstant[3]) ) ;
    NOR2_X1 calcRCon_U41 ( .A1 (calcRCon_n12), .A2 (calcRCon_n38), .ZN (roundConstant[2]) ) ;
    NOR2_X1 calcRCon_U40 ( .A1 (calcRCon_n14), .A2 (calcRCon_n38), .ZN (roundConstant[1]) ) ;
    NOR2_X1 calcRCon_U39 ( .A1 (calcRCon_n13), .A2 (calcRCon_n38), .ZN (roundConstant[0]) ) ;
    INV_X1 calcRCon_U38 ( .A (enRCon), .ZN (calcRCon_n38) ) ;
    NAND2_X1 calcRCon_U37 ( .A1 (calcRCon_n37), .A2 (calcRCon_n36), .ZN (notFirst) ) ;
    NOR2_X1 calcRCon_U36 ( .A1 (calcRCon_n35), .A2 (calcRCon_n34), .ZN (calcRCon_n36) ) ;
    NAND2_X1 calcRCon_U35 ( .A1 (calcRCon_n33), .A2 (calcRCon_n32), .ZN (calcRCon_n34) ) ;
    NOR2_X1 calcRCon_U34 ( .A1 (calcRCon_s_current_state_1_), .A2 (calcRCon_n15), .ZN (calcRCon_n32) ) ;
    NOR2_X1 calcRCon_U33 ( .A1 (calcRCon_s_current_state_6_), .A2 (calcRCon_n13), .ZN (calcRCon_n33) ) ;
    NAND2_X1 calcRCon_U32 ( .A1 (calcRCon_s_current_state_2_), .A2 (calcRCon_n3), .ZN (calcRCon_n35) ) ;
    NOR2_X1 calcRCon_U31 ( .A1 (calcRCon_s_current_state_4_), .A2 (calcRCon_s_current_state_5_), .ZN (calcRCon_n37) ) ;
    NAND2_X1 calcRCon_U30 ( .A1 (nReset), .A2 (calcRCon_n31), .ZN (calcRCon_n51) ) ;
    MUX2_X1 calcRCon_U29 ( .S (calcRCon_n5), .A (calcRCon_n11), .B (calcRCon_n13), .Z (calcRCon_n31) ) ;
    NAND2_X1 calcRCon_U28 ( .A1 (calcRCon_n30), .A2 (calcRCon_n29), .ZN (calcRCon_n50) ) ;
    NAND2_X1 calcRCon_U27 ( .A1 (calcRCon_n28), .A2 (calcRCon_s_current_state_1_), .ZN (calcRCon_n29) ) ;
    NAND2_X1 calcRCon_U26 ( .A1 (calcRCon_n27), .A2 (calcRCon_n26), .ZN (calcRCon_n30) ) ;
    XOR2_X1 calcRCon_U25 ( .A (calcRCon_s_current_state_0_), .B (calcRCon_n3), .Z (calcRCon_n27) ) ;
    NAND2_X1 calcRCon_U24 ( .A1 (nReset), .A2 (calcRCon_n25), .ZN (calcRCon_n49) ) ;
    MUX2_X1 calcRCon_U23 ( .S (calcRCon_n5), .A (calcRCon_n14), .B (calcRCon_n12), .Z (calcRCon_n25) ) ;
    NAND2_X1 calcRCon_U22 ( .A1 (nReset), .A2 (calcRCon_n24), .ZN (calcRCon_n48) ) ;
    MUX2_X1 calcRCon_U21 ( .S (calcRCon_n5), .A (calcRCon_n23), .B (calcRCon_n15), .Z (calcRCon_n24) ) ;
    XNOR2_X1 calcRCon_U20 ( .A (calcRCon_n3), .B (calcRCon_s_current_state_2_), .ZN (calcRCon_n23) ) ;
    NAND2_X1 calcRCon_U19 ( .A1 (calcRCon_n22), .A2 (calcRCon_n21), .ZN (calcRCon_n47) ) ;
    NAND2_X1 calcRCon_U18 ( .A1 (calcRCon_s_current_state_4_), .A2 (calcRCon_n28), .ZN (calcRCon_n21) ) ;
    NAND2_X1 calcRCon_U17 ( .A1 (calcRCon_n20), .A2 (calcRCon_n26), .ZN (calcRCon_n22) ) ;
    XOR2_X1 calcRCon_U16 ( .A (calcRCon_n15), .B (calcRCon_n11), .Z (calcRCon_n20) ) ;
    NAND2_X1 calcRCon_U15 ( .A1 (calcRCon_n19), .A2 (calcRCon_n18), .ZN (calcRCon_n46) ) ;
    NAND2_X1 calcRCon_U14 ( .A1 (calcRCon_s_current_state_4_), .A2 (calcRCon_n26), .ZN (calcRCon_n18) ) ;
    NAND2_X1 calcRCon_U13 ( .A1 (calcRCon_s_current_state_5_), .A2 (calcRCon_n28), .ZN (calcRCon_n19) ) ;
    NAND2_X1 calcRCon_U12 ( .A1 (calcRCon_n17), .A2 (calcRCon_n10), .ZN (calcRCon_n45) ) ;
    NAND2_X1 calcRCon_U11 ( .A1 (calcRCon_s_current_state_5_), .A2 (calcRCon_n26), .ZN (calcRCon_n10) ) ;
    NOR2_X1 calcRCon_U10 ( .A1 (calcRCon_n5), .A2 (calcRCon_n6), .ZN (calcRCon_n26) ) ;
    NAND2_X1 calcRCon_U9 ( .A1 (calcRCon_s_current_state_6_), .A2 (calcRCon_n28), .ZN (calcRCon_n17) ) ;
    NOR2_X1 calcRCon_U8 ( .A1 (selSR), .A2 (calcRCon_n6), .ZN (calcRCon_n28) ) ;
    NAND2_X1 calcRCon_U7 ( .A1 (nReset), .A2 (calcRCon_n9), .ZN (calcRCon_n44) ) ;
    MUX2_X1 calcRCon_U6 ( .S (calcRCon_n5), .A (calcRCon_n16), .B (calcRCon_n11), .Z (calcRCon_n9) ) ;
    NAND2_X1 calcRCon_U5 ( .A1 (calcRCon_s_current_state_4_), .A2 (calcRCon_s_current_state_2_), .ZN (calcRCon_n7) ) ;
    NAND2_X1 calcRCon_U4 ( .A1 (calcRCon_s_current_state_1_), .A2 (calcRCon_s_current_state_5_), .ZN (calcRCon_n8) ) ;
    INV_X1 calcRCon_U3 ( .A (nReset), .ZN (calcRCon_n6) ) ;
    INV_X1 calcRCon_U2 ( .A (selSR), .ZN (calcRCon_n5) ) ;
    NOR2_X1 calcRCon_U1 ( .A1 (calcRCon_n8), .A2 (calcRCon_n7), .ZN (intFinal) ) ;
    INV_X1 calcRCon_s_current_state_reg_0__U1 ( .A (calcRCon_s_current_state_0_), .ZN (calcRCon_n13) ) ;
    INV_X1 calcRCon_s_current_state_reg_1__U1 ( .A (calcRCon_s_current_state_1_), .ZN (calcRCon_n14) ) ;
    INV_X1 calcRCon_s_current_state_reg_2__U1 ( .A (calcRCon_s_current_state_2_), .ZN (calcRCon_n12) ) ;
    INV_X1 calcRCon_s_current_state_reg_3__U1 ( .A (calcRCon_s_current_state_3_), .ZN (calcRCon_n15) ) ;
    INV_X1 calcRCon_s_current_state_reg_6__U1 ( .A (calcRCon_s_current_state_6_), .ZN (calcRCon_n16) ) ;
    INV_X1 calcRCon_s_current_state_reg_7__U1 ( .A (calcRCon_n3), .ZN (calcRCon_n11) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_SboxIn_mux_inst_0_U1 ( .s (selMC), .b ({new_AGEMA_signal_1990, new_AGEMA_signal_1989, new_AGEMA_signal_1988, StateOutXORroundKey[0]}), .a ({new_AGEMA_signal_3727, new_AGEMA_signal_3726, new_AGEMA_signal_3725, keySBIn[0]}), .c ({new_AGEMA_signal_4516, new_AGEMA_signal_4515, new_AGEMA_signal_4514, SboxIn[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_SboxIn_mux_inst_1_U1 ( .s (selMC), .b ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, new_AGEMA_signal_1997, StateOutXORroundKey[1]}), .a ({new_AGEMA_signal_3736, new_AGEMA_signal_3735, new_AGEMA_signal_3734, keySBIn[1]}), .c ({new_AGEMA_signal_4519, new_AGEMA_signal_4518, new_AGEMA_signal_4517, SboxIn[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_SboxIn_mux_inst_2_U1 ( .s (selMC), .b ({new_AGEMA_signal_2008, new_AGEMA_signal_2007, new_AGEMA_signal_2006, StateOutXORroundKey[2]}), .a ({new_AGEMA_signal_3745, new_AGEMA_signal_3744, new_AGEMA_signal_3743, keySBIn[2]}), .c ({new_AGEMA_signal_4522, new_AGEMA_signal_4521, new_AGEMA_signal_4520, SboxIn[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_SboxIn_mux_inst_3_U1 ( .s (selMC), .b ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, new_AGEMA_signal_2015, StateOutXORroundKey[3]}), .a ({new_AGEMA_signal_3754, new_AGEMA_signal_3753, new_AGEMA_signal_3752, keySBIn[3]}), .c ({new_AGEMA_signal_4525, new_AGEMA_signal_4524, new_AGEMA_signal_4523, SboxIn[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_SboxIn_mux_inst_4_U1 ( .s (selMC), .b ({new_AGEMA_signal_2026, new_AGEMA_signal_2025, new_AGEMA_signal_2024, StateOutXORroundKey[4]}), .a ({new_AGEMA_signal_3763, new_AGEMA_signal_3762, new_AGEMA_signal_3761, keySBIn[4]}), .c ({new_AGEMA_signal_4528, new_AGEMA_signal_4527, new_AGEMA_signal_4526, SboxIn[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_SboxIn_mux_inst_5_U1 ( .s (selMC), .b ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, new_AGEMA_signal_2033, StateOutXORroundKey[5]}), .a ({new_AGEMA_signal_3772, new_AGEMA_signal_3771, new_AGEMA_signal_3770, keySBIn[5]}), .c ({new_AGEMA_signal_4531, new_AGEMA_signal_4530, new_AGEMA_signal_4529, SboxIn[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_SboxIn_mux_inst_6_U1 ( .s (selMC), .b ({new_AGEMA_signal_2044, new_AGEMA_signal_2043, new_AGEMA_signal_2042, StateOutXORroundKey[6]}), .a ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, new_AGEMA_signal_3779, keySBIn[6]}), .c ({new_AGEMA_signal_4534, new_AGEMA_signal_4533, new_AGEMA_signal_4532, SboxIn[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_SboxIn_mux_inst_7_U1 ( .s (selMC), .b ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, new_AGEMA_signal_2051, StateOutXORroundKey[7]}), .a ({new_AGEMA_signal_3790, new_AGEMA_signal_3789, new_AGEMA_signal_3788, keySBIn[7]}), .c ({new_AGEMA_signal_4537, new_AGEMA_signal_4536, new_AGEMA_signal_4535, SboxIn[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T1_U1 ( .a ({new_AGEMA_signal_4537, new_AGEMA_signal_4536, new_AGEMA_signal_4535, SboxIn[7]}), .b ({new_AGEMA_signal_4528, new_AGEMA_signal_4527, new_AGEMA_signal_4526, SboxIn[4]}), .c ({new_AGEMA_signal_4588, new_AGEMA_signal_4587, new_AGEMA_signal_4586, Inst_bSbox_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T2_U1 ( .a ({new_AGEMA_signal_4537, new_AGEMA_signal_4536, new_AGEMA_signal_4535, SboxIn[7]}), .b ({new_AGEMA_signal_4522, new_AGEMA_signal_4521, new_AGEMA_signal_4520, SboxIn[2]}), .c ({new_AGEMA_signal_4591, new_AGEMA_signal_4590, new_AGEMA_signal_4589, Inst_bSbox_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T3_U1 ( .a ({new_AGEMA_signal_4537, new_AGEMA_signal_4536, new_AGEMA_signal_4535, SboxIn[7]}), .b ({new_AGEMA_signal_4519, new_AGEMA_signal_4518, new_AGEMA_signal_4517, SboxIn[1]}), .c ({new_AGEMA_signal_4594, new_AGEMA_signal_4593, new_AGEMA_signal_4592, Inst_bSbox_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T4_U1 ( .a ({new_AGEMA_signal_4528, new_AGEMA_signal_4527, new_AGEMA_signal_4526, SboxIn[4]}), .b ({new_AGEMA_signal_4522, new_AGEMA_signal_4521, new_AGEMA_signal_4520, SboxIn[2]}), .c ({new_AGEMA_signal_4597, new_AGEMA_signal_4596, new_AGEMA_signal_4595, Inst_bSbox_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T5_U1 ( .a ({new_AGEMA_signal_4525, new_AGEMA_signal_4524, new_AGEMA_signal_4523, SboxIn[3]}), .b ({new_AGEMA_signal_4519, new_AGEMA_signal_4518, new_AGEMA_signal_4517, SboxIn[1]}), .c ({new_AGEMA_signal_4600, new_AGEMA_signal_4599, new_AGEMA_signal_4598, Inst_bSbox_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T6_U1 ( .a ({new_AGEMA_signal_4588, new_AGEMA_signal_4587, new_AGEMA_signal_4586, Inst_bSbox_T1}), .b ({new_AGEMA_signal_4600, new_AGEMA_signal_4599, new_AGEMA_signal_4598, Inst_bSbox_T5}), .c ({new_AGEMA_signal_5038, new_AGEMA_signal_5037, new_AGEMA_signal_5036, Inst_bSbox_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T7_U1 ( .a ({new_AGEMA_signal_4534, new_AGEMA_signal_4533, new_AGEMA_signal_4532, SboxIn[6]}), .b ({new_AGEMA_signal_4531, new_AGEMA_signal_4530, new_AGEMA_signal_4529, SboxIn[5]}), .c ({new_AGEMA_signal_4603, new_AGEMA_signal_4602, new_AGEMA_signal_4601, Inst_bSbox_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T8_U1 ( .a ({new_AGEMA_signal_4516, new_AGEMA_signal_4515, new_AGEMA_signal_4514, SboxIn[0]}), .b ({new_AGEMA_signal_5038, new_AGEMA_signal_5037, new_AGEMA_signal_5036, Inst_bSbox_T6}), .c ({new_AGEMA_signal_5134, new_AGEMA_signal_5133, new_AGEMA_signal_5132, Inst_bSbox_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T9_U1 ( .a ({new_AGEMA_signal_4516, new_AGEMA_signal_4515, new_AGEMA_signal_4514, SboxIn[0]}), .b ({new_AGEMA_signal_4603, new_AGEMA_signal_4602, new_AGEMA_signal_4601, Inst_bSbox_T7}), .c ({new_AGEMA_signal_5041, new_AGEMA_signal_5040, new_AGEMA_signal_5039, Inst_bSbox_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T10_U1 ( .a ({new_AGEMA_signal_5038, new_AGEMA_signal_5037, new_AGEMA_signal_5036, Inst_bSbox_T6}), .b ({new_AGEMA_signal_4603, new_AGEMA_signal_4602, new_AGEMA_signal_4601, Inst_bSbox_T7}), .c ({new_AGEMA_signal_5137, new_AGEMA_signal_5136, new_AGEMA_signal_5135, Inst_bSbox_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T11_U1 ( .a ({new_AGEMA_signal_4534, new_AGEMA_signal_4533, new_AGEMA_signal_4532, SboxIn[6]}), .b ({new_AGEMA_signal_4522, new_AGEMA_signal_4521, new_AGEMA_signal_4520, SboxIn[2]}), .c ({new_AGEMA_signal_4606, new_AGEMA_signal_4605, new_AGEMA_signal_4604, Inst_bSbox_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T12_U1 ( .a ({new_AGEMA_signal_4531, new_AGEMA_signal_4530, new_AGEMA_signal_4529, SboxIn[5]}), .b ({new_AGEMA_signal_4522, new_AGEMA_signal_4521, new_AGEMA_signal_4520, SboxIn[2]}), .c ({new_AGEMA_signal_4609, new_AGEMA_signal_4608, new_AGEMA_signal_4607, Inst_bSbox_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T13_U1 ( .a ({new_AGEMA_signal_4594, new_AGEMA_signal_4593, new_AGEMA_signal_4592, Inst_bSbox_T3}), .b ({new_AGEMA_signal_4597, new_AGEMA_signal_4596, new_AGEMA_signal_4595, Inst_bSbox_T4}), .c ({new_AGEMA_signal_5044, new_AGEMA_signal_5043, new_AGEMA_signal_5042, Inst_bSbox_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T14_U1 ( .a ({new_AGEMA_signal_5038, new_AGEMA_signal_5037, new_AGEMA_signal_5036, Inst_bSbox_T6}), .b ({new_AGEMA_signal_4606, new_AGEMA_signal_4605, new_AGEMA_signal_4604, Inst_bSbox_T11}), .c ({new_AGEMA_signal_5140, new_AGEMA_signal_5139, new_AGEMA_signal_5138, Inst_bSbox_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T15_U1 ( .a ({new_AGEMA_signal_4600, new_AGEMA_signal_4599, new_AGEMA_signal_4598, Inst_bSbox_T5}), .b ({new_AGEMA_signal_4606, new_AGEMA_signal_4605, new_AGEMA_signal_4604, Inst_bSbox_T11}), .c ({new_AGEMA_signal_5047, new_AGEMA_signal_5046, new_AGEMA_signal_5045, Inst_bSbox_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T16_U1 ( .a ({new_AGEMA_signal_4600, new_AGEMA_signal_4599, new_AGEMA_signal_4598, Inst_bSbox_T5}), .b ({new_AGEMA_signal_4609, new_AGEMA_signal_4608, new_AGEMA_signal_4607, Inst_bSbox_T12}), .c ({new_AGEMA_signal_5050, new_AGEMA_signal_5049, new_AGEMA_signal_5048, Inst_bSbox_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T17_U1 ( .a ({new_AGEMA_signal_5041, new_AGEMA_signal_5040, new_AGEMA_signal_5039, Inst_bSbox_T9}), .b ({new_AGEMA_signal_5050, new_AGEMA_signal_5049, new_AGEMA_signal_5048, Inst_bSbox_T16}), .c ({new_AGEMA_signal_5143, new_AGEMA_signal_5142, new_AGEMA_signal_5141, Inst_bSbox_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T18_U1 ( .a ({new_AGEMA_signal_4528, new_AGEMA_signal_4527, new_AGEMA_signal_4526, SboxIn[4]}), .b ({new_AGEMA_signal_4516, new_AGEMA_signal_4515, new_AGEMA_signal_4514, SboxIn[0]}), .c ({new_AGEMA_signal_4612, new_AGEMA_signal_4611, new_AGEMA_signal_4610, Inst_bSbox_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T19_U1 ( .a ({new_AGEMA_signal_4603, new_AGEMA_signal_4602, new_AGEMA_signal_4601, Inst_bSbox_T7}), .b ({new_AGEMA_signal_4612, new_AGEMA_signal_4611, new_AGEMA_signal_4610, Inst_bSbox_T18}), .c ({new_AGEMA_signal_5053, new_AGEMA_signal_5052, new_AGEMA_signal_5051, Inst_bSbox_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T20_U1 ( .a ({new_AGEMA_signal_4588, new_AGEMA_signal_4587, new_AGEMA_signal_4586, Inst_bSbox_T1}), .b ({new_AGEMA_signal_5053, new_AGEMA_signal_5052, new_AGEMA_signal_5051, Inst_bSbox_T19}), .c ({new_AGEMA_signal_5146, new_AGEMA_signal_5145, new_AGEMA_signal_5144, Inst_bSbox_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T21_U1 ( .a ({new_AGEMA_signal_4519, new_AGEMA_signal_4518, new_AGEMA_signal_4517, SboxIn[1]}), .b ({new_AGEMA_signal_4516, new_AGEMA_signal_4515, new_AGEMA_signal_4514, SboxIn[0]}), .c ({new_AGEMA_signal_4615, new_AGEMA_signal_4614, new_AGEMA_signal_4613, Inst_bSbox_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T22_U1 ( .a ({new_AGEMA_signal_4603, new_AGEMA_signal_4602, new_AGEMA_signal_4601, Inst_bSbox_T7}), .b ({new_AGEMA_signal_4615, new_AGEMA_signal_4614, new_AGEMA_signal_4613, Inst_bSbox_T21}), .c ({new_AGEMA_signal_5056, new_AGEMA_signal_5055, new_AGEMA_signal_5054, Inst_bSbox_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T23_U1 ( .a ({new_AGEMA_signal_4591, new_AGEMA_signal_4590, new_AGEMA_signal_4589, Inst_bSbox_T2}), .b ({new_AGEMA_signal_5056, new_AGEMA_signal_5055, new_AGEMA_signal_5054, Inst_bSbox_T22}), .c ({new_AGEMA_signal_5149, new_AGEMA_signal_5148, new_AGEMA_signal_5147, Inst_bSbox_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T24_U1 ( .a ({new_AGEMA_signal_4591, new_AGEMA_signal_4590, new_AGEMA_signal_4589, Inst_bSbox_T2}), .b ({new_AGEMA_signal_5137, new_AGEMA_signal_5136, new_AGEMA_signal_5135, Inst_bSbox_T10}), .c ({new_AGEMA_signal_5389, new_AGEMA_signal_5388, new_AGEMA_signal_5387, Inst_bSbox_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T25_U1 ( .a ({new_AGEMA_signal_5146, new_AGEMA_signal_5145, new_AGEMA_signal_5144, Inst_bSbox_T20}), .b ({new_AGEMA_signal_5143, new_AGEMA_signal_5142, new_AGEMA_signal_5141, Inst_bSbox_T17}), .c ({new_AGEMA_signal_5392, new_AGEMA_signal_5391, new_AGEMA_signal_5390, Inst_bSbox_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T26_U1 ( .a ({new_AGEMA_signal_4594, new_AGEMA_signal_4593, new_AGEMA_signal_4592, Inst_bSbox_T3}), .b ({new_AGEMA_signal_5050, new_AGEMA_signal_5049, new_AGEMA_signal_5048, Inst_bSbox_T16}), .c ({new_AGEMA_signal_5152, new_AGEMA_signal_5151, new_AGEMA_signal_5150, Inst_bSbox_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_T27_U1 ( .a ({new_AGEMA_signal_4588, new_AGEMA_signal_4587, new_AGEMA_signal_4586, Inst_bSbox_T1}), .b ({new_AGEMA_signal_4609, new_AGEMA_signal_4608, new_AGEMA_signal_4607, Inst_bSbox_T12}), .c ({new_AGEMA_signal_5059, new_AGEMA_signal_5058, new_AGEMA_signal_5057, Inst_bSbox_T27}) ) ;
    INV_X1 nReset_reg_U1 ( .A (nReset), .ZN (n10) ) ;
    ClockGatingController #(9) ClockGatingInst ( .clk (clk), .rst (start), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M1_U1 ( .a ({new_AGEMA_signal_5044, new_AGEMA_signal_5043, new_AGEMA_signal_5042, Inst_bSbox_T13}), .b ({new_AGEMA_signal_5038, new_AGEMA_signal_5037, new_AGEMA_signal_5036, Inst_bSbox_T6}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_5155, new_AGEMA_signal_5154, new_AGEMA_signal_5153, Inst_bSbox_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M2_U1 ( .a ({new_AGEMA_signal_5149, new_AGEMA_signal_5148, new_AGEMA_signal_5147, Inst_bSbox_T23}), .b ({new_AGEMA_signal_5134, new_AGEMA_signal_5133, new_AGEMA_signal_5132, Inst_bSbox_T8}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_5395, new_AGEMA_signal_5394, new_AGEMA_signal_5393, Inst_bSbox_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M3_U1 ( .a ({new_AGEMA_signal_5140, new_AGEMA_signal_5139, new_AGEMA_signal_5138, Inst_bSbox_T14}), .b ({new_AGEMA_signal_5155, new_AGEMA_signal_5154, new_AGEMA_signal_5153, Inst_bSbox_M1}), .c ({new_AGEMA_signal_5398, new_AGEMA_signal_5397, new_AGEMA_signal_5396, Inst_bSbox_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M4_U1 ( .a ({new_AGEMA_signal_5053, new_AGEMA_signal_5052, new_AGEMA_signal_5051, Inst_bSbox_T19}), .b ({new_AGEMA_signal_4516, new_AGEMA_signal_4515, new_AGEMA_signal_4514, SboxIn[0]}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_5158, new_AGEMA_signal_5157, new_AGEMA_signal_5156, Inst_bSbox_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M5_U1 ( .a ({new_AGEMA_signal_5158, new_AGEMA_signal_5157, new_AGEMA_signal_5156, Inst_bSbox_M4}), .b ({new_AGEMA_signal_5155, new_AGEMA_signal_5154, new_AGEMA_signal_5153, Inst_bSbox_M1}), .c ({new_AGEMA_signal_5401, new_AGEMA_signal_5400, new_AGEMA_signal_5399, Inst_bSbox_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M6_U1 ( .a ({new_AGEMA_signal_4594, new_AGEMA_signal_4593, new_AGEMA_signal_4592, Inst_bSbox_T3}), .b ({new_AGEMA_signal_5050, new_AGEMA_signal_5049, new_AGEMA_signal_5048, Inst_bSbox_T16}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_5161, new_AGEMA_signal_5160, new_AGEMA_signal_5159, Inst_bSbox_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M7_U1 ( .a ({new_AGEMA_signal_5056, new_AGEMA_signal_5055, new_AGEMA_signal_5054, Inst_bSbox_T22}), .b ({new_AGEMA_signal_5041, new_AGEMA_signal_5040, new_AGEMA_signal_5039, Inst_bSbox_T9}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_5164, new_AGEMA_signal_5163, new_AGEMA_signal_5162, Inst_bSbox_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M8_U1 ( .a ({new_AGEMA_signal_5152, new_AGEMA_signal_5151, new_AGEMA_signal_5150, Inst_bSbox_T26}), .b ({new_AGEMA_signal_5161, new_AGEMA_signal_5160, new_AGEMA_signal_5159, Inst_bSbox_M6}), .c ({new_AGEMA_signal_5404, new_AGEMA_signal_5403, new_AGEMA_signal_5402, Inst_bSbox_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M9_U1 ( .a ({new_AGEMA_signal_5146, new_AGEMA_signal_5145, new_AGEMA_signal_5144, Inst_bSbox_T20}), .b ({new_AGEMA_signal_5143, new_AGEMA_signal_5142, new_AGEMA_signal_5141, Inst_bSbox_T17}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_5407, new_AGEMA_signal_5406, new_AGEMA_signal_5405, Inst_bSbox_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M10_U1 ( .a ({new_AGEMA_signal_5407, new_AGEMA_signal_5406, new_AGEMA_signal_5405, Inst_bSbox_M9}), .b ({new_AGEMA_signal_5161, new_AGEMA_signal_5160, new_AGEMA_signal_5159, Inst_bSbox_M6}), .c ({new_AGEMA_signal_5824, new_AGEMA_signal_5823, new_AGEMA_signal_5822, Inst_bSbox_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M11_U1 ( .a ({new_AGEMA_signal_4588, new_AGEMA_signal_4587, new_AGEMA_signal_4586, Inst_bSbox_T1}), .b ({new_AGEMA_signal_5047, new_AGEMA_signal_5046, new_AGEMA_signal_5045, Inst_bSbox_T15}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_5167, new_AGEMA_signal_5166, new_AGEMA_signal_5165, Inst_bSbox_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M12_U1 ( .a ({new_AGEMA_signal_4597, new_AGEMA_signal_4596, new_AGEMA_signal_4595, Inst_bSbox_T4}), .b ({new_AGEMA_signal_5059, new_AGEMA_signal_5058, new_AGEMA_signal_5057, Inst_bSbox_T27}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_5170, new_AGEMA_signal_5169, new_AGEMA_signal_5168, Inst_bSbox_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M13_U1 ( .a ({new_AGEMA_signal_5170, new_AGEMA_signal_5169, new_AGEMA_signal_5168, Inst_bSbox_M12}), .b ({new_AGEMA_signal_5167, new_AGEMA_signal_5166, new_AGEMA_signal_5165, Inst_bSbox_M11}), .c ({new_AGEMA_signal_5410, new_AGEMA_signal_5409, new_AGEMA_signal_5408, Inst_bSbox_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M14_U1 ( .a ({new_AGEMA_signal_4591, new_AGEMA_signal_4590, new_AGEMA_signal_4589, Inst_bSbox_T2}), .b ({new_AGEMA_signal_5137, new_AGEMA_signal_5136, new_AGEMA_signal_5135, Inst_bSbox_T10}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_5413, new_AGEMA_signal_5412, new_AGEMA_signal_5411, Inst_bSbox_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M15_U1 ( .a ({new_AGEMA_signal_5413, new_AGEMA_signal_5412, new_AGEMA_signal_5411, Inst_bSbox_M14}), .b ({new_AGEMA_signal_5167, new_AGEMA_signal_5166, new_AGEMA_signal_5165, Inst_bSbox_M11}), .c ({new_AGEMA_signal_5827, new_AGEMA_signal_5826, new_AGEMA_signal_5825, Inst_bSbox_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M16_U1 ( .a ({new_AGEMA_signal_5398, new_AGEMA_signal_5397, new_AGEMA_signal_5396, Inst_bSbox_M3}), .b ({new_AGEMA_signal_5395, new_AGEMA_signal_5394, new_AGEMA_signal_5393, Inst_bSbox_M2}), .c ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, new_AGEMA_signal_5828, Inst_bSbox_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M17_U1 ( .a ({new_AGEMA_signal_5401, new_AGEMA_signal_5400, new_AGEMA_signal_5399, Inst_bSbox_M5}), .b ({new_AGEMA_signal_5389, new_AGEMA_signal_5388, new_AGEMA_signal_5387, Inst_bSbox_T24}), .c ({new_AGEMA_signal_5833, new_AGEMA_signal_5832, new_AGEMA_signal_5831, Inst_bSbox_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M18_U1 ( .a ({new_AGEMA_signal_5404, new_AGEMA_signal_5403, new_AGEMA_signal_5402, Inst_bSbox_M8}), .b ({new_AGEMA_signal_5164, new_AGEMA_signal_5163, new_AGEMA_signal_5162, Inst_bSbox_M7}), .c ({new_AGEMA_signal_5836, new_AGEMA_signal_5835, new_AGEMA_signal_5834, Inst_bSbox_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M19_U1 ( .a ({new_AGEMA_signal_5824, new_AGEMA_signal_5823, new_AGEMA_signal_5822, Inst_bSbox_M10}), .b ({new_AGEMA_signal_5827, new_AGEMA_signal_5826, new_AGEMA_signal_5825, Inst_bSbox_M15}), .c ({new_AGEMA_signal_6151, new_AGEMA_signal_6150, new_AGEMA_signal_6149, Inst_bSbox_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M20_U1 ( .a ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, new_AGEMA_signal_5828, Inst_bSbox_M16}), .b ({new_AGEMA_signal_5410, new_AGEMA_signal_5409, new_AGEMA_signal_5408, Inst_bSbox_M13}), .c ({new_AGEMA_signal_6154, new_AGEMA_signal_6153, new_AGEMA_signal_6152, Inst_bSbox_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M21_U1 ( .a ({new_AGEMA_signal_5833, new_AGEMA_signal_5832, new_AGEMA_signal_5831, Inst_bSbox_M17}), .b ({new_AGEMA_signal_5827, new_AGEMA_signal_5826, new_AGEMA_signal_5825, Inst_bSbox_M15}), .c ({new_AGEMA_signal_6157, new_AGEMA_signal_6156, new_AGEMA_signal_6155, Inst_bSbox_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M22_U1 ( .a ({new_AGEMA_signal_5836, new_AGEMA_signal_5835, new_AGEMA_signal_5834, Inst_bSbox_M18}), .b ({new_AGEMA_signal_5410, new_AGEMA_signal_5409, new_AGEMA_signal_5408, Inst_bSbox_M13}), .c ({new_AGEMA_signal_6160, new_AGEMA_signal_6159, new_AGEMA_signal_6158, Inst_bSbox_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M23_U1 ( .a ({new_AGEMA_signal_6151, new_AGEMA_signal_6150, new_AGEMA_signal_6149, Inst_bSbox_M19}), .b ({new_AGEMA_signal_5392, new_AGEMA_signal_5391, new_AGEMA_signal_5390, Inst_bSbox_T25}), .c ({new_AGEMA_signal_6187, new_AGEMA_signal_6186, new_AGEMA_signal_6185, Inst_bSbox_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M24_U1 ( .a ({new_AGEMA_signal_6160, new_AGEMA_signal_6159, new_AGEMA_signal_6158, Inst_bSbox_M22}), .b ({new_AGEMA_signal_6187, new_AGEMA_signal_6186, new_AGEMA_signal_6185, Inst_bSbox_M23}), .c ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, new_AGEMA_signal_6197, Inst_bSbox_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M27_U1 ( .a ({new_AGEMA_signal_6154, new_AGEMA_signal_6153, new_AGEMA_signal_6152, Inst_bSbox_M20}), .b ({new_AGEMA_signal_6157, new_AGEMA_signal_6156, new_AGEMA_signal_6155, Inst_bSbox_M21}), .c ({new_AGEMA_signal_6193, new_AGEMA_signal_6192, new_AGEMA_signal_6191, Inst_bSbox_M27}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M25_U1 ( .a ({new_AGEMA_signal_6160, new_AGEMA_signal_6159, new_AGEMA_signal_6158, Inst_bSbox_M22}), .b ({new_AGEMA_signal_6154, new_AGEMA_signal_6153, new_AGEMA_signal_6152, Inst_bSbox_M20}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_6190, new_AGEMA_signal_6189, new_AGEMA_signal_6188, Inst_bSbox_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M26_U1 ( .a ({new_AGEMA_signal_6157, new_AGEMA_signal_6156, new_AGEMA_signal_6155, Inst_bSbox_M21}), .b ({new_AGEMA_signal_6190, new_AGEMA_signal_6189, new_AGEMA_signal_6188, Inst_bSbox_M25}), .c ({new_AGEMA_signal_6202, new_AGEMA_signal_6201, new_AGEMA_signal_6200, Inst_bSbox_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M28_U1 ( .a ({new_AGEMA_signal_6187, new_AGEMA_signal_6186, new_AGEMA_signal_6185, Inst_bSbox_M23}), .b ({new_AGEMA_signal_6190, new_AGEMA_signal_6189, new_AGEMA_signal_6188, Inst_bSbox_M25}), .c ({new_AGEMA_signal_6205, new_AGEMA_signal_6204, new_AGEMA_signal_6203, Inst_bSbox_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M31_U1 ( .a ({new_AGEMA_signal_6154, new_AGEMA_signal_6153, new_AGEMA_signal_6152, Inst_bSbox_M20}), .b ({new_AGEMA_signal_6187, new_AGEMA_signal_6186, new_AGEMA_signal_6185, Inst_bSbox_M23}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_6208, new_AGEMA_signal_6207, new_AGEMA_signal_6206, Inst_bSbox_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M33_U1 ( .a ({new_AGEMA_signal_6193, new_AGEMA_signal_6192, new_AGEMA_signal_6191, Inst_bSbox_M27}), .b ({new_AGEMA_signal_6190, new_AGEMA_signal_6189, new_AGEMA_signal_6188, Inst_bSbox_M25}), .c ({new_AGEMA_signal_6211, new_AGEMA_signal_6210, new_AGEMA_signal_6209, Inst_bSbox_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M34_U1 ( .a ({new_AGEMA_signal_6157, new_AGEMA_signal_6156, new_AGEMA_signal_6155, Inst_bSbox_M21}), .b ({new_AGEMA_signal_6160, new_AGEMA_signal_6159, new_AGEMA_signal_6158, Inst_bSbox_M22}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_6196, new_AGEMA_signal_6195, new_AGEMA_signal_6194, Inst_bSbox_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M36_U1 ( .a ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, new_AGEMA_signal_6197, Inst_bSbox_M24}), .b ({new_AGEMA_signal_6190, new_AGEMA_signal_6189, new_AGEMA_signal_6188, Inst_bSbox_M25}), .c ({new_AGEMA_signal_6226, new_AGEMA_signal_6225, new_AGEMA_signal_6224, Inst_bSbox_M36}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M29_U1 ( .a ({new_AGEMA_signal_6205, new_AGEMA_signal_6204, new_AGEMA_signal_6203, Inst_bSbox_M28}), .b ({new_AGEMA_signal_6193, new_AGEMA_signal_6192, new_AGEMA_signal_6191, Inst_bSbox_M27}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_6214, new_AGEMA_signal_6213, new_AGEMA_signal_6212, Inst_bSbox_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M30_U1 ( .a ({new_AGEMA_signal_6202, new_AGEMA_signal_6201, new_AGEMA_signal_6200, Inst_bSbox_M26}), .b ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, new_AGEMA_signal_6197, Inst_bSbox_M24}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_6217, new_AGEMA_signal_6216, new_AGEMA_signal_6215, Inst_bSbox_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M32_U1 ( .a ({new_AGEMA_signal_6193, new_AGEMA_signal_6192, new_AGEMA_signal_6191, Inst_bSbox_M27}), .b ({new_AGEMA_signal_6208, new_AGEMA_signal_6207, new_AGEMA_signal_6206, Inst_bSbox_M31}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_6220, new_AGEMA_signal_6219, new_AGEMA_signal_6218, Inst_bSbox_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M35_U1 ( .a ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, new_AGEMA_signal_6197, Inst_bSbox_M24}), .b ({new_AGEMA_signal_6196, new_AGEMA_signal_6195, new_AGEMA_signal_6194, Inst_bSbox_M34}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_6223, new_AGEMA_signal_6222, new_AGEMA_signal_6221, Inst_bSbox_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M37_U1 ( .a ({new_AGEMA_signal_6157, new_AGEMA_signal_6156, new_AGEMA_signal_6155, Inst_bSbox_M21}), .b ({new_AGEMA_signal_6214, new_AGEMA_signal_6213, new_AGEMA_signal_6212, Inst_bSbox_M29}), .c ({new_AGEMA_signal_6229, new_AGEMA_signal_6228, new_AGEMA_signal_6227, Inst_bSbox_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M38_U1 ( .a ({new_AGEMA_signal_6220, new_AGEMA_signal_6219, new_AGEMA_signal_6218, Inst_bSbox_M32}), .b ({new_AGEMA_signal_6211, new_AGEMA_signal_6210, new_AGEMA_signal_6209, Inst_bSbox_M33}), .c ({new_AGEMA_signal_6232, new_AGEMA_signal_6231, new_AGEMA_signal_6230, Inst_bSbox_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M39_U1 ( .a ({new_AGEMA_signal_6187, new_AGEMA_signal_6186, new_AGEMA_signal_6185, Inst_bSbox_M23}), .b ({new_AGEMA_signal_6217, new_AGEMA_signal_6216, new_AGEMA_signal_6215, Inst_bSbox_M30}), .c ({new_AGEMA_signal_6235, new_AGEMA_signal_6234, new_AGEMA_signal_6233, Inst_bSbox_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M40_U1 ( .a ({new_AGEMA_signal_6223, new_AGEMA_signal_6222, new_AGEMA_signal_6221, Inst_bSbox_M35}), .b ({new_AGEMA_signal_6226, new_AGEMA_signal_6225, new_AGEMA_signal_6224, Inst_bSbox_M36}), .c ({new_AGEMA_signal_6238, new_AGEMA_signal_6237, new_AGEMA_signal_6236, Inst_bSbox_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M41_U1 ( .a ({new_AGEMA_signal_6232, new_AGEMA_signal_6231, new_AGEMA_signal_6230, Inst_bSbox_M38}), .b ({new_AGEMA_signal_6238, new_AGEMA_signal_6237, new_AGEMA_signal_6236, Inst_bSbox_M40}), .c ({new_AGEMA_signal_6241, new_AGEMA_signal_6240, new_AGEMA_signal_6239, Inst_bSbox_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M42_U1 ( .a ({new_AGEMA_signal_6229, new_AGEMA_signal_6228, new_AGEMA_signal_6227, Inst_bSbox_M37}), .b ({new_AGEMA_signal_6235, new_AGEMA_signal_6234, new_AGEMA_signal_6233, Inst_bSbox_M39}), .c ({new_AGEMA_signal_6244, new_AGEMA_signal_6243, new_AGEMA_signal_6242, Inst_bSbox_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M43_U1 ( .a ({new_AGEMA_signal_6229, new_AGEMA_signal_6228, new_AGEMA_signal_6227, Inst_bSbox_M37}), .b ({new_AGEMA_signal_6232, new_AGEMA_signal_6231, new_AGEMA_signal_6230, Inst_bSbox_M38}), .c ({new_AGEMA_signal_6247, new_AGEMA_signal_6246, new_AGEMA_signal_6245, Inst_bSbox_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M44_U1 ( .a ({new_AGEMA_signal_6235, new_AGEMA_signal_6234, new_AGEMA_signal_6233, Inst_bSbox_M39}), .b ({new_AGEMA_signal_6238, new_AGEMA_signal_6237, new_AGEMA_signal_6236, Inst_bSbox_M40}), .c ({new_AGEMA_signal_6250, new_AGEMA_signal_6249, new_AGEMA_signal_6248, Inst_bSbox_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_M45_U1 ( .a ({new_AGEMA_signal_6244, new_AGEMA_signal_6243, new_AGEMA_signal_6242, Inst_bSbox_M42}), .b ({new_AGEMA_signal_6241, new_AGEMA_signal_6240, new_AGEMA_signal_6239, Inst_bSbox_M41}), .c ({new_AGEMA_signal_6277, new_AGEMA_signal_6276, new_AGEMA_signal_6275, Inst_bSbox_M45}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateIn_mux_inst_0_U1 ( .s (intFinal), .b ({new_AGEMA_signal_6400, new_AGEMA_signal_6399, new_AGEMA_signal_6398, SboxOut[0]}), .a ({new_AGEMA_signal_1990, new_AGEMA_signal_1989, new_AGEMA_signal_1988, StateOutXORroundKey[0]}), .c ({new_AGEMA_signal_6403, new_AGEMA_signal_6402, new_AGEMA_signal_6401, StateIn[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateIn_mux_inst_1_U1 ( .s (intFinal), .b ({new_AGEMA_signal_6427, new_AGEMA_signal_6426, new_AGEMA_signal_6425, SboxOut[1]}), .a ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, new_AGEMA_signal_1997, StateOutXORroundKey[1]}), .c ({new_AGEMA_signal_6430, new_AGEMA_signal_6429, new_AGEMA_signal_6428, StateIn[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateIn_mux_inst_2_U1 ( .s (intFinal), .b ({new_AGEMA_signal_6424, new_AGEMA_signal_6423, new_AGEMA_signal_6422, SboxOut[2]}), .a ({new_AGEMA_signal_2008, new_AGEMA_signal_2007, new_AGEMA_signal_2006, StateOutXORroundKey[2]}), .c ({new_AGEMA_signal_6433, new_AGEMA_signal_6432, new_AGEMA_signal_6431, StateIn[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateIn_mux_inst_3_U1 ( .s (intFinal), .b ({new_AGEMA_signal_6421, new_AGEMA_signal_6420, new_AGEMA_signal_6419, SboxOut[3]}), .a ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, new_AGEMA_signal_2015, StateOutXORroundKey[3]}), .c ({new_AGEMA_signal_6436, new_AGEMA_signal_6435, new_AGEMA_signal_6434, StateIn[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateIn_mux_inst_4_U1 ( .s (intFinal), .b ({new_AGEMA_signal_6418, new_AGEMA_signal_6417, new_AGEMA_signal_6416, SboxOut[4]}), .a ({new_AGEMA_signal_2026, new_AGEMA_signal_2025, new_AGEMA_signal_2024, StateOutXORroundKey[4]}), .c ({new_AGEMA_signal_6439, new_AGEMA_signal_6438, new_AGEMA_signal_6437, StateIn[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateIn_mux_inst_5_U1 ( .s (intFinal), .b ({new_AGEMA_signal_6415, new_AGEMA_signal_6414, new_AGEMA_signal_6413, SboxOut[5]}), .a ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, new_AGEMA_signal_2033, StateOutXORroundKey[5]}), .c ({new_AGEMA_signal_6442, new_AGEMA_signal_6441, new_AGEMA_signal_6440, StateIn[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateIn_mux_inst_6_U1 ( .s (intFinal), .b ({new_AGEMA_signal_6412, new_AGEMA_signal_6411, new_AGEMA_signal_6410, SboxOut[6]}), .a ({new_AGEMA_signal_2044, new_AGEMA_signal_2043, new_AGEMA_signal_2042, StateOutXORroundKey[6]}), .c ({new_AGEMA_signal_6445, new_AGEMA_signal_6444, new_AGEMA_signal_6443, StateIn[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_StateIn_mux_inst_7_U1 ( .s (intFinal), .b ({new_AGEMA_signal_6409, new_AGEMA_signal_6408, new_AGEMA_signal_6407, SboxOut[7]}), .a ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, new_AGEMA_signal_2051, StateOutXORroundKey[7]}), .c ({new_AGEMA_signal_6448, new_AGEMA_signal_6447, new_AGEMA_signal_6446, StateIn[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S33reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_6502, new_AGEMA_signal_6501, new_AGEMA_signal_6500, stateArray_inS33ser[0]}), .a ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .c ({new_AGEMA_signal_6529, new_AGEMA_signal_6528, new_AGEMA_signal_6527, stateArray_S33reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S33reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_6535, new_AGEMA_signal_6534, new_AGEMA_signal_6533, stateArray_inS33ser[1]}), .a ({ciphertext_s3[9], ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .c ({new_AGEMA_signal_6598, new_AGEMA_signal_6597, new_AGEMA_signal_6596, stateArray_S33reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S33reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_6541, new_AGEMA_signal_6540, new_AGEMA_signal_6539, stateArray_inS33ser[2]}), .a ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_6601, new_AGEMA_signal_6600, new_AGEMA_signal_6599, stateArray_S33reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S33reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_6547, new_AGEMA_signal_6546, new_AGEMA_signal_6545, stateArray_inS33ser[3]}), .a ({ciphertext_s3[11], ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .c ({new_AGEMA_signal_6604, new_AGEMA_signal_6603, new_AGEMA_signal_6602, stateArray_S33reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S33reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_6553, new_AGEMA_signal_6552, new_AGEMA_signal_6551, stateArray_inS33ser[4]}), .a ({ciphertext_s3[12], ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .c ({new_AGEMA_signal_6607, new_AGEMA_signal_6606, new_AGEMA_signal_6605, stateArray_S33reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S33reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_6559, new_AGEMA_signal_6558, new_AGEMA_signal_6557, stateArray_inS33ser[5]}), .a ({ciphertext_s3[13], ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .c ({new_AGEMA_signal_6610, new_AGEMA_signal_6609, new_AGEMA_signal_6608, stateArray_S33reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S33reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_6565, new_AGEMA_signal_6564, new_AGEMA_signal_6563, stateArray_inS33ser[6]}), .a ({ciphertext_s3[14], ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .c ({new_AGEMA_signal_6613, new_AGEMA_signal_6612, new_AGEMA_signal_6611, stateArray_S33reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_S33reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_6571, new_AGEMA_signal_6570, new_AGEMA_signal_6569, stateArray_inS33ser[7]}), .a ({ciphertext_s3[15], ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .c ({new_AGEMA_signal_6616, new_AGEMA_signal_6615, new_AGEMA_signal_6614, stateArray_S33reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_input_MC_mux_inst_0_U1 ( .s (stateArray_n22), .b ({new_AGEMA_signal_6403, new_AGEMA_signal_6402, new_AGEMA_signal_6401, StateIn[0]}), .a ({new_AGEMA_signal_4618, new_AGEMA_signal_4617, new_AGEMA_signal_4616, StateInMC[0]}), .c ({new_AGEMA_signal_6451, new_AGEMA_signal_6450, new_AGEMA_signal_6449, stateArray_input_MC[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_input_MC_mux_inst_1_U1 ( .s (stateArray_n22), .b ({new_AGEMA_signal_6430, new_AGEMA_signal_6429, new_AGEMA_signal_6428, StateIn[1]}), .a ({new_AGEMA_signal_4621, new_AGEMA_signal_4620, new_AGEMA_signal_4619, StateInMC[1]}), .c ({new_AGEMA_signal_6478, new_AGEMA_signal_6477, new_AGEMA_signal_6476, stateArray_input_MC[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_input_MC_mux_inst_2_U1 ( .s (stateArray_n22), .b ({new_AGEMA_signal_6433, new_AGEMA_signal_6432, new_AGEMA_signal_6431, StateIn[2]}), .a ({new_AGEMA_signal_4540, new_AGEMA_signal_4539, new_AGEMA_signal_4538, StateInMC[2]}), .c ({new_AGEMA_signal_6481, new_AGEMA_signal_6480, new_AGEMA_signal_6479, stateArray_input_MC[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_input_MC_mux_inst_3_U1 ( .s (stateArray_n22), .b ({new_AGEMA_signal_6436, new_AGEMA_signal_6435, new_AGEMA_signal_6434, StateIn[3]}), .a ({new_AGEMA_signal_4624, new_AGEMA_signal_4623, new_AGEMA_signal_4622, StateInMC[3]}), .c ({new_AGEMA_signal_6484, new_AGEMA_signal_6483, new_AGEMA_signal_6482, stateArray_input_MC[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_input_MC_mux_inst_4_U1 ( .s (stateArray_n22), .b ({new_AGEMA_signal_6439, new_AGEMA_signal_6438, new_AGEMA_signal_6437, StateIn[4]}), .a ({new_AGEMA_signal_4627, new_AGEMA_signal_4626, new_AGEMA_signal_4625, StateInMC[4]}), .c ({new_AGEMA_signal_6487, new_AGEMA_signal_6486, new_AGEMA_signal_6485, stateArray_input_MC[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_input_MC_mux_inst_5_U1 ( .s (stateArray_n22), .b ({new_AGEMA_signal_6442, new_AGEMA_signal_6441, new_AGEMA_signal_6440, StateIn[5]}), .a ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, new_AGEMA_signal_4541, StateInMC[5]}), .c ({new_AGEMA_signal_6490, new_AGEMA_signal_6489, new_AGEMA_signal_6488, stateArray_input_MC[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_input_MC_mux_inst_6_U1 ( .s (stateArray_n22), .b ({new_AGEMA_signal_6445, new_AGEMA_signal_6444, new_AGEMA_signal_6443, StateIn[6]}), .a ({new_AGEMA_signal_4546, new_AGEMA_signal_4545, new_AGEMA_signal_4544, StateInMC[6]}), .c ({new_AGEMA_signal_6493, new_AGEMA_signal_6492, new_AGEMA_signal_6491, stateArray_input_MC[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_input_MC_mux_inst_7_U1 ( .s (stateArray_n22), .b ({new_AGEMA_signal_6448, new_AGEMA_signal_6447, new_AGEMA_signal_6446, StateIn[7]}), .a ({new_AGEMA_signal_4549, new_AGEMA_signal_4548, new_AGEMA_signal_4547, StateInMC[7]}), .c ({new_AGEMA_signal_6496, new_AGEMA_signal_6495, new_AGEMA_signal_6494, stateArray_input_MC[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS33ser_mux_inst_0_U1 ( .s (stateArray_n25), .b ({plaintext_s3[0], plaintext_s2[0], plaintext_s1[0], plaintext_s0[0]}), .a ({new_AGEMA_signal_6451, new_AGEMA_signal_6450, new_AGEMA_signal_6449, stateArray_input_MC[0]}), .c ({new_AGEMA_signal_6502, new_AGEMA_signal_6501, new_AGEMA_signal_6500, stateArray_inS33ser[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS33ser_mux_inst_1_U1 ( .s (stateArray_n25), .b ({plaintext_s3[1], plaintext_s2[1], plaintext_s1[1], plaintext_s0[1]}), .a ({new_AGEMA_signal_6478, new_AGEMA_signal_6477, new_AGEMA_signal_6476, stateArray_input_MC[1]}), .c ({new_AGEMA_signal_6535, new_AGEMA_signal_6534, new_AGEMA_signal_6533, stateArray_inS33ser[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS33ser_mux_inst_2_U1 ( .s (stateArray_n25), .b ({plaintext_s3[2], plaintext_s2[2], plaintext_s1[2], plaintext_s0[2]}), .a ({new_AGEMA_signal_6481, new_AGEMA_signal_6480, new_AGEMA_signal_6479, stateArray_input_MC[2]}), .c ({new_AGEMA_signal_6541, new_AGEMA_signal_6540, new_AGEMA_signal_6539, stateArray_inS33ser[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS33ser_mux_inst_3_U1 ( .s (stateArray_n25), .b ({plaintext_s3[3], plaintext_s2[3], plaintext_s1[3], plaintext_s0[3]}), .a ({new_AGEMA_signal_6484, new_AGEMA_signal_6483, new_AGEMA_signal_6482, stateArray_input_MC[3]}), .c ({new_AGEMA_signal_6547, new_AGEMA_signal_6546, new_AGEMA_signal_6545, stateArray_inS33ser[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS33ser_mux_inst_4_U1 ( .s (stateArray_n25), .b ({plaintext_s3[4], plaintext_s2[4], plaintext_s1[4], plaintext_s0[4]}), .a ({new_AGEMA_signal_6487, new_AGEMA_signal_6486, new_AGEMA_signal_6485, stateArray_input_MC[4]}), .c ({new_AGEMA_signal_6553, new_AGEMA_signal_6552, new_AGEMA_signal_6551, stateArray_inS33ser[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS33ser_mux_inst_5_U1 ( .s (stateArray_n25), .b ({plaintext_s3[5], plaintext_s2[5], plaintext_s1[5], plaintext_s0[5]}), .a ({new_AGEMA_signal_6490, new_AGEMA_signal_6489, new_AGEMA_signal_6488, stateArray_input_MC[5]}), .c ({new_AGEMA_signal_6559, new_AGEMA_signal_6558, new_AGEMA_signal_6557, stateArray_inS33ser[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS33ser_mux_inst_6_U1 ( .s (stateArray_n25), .b ({plaintext_s3[6], plaintext_s2[6], plaintext_s1[6], plaintext_s0[6]}), .a ({new_AGEMA_signal_6493, new_AGEMA_signal_6492, new_AGEMA_signal_6491, stateArray_input_MC[6]}), .c ({new_AGEMA_signal_6565, new_AGEMA_signal_6564, new_AGEMA_signal_6563, stateArray_inS33ser[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateArray_MUX_inS33ser_mux_inst_7_U1 ( .s (stateArray_n25), .b ({plaintext_s3[7], plaintext_s2[7], plaintext_s1[7], plaintext_s0[7]}), .a ({new_AGEMA_signal_6496, new_AGEMA_signal_6495, new_AGEMA_signal_6494, stateArray_input_MC[7]}), .c ({new_AGEMA_signal_6571, new_AGEMA_signal_6570, new_AGEMA_signal_6569, stateArray_inS33ser[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U42 ( .a ({new_AGEMA_signal_6454, new_AGEMA_signal_6453, new_AGEMA_signal_6452, KeyArray_n55}), .b ({new_AGEMA_signal_2050, new_AGEMA_signal_2049, new_AGEMA_signal_2048, keyStateIn[7]}), .c ({new_AGEMA_signal_6505, new_AGEMA_signal_6504, new_AGEMA_signal_6503, KeyArray_inS30par[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U41 ( .a ({1'b0, 1'b0, 1'b0, roundConstant[7]}), .b ({new_AGEMA_signal_6409, new_AGEMA_signal_6408, new_AGEMA_signal_6407, SboxOut[7]}), .c ({new_AGEMA_signal_6454, new_AGEMA_signal_6453, new_AGEMA_signal_6452, KeyArray_n55}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U40 ( .a ({new_AGEMA_signal_6457, new_AGEMA_signal_6456, new_AGEMA_signal_6455, KeyArray_n54}), .b ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, new_AGEMA_signal_2039, keyStateIn[6]}), .c ({new_AGEMA_signal_6508, new_AGEMA_signal_6507, new_AGEMA_signal_6506, KeyArray_inS30par[6]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U39 ( .a ({1'b0, 1'b0, 1'b0, roundConstant[6]}), .b ({new_AGEMA_signal_6412, new_AGEMA_signal_6411, new_AGEMA_signal_6410, SboxOut[6]}), .c ({new_AGEMA_signal_6457, new_AGEMA_signal_6456, new_AGEMA_signal_6455, KeyArray_n54}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U38 ( .a ({new_AGEMA_signal_6460, new_AGEMA_signal_6459, new_AGEMA_signal_6458, KeyArray_n53}), .b ({new_AGEMA_signal_2032, new_AGEMA_signal_2031, new_AGEMA_signal_2030, keyStateIn[5]}), .c ({new_AGEMA_signal_6511, new_AGEMA_signal_6510, new_AGEMA_signal_6509, KeyArray_inS30par[5]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U37 ( .a ({1'b0, 1'b0, 1'b0, roundConstant[5]}), .b ({new_AGEMA_signal_6415, new_AGEMA_signal_6414, new_AGEMA_signal_6413, SboxOut[5]}), .c ({new_AGEMA_signal_6460, new_AGEMA_signal_6459, new_AGEMA_signal_6458, KeyArray_n53}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U36 ( .a ({new_AGEMA_signal_6463, new_AGEMA_signal_6462, new_AGEMA_signal_6461, KeyArray_n52}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, new_AGEMA_signal_2021, keyStateIn[4]}), .c ({new_AGEMA_signal_6514, new_AGEMA_signal_6513, new_AGEMA_signal_6512, KeyArray_inS30par[4]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U35 ( .a ({1'b0, 1'b0, 1'b0, roundConstant[4]}), .b ({new_AGEMA_signal_6418, new_AGEMA_signal_6417, new_AGEMA_signal_6416, SboxOut[4]}), .c ({new_AGEMA_signal_6463, new_AGEMA_signal_6462, new_AGEMA_signal_6461, KeyArray_n52}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U34 ( .a ({new_AGEMA_signal_6466, new_AGEMA_signal_6465, new_AGEMA_signal_6464, KeyArray_n51}), .b ({new_AGEMA_signal_2014, new_AGEMA_signal_2013, new_AGEMA_signal_2012, keyStateIn[3]}), .c ({new_AGEMA_signal_6517, new_AGEMA_signal_6516, new_AGEMA_signal_6515, KeyArray_inS30par[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U33 ( .a ({1'b0, 1'b0, 1'b0, roundConstant[3]}), .b ({new_AGEMA_signal_6421, new_AGEMA_signal_6420, new_AGEMA_signal_6419, SboxOut[3]}), .c ({new_AGEMA_signal_6466, new_AGEMA_signal_6465, new_AGEMA_signal_6464, KeyArray_n51}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U32 ( .a ({new_AGEMA_signal_6469, new_AGEMA_signal_6468, new_AGEMA_signal_6467, KeyArray_n50}), .b ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, new_AGEMA_signal_2003, keyStateIn[2]}), .c ({new_AGEMA_signal_6520, new_AGEMA_signal_6519, new_AGEMA_signal_6518, KeyArray_inS30par[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U31 ( .a ({1'b0, 1'b0, 1'b0, roundConstant[2]}), .b ({new_AGEMA_signal_6424, new_AGEMA_signal_6423, new_AGEMA_signal_6422, SboxOut[2]}), .c ({new_AGEMA_signal_6469, new_AGEMA_signal_6468, new_AGEMA_signal_6467, KeyArray_n50}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U30 ( .a ({new_AGEMA_signal_6472, new_AGEMA_signal_6471, new_AGEMA_signal_6470, KeyArray_n49}), .b ({new_AGEMA_signal_1996, new_AGEMA_signal_1995, new_AGEMA_signal_1994, keyStateIn[1]}), .c ({new_AGEMA_signal_6523, new_AGEMA_signal_6522, new_AGEMA_signal_6521, KeyArray_inS30par[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U29 ( .a ({1'b0, 1'b0, 1'b0, roundConstant[1]}), .b ({new_AGEMA_signal_6427, new_AGEMA_signal_6426, new_AGEMA_signal_6425, SboxOut[1]}), .c ({new_AGEMA_signal_6472, new_AGEMA_signal_6471, new_AGEMA_signal_6470, KeyArray_n49}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U28 ( .a ({new_AGEMA_signal_6406, new_AGEMA_signal_6405, new_AGEMA_signal_6404, KeyArray_n48}), .b ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, new_AGEMA_signal_1985, keyStateIn[0]}), .c ({new_AGEMA_signal_6475, new_AGEMA_signal_6474, new_AGEMA_signal_6473, KeyArray_inS30par[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyArray_U27 ( .a ({1'b0, 1'b0, 1'b0, roundConstant[0]}), .b ({new_AGEMA_signal_6400, new_AGEMA_signal_6399, new_AGEMA_signal_6398, SboxOut[0]}), .c ({new_AGEMA_signal_6406, new_AGEMA_signal_6405, new_AGEMA_signal_6404, KeyArray_n48}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_0_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_4087, new_AGEMA_signal_4086, new_AGEMA_signal_4085, KeyArray_outS30ser[0]}), .a ({new_AGEMA_signal_6526, new_AGEMA_signal_6525, new_AGEMA_signal_6524, KeyArray_S30reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_6574, new_AGEMA_signal_6573, new_AGEMA_signal_6572, KeyArray_S30reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_4162, new_AGEMA_signal_4161, new_AGEMA_signal_4160, KeyArray_inS30ser[0]}), .a ({new_AGEMA_signal_6475, new_AGEMA_signal_6474, new_AGEMA_signal_6473, KeyArray_inS30par[0]}), .c ({new_AGEMA_signal_6526, new_AGEMA_signal_6525, new_AGEMA_signal_6524, KeyArray_S30reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_1_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_4096, new_AGEMA_signal_4095, new_AGEMA_signal_4094, KeyArray_outS30ser[1]}), .a ({new_AGEMA_signal_6577, new_AGEMA_signal_6576, new_AGEMA_signal_6575, KeyArray_S30reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_6619, new_AGEMA_signal_6618, new_AGEMA_signal_6617, KeyArray_S30reg_gff_1_SFF_1_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_4171, new_AGEMA_signal_4170, new_AGEMA_signal_4169, KeyArray_inS30ser[1]}), .a ({new_AGEMA_signal_6523, new_AGEMA_signal_6522, new_AGEMA_signal_6521, KeyArray_inS30par[1]}), .c ({new_AGEMA_signal_6577, new_AGEMA_signal_6576, new_AGEMA_signal_6575, KeyArray_S30reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_2_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_4105, new_AGEMA_signal_4104, new_AGEMA_signal_4103, KeyArray_outS30ser[2]}), .a ({new_AGEMA_signal_6580, new_AGEMA_signal_6579, new_AGEMA_signal_6578, KeyArray_S30reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_6622, new_AGEMA_signal_6621, new_AGEMA_signal_6620, KeyArray_S30reg_gff_1_SFF_2_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_4180, new_AGEMA_signal_4179, new_AGEMA_signal_4178, KeyArray_inS30ser[2]}), .a ({new_AGEMA_signal_6520, new_AGEMA_signal_6519, new_AGEMA_signal_6518, KeyArray_inS30par[2]}), .c ({new_AGEMA_signal_6580, new_AGEMA_signal_6579, new_AGEMA_signal_6578, KeyArray_S30reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_3_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_4114, new_AGEMA_signal_4113, new_AGEMA_signal_4112, KeyArray_outS30ser[3]}), .a ({new_AGEMA_signal_6583, new_AGEMA_signal_6582, new_AGEMA_signal_6581, KeyArray_S30reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_6625, new_AGEMA_signal_6624, new_AGEMA_signal_6623, KeyArray_S30reg_gff_1_SFF_3_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_4189, new_AGEMA_signal_4188, new_AGEMA_signal_4187, KeyArray_inS30ser[3]}), .a ({new_AGEMA_signal_6517, new_AGEMA_signal_6516, new_AGEMA_signal_6515, KeyArray_inS30par[3]}), .c ({new_AGEMA_signal_6583, new_AGEMA_signal_6582, new_AGEMA_signal_6581, KeyArray_S30reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_4_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_4123, new_AGEMA_signal_4122, new_AGEMA_signal_4121, KeyArray_outS30ser[4]}), .a ({new_AGEMA_signal_6586, new_AGEMA_signal_6585, new_AGEMA_signal_6584, KeyArray_S30reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_6628, new_AGEMA_signal_6627, new_AGEMA_signal_6626, KeyArray_S30reg_gff_1_SFF_4_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_4198, new_AGEMA_signal_4197, new_AGEMA_signal_4196, KeyArray_inS30ser[4]}), .a ({new_AGEMA_signal_6514, new_AGEMA_signal_6513, new_AGEMA_signal_6512, KeyArray_inS30par[4]}), .c ({new_AGEMA_signal_6586, new_AGEMA_signal_6585, new_AGEMA_signal_6584, KeyArray_S30reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_5_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_4132, new_AGEMA_signal_4131, new_AGEMA_signal_4130, KeyArray_outS30ser[5]}), .a ({new_AGEMA_signal_6589, new_AGEMA_signal_6588, new_AGEMA_signal_6587, KeyArray_S30reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_6631, new_AGEMA_signal_6630, new_AGEMA_signal_6629, KeyArray_S30reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_4207, new_AGEMA_signal_4206, new_AGEMA_signal_4205, KeyArray_inS30ser[5]}), .a ({new_AGEMA_signal_6511, new_AGEMA_signal_6510, new_AGEMA_signal_6509, KeyArray_inS30par[5]}), .c ({new_AGEMA_signal_6589, new_AGEMA_signal_6588, new_AGEMA_signal_6587, KeyArray_S30reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_6_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_4141, new_AGEMA_signal_4140, new_AGEMA_signal_4139, KeyArray_outS30ser[6]}), .a ({new_AGEMA_signal_6592, new_AGEMA_signal_6591, new_AGEMA_signal_6590, KeyArray_S30reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_6634, new_AGEMA_signal_6633, new_AGEMA_signal_6632, KeyArray_S30reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_4216, new_AGEMA_signal_4215, new_AGEMA_signal_4214, KeyArray_inS30ser[6]}), .a ({new_AGEMA_signal_6508, new_AGEMA_signal_6507, new_AGEMA_signal_6506, KeyArray_inS30par[6]}), .c ({new_AGEMA_signal_6592, new_AGEMA_signal_6591, new_AGEMA_signal_6590, KeyArray_S30reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_7_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_4150, new_AGEMA_signal_4149, new_AGEMA_signal_4148, KeyArray_outS30ser[7]}), .a ({new_AGEMA_signal_6595, new_AGEMA_signal_6594, new_AGEMA_signal_6593, KeyArray_S30reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_6637, new_AGEMA_signal_6636, new_AGEMA_signal_6635, KeyArray_S30reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_4225, new_AGEMA_signal_4224, new_AGEMA_signal_4223, KeyArray_inS30ser[7]}), .a ({new_AGEMA_signal_6505, new_AGEMA_signal_6504, new_AGEMA_signal_6503, KeyArray_inS30par[7]}), .c ({new_AGEMA_signal_6595, new_AGEMA_signal_6594, new_AGEMA_signal_6593, KeyArray_S30reg_gff_1_SFF_7_QD}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M46_U1 ( .a ({new_AGEMA_signal_6250, new_AGEMA_signal_6249, new_AGEMA_signal_6248, Inst_bSbox_M44}), .b ({new_AGEMA_signal_5038, new_AGEMA_signal_5037, new_AGEMA_signal_5036, Inst_bSbox_T6}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_6280, new_AGEMA_signal_6279, new_AGEMA_signal_6278, Inst_bSbox_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M47_U1 ( .a ({new_AGEMA_signal_6238, new_AGEMA_signal_6237, new_AGEMA_signal_6236, Inst_bSbox_M40}), .b ({new_AGEMA_signal_5134, new_AGEMA_signal_5133, new_AGEMA_signal_5132, Inst_bSbox_T8}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_6253, new_AGEMA_signal_6252, new_AGEMA_signal_6251, Inst_bSbox_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M48_U1 ( .a ({new_AGEMA_signal_6235, new_AGEMA_signal_6234, new_AGEMA_signal_6233, Inst_bSbox_M39}), .b ({new_AGEMA_signal_4516, new_AGEMA_signal_4515, new_AGEMA_signal_4514, SboxIn[0]}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_6256, new_AGEMA_signal_6255, new_AGEMA_signal_6254, Inst_bSbox_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M49_U1 ( .a ({new_AGEMA_signal_6247, new_AGEMA_signal_6246, new_AGEMA_signal_6245, Inst_bSbox_M43}), .b ({new_AGEMA_signal_5050, new_AGEMA_signal_5049, new_AGEMA_signal_5048, Inst_bSbox_T16}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_6283, new_AGEMA_signal_6282, new_AGEMA_signal_6281, Inst_bSbox_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M50_U1 ( .a ({new_AGEMA_signal_6232, new_AGEMA_signal_6231, new_AGEMA_signal_6230, Inst_bSbox_M38}), .b ({new_AGEMA_signal_5041, new_AGEMA_signal_5040, new_AGEMA_signal_5039, Inst_bSbox_T9}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_6259, new_AGEMA_signal_6258, new_AGEMA_signal_6257, Inst_bSbox_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M51_U1 ( .a ({new_AGEMA_signal_6229, new_AGEMA_signal_6228, new_AGEMA_signal_6227, Inst_bSbox_M37}), .b ({new_AGEMA_signal_5143, new_AGEMA_signal_5142, new_AGEMA_signal_5141, Inst_bSbox_T17}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_6262, new_AGEMA_signal_6261, new_AGEMA_signal_6260, Inst_bSbox_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M52_U1 ( .a ({new_AGEMA_signal_6244, new_AGEMA_signal_6243, new_AGEMA_signal_6242, Inst_bSbox_M42}), .b ({new_AGEMA_signal_5047, new_AGEMA_signal_5046, new_AGEMA_signal_5045, Inst_bSbox_T15}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_6286, new_AGEMA_signal_6285, new_AGEMA_signal_6284, Inst_bSbox_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M53_U1 ( .a ({new_AGEMA_signal_6277, new_AGEMA_signal_6276, new_AGEMA_signal_6275, Inst_bSbox_M45}), .b ({new_AGEMA_signal_5059, new_AGEMA_signal_5058, new_AGEMA_signal_5057, Inst_bSbox_T27}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_6313, new_AGEMA_signal_6312, new_AGEMA_signal_6311, Inst_bSbox_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M54_U1 ( .a ({new_AGEMA_signal_6241, new_AGEMA_signal_6240, new_AGEMA_signal_6239, Inst_bSbox_M41}), .b ({new_AGEMA_signal_5137, new_AGEMA_signal_5136, new_AGEMA_signal_5135, Inst_bSbox_T10}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_6289, new_AGEMA_signal_6288, new_AGEMA_signal_6287, Inst_bSbox_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M55_U1 ( .a ({new_AGEMA_signal_6250, new_AGEMA_signal_6249, new_AGEMA_signal_6248, Inst_bSbox_M44}), .b ({new_AGEMA_signal_5044, new_AGEMA_signal_5043, new_AGEMA_signal_5042, Inst_bSbox_T13}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_6292, new_AGEMA_signal_6291, new_AGEMA_signal_6290, Inst_bSbox_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M56_U1 ( .a ({new_AGEMA_signal_6238, new_AGEMA_signal_6237, new_AGEMA_signal_6236, Inst_bSbox_M40}), .b ({new_AGEMA_signal_5149, new_AGEMA_signal_5148, new_AGEMA_signal_5147, Inst_bSbox_T23}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_6265, new_AGEMA_signal_6264, new_AGEMA_signal_6263, Inst_bSbox_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M57_U1 ( .a ({new_AGEMA_signal_6235, new_AGEMA_signal_6234, new_AGEMA_signal_6233, Inst_bSbox_M39}), .b ({new_AGEMA_signal_5053, new_AGEMA_signal_5052, new_AGEMA_signal_5051, Inst_bSbox_T19}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_6268, new_AGEMA_signal_6267, new_AGEMA_signal_6266, Inst_bSbox_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M58_U1 ( .a ({new_AGEMA_signal_6247, new_AGEMA_signal_6246, new_AGEMA_signal_6245, Inst_bSbox_M43}), .b ({new_AGEMA_signal_4594, new_AGEMA_signal_4593, new_AGEMA_signal_4592, Inst_bSbox_T3}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_6295, new_AGEMA_signal_6294, new_AGEMA_signal_6293, Inst_bSbox_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M59_U1 ( .a ({new_AGEMA_signal_6232, new_AGEMA_signal_6231, new_AGEMA_signal_6230, Inst_bSbox_M38}), .b ({new_AGEMA_signal_5056, new_AGEMA_signal_5055, new_AGEMA_signal_5054, Inst_bSbox_T22}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_6271, new_AGEMA_signal_6270, new_AGEMA_signal_6269, Inst_bSbox_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M60_U1 ( .a ({new_AGEMA_signal_6229, new_AGEMA_signal_6228, new_AGEMA_signal_6227, Inst_bSbox_M37}), .b ({new_AGEMA_signal_5146, new_AGEMA_signal_5145, new_AGEMA_signal_5144, Inst_bSbox_T20}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_6274, new_AGEMA_signal_6273, new_AGEMA_signal_6272, Inst_bSbox_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M61_U1 ( .a ({new_AGEMA_signal_6244, new_AGEMA_signal_6243, new_AGEMA_signal_6242, Inst_bSbox_M42}), .b ({new_AGEMA_signal_4588, new_AGEMA_signal_4587, new_AGEMA_signal_4586, Inst_bSbox_T1}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_6298, new_AGEMA_signal_6297, new_AGEMA_signal_6296, Inst_bSbox_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M62_U1 ( .a ({new_AGEMA_signal_6277, new_AGEMA_signal_6276, new_AGEMA_signal_6275, Inst_bSbox_M45}), .b ({new_AGEMA_signal_4597, new_AGEMA_signal_4596, new_AGEMA_signal_4595, Inst_bSbox_T4}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_6316, new_AGEMA_signal_6315, new_AGEMA_signal_6314, Inst_bSbox_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_AND_M63_U1 ( .a ({new_AGEMA_signal_6241, new_AGEMA_signal_6240, new_AGEMA_signal_6239, Inst_bSbox_M41}), .b ({new_AGEMA_signal_4591, new_AGEMA_signal_4590, new_AGEMA_signal_4589, Inst_bSbox_T2}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_6301, new_AGEMA_signal_6300, new_AGEMA_signal_6299, Inst_bSbox_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L0_U1 ( .a ({new_AGEMA_signal_6298, new_AGEMA_signal_6297, new_AGEMA_signal_6296, Inst_bSbox_M61}), .b ({new_AGEMA_signal_6316, new_AGEMA_signal_6315, new_AGEMA_signal_6314, Inst_bSbox_M62}), .c ({new_AGEMA_signal_6343, new_AGEMA_signal_6342, new_AGEMA_signal_6341, Inst_bSbox_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L1_U1 ( .a ({new_AGEMA_signal_6259, new_AGEMA_signal_6258, new_AGEMA_signal_6257, Inst_bSbox_M50}), .b ({new_AGEMA_signal_6265, new_AGEMA_signal_6264, new_AGEMA_signal_6263, Inst_bSbox_M56}), .c ({new_AGEMA_signal_6304, new_AGEMA_signal_6303, new_AGEMA_signal_6302, Inst_bSbox_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L2_U1 ( .a ({new_AGEMA_signal_6280, new_AGEMA_signal_6279, new_AGEMA_signal_6278, Inst_bSbox_M46}), .b ({new_AGEMA_signal_6256, new_AGEMA_signal_6255, new_AGEMA_signal_6254, Inst_bSbox_M48}), .c ({new_AGEMA_signal_6319, new_AGEMA_signal_6318, new_AGEMA_signal_6317, Inst_bSbox_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L3_U1 ( .a ({new_AGEMA_signal_6253, new_AGEMA_signal_6252, new_AGEMA_signal_6251, Inst_bSbox_M47}), .b ({new_AGEMA_signal_6292, new_AGEMA_signal_6291, new_AGEMA_signal_6290, Inst_bSbox_M55}), .c ({new_AGEMA_signal_6322, new_AGEMA_signal_6321, new_AGEMA_signal_6320, Inst_bSbox_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L4_U1 ( .a ({new_AGEMA_signal_6289, new_AGEMA_signal_6288, new_AGEMA_signal_6287, Inst_bSbox_M54}), .b ({new_AGEMA_signal_6295, new_AGEMA_signal_6294, new_AGEMA_signal_6293, Inst_bSbox_M58}), .c ({new_AGEMA_signal_6325, new_AGEMA_signal_6324, new_AGEMA_signal_6323, Inst_bSbox_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L5_U1 ( .a ({new_AGEMA_signal_6283, new_AGEMA_signal_6282, new_AGEMA_signal_6281, Inst_bSbox_M49}), .b ({new_AGEMA_signal_6298, new_AGEMA_signal_6297, new_AGEMA_signal_6296, Inst_bSbox_M61}), .c ({new_AGEMA_signal_6328, new_AGEMA_signal_6327, new_AGEMA_signal_6326, Inst_bSbox_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L6_U1 ( .a ({new_AGEMA_signal_6316, new_AGEMA_signal_6315, new_AGEMA_signal_6314, Inst_bSbox_M62}), .b ({new_AGEMA_signal_6328, new_AGEMA_signal_6327, new_AGEMA_signal_6326, Inst_bSbox_L5}), .c ({new_AGEMA_signal_6346, new_AGEMA_signal_6345, new_AGEMA_signal_6344, Inst_bSbox_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L7_U1 ( .a ({new_AGEMA_signal_6280, new_AGEMA_signal_6279, new_AGEMA_signal_6278, Inst_bSbox_M46}), .b ({new_AGEMA_signal_6322, new_AGEMA_signal_6321, new_AGEMA_signal_6320, Inst_bSbox_L3}), .c ({new_AGEMA_signal_6349, new_AGEMA_signal_6348, new_AGEMA_signal_6347, Inst_bSbox_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L8_U1 ( .a ({new_AGEMA_signal_6262, new_AGEMA_signal_6261, new_AGEMA_signal_6260, Inst_bSbox_M51}), .b ({new_AGEMA_signal_6271, new_AGEMA_signal_6270, new_AGEMA_signal_6269, Inst_bSbox_M59}), .c ({new_AGEMA_signal_6307, new_AGEMA_signal_6306, new_AGEMA_signal_6305, Inst_bSbox_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L9_U1 ( .a ({new_AGEMA_signal_6286, new_AGEMA_signal_6285, new_AGEMA_signal_6284, Inst_bSbox_M52}), .b ({new_AGEMA_signal_6313, new_AGEMA_signal_6312, new_AGEMA_signal_6311, Inst_bSbox_M53}), .c ({new_AGEMA_signal_6352, new_AGEMA_signal_6351, new_AGEMA_signal_6350, Inst_bSbox_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L10_U1 ( .a ({new_AGEMA_signal_6313, new_AGEMA_signal_6312, new_AGEMA_signal_6311, Inst_bSbox_M53}), .b ({new_AGEMA_signal_6325, new_AGEMA_signal_6324, new_AGEMA_signal_6323, Inst_bSbox_L4}), .c ({new_AGEMA_signal_6355, new_AGEMA_signal_6354, new_AGEMA_signal_6353, Inst_bSbox_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L11_U1 ( .a ({new_AGEMA_signal_6274, new_AGEMA_signal_6273, new_AGEMA_signal_6272, Inst_bSbox_M60}), .b ({new_AGEMA_signal_6319, new_AGEMA_signal_6318, new_AGEMA_signal_6317, Inst_bSbox_L2}), .c ({new_AGEMA_signal_6358, new_AGEMA_signal_6357, new_AGEMA_signal_6356, Inst_bSbox_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L12_U1 ( .a ({new_AGEMA_signal_6256, new_AGEMA_signal_6255, new_AGEMA_signal_6254, Inst_bSbox_M48}), .b ({new_AGEMA_signal_6262, new_AGEMA_signal_6261, new_AGEMA_signal_6260, Inst_bSbox_M51}), .c ({new_AGEMA_signal_6310, new_AGEMA_signal_6309, new_AGEMA_signal_6308, Inst_bSbox_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L13_U1 ( .a ({new_AGEMA_signal_6259, new_AGEMA_signal_6258, new_AGEMA_signal_6257, Inst_bSbox_M50}), .b ({new_AGEMA_signal_6343, new_AGEMA_signal_6342, new_AGEMA_signal_6341, Inst_bSbox_L0}), .c ({new_AGEMA_signal_6370, new_AGEMA_signal_6369, new_AGEMA_signal_6368, Inst_bSbox_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L14_U1 ( .a ({new_AGEMA_signal_6286, new_AGEMA_signal_6285, new_AGEMA_signal_6284, Inst_bSbox_M52}), .b ({new_AGEMA_signal_6298, new_AGEMA_signal_6297, new_AGEMA_signal_6296, Inst_bSbox_M61}), .c ({new_AGEMA_signal_6331, new_AGEMA_signal_6330, new_AGEMA_signal_6329, Inst_bSbox_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L15_U1 ( .a ({new_AGEMA_signal_6292, new_AGEMA_signal_6291, new_AGEMA_signal_6290, Inst_bSbox_M55}), .b ({new_AGEMA_signal_6304, new_AGEMA_signal_6303, new_AGEMA_signal_6302, Inst_bSbox_L1}), .c ({new_AGEMA_signal_6334, new_AGEMA_signal_6333, new_AGEMA_signal_6332, Inst_bSbox_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L16_U1 ( .a ({new_AGEMA_signal_6265, new_AGEMA_signal_6264, new_AGEMA_signal_6263, Inst_bSbox_M56}), .b ({new_AGEMA_signal_6343, new_AGEMA_signal_6342, new_AGEMA_signal_6341, Inst_bSbox_L0}), .c ({new_AGEMA_signal_6373, new_AGEMA_signal_6372, new_AGEMA_signal_6371, Inst_bSbox_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L17_U1 ( .a ({new_AGEMA_signal_6268, new_AGEMA_signal_6267, new_AGEMA_signal_6266, Inst_bSbox_M57}), .b ({new_AGEMA_signal_6304, new_AGEMA_signal_6303, new_AGEMA_signal_6302, Inst_bSbox_L1}), .c ({new_AGEMA_signal_6337, new_AGEMA_signal_6336, new_AGEMA_signal_6335, Inst_bSbox_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L18_U1 ( .a ({new_AGEMA_signal_6295, new_AGEMA_signal_6294, new_AGEMA_signal_6293, Inst_bSbox_M58}), .b ({new_AGEMA_signal_6307, new_AGEMA_signal_6306, new_AGEMA_signal_6305, Inst_bSbox_L8}), .c ({new_AGEMA_signal_6340, new_AGEMA_signal_6339, new_AGEMA_signal_6338, Inst_bSbox_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L19_U1 ( .a ({new_AGEMA_signal_6301, new_AGEMA_signal_6300, new_AGEMA_signal_6299, Inst_bSbox_M63}), .b ({new_AGEMA_signal_6325, new_AGEMA_signal_6324, new_AGEMA_signal_6323, Inst_bSbox_L4}), .c ({new_AGEMA_signal_6361, new_AGEMA_signal_6360, new_AGEMA_signal_6359, Inst_bSbox_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L20_U1 ( .a ({new_AGEMA_signal_6343, new_AGEMA_signal_6342, new_AGEMA_signal_6341, Inst_bSbox_L0}), .b ({new_AGEMA_signal_6304, new_AGEMA_signal_6303, new_AGEMA_signal_6302, Inst_bSbox_L1}), .c ({new_AGEMA_signal_6376, new_AGEMA_signal_6375, new_AGEMA_signal_6374, Inst_bSbox_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L21_U1 ( .a ({new_AGEMA_signal_6304, new_AGEMA_signal_6303, new_AGEMA_signal_6302, Inst_bSbox_L1}), .b ({new_AGEMA_signal_6349, new_AGEMA_signal_6348, new_AGEMA_signal_6347, Inst_bSbox_L7}), .c ({new_AGEMA_signal_6379, new_AGEMA_signal_6378, new_AGEMA_signal_6377, Inst_bSbox_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L22_U1 ( .a ({new_AGEMA_signal_6322, new_AGEMA_signal_6321, new_AGEMA_signal_6320, Inst_bSbox_L3}), .b ({new_AGEMA_signal_6310, new_AGEMA_signal_6309, new_AGEMA_signal_6308, Inst_bSbox_L12}), .c ({new_AGEMA_signal_6364, new_AGEMA_signal_6363, new_AGEMA_signal_6362, Inst_bSbox_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L23_U1 ( .a ({new_AGEMA_signal_6340, new_AGEMA_signal_6339, new_AGEMA_signal_6338, Inst_bSbox_L18}), .b ({new_AGEMA_signal_6319, new_AGEMA_signal_6318, new_AGEMA_signal_6317, Inst_bSbox_L2}), .c ({new_AGEMA_signal_6367, new_AGEMA_signal_6366, new_AGEMA_signal_6365, Inst_bSbox_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L24_U1 ( .a ({new_AGEMA_signal_6334, new_AGEMA_signal_6333, new_AGEMA_signal_6332, Inst_bSbox_L15}), .b ({new_AGEMA_signal_6352, new_AGEMA_signal_6351, new_AGEMA_signal_6350, Inst_bSbox_L9}), .c ({new_AGEMA_signal_6382, new_AGEMA_signal_6381, new_AGEMA_signal_6380, Inst_bSbox_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L25_U1 ( .a ({new_AGEMA_signal_6346, new_AGEMA_signal_6345, new_AGEMA_signal_6344, Inst_bSbox_L6}), .b ({new_AGEMA_signal_6355, new_AGEMA_signal_6354, new_AGEMA_signal_6353, Inst_bSbox_L10}), .c ({new_AGEMA_signal_6385, new_AGEMA_signal_6384, new_AGEMA_signal_6383, Inst_bSbox_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L26_U1 ( .a ({new_AGEMA_signal_6349, new_AGEMA_signal_6348, new_AGEMA_signal_6347, Inst_bSbox_L7}), .b ({new_AGEMA_signal_6352, new_AGEMA_signal_6351, new_AGEMA_signal_6350, Inst_bSbox_L9}), .c ({new_AGEMA_signal_6388, new_AGEMA_signal_6387, new_AGEMA_signal_6386, Inst_bSbox_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L27_U1 ( .a ({new_AGEMA_signal_6307, new_AGEMA_signal_6306, new_AGEMA_signal_6305, Inst_bSbox_L8}), .b ({new_AGEMA_signal_6355, new_AGEMA_signal_6354, new_AGEMA_signal_6353, Inst_bSbox_L10}), .c ({new_AGEMA_signal_6391, new_AGEMA_signal_6390, new_AGEMA_signal_6389, Inst_bSbox_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L28_U1 ( .a ({new_AGEMA_signal_6358, new_AGEMA_signal_6357, new_AGEMA_signal_6356, Inst_bSbox_L11}), .b ({new_AGEMA_signal_6331, new_AGEMA_signal_6330, new_AGEMA_signal_6329, Inst_bSbox_L14}), .c ({new_AGEMA_signal_6394, new_AGEMA_signal_6393, new_AGEMA_signal_6392, Inst_bSbox_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_L29_U1 ( .a ({new_AGEMA_signal_6358, new_AGEMA_signal_6357, new_AGEMA_signal_6356, Inst_bSbox_L11}), .b ({new_AGEMA_signal_6337, new_AGEMA_signal_6336, new_AGEMA_signal_6335, Inst_bSbox_L17}), .c ({new_AGEMA_signal_6397, new_AGEMA_signal_6396, new_AGEMA_signal_6395, Inst_bSbox_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_S0_U1 ( .a ({new_AGEMA_signal_6346, new_AGEMA_signal_6345, new_AGEMA_signal_6344, Inst_bSbox_L6}), .b ({new_AGEMA_signal_6382, new_AGEMA_signal_6381, new_AGEMA_signal_6380, Inst_bSbox_L24}), .c ({new_AGEMA_signal_6409, new_AGEMA_signal_6408, new_AGEMA_signal_6407, SboxOut[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_S1_U1 ( .a ({new_AGEMA_signal_6373, new_AGEMA_signal_6372, new_AGEMA_signal_6371, Inst_bSbox_L16}), .b ({new_AGEMA_signal_6388, new_AGEMA_signal_6387, new_AGEMA_signal_6386, Inst_bSbox_L26}), .c ({new_AGEMA_signal_6412, new_AGEMA_signal_6411, new_AGEMA_signal_6410, SboxOut[6]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_S2_U1 ( .a ({new_AGEMA_signal_6361, new_AGEMA_signal_6360, new_AGEMA_signal_6359, Inst_bSbox_L19}), .b ({new_AGEMA_signal_6394, new_AGEMA_signal_6393, new_AGEMA_signal_6392, Inst_bSbox_L28}), .c ({new_AGEMA_signal_6415, new_AGEMA_signal_6414, new_AGEMA_signal_6413, SboxOut[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_S3_U1 ( .a ({new_AGEMA_signal_6346, new_AGEMA_signal_6345, new_AGEMA_signal_6344, Inst_bSbox_L6}), .b ({new_AGEMA_signal_6379, new_AGEMA_signal_6378, new_AGEMA_signal_6377, Inst_bSbox_L21}), .c ({new_AGEMA_signal_6418, new_AGEMA_signal_6417, new_AGEMA_signal_6416, SboxOut[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_S4_U1 ( .a ({new_AGEMA_signal_6376, new_AGEMA_signal_6375, new_AGEMA_signal_6374, Inst_bSbox_L20}), .b ({new_AGEMA_signal_6364, new_AGEMA_signal_6363, new_AGEMA_signal_6362, Inst_bSbox_L22}), .c ({new_AGEMA_signal_6421, new_AGEMA_signal_6420, new_AGEMA_signal_6419, SboxOut[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_S5_U1 ( .a ({new_AGEMA_signal_6385, new_AGEMA_signal_6384, new_AGEMA_signal_6383, Inst_bSbox_L25}), .b ({new_AGEMA_signal_6397, new_AGEMA_signal_6396, new_AGEMA_signal_6395, Inst_bSbox_L29}), .c ({new_AGEMA_signal_6424, new_AGEMA_signal_6423, new_AGEMA_signal_6422, SboxOut[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_S6_U1 ( .a ({new_AGEMA_signal_6370, new_AGEMA_signal_6369, new_AGEMA_signal_6368, Inst_bSbox_L13}), .b ({new_AGEMA_signal_6391, new_AGEMA_signal_6390, new_AGEMA_signal_6389, Inst_bSbox_L27}), .c ({new_AGEMA_signal_6427, new_AGEMA_signal_6426, new_AGEMA_signal_6425, SboxOut[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Inst_bSbox_XOR_S7_U1 ( .a ({new_AGEMA_signal_6346, new_AGEMA_signal_6345, new_AGEMA_signal_6344, Inst_bSbox_L6}), .b ({new_AGEMA_signal_6367, new_AGEMA_signal_6366, new_AGEMA_signal_6365, Inst_bSbox_L23}), .c ({new_AGEMA_signal_6400, new_AGEMA_signal_6399, new_AGEMA_signal_6398, SboxOut[0]}) ) ;

    /* register cells */
    DFF_X1 ctrl_seq6_SFF_0_Q_reg_FF_FF ( .CK (clk_gated), .D (ctrl_seq6_SFF_0_QD), .Q (ctrl_seq6In_1_), .QN () ) ;
    DFF_X1 ctrl_seq6_SFF_1_Q_reg_FF_FF ( .CK (clk_gated), .D (ctrl_seq6_SFF_1_QD), .Q (ctrl_seq6In_2_), .QN () ) ;
    DFF_X1 ctrl_seq6_SFF_2_Q_reg_FF_FF ( .CK (clk_gated), .D (ctrl_seq6_SFF_2_QD), .Q (ctrl_seq6In_3_), .QN () ) ;
    DFF_X1 ctrl_seq6_SFF_3_Q_reg_FF_FF ( .CK (clk_gated), .D (ctrl_seq6_SFF_3_QD), .Q (ctrl_seq6In_4_), .QN () ) ;
    DFF_X1 ctrl_seq6_SFF_4_Q_reg_FF_FF ( .CK (clk_gated), .D (ctrl_seq6_SFF_4_QD), .Q (ctrl_seq6Out_4_), .QN () ) ;
    DFF_X1 ctrl_seq4_SFF_0_Q_reg_FF_FF ( .CK (clk_gated), .D (ctrl_seq4_SFF_0_QD), .Q (ctrl_seq4In_1_), .QN () ) ;
    DFF_X1 ctrl_seq4_SFF_1_Q_reg_FF_FF ( .CK (clk_gated), .D (ctrl_seq4_SFF_1_QD), .Q (ctrl_seq4Out_1_), .QN () ) ;
    DFF_X1 ctrl_CSselMC_reg_FF_FF ( .CK (clk_gated), .D (ctrl_N14), .Q (ctrl_n6), .QN () ) ;
    DFF_X1 ctrl_CSenRC_reg_FF_FF ( .CK (clk_gated), .D (selSR), .Q (enRCon), .QN () ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5416, new_AGEMA_signal_5415, new_AGEMA_signal_5414, stateArray_S00reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5419, new_AGEMA_signal_5418, new_AGEMA_signal_5417, stateArray_S00reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5422, new_AGEMA_signal_5421, new_AGEMA_signal_5420, stateArray_S00reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5425, new_AGEMA_signal_5424, new_AGEMA_signal_5423, stateArray_S00reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s3[123], ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5428, new_AGEMA_signal_5427, new_AGEMA_signal_5426, stateArray_S00reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5431, new_AGEMA_signal_5430, new_AGEMA_signal_5429, stateArray_S00reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s3[125], ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5434, new_AGEMA_signal_5433, new_AGEMA_signal_5432, stateArray_S00reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s3[126], ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5437, new_AGEMA_signal_5436, new_AGEMA_signal_5435, stateArray_S00reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5440, new_AGEMA_signal_5439, new_AGEMA_signal_5438, stateArray_S01reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s3[112], ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5443, new_AGEMA_signal_5442, new_AGEMA_signal_5441, stateArray_S01reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s3[113], ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5446, new_AGEMA_signal_5445, new_AGEMA_signal_5444, stateArray_S01reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s3[114], ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5449, new_AGEMA_signal_5448, new_AGEMA_signal_5447, stateArray_S01reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s3[115], ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5452, new_AGEMA_signal_5451, new_AGEMA_signal_5450, stateArray_S01reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s3[116], ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5455, new_AGEMA_signal_5454, new_AGEMA_signal_5453, stateArray_S01reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s3[117], ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5458, new_AGEMA_signal_5457, new_AGEMA_signal_5456, stateArray_S01reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s3[118], ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5461, new_AGEMA_signal_5460, new_AGEMA_signal_5459, stateArray_S01reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s3[119], ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5464, new_AGEMA_signal_5463, new_AGEMA_signal_5462, stateArray_S02reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s3[104], ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5467, new_AGEMA_signal_5466, new_AGEMA_signal_5465, stateArray_S02reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s3[105], ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5470, new_AGEMA_signal_5469, new_AGEMA_signal_5468, stateArray_S02reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s3[106], ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5473, new_AGEMA_signal_5472, new_AGEMA_signal_5471, stateArray_S02reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s3[107], ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5476, new_AGEMA_signal_5475, new_AGEMA_signal_5474, stateArray_S02reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s3[108], ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5479, new_AGEMA_signal_5478, new_AGEMA_signal_5477, stateArray_S02reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s3[109], ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5482, new_AGEMA_signal_5481, new_AGEMA_signal_5480, stateArray_S02reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s3[110], ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5485, new_AGEMA_signal_5484, new_AGEMA_signal_5483, stateArray_S02reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s3[111], ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5488, new_AGEMA_signal_5487, new_AGEMA_signal_5486, stateArray_S03reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s3[96], ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5491, new_AGEMA_signal_5490, new_AGEMA_signal_5489, stateArray_S03reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s3[97], ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5494, new_AGEMA_signal_5493, new_AGEMA_signal_5492, stateArray_S03reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s3[98], ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5497, new_AGEMA_signal_5496, new_AGEMA_signal_5495, stateArray_S03reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s3[99], ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5500, new_AGEMA_signal_5499, new_AGEMA_signal_5498, stateArray_S03reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s3[100], ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5503, new_AGEMA_signal_5502, new_AGEMA_signal_5501, stateArray_S03reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s3[101], ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5506, new_AGEMA_signal_5505, new_AGEMA_signal_5504, stateArray_S03reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s3[102], ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5509, new_AGEMA_signal_5508, new_AGEMA_signal_5507, stateArray_S03reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s3[103], ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5512, new_AGEMA_signal_5511, new_AGEMA_signal_5510, stateArray_S10reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5515, new_AGEMA_signal_5514, new_AGEMA_signal_5513, stateArray_S10reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5518, new_AGEMA_signal_5517, new_AGEMA_signal_5516, stateArray_S10reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5521, new_AGEMA_signal_5520, new_AGEMA_signal_5519, stateArray_S10reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s3[91], ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5524, new_AGEMA_signal_5523, new_AGEMA_signal_5522, stateArray_S10reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5527, new_AGEMA_signal_5526, new_AGEMA_signal_5525, stateArray_S10reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s3[93], ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5530, new_AGEMA_signal_5529, new_AGEMA_signal_5528, stateArray_S10reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s3[94], ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5533, new_AGEMA_signal_5532, new_AGEMA_signal_5531, stateArray_S10reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5536, new_AGEMA_signal_5535, new_AGEMA_signal_5534, stateArray_S11reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s3[80], ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5539, new_AGEMA_signal_5538, new_AGEMA_signal_5537, stateArray_S11reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s3[81], ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5542, new_AGEMA_signal_5541, new_AGEMA_signal_5540, stateArray_S11reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s3[82], ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5545, new_AGEMA_signal_5544, new_AGEMA_signal_5543, stateArray_S11reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s3[83], ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5548, new_AGEMA_signal_5547, new_AGEMA_signal_5546, stateArray_S11reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s3[84], ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5551, new_AGEMA_signal_5550, new_AGEMA_signal_5549, stateArray_S11reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s3[85], ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5554, new_AGEMA_signal_5553, new_AGEMA_signal_5552, stateArray_S11reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s3[86], ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5557, new_AGEMA_signal_5556, new_AGEMA_signal_5555, stateArray_S11reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s3[87], ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5560, new_AGEMA_signal_5559, new_AGEMA_signal_5558, stateArray_S12reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s3[72], ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5563, new_AGEMA_signal_5562, new_AGEMA_signal_5561, stateArray_S12reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s3[73], ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5566, new_AGEMA_signal_5565, new_AGEMA_signal_5564, stateArray_S12reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s3[74], ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5569, new_AGEMA_signal_5568, new_AGEMA_signal_5567, stateArray_S12reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s3[75], ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5572, new_AGEMA_signal_5571, new_AGEMA_signal_5570, stateArray_S12reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s3[76], ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5575, new_AGEMA_signal_5574, new_AGEMA_signal_5573, stateArray_S12reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s3[77], ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5578, new_AGEMA_signal_5577, new_AGEMA_signal_5576, stateArray_S12reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s3[78], ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5581, new_AGEMA_signal_5580, new_AGEMA_signal_5579, stateArray_S12reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s3[79], ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5584, new_AGEMA_signal_5583, new_AGEMA_signal_5582, stateArray_S13reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s3[64], ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5587, new_AGEMA_signal_5586, new_AGEMA_signal_5585, stateArray_S13reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s3[65], ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5590, new_AGEMA_signal_5589, new_AGEMA_signal_5588, stateArray_S13reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s3[66], ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5593, new_AGEMA_signal_5592, new_AGEMA_signal_5591, stateArray_S13reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s3[67], ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5596, new_AGEMA_signal_5595, new_AGEMA_signal_5594, stateArray_S13reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s3[68], ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5599, new_AGEMA_signal_5598, new_AGEMA_signal_5597, stateArray_S13reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s3[69], ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5602, new_AGEMA_signal_5601, new_AGEMA_signal_5600, stateArray_S13reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s3[70], ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5605, new_AGEMA_signal_5604, new_AGEMA_signal_5603, stateArray_S13reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s3[71], ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5608, new_AGEMA_signal_5607, new_AGEMA_signal_5606, stateArray_S20reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5611, new_AGEMA_signal_5610, new_AGEMA_signal_5609, stateArray_S20reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5614, new_AGEMA_signal_5613, new_AGEMA_signal_5612, stateArray_S20reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5617, new_AGEMA_signal_5616, new_AGEMA_signal_5615, stateArray_S20reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5620, new_AGEMA_signal_5619, new_AGEMA_signal_5618, stateArray_S20reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5623, new_AGEMA_signal_5622, new_AGEMA_signal_5621, stateArray_S20reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5626, new_AGEMA_signal_5625, new_AGEMA_signal_5624, stateArray_S20reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5629, new_AGEMA_signal_5628, new_AGEMA_signal_5627, stateArray_S20reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5632, new_AGEMA_signal_5631, new_AGEMA_signal_5630, stateArray_S21reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5635, new_AGEMA_signal_5634, new_AGEMA_signal_5633, stateArray_S21reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s3[49], ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5638, new_AGEMA_signal_5637, new_AGEMA_signal_5636, stateArray_S21reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5641, new_AGEMA_signal_5640, new_AGEMA_signal_5639, stateArray_S21reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s3[51], ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5644, new_AGEMA_signal_5643, new_AGEMA_signal_5642, stateArray_S21reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s3[52], ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5647, new_AGEMA_signal_5646, new_AGEMA_signal_5645, stateArray_S21reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s3[53], ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5650, new_AGEMA_signal_5649, new_AGEMA_signal_5648, stateArray_S21reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s3[54], ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5653, new_AGEMA_signal_5652, new_AGEMA_signal_5651, stateArray_S21reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s3[55], ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5656, new_AGEMA_signal_5655, new_AGEMA_signal_5654, stateArray_S22reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5659, new_AGEMA_signal_5658, new_AGEMA_signal_5657, stateArray_S22reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s3[41], ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5662, new_AGEMA_signal_5661, new_AGEMA_signal_5660, stateArray_S22reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5665, new_AGEMA_signal_5664, new_AGEMA_signal_5663, stateArray_S22reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s3[43], ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5668, new_AGEMA_signal_5667, new_AGEMA_signal_5666, stateArray_S22reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s3[44], ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5671, new_AGEMA_signal_5670, new_AGEMA_signal_5669, stateArray_S22reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s3[45], ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5674, new_AGEMA_signal_5673, new_AGEMA_signal_5672, stateArray_S22reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s3[46], ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5677, new_AGEMA_signal_5676, new_AGEMA_signal_5675, stateArray_S22reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s3[47], ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5680, new_AGEMA_signal_5679, new_AGEMA_signal_5678, stateArray_S23reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5683, new_AGEMA_signal_5682, new_AGEMA_signal_5681, stateArray_S23reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s3[33], ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5686, new_AGEMA_signal_5685, new_AGEMA_signal_5684, stateArray_S23reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5689, new_AGEMA_signal_5688, new_AGEMA_signal_5687, stateArray_S23reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s3[35], ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5692, new_AGEMA_signal_5691, new_AGEMA_signal_5690, stateArray_S23reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s3[36], ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5695, new_AGEMA_signal_5694, new_AGEMA_signal_5693, stateArray_S23reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s3[37], ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5698, new_AGEMA_signal_5697, new_AGEMA_signal_5696, stateArray_S23reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s3[38], ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5701, new_AGEMA_signal_5700, new_AGEMA_signal_5699, stateArray_S23reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s3[39], ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5704, new_AGEMA_signal_5703, new_AGEMA_signal_5702, stateArray_S30reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5707, new_AGEMA_signal_5706, new_AGEMA_signal_5705, stateArray_S30reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5710, new_AGEMA_signal_5709, new_AGEMA_signal_5708, stateArray_S30reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5713, new_AGEMA_signal_5712, new_AGEMA_signal_5711, stateArray_S30reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5716, new_AGEMA_signal_5715, new_AGEMA_signal_5714, stateArray_S30reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5719, new_AGEMA_signal_5718, new_AGEMA_signal_5717, stateArray_S30reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5722, new_AGEMA_signal_5721, new_AGEMA_signal_5720, stateArray_S30reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5725, new_AGEMA_signal_5724, new_AGEMA_signal_5723, stateArray_S30reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5728, new_AGEMA_signal_5727, new_AGEMA_signal_5726, stateArray_S31reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5731, new_AGEMA_signal_5730, new_AGEMA_signal_5729, stateArray_S31reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s3[17], ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5734, new_AGEMA_signal_5733, new_AGEMA_signal_5732, stateArray_S31reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5737, new_AGEMA_signal_5736, new_AGEMA_signal_5735, stateArray_S31reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s3[19], ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5740, new_AGEMA_signal_5739, new_AGEMA_signal_5738, stateArray_S31reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s3[20], ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5743, new_AGEMA_signal_5742, new_AGEMA_signal_5741, stateArray_S31reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s3[21], ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5746, new_AGEMA_signal_5745, new_AGEMA_signal_5744, stateArray_S31reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s3[22], ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5749, new_AGEMA_signal_5748, new_AGEMA_signal_5747, stateArray_S31reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s3[23], ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5752, new_AGEMA_signal_5751, new_AGEMA_signal_5750, stateArray_S32reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5755, new_AGEMA_signal_5754, new_AGEMA_signal_5753, stateArray_S32reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s3[9], ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5758, new_AGEMA_signal_5757, new_AGEMA_signal_5756, stateArray_S32reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5761, new_AGEMA_signal_5760, new_AGEMA_signal_5759, stateArray_S32reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s3[11], ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5764, new_AGEMA_signal_5763, new_AGEMA_signal_5762, stateArray_S32reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s3[12], ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5767, new_AGEMA_signal_5766, new_AGEMA_signal_5765, stateArray_S32reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s3[13], ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5770, new_AGEMA_signal_5769, new_AGEMA_signal_5768, stateArray_S32reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s3[14], ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5773, new_AGEMA_signal_5772, new_AGEMA_signal_5771, stateArray_S32reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s3[15], ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6529, new_AGEMA_signal_6528, new_AGEMA_signal_6527, stateArray_S33reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6598, new_AGEMA_signal_6597, new_AGEMA_signal_6596, stateArray_S33reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s3[1], ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6601, new_AGEMA_signal_6600, new_AGEMA_signal_6599, stateArray_S33reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6604, new_AGEMA_signal_6603, new_AGEMA_signal_6602, stateArray_S33reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s3[3], ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6607, new_AGEMA_signal_6606, new_AGEMA_signal_6605, stateArray_S33reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s3[4], ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6610, new_AGEMA_signal_6609, new_AGEMA_signal_6608, stateArray_S33reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s3[5], ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6613, new_AGEMA_signal_6612, new_AGEMA_signal_6611, stateArray_S33reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s3[6], ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6616, new_AGEMA_signal_6615, new_AGEMA_signal_6614, stateArray_S33reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s3[7], ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6163, new_AGEMA_signal_6162, new_AGEMA_signal_6161, KeyArray_S00reg_gff_1_SFF_0_n5}), .Q ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, new_AGEMA_signal_1985, keyStateIn[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6166, new_AGEMA_signal_6165, new_AGEMA_signal_6164, KeyArray_S00reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_1996, new_AGEMA_signal_1995, new_AGEMA_signal_1994, keyStateIn[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6169, new_AGEMA_signal_6168, new_AGEMA_signal_6167, KeyArray_S00reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, new_AGEMA_signal_2003, keyStateIn[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6172, new_AGEMA_signal_6171, new_AGEMA_signal_6170, KeyArray_S00reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_2014, new_AGEMA_signal_2013, new_AGEMA_signal_2012, keyStateIn[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6175, new_AGEMA_signal_6174, new_AGEMA_signal_6173, KeyArray_S00reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, new_AGEMA_signal_2021, keyStateIn[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6178, new_AGEMA_signal_6177, new_AGEMA_signal_6176, KeyArray_S00reg_gff_1_SFF_5_n6}), .Q ({new_AGEMA_signal_2032, new_AGEMA_signal_2031, new_AGEMA_signal_2030, keyStateIn[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6181, new_AGEMA_signal_6180, new_AGEMA_signal_6179, KeyArray_S00reg_gff_1_SFF_6_n6}), .Q ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, new_AGEMA_signal_2039, keyStateIn[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6184, new_AGEMA_signal_6183, new_AGEMA_signal_6182, KeyArray_S00reg_gff_1_SFF_7_n6}), .Q ({new_AGEMA_signal_2050, new_AGEMA_signal_2049, new_AGEMA_signal_2048, keyStateIn[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5863, new_AGEMA_signal_5862, new_AGEMA_signal_5861, KeyArray_S01reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_2098, new_AGEMA_signal_2097, new_AGEMA_signal_2096, KeyArray_outS01ser_0_}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5866, new_AGEMA_signal_5865, new_AGEMA_signal_5864, KeyArray_S01reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_2092, new_AGEMA_signal_2091, new_AGEMA_signal_2090, KeyArray_outS01ser_1_}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5869, new_AGEMA_signal_5868, new_AGEMA_signal_5867, KeyArray_S01reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_2086, new_AGEMA_signal_2085, new_AGEMA_signal_2084, KeyArray_outS01ser_2_}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5872, new_AGEMA_signal_5871, new_AGEMA_signal_5870, KeyArray_S01reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_2080, new_AGEMA_signal_2079, new_AGEMA_signal_2078, KeyArray_outS01ser_3_}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5875, new_AGEMA_signal_5874, new_AGEMA_signal_5873, KeyArray_S01reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_2074, new_AGEMA_signal_2073, new_AGEMA_signal_2072, KeyArray_outS01ser_4_}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5878, new_AGEMA_signal_5877, new_AGEMA_signal_5876, KeyArray_S01reg_gff_1_SFF_5_n6}), .Q ({new_AGEMA_signal_2068, new_AGEMA_signal_2067, new_AGEMA_signal_2066, KeyArray_outS01ser_5_}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5881, new_AGEMA_signal_5880, new_AGEMA_signal_5879, KeyArray_S01reg_gff_1_SFF_6_n6}), .Q ({new_AGEMA_signal_2062, new_AGEMA_signal_2061, new_AGEMA_signal_2060, KeyArray_outS01ser_6_}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5884, new_AGEMA_signal_5883, new_AGEMA_signal_5882, KeyArray_S01reg_gff_1_SFF_7_n6}), .Q ({new_AGEMA_signal_2056, new_AGEMA_signal_2055, new_AGEMA_signal_2054, KeyArray_outS01ser_7_}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5887, new_AGEMA_signal_5886, new_AGEMA_signal_5885, KeyArray_S02reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, new_AGEMA_signal_3365, KeyArray_outS02ser[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5890, new_AGEMA_signal_5889, new_AGEMA_signal_5888, KeyArray_S02reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_3376, new_AGEMA_signal_3375, new_AGEMA_signal_3374, KeyArray_outS02ser[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5893, new_AGEMA_signal_5892, new_AGEMA_signal_5891, KeyArray_S02reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, new_AGEMA_signal_3383, KeyArray_outS02ser[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5896, new_AGEMA_signal_5895, new_AGEMA_signal_5894, KeyArray_S02reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_3394, new_AGEMA_signal_3393, new_AGEMA_signal_3392, KeyArray_outS02ser[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5899, new_AGEMA_signal_5898, new_AGEMA_signal_5897, KeyArray_S02reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, new_AGEMA_signal_3401, KeyArray_outS02ser[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5902, new_AGEMA_signal_5901, new_AGEMA_signal_5900, KeyArray_S02reg_gff_1_SFF_5_n6}), .Q ({new_AGEMA_signal_3412, new_AGEMA_signal_3411, new_AGEMA_signal_3410, KeyArray_outS02ser[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5905, new_AGEMA_signal_5904, new_AGEMA_signal_5903, KeyArray_S02reg_gff_1_SFF_6_n6}), .Q ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, new_AGEMA_signal_3419, KeyArray_outS02ser[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5908, new_AGEMA_signal_5907, new_AGEMA_signal_5906, KeyArray_S02reg_gff_1_SFF_7_n6}), .Q ({new_AGEMA_signal_3430, new_AGEMA_signal_3429, new_AGEMA_signal_3428, KeyArray_outS02ser[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5911, new_AGEMA_signal_5910, new_AGEMA_signal_5909, KeyArray_S03reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_3439, new_AGEMA_signal_3438, new_AGEMA_signal_3437, KeyArray_outS03ser[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5914, new_AGEMA_signal_5913, new_AGEMA_signal_5912, KeyArray_S03reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_3448, new_AGEMA_signal_3447, new_AGEMA_signal_3446, KeyArray_outS03ser[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5917, new_AGEMA_signal_5916, new_AGEMA_signal_5915, KeyArray_S03reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, new_AGEMA_signal_3455, KeyArray_outS03ser[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5920, new_AGEMA_signal_5919, new_AGEMA_signal_5918, KeyArray_S03reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_3466, new_AGEMA_signal_3465, new_AGEMA_signal_3464, KeyArray_outS03ser[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5923, new_AGEMA_signal_5922, new_AGEMA_signal_5921, KeyArray_S03reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, new_AGEMA_signal_3473, KeyArray_outS03ser[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5926, new_AGEMA_signal_5925, new_AGEMA_signal_5924, KeyArray_S03reg_gff_1_SFF_5_n5}), .Q ({new_AGEMA_signal_3484, new_AGEMA_signal_3483, new_AGEMA_signal_3482, KeyArray_outS03ser[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5929, new_AGEMA_signal_5928, new_AGEMA_signal_5927, KeyArray_S03reg_gff_1_SFF_6_n5}), .Q ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, new_AGEMA_signal_3491, KeyArray_outS03ser[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5932, new_AGEMA_signal_5931, new_AGEMA_signal_5930, KeyArray_S03reg_gff_1_SFF_7_n5}), .Q ({new_AGEMA_signal_3502, new_AGEMA_signal_3501, new_AGEMA_signal_3500, KeyArray_outS03ser[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5935, new_AGEMA_signal_5934, new_AGEMA_signal_5933, KeyArray_S10reg_gff_1_SFF_0_n5}), .Q ({new_AGEMA_signal_3511, new_AGEMA_signal_3510, new_AGEMA_signal_3509, KeyArray_outS10ser[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5938, new_AGEMA_signal_5937, new_AGEMA_signal_5936, KeyArray_S10reg_gff_1_SFF_1_n5}), .Q ({new_AGEMA_signal_3520, new_AGEMA_signal_3519, new_AGEMA_signal_3518, KeyArray_outS10ser[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5941, new_AGEMA_signal_5940, new_AGEMA_signal_5939, KeyArray_S10reg_gff_1_SFF_2_n5}), .Q ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, new_AGEMA_signal_3527, KeyArray_outS10ser[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5944, new_AGEMA_signal_5943, new_AGEMA_signal_5942, KeyArray_S10reg_gff_1_SFF_3_n5}), .Q ({new_AGEMA_signal_3538, new_AGEMA_signal_3537, new_AGEMA_signal_3536, KeyArray_outS10ser[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5947, new_AGEMA_signal_5946, new_AGEMA_signal_5945, KeyArray_S10reg_gff_1_SFF_4_n5}), .Q ({new_AGEMA_signal_3547, new_AGEMA_signal_3546, new_AGEMA_signal_3545, KeyArray_outS10ser[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5950, new_AGEMA_signal_5949, new_AGEMA_signal_5948, KeyArray_S10reg_gff_1_SFF_5_n5}), .Q ({new_AGEMA_signal_3556, new_AGEMA_signal_3555, new_AGEMA_signal_3554, KeyArray_outS10ser[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5953, new_AGEMA_signal_5952, new_AGEMA_signal_5951, KeyArray_S10reg_gff_1_SFF_6_n5}), .Q ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, new_AGEMA_signal_3563, KeyArray_outS10ser[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5956, new_AGEMA_signal_5955, new_AGEMA_signal_5954, KeyArray_S10reg_gff_1_SFF_7_n5}), .Q ({new_AGEMA_signal_3574, new_AGEMA_signal_3573, new_AGEMA_signal_3572, KeyArray_outS10ser[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5959, new_AGEMA_signal_5958, new_AGEMA_signal_5957, KeyArray_S11reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, new_AGEMA_signal_3581, KeyArray_outS11ser[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5962, new_AGEMA_signal_5961, new_AGEMA_signal_5960, KeyArray_S11reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_3592, new_AGEMA_signal_3591, new_AGEMA_signal_3590, KeyArray_outS11ser[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5965, new_AGEMA_signal_5964, new_AGEMA_signal_5963, KeyArray_S11reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, new_AGEMA_signal_3599, KeyArray_outS11ser[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5968, new_AGEMA_signal_5967, new_AGEMA_signal_5966, KeyArray_S11reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_3610, new_AGEMA_signal_3609, new_AGEMA_signal_3608, KeyArray_outS11ser[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5971, new_AGEMA_signal_5970, new_AGEMA_signal_5969, KeyArray_S11reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_3619, new_AGEMA_signal_3618, new_AGEMA_signal_3617, KeyArray_outS11ser[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5974, new_AGEMA_signal_5973, new_AGEMA_signal_5972, KeyArray_S11reg_gff_1_SFF_5_n6}), .Q ({new_AGEMA_signal_3628, new_AGEMA_signal_3627, new_AGEMA_signal_3626, KeyArray_outS11ser[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5977, new_AGEMA_signal_5976, new_AGEMA_signal_5975, KeyArray_S11reg_gff_1_SFF_6_n6}), .Q ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, new_AGEMA_signal_3635, KeyArray_outS11ser[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5980, new_AGEMA_signal_5979, new_AGEMA_signal_5978, KeyArray_S11reg_gff_1_SFF_7_n6}), .Q ({new_AGEMA_signal_3646, new_AGEMA_signal_3645, new_AGEMA_signal_3644, KeyArray_outS11ser[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5317, new_AGEMA_signal_5316, new_AGEMA_signal_5315, KeyArray_S12reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_3655, new_AGEMA_signal_3654, new_AGEMA_signal_3653, KeyArray_outS12ser[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5320, new_AGEMA_signal_5319, new_AGEMA_signal_5318, KeyArray_S12reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_3664, new_AGEMA_signal_3663, new_AGEMA_signal_3662, KeyArray_outS12ser[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5323, new_AGEMA_signal_5322, new_AGEMA_signal_5321, KeyArray_S12reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, new_AGEMA_signal_3671, KeyArray_outS12ser[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5326, new_AGEMA_signal_5325, new_AGEMA_signal_5324, KeyArray_S12reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_3682, new_AGEMA_signal_3681, new_AGEMA_signal_3680, KeyArray_outS12ser[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5329, new_AGEMA_signal_5328, new_AGEMA_signal_5327, KeyArray_S12reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_3691, new_AGEMA_signal_3690, new_AGEMA_signal_3689, KeyArray_outS12ser[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5332, new_AGEMA_signal_5331, new_AGEMA_signal_5330, KeyArray_S12reg_gff_1_SFF_5_n6}), .Q ({new_AGEMA_signal_3700, new_AGEMA_signal_3699, new_AGEMA_signal_3698, KeyArray_outS12ser[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5335, new_AGEMA_signal_5334, new_AGEMA_signal_5333, KeyArray_S12reg_gff_1_SFF_6_n6}), .Q ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, new_AGEMA_signal_3707, KeyArray_outS12ser[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5338, new_AGEMA_signal_5337, new_AGEMA_signal_5336, KeyArray_S12reg_gff_1_SFF_7_n6}), .Q ({new_AGEMA_signal_3718, new_AGEMA_signal_3717, new_AGEMA_signal_3716, KeyArray_outS12ser[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5341, new_AGEMA_signal_5340, new_AGEMA_signal_5339, KeyArray_S13reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_3727, new_AGEMA_signal_3726, new_AGEMA_signal_3725, keySBIn[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5344, new_AGEMA_signal_5343, new_AGEMA_signal_5342, KeyArray_S13reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_3736, new_AGEMA_signal_3735, new_AGEMA_signal_3734, keySBIn[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5347, new_AGEMA_signal_5346, new_AGEMA_signal_5345, KeyArray_S13reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_3745, new_AGEMA_signal_3744, new_AGEMA_signal_3743, keySBIn[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5350, new_AGEMA_signal_5349, new_AGEMA_signal_5348, KeyArray_S13reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_3754, new_AGEMA_signal_3753, new_AGEMA_signal_3752, keySBIn[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5353, new_AGEMA_signal_5352, new_AGEMA_signal_5351, KeyArray_S13reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_3763, new_AGEMA_signal_3762, new_AGEMA_signal_3761, keySBIn[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5356, new_AGEMA_signal_5355, new_AGEMA_signal_5354, KeyArray_S13reg_gff_1_SFF_5_n5}), .Q ({new_AGEMA_signal_3772, new_AGEMA_signal_3771, new_AGEMA_signal_3770, keySBIn[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5359, new_AGEMA_signal_5358, new_AGEMA_signal_5357, KeyArray_S13reg_gff_1_SFF_6_n5}), .Q ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, new_AGEMA_signal_3779, keySBIn[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5362, new_AGEMA_signal_5361, new_AGEMA_signal_5360, KeyArray_S13reg_gff_1_SFF_7_n5}), .Q ({new_AGEMA_signal_3790, new_AGEMA_signal_3789, new_AGEMA_signal_3788, keySBIn[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5983, new_AGEMA_signal_5982, new_AGEMA_signal_5981, KeyArray_S20reg_gff_1_SFF_0_n5}), .Q ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, new_AGEMA_signal_3797, KeyArray_outS20ser[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5986, new_AGEMA_signal_5985, new_AGEMA_signal_5984, KeyArray_S20reg_gff_1_SFF_1_n5}), .Q ({new_AGEMA_signal_3808, new_AGEMA_signal_3807, new_AGEMA_signal_3806, KeyArray_outS20ser[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5989, new_AGEMA_signal_5988, new_AGEMA_signal_5987, KeyArray_S20reg_gff_1_SFF_2_n5}), .Q ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, new_AGEMA_signal_3815, KeyArray_outS20ser[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5992, new_AGEMA_signal_5991, new_AGEMA_signal_5990, KeyArray_S20reg_gff_1_SFF_3_n5}), .Q ({new_AGEMA_signal_3826, new_AGEMA_signal_3825, new_AGEMA_signal_3824, KeyArray_outS20ser[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5995, new_AGEMA_signal_5994, new_AGEMA_signal_5993, KeyArray_S20reg_gff_1_SFF_4_n5}), .Q ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, new_AGEMA_signal_3833, KeyArray_outS20ser[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5998, new_AGEMA_signal_5997, new_AGEMA_signal_5996, KeyArray_S20reg_gff_1_SFF_5_n5}), .Q ({new_AGEMA_signal_3844, new_AGEMA_signal_3843, new_AGEMA_signal_3842, KeyArray_outS20ser[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6001, new_AGEMA_signal_6000, new_AGEMA_signal_5999, KeyArray_S20reg_gff_1_SFF_6_n5}), .Q ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, new_AGEMA_signal_3851, KeyArray_outS20ser[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6004, new_AGEMA_signal_6003, new_AGEMA_signal_6002, KeyArray_S20reg_gff_1_SFF_7_n5}), .Q ({new_AGEMA_signal_3862, new_AGEMA_signal_3861, new_AGEMA_signal_3860, KeyArray_outS20ser[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6007, new_AGEMA_signal_6006, new_AGEMA_signal_6005, KeyArray_S21reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, new_AGEMA_signal_3869, KeyArray_outS21ser[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6010, new_AGEMA_signal_6009, new_AGEMA_signal_6008, KeyArray_S21reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_3880, new_AGEMA_signal_3879, new_AGEMA_signal_3878, KeyArray_outS21ser[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6013, new_AGEMA_signal_6012, new_AGEMA_signal_6011, KeyArray_S21reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_3889, new_AGEMA_signal_3888, new_AGEMA_signal_3887, KeyArray_outS21ser[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6016, new_AGEMA_signal_6015, new_AGEMA_signal_6014, KeyArray_S21reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_3898, new_AGEMA_signal_3897, new_AGEMA_signal_3896, KeyArray_outS21ser[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6019, new_AGEMA_signal_6018, new_AGEMA_signal_6017, KeyArray_S21reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_3907, new_AGEMA_signal_3906, new_AGEMA_signal_3905, KeyArray_outS21ser[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6022, new_AGEMA_signal_6021, new_AGEMA_signal_6020, KeyArray_S21reg_gff_1_SFF_5_n6}), .Q ({new_AGEMA_signal_3916, new_AGEMA_signal_3915, new_AGEMA_signal_3914, KeyArray_outS21ser[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6025, new_AGEMA_signal_6024, new_AGEMA_signal_6023, KeyArray_S21reg_gff_1_SFF_6_n6}), .Q ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, new_AGEMA_signal_3923, KeyArray_outS21ser[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6028, new_AGEMA_signal_6027, new_AGEMA_signal_6026, KeyArray_S21reg_gff_1_SFF_7_n6}), .Q ({new_AGEMA_signal_3934, new_AGEMA_signal_3933, new_AGEMA_signal_3932, KeyArray_outS21ser[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6031, new_AGEMA_signal_6030, new_AGEMA_signal_6029, KeyArray_S22reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_3943, new_AGEMA_signal_3942, new_AGEMA_signal_3941, KeyArray_outS22ser[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6034, new_AGEMA_signal_6033, new_AGEMA_signal_6032, KeyArray_S22reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_3952, new_AGEMA_signal_3951, new_AGEMA_signal_3950, KeyArray_outS22ser[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6037, new_AGEMA_signal_6036, new_AGEMA_signal_6035, KeyArray_S22reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_3961, new_AGEMA_signal_3960, new_AGEMA_signal_3959, KeyArray_outS22ser[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6040, new_AGEMA_signal_6039, new_AGEMA_signal_6038, KeyArray_S22reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_3970, new_AGEMA_signal_3969, new_AGEMA_signal_3968, KeyArray_outS22ser[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6043, new_AGEMA_signal_6042, new_AGEMA_signal_6041, KeyArray_S22reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_3979, new_AGEMA_signal_3978, new_AGEMA_signal_3977, KeyArray_outS22ser[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6046, new_AGEMA_signal_6045, new_AGEMA_signal_6044, KeyArray_S22reg_gff_1_SFF_5_n6}), .Q ({new_AGEMA_signal_3988, new_AGEMA_signal_3987, new_AGEMA_signal_3986, KeyArray_outS22ser[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6049, new_AGEMA_signal_6048, new_AGEMA_signal_6047, KeyArray_S22reg_gff_1_SFF_6_n6}), .Q ({new_AGEMA_signal_3997, new_AGEMA_signal_3996, new_AGEMA_signal_3995, KeyArray_outS22ser[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6052, new_AGEMA_signal_6051, new_AGEMA_signal_6050, KeyArray_S22reg_gff_1_SFF_7_n6}), .Q ({new_AGEMA_signal_4006, new_AGEMA_signal_4005, new_AGEMA_signal_4004, KeyArray_outS22ser[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6055, new_AGEMA_signal_6054, new_AGEMA_signal_6053, KeyArray_S23reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_4015, new_AGEMA_signal_4014, new_AGEMA_signal_4013, KeyArray_outS23ser[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6058, new_AGEMA_signal_6057, new_AGEMA_signal_6056, KeyArray_S23reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_4024, new_AGEMA_signal_4023, new_AGEMA_signal_4022, KeyArray_outS23ser[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6061, new_AGEMA_signal_6060, new_AGEMA_signal_6059, KeyArray_S23reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_4033, new_AGEMA_signal_4032, new_AGEMA_signal_4031, KeyArray_outS23ser[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6064, new_AGEMA_signal_6063, new_AGEMA_signal_6062, KeyArray_S23reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_4042, new_AGEMA_signal_4041, new_AGEMA_signal_4040, KeyArray_outS23ser[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6067, new_AGEMA_signal_6066, new_AGEMA_signal_6065, KeyArray_S23reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_4051, new_AGEMA_signal_4050, new_AGEMA_signal_4049, KeyArray_outS23ser[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6070, new_AGEMA_signal_6069, new_AGEMA_signal_6068, KeyArray_S23reg_gff_1_SFF_5_n5}), .Q ({new_AGEMA_signal_4060, new_AGEMA_signal_4059, new_AGEMA_signal_4058, KeyArray_outS23ser[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6073, new_AGEMA_signal_6072, new_AGEMA_signal_6071, KeyArray_S23reg_gff_1_SFF_6_n5}), .Q ({new_AGEMA_signal_4069, new_AGEMA_signal_4068, new_AGEMA_signal_4067, KeyArray_outS23ser[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6076, new_AGEMA_signal_6075, new_AGEMA_signal_6074, KeyArray_S23reg_gff_1_SFF_7_n5}), .Q ({new_AGEMA_signal_4078, new_AGEMA_signal_4077, new_AGEMA_signal_4076, KeyArray_outS23ser[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6574, new_AGEMA_signal_6573, new_AGEMA_signal_6572, KeyArray_S30reg_gff_1_SFF_0_n5}), .Q ({new_AGEMA_signal_4087, new_AGEMA_signal_4086, new_AGEMA_signal_4085, KeyArray_outS30ser[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6619, new_AGEMA_signal_6618, new_AGEMA_signal_6617, KeyArray_S30reg_gff_1_SFF_1_n5}), .Q ({new_AGEMA_signal_4096, new_AGEMA_signal_4095, new_AGEMA_signal_4094, KeyArray_outS30ser[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6622, new_AGEMA_signal_6621, new_AGEMA_signal_6620, KeyArray_S30reg_gff_1_SFF_2_n5}), .Q ({new_AGEMA_signal_4105, new_AGEMA_signal_4104, new_AGEMA_signal_4103, KeyArray_outS30ser[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6625, new_AGEMA_signal_6624, new_AGEMA_signal_6623, KeyArray_S30reg_gff_1_SFF_3_n5}), .Q ({new_AGEMA_signal_4114, new_AGEMA_signal_4113, new_AGEMA_signal_4112, KeyArray_outS30ser[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6628, new_AGEMA_signal_6627, new_AGEMA_signal_6626, KeyArray_S30reg_gff_1_SFF_4_n5}), .Q ({new_AGEMA_signal_4123, new_AGEMA_signal_4122, new_AGEMA_signal_4121, KeyArray_outS30ser[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6631, new_AGEMA_signal_6630, new_AGEMA_signal_6629, KeyArray_S30reg_gff_1_SFF_5_n5}), .Q ({new_AGEMA_signal_4132, new_AGEMA_signal_4131, new_AGEMA_signal_4130, KeyArray_outS30ser[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6634, new_AGEMA_signal_6633, new_AGEMA_signal_6632, KeyArray_S30reg_gff_1_SFF_6_n5}), .Q ({new_AGEMA_signal_4141, new_AGEMA_signal_4140, new_AGEMA_signal_4139, KeyArray_outS30ser[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6637, new_AGEMA_signal_6636, new_AGEMA_signal_6635, KeyArray_S30reg_gff_1_SFF_7_n5}), .Q ({new_AGEMA_signal_4150, new_AGEMA_signal_4149, new_AGEMA_signal_4148, KeyArray_outS30ser[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6079, new_AGEMA_signal_6078, new_AGEMA_signal_6077, KeyArray_S31reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_4159, new_AGEMA_signal_4158, new_AGEMA_signal_4157, KeyArray_outS31ser[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6082, new_AGEMA_signal_6081, new_AGEMA_signal_6080, KeyArray_S31reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_4168, new_AGEMA_signal_4167, new_AGEMA_signal_4166, KeyArray_outS31ser[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6085, new_AGEMA_signal_6084, new_AGEMA_signal_6083, KeyArray_S31reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_4177, new_AGEMA_signal_4176, new_AGEMA_signal_4175, KeyArray_outS31ser[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6088, new_AGEMA_signal_6087, new_AGEMA_signal_6086, KeyArray_S31reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_4186, new_AGEMA_signal_4185, new_AGEMA_signal_4184, KeyArray_outS31ser[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6091, new_AGEMA_signal_6090, new_AGEMA_signal_6089, KeyArray_S31reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_4195, new_AGEMA_signal_4194, new_AGEMA_signal_4193, KeyArray_outS31ser[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6094, new_AGEMA_signal_6093, new_AGEMA_signal_6092, KeyArray_S31reg_gff_1_SFF_5_n6}), .Q ({new_AGEMA_signal_4204, new_AGEMA_signal_4203, new_AGEMA_signal_4202, KeyArray_outS31ser[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6097, new_AGEMA_signal_6096, new_AGEMA_signal_6095, KeyArray_S31reg_gff_1_SFF_6_n6}), .Q ({new_AGEMA_signal_4213, new_AGEMA_signal_4212, new_AGEMA_signal_4211, KeyArray_outS31ser[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6100, new_AGEMA_signal_6099, new_AGEMA_signal_6098, KeyArray_S31reg_gff_1_SFF_7_n6}), .Q ({new_AGEMA_signal_4222, new_AGEMA_signal_4221, new_AGEMA_signal_4220, KeyArray_outS31ser[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6103, new_AGEMA_signal_6102, new_AGEMA_signal_6101, KeyArray_S32reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_4231, new_AGEMA_signal_4230, new_AGEMA_signal_4229, KeyArray_outS32ser[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6106, new_AGEMA_signal_6105, new_AGEMA_signal_6104, KeyArray_S32reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_4240, new_AGEMA_signal_4239, new_AGEMA_signal_4238, KeyArray_outS32ser[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6109, new_AGEMA_signal_6108, new_AGEMA_signal_6107, KeyArray_S32reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_4249, new_AGEMA_signal_4248, new_AGEMA_signal_4247, KeyArray_outS32ser[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6112, new_AGEMA_signal_6111, new_AGEMA_signal_6110, KeyArray_S32reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_4258, new_AGEMA_signal_4257, new_AGEMA_signal_4256, KeyArray_outS32ser[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6115, new_AGEMA_signal_6114, new_AGEMA_signal_6113, KeyArray_S32reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_4267, new_AGEMA_signal_4266, new_AGEMA_signal_4265, KeyArray_outS32ser[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6118, new_AGEMA_signal_6117, new_AGEMA_signal_6116, KeyArray_S32reg_gff_1_SFF_5_n6}), .Q ({new_AGEMA_signal_4276, new_AGEMA_signal_4275, new_AGEMA_signal_4274, KeyArray_outS32ser[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6121, new_AGEMA_signal_6120, new_AGEMA_signal_6119, KeyArray_S32reg_gff_1_SFF_6_n5}), .Q ({new_AGEMA_signal_4285, new_AGEMA_signal_4284, new_AGEMA_signal_4283, KeyArray_outS32ser[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6124, new_AGEMA_signal_6123, new_AGEMA_signal_6122, KeyArray_S32reg_gff_1_SFF_7_n5}), .Q ({new_AGEMA_signal_4294, new_AGEMA_signal_4293, new_AGEMA_signal_4292, KeyArray_outS32ser[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6127, new_AGEMA_signal_6126, new_AGEMA_signal_6125, KeyArray_S33reg_gff_1_SFF_0_n5}), .Q ({new_AGEMA_signal_4303, new_AGEMA_signal_4302, new_AGEMA_signal_4301, KeyArray_outS33ser[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6130, new_AGEMA_signal_6129, new_AGEMA_signal_6128, KeyArray_S33reg_gff_1_SFF_1_n5}), .Q ({new_AGEMA_signal_4312, new_AGEMA_signal_4311, new_AGEMA_signal_4310, KeyArray_outS33ser[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6133, new_AGEMA_signal_6132, new_AGEMA_signal_6131, KeyArray_S33reg_gff_1_SFF_2_n5}), .Q ({new_AGEMA_signal_4321, new_AGEMA_signal_4320, new_AGEMA_signal_4319, KeyArray_outS33ser[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6136, new_AGEMA_signal_6135, new_AGEMA_signal_6134, KeyArray_S33reg_gff_1_SFF_3_n5}), .Q ({new_AGEMA_signal_4330, new_AGEMA_signal_4329, new_AGEMA_signal_4328, KeyArray_outS33ser[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6139, new_AGEMA_signal_6138, new_AGEMA_signal_6137, KeyArray_S33reg_gff_1_SFF_4_n5}), .Q ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, new_AGEMA_signal_4337, KeyArray_outS33ser[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6142, new_AGEMA_signal_6141, new_AGEMA_signal_6140, KeyArray_S33reg_gff_1_SFF_5_n5}), .Q ({new_AGEMA_signal_4348, new_AGEMA_signal_4347, new_AGEMA_signal_4346, KeyArray_outS33ser[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6145, new_AGEMA_signal_6144, new_AGEMA_signal_6143, KeyArray_S33reg_gff_1_SFF_6_n5}), .Q ({new_AGEMA_signal_4357, new_AGEMA_signal_4356, new_AGEMA_signal_4355, KeyArray_outS33ser[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_6148, new_AGEMA_signal_6147, new_AGEMA_signal_6146, KeyArray_S33reg_gff_1_SFF_7_n5}), .Q ({new_AGEMA_signal_4366, new_AGEMA_signal_4365, new_AGEMA_signal_4364, KeyArray_outS33ser[7]}) ) ;
    DFF_X1 calcRCon_s_current_state_reg_0__FF_FF ( .CK (clk_gated), .D (calcRCon_n51), .Q (calcRCon_s_current_state_0_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_1__FF_FF ( .CK (clk_gated), .D (calcRCon_n50), .Q (calcRCon_s_current_state_1_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_2__FF_FF ( .CK (clk_gated), .D (calcRCon_n49), .Q (calcRCon_s_current_state_2_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_3__FF_FF ( .CK (clk_gated), .D (calcRCon_n48), .Q (calcRCon_s_current_state_3_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_4__FF_FF ( .CK (clk_gated), .D (calcRCon_n47), .Q (calcRCon_s_current_state_4_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_5__FF_FF ( .CK (clk_gated), .D (calcRCon_n46), .Q (calcRCon_s_current_state_5_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_6__FF_FF ( .CK (clk_gated), .D (calcRCon_n45), .Q (calcRCon_s_current_state_6_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_7__FF_FF ( .CK (clk_gated), .D (calcRCon_n44), .Q (calcRCon_n3), .QN () ) ;
    DFF_X1 nReset_reg_FF_FF ( .CK (clk_gated), .D (n9), .Q (nReset), .QN () ) ;
endmodule
