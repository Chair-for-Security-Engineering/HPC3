////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module sbox in file Designs/AESSbox/optBP2/AGEMA/sbox.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module sbox_HPC2_ClockGating_d3 (X_s0, clk, X_s1, X_s2, X_s3, Fresh, rst, Y_s0, Y_s1, Y_s2, Y_s3, Synch);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input [7:0] X_s3 ;
    input rst ;
    input [203:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    output [7:0] Y_s3 ;
    output Synch ;
    wire T1 ;
    wire T2 ;
    wire T3 ;
    wire T4 ;
    wire T5 ;
    wire T6 ;
    wire T7 ;
    wire T8 ;
    wire T9 ;
    wire T10 ;
    wire T11 ;
    wire T12 ;
    wire T13 ;
    wire T14 ;
    wire T15 ;
    wire T16 ;
    wire T17 ;
    wire T18 ;
    wire T19 ;
    wire T20 ;
    wire T21 ;
    wire T22 ;
    wire T23 ;
    wire T24 ;
    wire T25 ;
    wire T26 ;
    wire T27 ;
    wire M1 ;
    wire M2 ;
    wire M3 ;
    wire M4 ;
    wire M5 ;
    wire M6 ;
    wire M7 ;
    wire M8 ;
    wire M9 ;
    wire M10 ;
    wire M11 ;
    wire M12 ;
    wire M13 ;
    wire M14 ;
    wire M15 ;
    wire M16 ;
    wire M17 ;
    wire M18 ;
    wire M19 ;
    wire M20 ;
    wire M21 ;
    wire M22 ;
    wire M23 ;
    wire M24 ;
    wire M25 ;
    wire M26 ;
    wire M27 ;
    wire M28 ;
    wire M29 ;
    wire M30 ;
    wire M31 ;
    wire M32 ;
    wire M33 ;
    wire M34 ;
    wire M35 ;
    wire M36 ;
    wire M37 ;
    wire M38 ;
    wire M39 ;
    wire M40 ;
    wire M41 ;
    wire M42 ;
    wire M43 ;
    wire M44 ;
    wire M45 ;
    wire M46 ;
    wire M47 ;
    wire M48 ;
    wire M49 ;
    wire M50 ;
    wire M51 ;
    wire M52 ;
    wire M53 ;
    wire M54 ;
    wire M55 ;
    wire M56 ;
    wire M57 ;
    wire M58 ;
    wire M59 ;
    wire M60 ;
    wire M61 ;
    wire M62 ;
    wire M63 ;
    wire L0 ;
    wire L1 ;
    wire L2 ;
    wire L3 ;
    wire L4 ;
    wire L5 ;
    wire L6 ;
    wire L7 ;
    wire L8 ;
    wire L9 ;
    wire L10 ;
    wire L11 ;
    wire L12 ;
    wire L13 ;
    wire L14 ;
    wire L15 ;
    wire L16 ;
    wire L17 ;
    wire L18 ;
    wire L19 ;
    wire L20 ;
    wire L21 ;
    wire L22 ;
    wire L23 ;
    wire L24 ;
    wire L25 ;
    wire L26 ;
    wire L27 ;
    wire L28 ;
    wire L29 ;
    wire [7:0] O ;
    wire new_AGEMA_signal_157 ;
    wire new_AGEMA_signal_158 ;
    wire new_AGEMA_signal_159 ;
    wire new_AGEMA_signal_163 ;
    wire new_AGEMA_signal_164 ;
    wire new_AGEMA_signal_165 ;
    wire new_AGEMA_signal_169 ;
    wire new_AGEMA_signal_170 ;
    wire new_AGEMA_signal_171 ;
    wire new_AGEMA_signal_172 ;
    wire new_AGEMA_signal_173 ;
    wire new_AGEMA_signal_174 ;
    wire new_AGEMA_signal_178 ;
    wire new_AGEMA_signal_179 ;
    wire new_AGEMA_signal_180 ;
    wire new_AGEMA_signal_187 ;
    wire new_AGEMA_signal_188 ;
    wire new_AGEMA_signal_189 ;
    wire new_AGEMA_signal_190 ;
    wire new_AGEMA_signal_191 ;
    wire new_AGEMA_signal_192 ;
    wire new_AGEMA_signal_193 ;
    wire new_AGEMA_signal_194 ;
    wire new_AGEMA_signal_195 ;
    wire new_AGEMA_signal_199 ;
    wire new_AGEMA_signal_200 ;
    wire new_AGEMA_signal_201 ;
    wire new_AGEMA_signal_202 ;
    wire new_AGEMA_signal_203 ;
    wire new_AGEMA_signal_204 ;
    wire new_AGEMA_signal_205 ;
    wire new_AGEMA_signal_206 ;
    wire new_AGEMA_signal_207 ;
    wire new_AGEMA_signal_208 ;
    wire new_AGEMA_signal_209 ;
    wire new_AGEMA_signal_210 ;
    wire new_AGEMA_signal_211 ;
    wire new_AGEMA_signal_212 ;
    wire new_AGEMA_signal_213 ;
    wire new_AGEMA_signal_214 ;
    wire new_AGEMA_signal_215 ;
    wire new_AGEMA_signal_216 ;
    wire new_AGEMA_signal_217 ;
    wire new_AGEMA_signal_218 ;
    wire new_AGEMA_signal_219 ;
    wire new_AGEMA_signal_220 ;
    wire new_AGEMA_signal_221 ;
    wire new_AGEMA_signal_222 ;
    wire new_AGEMA_signal_223 ;
    wire new_AGEMA_signal_224 ;
    wire new_AGEMA_signal_225 ;
    wire new_AGEMA_signal_226 ;
    wire new_AGEMA_signal_227 ;
    wire new_AGEMA_signal_228 ;
    wire new_AGEMA_signal_229 ;
    wire new_AGEMA_signal_230 ;
    wire new_AGEMA_signal_231 ;
    wire new_AGEMA_signal_232 ;
    wire new_AGEMA_signal_233 ;
    wire new_AGEMA_signal_234 ;
    wire new_AGEMA_signal_235 ;
    wire new_AGEMA_signal_236 ;
    wire new_AGEMA_signal_237 ;
    wire new_AGEMA_signal_238 ;
    wire new_AGEMA_signal_239 ;
    wire new_AGEMA_signal_240 ;
    wire new_AGEMA_signal_241 ;
    wire new_AGEMA_signal_242 ;
    wire new_AGEMA_signal_243 ;
    wire new_AGEMA_signal_244 ;
    wire new_AGEMA_signal_245 ;
    wire new_AGEMA_signal_246 ;
    wire new_AGEMA_signal_247 ;
    wire new_AGEMA_signal_248 ;
    wire new_AGEMA_signal_249 ;
    wire new_AGEMA_signal_250 ;
    wire new_AGEMA_signal_251 ;
    wire new_AGEMA_signal_252 ;
    wire new_AGEMA_signal_253 ;
    wire new_AGEMA_signal_254 ;
    wire new_AGEMA_signal_255 ;
    wire new_AGEMA_signal_256 ;
    wire new_AGEMA_signal_257 ;
    wire new_AGEMA_signal_258 ;
    wire new_AGEMA_signal_259 ;
    wire new_AGEMA_signal_260 ;
    wire new_AGEMA_signal_261 ;
    wire new_AGEMA_signal_262 ;
    wire new_AGEMA_signal_263 ;
    wire new_AGEMA_signal_264 ;
    wire new_AGEMA_signal_265 ;
    wire new_AGEMA_signal_266 ;
    wire new_AGEMA_signal_267 ;
    wire new_AGEMA_signal_268 ;
    wire new_AGEMA_signal_269 ;
    wire new_AGEMA_signal_270 ;
    wire new_AGEMA_signal_271 ;
    wire new_AGEMA_signal_272 ;
    wire new_AGEMA_signal_273 ;
    wire new_AGEMA_signal_274 ;
    wire new_AGEMA_signal_275 ;
    wire new_AGEMA_signal_276 ;
    wire new_AGEMA_signal_277 ;
    wire new_AGEMA_signal_278 ;
    wire new_AGEMA_signal_279 ;
    wire new_AGEMA_signal_280 ;
    wire new_AGEMA_signal_281 ;
    wire new_AGEMA_signal_282 ;
    wire new_AGEMA_signal_283 ;
    wire new_AGEMA_signal_284 ;
    wire new_AGEMA_signal_285 ;
    wire new_AGEMA_signal_286 ;
    wire new_AGEMA_signal_287 ;
    wire new_AGEMA_signal_288 ;
    wire new_AGEMA_signal_289 ;
    wire new_AGEMA_signal_290 ;
    wire new_AGEMA_signal_291 ;
    wire new_AGEMA_signal_292 ;
    wire new_AGEMA_signal_293 ;
    wire new_AGEMA_signal_294 ;
    wire new_AGEMA_signal_295 ;
    wire new_AGEMA_signal_296 ;
    wire new_AGEMA_signal_297 ;
    wire new_AGEMA_signal_298 ;
    wire new_AGEMA_signal_299 ;
    wire new_AGEMA_signal_300 ;
    wire new_AGEMA_signal_301 ;
    wire new_AGEMA_signal_302 ;
    wire new_AGEMA_signal_303 ;
    wire new_AGEMA_signal_304 ;
    wire new_AGEMA_signal_305 ;
    wire new_AGEMA_signal_306 ;
    wire new_AGEMA_signal_307 ;
    wire new_AGEMA_signal_308 ;
    wire new_AGEMA_signal_309 ;
    wire new_AGEMA_signal_310 ;
    wire new_AGEMA_signal_311 ;
    wire new_AGEMA_signal_312 ;
    wire new_AGEMA_signal_313 ;
    wire new_AGEMA_signal_314 ;
    wire new_AGEMA_signal_315 ;
    wire new_AGEMA_signal_316 ;
    wire new_AGEMA_signal_317 ;
    wire new_AGEMA_signal_318 ;
    wire new_AGEMA_signal_319 ;
    wire new_AGEMA_signal_320 ;
    wire new_AGEMA_signal_321 ;
    wire new_AGEMA_signal_322 ;
    wire new_AGEMA_signal_323 ;
    wire new_AGEMA_signal_324 ;
    wire new_AGEMA_signal_325 ;
    wire new_AGEMA_signal_326 ;
    wire new_AGEMA_signal_327 ;
    wire new_AGEMA_signal_328 ;
    wire new_AGEMA_signal_329 ;
    wire new_AGEMA_signal_330 ;
    wire new_AGEMA_signal_331 ;
    wire new_AGEMA_signal_332 ;
    wire new_AGEMA_signal_333 ;
    wire new_AGEMA_signal_334 ;
    wire new_AGEMA_signal_335 ;
    wire new_AGEMA_signal_336 ;
    wire new_AGEMA_signal_337 ;
    wire new_AGEMA_signal_338 ;
    wire new_AGEMA_signal_339 ;
    wire new_AGEMA_signal_340 ;
    wire new_AGEMA_signal_341 ;
    wire new_AGEMA_signal_342 ;
    wire new_AGEMA_signal_343 ;
    wire new_AGEMA_signal_344 ;
    wire new_AGEMA_signal_345 ;
    wire new_AGEMA_signal_346 ;
    wire new_AGEMA_signal_347 ;
    wire new_AGEMA_signal_348 ;
    wire new_AGEMA_signal_349 ;
    wire new_AGEMA_signal_350 ;
    wire new_AGEMA_signal_351 ;
    wire new_AGEMA_signal_352 ;
    wire new_AGEMA_signal_353 ;
    wire new_AGEMA_signal_354 ;
    wire new_AGEMA_signal_355 ;
    wire new_AGEMA_signal_356 ;
    wire new_AGEMA_signal_357 ;
    wire new_AGEMA_signal_358 ;
    wire new_AGEMA_signal_359 ;
    wire new_AGEMA_signal_360 ;
    wire new_AGEMA_signal_361 ;
    wire new_AGEMA_signal_362 ;
    wire new_AGEMA_signal_363 ;
    wire new_AGEMA_signal_364 ;
    wire new_AGEMA_signal_365 ;
    wire new_AGEMA_signal_366 ;
    wire new_AGEMA_signal_367 ;
    wire new_AGEMA_signal_368 ;
    wire new_AGEMA_signal_369 ;
    wire new_AGEMA_signal_370 ;
    wire new_AGEMA_signal_371 ;
    wire new_AGEMA_signal_372 ;
    wire new_AGEMA_signal_373 ;
    wire new_AGEMA_signal_374 ;
    wire new_AGEMA_signal_375 ;
    wire new_AGEMA_signal_376 ;
    wire new_AGEMA_signal_377 ;
    wire new_AGEMA_signal_378 ;
    wire new_AGEMA_signal_379 ;
    wire new_AGEMA_signal_380 ;
    wire new_AGEMA_signal_381 ;
    wire new_AGEMA_signal_382 ;
    wire new_AGEMA_signal_383 ;
    wire new_AGEMA_signal_384 ;
    wire new_AGEMA_signal_385 ;
    wire new_AGEMA_signal_386 ;
    wire new_AGEMA_signal_387 ;
    wire new_AGEMA_signal_388 ;
    wire new_AGEMA_signal_389 ;
    wire new_AGEMA_signal_390 ;
    wire new_AGEMA_signal_391 ;
    wire new_AGEMA_signal_392 ;
    wire new_AGEMA_signal_393 ;
    wire new_AGEMA_signal_394 ;
    wire new_AGEMA_signal_395 ;
    wire new_AGEMA_signal_396 ;
    wire new_AGEMA_signal_397 ;
    wire new_AGEMA_signal_398 ;
    wire new_AGEMA_signal_399 ;
    wire new_AGEMA_signal_400 ;
    wire new_AGEMA_signal_401 ;
    wire new_AGEMA_signal_402 ;
    wire new_AGEMA_signal_403 ;
    wire new_AGEMA_signal_404 ;
    wire new_AGEMA_signal_405 ;
    wire new_AGEMA_signal_406 ;
    wire new_AGEMA_signal_407 ;
    wire new_AGEMA_signal_408 ;
    wire new_AGEMA_signal_409 ;
    wire new_AGEMA_signal_410 ;
    wire new_AGEMA_signal_411 ;
    wire new_AGEMA_signal_412 ;
    wire new_AGEMA_signal_413 ;
    wire new_AGEMA_signal_414 ;
    wire new_AGEMA_signal_415 ;
    wire new_AGEMA_signal_416 ;
    wire new_AGEMA_signal_417 ;
    wire new_AGEMA_signal_418 ;
    wire new_AGEMA_signal_419 ;
    wire new_AGEMA_signal_420 ;
    wire new_AGEMA_signal_421 ;
    wire new_AGEMA_signal_422 ;
    wire new_AGEMA_signal_423 ;
    wire new_AGEMA_signal_424 ;
    wire new_AGEMA_signal_425 ;
    wire new_AGEMA_signal_426 ;
    wire new_AGEMA_signal_427 ;
    wire new_AGEMA_signal_428 ;
    wire new_AGEMA_signal_429 ;
    wire new_AGEMA_signal_430 ;
    wire new_AGEMA_signal_431 ;
    wire new_AGEMA_signal_432 ;
    wire new_AGEMA_signal_433 ;
    wire new_AGEMA_signal_434 ;
    wire new_AGEMA_signal_435 ;
    wire new_AGEMA_signal_436 ;
    wire new_AGEMA_signal_437 ;
    wire new_AGEMA_signal_438 ;
    wire new_AGEMA_signal_439 ;
    wire new_AGEMA_signal_440 ;
    wire new_AGEMA_signal_441 ;
    wire new_AGEMA_signal_442 ;
    wire new_AGEMA_signal_443 ;
    wire new_AGEMA_signal_444 ;
    wire new_AGEMA_signal_445 ;
    wire new_AGEMA_signal_446 ;
    wire new_AGEMA_signal_447 ;
    wire new_AGEMA_signal_448 ;
    wire new_AGEMA_signal_449 ;
    wire new_AGEMA_signal_450 ;
    wire new_AGEMA_signal_451 ;
    wire new_AGEMA_signal_452 ;
    wire new_AGEMA_signal_453 ;
    wire new_AGEMA_signal_454 ;
    wire new_AGEMA_signal_455 ;
    wire new_AGEMA_signal_456 ;
    wire new_AGEMA_signal_457 ;
    wire new_AGEMA_signal_458 ;
    wire new_AGEMA_signal_459 ;
    wire new_AGEMA_signal_460 ;
    wire new_AGEMA_signal_461 ;
    wire new_AGEMA_signal_462 ;
    wire new_AGEMA_signal_463 ;
    wire new_AGEMA_signal_464 ;
    wire new_AGEMA_signal_465 ;
    wire new_AGEMA_signal_466 ;
    wire new_AGEMA_signal_467 ;
    wire new_AGEMA_signal_468 ;
    wire new_AGEMA_signal_469 ;
    wire new_AGEMA_signal_470 ;
    wire new_AGEMA_signal_471 ;
    wire new_AGEMA_signal_472 ;
    wire new_AGEMA_signal_473 ;
    wire new_AGEMA_signal_474 ;
    wire new_AGEMA_signal_475 ;
    wire new_AGEMA_signal_476 ;
    wire new_AGEMA_signal_477 ;
    wire new_AGEMA_signal_478 ;
    wire new_AGEMA_signal_479 ;
    wire new_AGEMA_signal_480 ;
    wire new_AGEMA_signal_481 ;
    wire new_AGEMA_signal_482 ;
    wire new_AGEMA_signal_483 ;
    wire new_AGEMA_signal_484 ;
    wire new_AGEMA_signal_485 ;
    wire new_AGEMA_signal_486 ;
    wire new_AGEMA_signal_487 ;
    wire new_AGEMA_signal_488 ;
    wire new_AGEMA_signal_489 ;
    wire new_AGEMA_signal_490 ;
    wire new_AGEMA_signal_491 ;
    wire new_AGEMA_signal_492 ;
    wire new_AGEMA_signal_493 ;
    wire new_AGEMA_signal_494 ;
    wire new_AGEMA_signal_495 ;
    wire new_AGEMA_signal_496 ;
    wire new_AGEMA_signal_497 ;
    wire new_AGEMA_signal_498 ;
    wire new_AGEMA_signal_499 ;
    wire new_AGEMA_signal_500 ;
    wire new_AGEMA_signal_501 ;
    wire new_AGEMA_signal_502 ;
    wire new_AGEMA_signal_503 ;
    wire new_AGEMA_signal_504 ;
    wire new_AGEMA_signal_505 ;
    wire new_AGEMA_signal_506 ;
    wire new_AGEMA_signal_507 ;
    wire new_AGEMA_signal_508 ;
    wire new_AGEMA_signal_509 ;
    wire new_AGEMA_signal_510 ;
    wire new_AGEMA_signal_511 ;
    wire new_AGEMA_signal_512 ;
    wire new_AGEMA_signal_513 ;
    wire new_AGEMA_signal_514 ;
    wire new_AGEMA_signal_515 ;
    wire new_AGEMA_signal_516 ;
    wire new_AGEMA_signal_517 ;
    wire new_AGEMA_signal_518 ;
    wire new_AGEMA_signal_519 ;
    wire new_AGEMA_signal_520 ;
    wire new_AGEMA_signal_521 ;
    wire new_AGEMA_signal_522 ;
    wire new_AGEMA_signal_523 ;
    wire new_AGEMA_signal_524 ;
    wire new_AGEMA_signal_525 ;
    wire new_AGEMA_signal_526 ;
    wire new_AGEMA_signal_527 ;
    wire new_AGEMA_signal_528 ;
    wire new_AGEMA_signal_529 ;
    wire new_AGEMA_signal_530 ;
    wire new_AGEMA_signal_531 ;
    wire new_AGEMA_signal_532 ;
    wire new_AGEMA_signal_533 ;
    wire new_AGEMA_signal_534 ;
    wire new_AGEMA_signal_535 ;
    wire new_AGEMA_signal_536 ;
    wire new_AGEMA_signal_537 ;
    wire new_AGEMA_signal_538 ;
    wire new_AGEMA_signal_539 ;
    wire new_AGEMA_signal_540 ;
    wire new_AGEMA_signal_541 ;
    wire new_AGEMA_signal_542 ;
    wire new_AGEMA_signal_543 ;
    wire new_AGEMA_signal_544 ;
    wire new_AGEMA_signal_545 ;
    wire new_AGEMA_signal_546 ;
    wire new_AGEMA_signal_547 ;
    wire new_AGEMA_signal_548 ;
    wire new_AGEMA_signal_549 ;
    wire new_AGEMA_signal_550 ;
    wire new_AGEMA_signal_551 ;
    wire new_AGEMA_signal_552 ;
    wire new_AGEMA_signal_553 ;
    wire new_AGEMA_signal_554 ;
    wire new_AGEMA_signal_555 ;
    wire new_AGEMA_signal_556 ;
    wire new_AGEMA_signal_557 ;
    wire new_AGEMA_signal_558 ;
    wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T1_U1 ( .a ({X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .c ({new_AGEMA_signal_159, new_AGEMA_signal_158, new_AGEMA_signal_157, T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T2_U1 ( .a ({X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_165, new_AGEMA_signal_164, new_AGEMA_signal_163, T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T3_U1 ( .a ({X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .c ({new_AGEMA_signal_171, new_AGEMA_signal_170, new_AGEMA_signal_169, T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T4_U1 ( .a ({X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_174, new_AGEMA_signal_173, new_AGEMA_signal_172, T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T5_U1 ( .a ({X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .c ({new_AGEMA_signal_180, new_AGEMA_signal_179, new_AGEMA_signal_178, T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T6_U1 ( .a ({new_AGEMA_signal_159, new_AGEMA_signal_158, new_AGEMA_signal_157, T1}), .b ({new_AGEMA_signal_180, new_AGEMA_signal_179, new_AGEMA_signal_178, T5}), .c ({new_AGEMA_signal_207, new_AGEMA_signal_206, new_AGEMA_signal_205, T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T7_U1 ( .a ({X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .c ({new_AGEMA_signal_189, new_AGEMA_signal_188, new_AGEMA_signal_187, T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T8_U1 ( .a ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({new_AGEMA_signal_207, new_AGEMA_signal_206, new_AGEMA_signal_205, T6}), .c ({new_AGEMA_signal_231, new_AGEMA_signal_230, new_AGEMA_signal_229, T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T9_U1 ( .a ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({new_AGEMA_signal_189, new_AGEMA_signal_188, new_AGEMA_signal_187, T7}), .c ({new_AGEMA_signal_210, new_AGEMA_signal_209, new_AGEMA_signal_208, T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T10_U1 ( .a ({new_AGEMA_signal_207, new_AGEMA_signal_206, new_AGEMA_signal_205, T6}), .b ({new_AGEMA_signal_189, new_AGEMA_signal_188, new_AGEMA_signal_187, T7}), .c ({new_AGEMA_signal_234, new_AGEMA_signal_233, new_AGEMA_signal_232, T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T11_U1 ( .a ({X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_192, new_AGEMA_signal_191, new_AGEMA_signal_190, T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T12_U1 ( .a ({X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_195, new_AGEMA_signal_194, new_AGEMA_signal_193, T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T13_U1 ( .a ({new_AGEMA_signal_171, new_AGEMA_signal_170, new_AGEMA_signal_169, T3}), .b ({new_AGEMA_signal_174, new_AGEMA_signal_173, new_AGEMA_signal_172, T4}), .c ({new_AGEMA_signal_213, new_AGEMA_signal_212, new_AGEMA_signal_211, T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T14_U1 ( .a ({new_AGEMA_signal_207, new_AGEMA_signal_206, new_AGEMA_signal_205, T6}), .b ({new_AGEMA_signal_192, new_AGEMA_signal_191, new_AGEMA_signal_190, T11}), .c ({new_AGEMA_signal_237, new_AGEMA_signal_236, new_AGEMA_signal_235, T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T15_U1 ( .a ({new_AGEMA_signal_180, new_AGEMA_signal_179, new_AGEMA_signal_178, T5}), .b ({new_AGEMA_signal_192, new_AGEMA_signal_191, new_AGEMA_signal_190, T11}), .c ({new_AGEMA_signal_216, new_AGEMA_signal_215, new_AGEMA_signal_214, T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T16_U1 ( .a ({new_AGEMA_signal_180, new_AGEMA_signal_179, new_AGEMA_signal_178, T5}), .b ({new_AGEMA_signal_195, new_AGEMA_signal_194, new_AGEMA_signal_193, T12}), .c ({new_AGEMA_signal_219, new_AGEMA_signal_218, new_AGEMA_signal_217, T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T17_U1 ( .a ({new_AGEMA_signal_210, new_AGEMA_signal_209, new_AGEMA_signal_208, T9}), .b ({new_AGEMA_signal_219, new_AGEMA_signal_218, new_AGEMA_signal_217, T16}), .c ({new_AGEMA_signal_240, new_AGEMA_signal_239, new_AGEMA_signal_238, T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T18_U1 ( .a ({X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({new_AGEMA_signal_201, new_AGEMA_signal_200, new_AGEMA_signal_199, T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T19_U1 ( .a ({new_AGEMA_signal_189, new_AGEMA_signal_188, new_AGEMA_signal_187, T7}), .b ({new_AGEMA_signal_201, new_AGEMA_signal_200, new_AGEMA_signal_199, T18}), .c ({new_AGEMA_signal_222, new_AGEMA_signal_221, new_AGEMA_signal_220, T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T20_U1 ( .a ({new_AGEMA_signal_159, new_AGEMA_signal_158, new_AGEMA_signal_157, T1}), .b ({new_AGEMA_signal_222, new_AGEMA_signal_221, new_AGEMA_signal_220, T19}), .c ({new_AGEMA_signal_243, new_AGEMA_signal_242, new_AGEMA_signal_241, T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T21_U1 ( .a ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({new_AGEMA_signal_204, new_AGEMA_signal_203, new_AGEMA_signal_202, T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T22_U1 ( .a ({new_AGEMA_signal_189, new_AGEMA_signal_188, new_AGEMA_signal_187, T7}), .b ({new_AGEMA_signal_204, new_AGEMA_signal_203, new_AGEMA_signal_202, T21}), .c ({new_AGEMA_signal_225, new_AGEMA_signal_224, new_AGEMA_signal_223, T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T23_U1 ( .a ({new_AGEMA_signal_165, new_AGEMA_signal_164, new_AGEMA_signal_163, T2}), .b ({new_AGEMA_signal_225, new_AGEMA_signal_224, new_AGEMA_signal_223, T22}), .c ({new_AGEMA_signal_246, new_AGEMA_signal_245, new_AGEMA_signal_244, T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T24_U1 ( .a ({new_AGEMA_signal_165, new_AGEMA_signal_164, new_AGEMA_signal_163, T2}), .b ({new_AGEMA_signal_234, new_AGEMA_signal_233, new_AGEMA_signal_232, T10}), .c ({new_AGEMA_signal_270, new_AGEMA_signal_269, new_AGEMA_signal_268, T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T25_U1 ( .a ({new_AGEMA_signal_243, new_AGEMA_signal_242, new_AGEMA_signal_241, T20}), .b ({new_AGEMA_signal_240, new_AGEMA_signal_239, new_AGEMA_signal_238, T17}), .c ({new_AGEMA_signal_273, new_AGEMA_signal_272, new_AGEMA_signal_271, T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T26_U1 ( .a ({new_AGEMA_signal_171, new_AGEMA_signal_170, new_AGEMA_signal_169, T3}), .b ({new_AGEMA_signal_219, new_AGEMA_signal_218, new_AGEMA_signal_217, T16}), .c ({new_AGEMA_signal_249, new_AGEMA_signal_248, new_AGEMA_signal_247, T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_T27_U1 ( .a ({new_AGEMA_signal_159, new_AGEMA_signal_158, new_AGEMA_signal_157, T1}), .b ({new_AGEMA_signal_195, new_AGEMA_signal_194, new_AGEMA_signal_193, T12}), .c ({new_AGEMA_signal_228, new_AGEMA_signal_227, new_AGEMA_signal_226, T27}) ) ;
    

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M1_U1 ( .a ({new_AGEMA_signal_213, new_AGEMA_signal_212, new_AGEMA_signal_211, T13}), .b ({new_AGEMA_signal_207, new_AGEMA_signal_206, new_AGEMA_signal_205, T6}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_252, new_AGEMA_signal_251, new_AGEMA_signal_250, M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M2_U1 ( .a ({new_AGEMA_signal_246, new_AGEMA_signal_245, new_AGEMA_signal_244, T23}), .b ({new_AGEMA_signal_231, new_AGEMA_signal_230, new_AGEMA_signal_229, T8}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_276, new_AGEMA_signal_275, new_AGEMA_signal_274, M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M3_U1 ( .a ({new_AGEMA_signal_237, new_AGEMA_signal_236, new_AGEMA_signal_235, T14}), .b ({new_AGEMA_signal_252, new_AGEMA_signal_251, new_AGEMA_signal_250, M1}), .c ({new_AGEMA_signal_279, new_AGEMA_signal_278, new_AGEMA_signal_277, M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M4_U1 ( .a ({new_AGEMA_signal_222, new_AGEMA_signal_221, new_AGEMA_signal_220, T19}), .b ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_255, new_AGEMA_signal_254, new_AGEMA_signal_253, M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M5_U1 ( .a ({new_AGEMA_signal_255, new_AGEMA_signal_254, new_AGEMA_signal_253, M4}), .b ({new_AGEMA_signal_252, new_AGEMA_signal_251, new_AGEMA_signal_250, M1}), .c ({new_AGEMA_signal_282, new_AGEMA_signal_281, new_AGEMA_signal_280, M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M6_U1 ( .a ({new_AGEMA_signal_171, new_AGEMA_signal_170, new_AGEMA_signal_169, T3}), .b ({new_AGEMA_signal_219, new_AGEMA_signal_218, new_AGEMA_signal_217, T16}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_258, new_AGEMA_signal_257, new_AGEMA_signal_256, M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M7_U1 ( .a ({new_AGEMA_signal_225, new_AGEMA_signal_224, new_AGEMA_signal_223, T22}), .b ({new_AGEMA_signal_210, new_AGEMA_signal_209, new_AGEMA_signal_208, T9}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_261, new_AGEMA_signal_260, new_AGEMA_signal_259, M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M8_U1 ( .a ({new_AGEMA_signal_249, new_AGEMA_signal_248, new_AGEMA_signal_247, T26}), .b ({new_AGEMA_signal_258, new_AGEMA_signal_257, new_AGEMA_signal_256, M6}), .c ({new_AGEMA_signal_285, new_AGEMA_signal_284, new_AGEMA_signal_283, M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M9_U1 ( .a ({new_AGEMA_signal_243, new_AGEMA_signal_242, new_AGEMA_signal_241, T20}), .b ({new_AGEMA_signal_240, new_AGEMA_signal_239, new_AGEMA_signal_238, T17}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_288, new_AGEMA_signal_287, new_AGEMA_signal_286, M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M10_U1 ( .a ({new_AGEMA_signal_288, new_AGEMA_signal_287, new_AGEMA_signal_286, M9}), .b ({new_AGEMA_signal_258, new_AGEMA_signal_257, new_AGEMA_signal_256, M6}), .c ({new_AGEMA_signal_297, new_AGEMA_signal_296, new_AGEMA_signal_295, M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M11_U1 ( .a ({new_AGEMA_signal_159, new_AGEMA_signal_158, new_AGEMA_signal_157, T1}), .b ({new_AGEMA_signal_216, new_AGEMA_signal_215, new_AGEMA_signal_214, T15}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_264, new_AGEMA_signal_263, new_AGEMA_signal_262, M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M12_U1 ( .a ({new_AGEMA_signal_174, new_AGEMA_signal_173, new_AGEMA_signal_172, T4}), .b ({new_AGEMA_signal_228, new_AGEMA_signal_227, new_AGEMA_signal_226, T27}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_267, new_AGEMA_signal_266, new_AGEMA_signal_265, M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M13_U1 ( .a ({new_AGEMA_signal_267, new_AGEMA_signal_266, new_AGEMA_signal_265, M12}), .b ({new_AGEMA_signal_264, new_AGEMA_signal_263, new_AGEMA_signal_262, M11}), .c ({new_AGEMA_signal_291, new_AGEMA_signal_290, new_AGEMA_signal_289, M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M14_U1 ( .a ({new_AGEMA_signal_165, new_AGEMA_signal_164, new_AGEMA_signal_163, T2}), .b ({new_AGEMA_signal_234, new_AGEMA_signal_233, new_AGEMA_signal_232, T10}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_294, new_AGEMA_signal_293, new_AGEMA_signal_292, M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M15_U1 ( .a ({new_AGEMA_signal_294, new_AGEMA_signal_293, new_AGEMA_signal_292, M14}), .b ({new_AGEMA_signal_264, new_AGEMA_signal_263, new_AGEMA_signal_262, M11}), .c ({new_AGEMA_signal_300, new_AGEMA_signal_299, new_AGEMA_signal_298, M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M16_U1 ( .a ({new_AGEMA_signal_279, new_AGEMA_signal_278, new_AGEMA_signal_277, M3}), .b ({new_AGEMA_signal_276, new_AGEMA_signal_275, new_AGEMA_signal_274, M2}), .c ({new_AGEMA_signal_303, new_AGEMA_signal_302, new_AGEMA_signal_301, M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M17_U1 ( .a ({new_AGEMA_signal_282, new_AGEMA_signal_281, new_AGEMA_signal_280, M5}), .b ({new_AGEMA_signal_270, new_AGEMA_signal_269, new_AGEMA_signal_268, T24}), .c ({new_AGEMA_signal_306, new_AGEMA_signal_305, new_AGEMA_signal_304, M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M18_U1 ( .a ({new_AGEMA_signal_285, new_AGEMA_signal_284, new_AGEMA_signal_283, M8}), .b ({new_AGEMA_signal_261, new_AGEMA_signal_260, new_AGEMA_signal_259, M7}), .c ({new_AGEMA_signal_309, new_AGEMA_signal_308, new_AGEMA_signal_307, M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M19_U1 ( .a ({new_AGEMA_signal_297, new_AGEMA_signal_296, new_AGEMA_signal_295, M10}), .b ({new_AGEMA_signal_300, new_AGEMA_signal_299, new_AGEMA_signal_298, M15}), .c ({new_AGEMA_signal_312, new_AGEMA_signal_311, new_AGEMA_signal_310, M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M20_U1 ( .a ({new_AGEMA_signal_303, new_AGEMA_signal_302, new_AGEMA_signal_301, M16}), .b ({new_AGEMA_signal_291, new_AGEMA_signal_290, new_AGEMA_signal_289, M13}), .c ({new_AGEMA_signal_315, new_AGEMA_signal_314, new_AGEMA_signal_313, M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M21_U1 ( .a ({new_AGEMA_signal_306, new_AGEMA_signal_305, new_AGEMA_signal_304, M17}), .b ({new_AGEMA_signal_300, new_AGEMA_signal_299, new_AGEMA_signal_298, M15}), .c ({new_AGEMA_signal_318, new_AGEMA_signal_317, new_AGEMA_signal_316, M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M22_U1 ( .a ({new_AGEMA_signal_309, new_AGEMA_signal_308, new_AGEMA_signal_307, M18}), .b ({new_AGEMA_signal_291, new_AGEMA_signal_290, new_AGEMA_signal_289, M13}), .c ({new_AGEMA_signal_321, new_AGEMA_signal_320, new_AGEMA_signal_319, M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M23_U1 ( .a ({new_AGEMA_signal_312, new_AGEMA_signal_311, new_AGEMA_signal_310, M19}), .b ({new_AGEMA_signal_273, new_AGEMA_signal_272, new_AGEMA_signal_271, T25}), .c ({new_AGEMA_signal_324, new_AGEMA_signal_323, new_AGEMA_signal_322, M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M24_U1 ( .a ({new_AGEMA_signal_321, new_AGEMA_signal_320, new_AGEMA_signal_319, M22}), .b ({new_AGEMA_signal_324, new_AGEMA_signal_323, new_AGEMA_signal_322, M23}), .c ({new_AGEMA_signal_336, new_AGEMA_signal_335, new_AGEMA_signal_334, M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M27_U1 ( .a ({new_AGEMA_signal_315, new_AGEMA_signal_314, new_AGEMA_signal_313, M20}), .b ({new_AGEMA_signal_318, new_AGEMA_signal_317, new_AGEMA_signal_316, M21}), .c ({new_AGEMA_signal_330, new_AGEMA_signal_329, new_AGEMA_signal_328, M27}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M25_U1 ( .a ({new_AGEMA_signal_321, new_AGEMA_signal_320, new_AGEMA_signal_319, M22}), .b ({new_AGEMA_signal_315, new_AGEMA_signal_314, new_AGEMA_signal_313, M20}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_327, new_AGEMA_signal_326, new_AGEMA_signal_325, M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M26_U1 ( .a ({new_AGEMA_signal_318, new_AGEMA_signal_317, new_AGEMA_signal_316, M21}), .b ({new_AGEMA_signal_327, new_AGEMA_signal_326, new_AGEMA_signal_325, M25}), .c ({new_AGEMA_signal_339, new_AGEMA_signal_338, new_AGEMA_signal_337, M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M28_U1 ( .a ({new_AGEMA_signal_324, new_AGEMA_signal_323, new_AGEMA_signal_322, M23}), .b ({new_AGEMA_signal_327, new_AGEMA_signal_326, new_AGEMA_signal_325, M25}), .c ({new_AGEMA_signal_342, new_AGEMA_signal_341, new_AGEMA_signal_340, M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M31_U1 ( .a ({new_AGEMA_signal_315, new_AGEMA_signal_314, new_AGEMA_signal_313, M20}), .b ({new_AGEMA_signal_324, new_AGEMA_signal_323, new_AGEMA_signal_322, M23}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_345, new_AGEMA_signal_344, new_AGEMA_signal_343, M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M33_U1 ( .a ({new_AGEMA_signal_330, new_AGEMA_signal_329, new_AGEMA_signal_328, M27}), .b ({new_AGEMA_signal_327, new_AGEMA_signal_326, new_AGEMA_signal_325, M25}), .c ({new_AGEMA_signal_348, new_AGEMA_signal_347, new_AGEMA_signal_346, M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M34_U1 ( .a ({new_AGEMA_signal_318, new_AGEMA_signal_317, new_AGEMA_signal_316, M21}), .b ({new_AGEMA_signal_321, new_AGEMA_signal_320, new_AGEMA_signal_319, M22}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_333, new_AGEMA_signal_332, new_AGEMA_signal_331, M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M36_U1 ( .a ({new_AGEMA_signal_336, new_AGEMA_signal_335, new_AGEMA_signal_334, M24}), .b ({new_AGEMA_signal_327, new_AGEMA_signal_326, new_AGEMA_signal_325, M25}), .c ({new_AGEMA_signal_363, new_AGEMA_signal_362, new_AGEMA_signal_361, M36}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M29_U1 ( .a ({new_AGEMA_signal_342, new_AGEMA_signal_341, new_AGEMA_signal_340, M28}), .b ({new_AGEMA_signal_330, new_AGEMA_signal_329, new_AGEMA_signal_328, M27}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_351, new_AGEMA_signal_350, new_AGEMA_signal_349, M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M30_U1 ( .a ({new_AGEMA_signal_339, new_AGEMA_signal_338, new_AGEMA_signal_337, M26}), .b ({new_AGEMA_signal_336, new_AGEMA_signal_335, new_AGEMA_signal_334, M24}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_354, new_AGEMA_signal_353, new_AGEMA_signal_352, M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M32_U1 ( .a ({new_AGEMA_signal_330, new_AGEMA_signal_329, new_AGEMA_signal_328, M27}), .b ({new_AGEMA_signal_345, new_AGEMA_signal_344, new_AGEMA_signal_343, M31}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_357, new_AGEMA_signal_356, new_AGEMA_signal_355, M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M35_U1 ( .a ({new_AGEMA_signal_336, new_AGEMA_signal_335, new_AGEMA_signal_334, M24}), .b ({new_AGEMA_signal_333, new_AGEMA_signal_332, new_AGEMA_signal_331, M34}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_360, new_AGEMA_signal_359, new_AGEMA_signal_358, M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M37_U1 ( .a ({new_AGEMA_signal_318, new_AGEMA_signal_317, new_AGEMA_signal_316, M21}), .b ({new_AGEMA_signal_351, new_AGEMA_signal_350, new_AGEMA_signal_349, M29}), .c ({new_AGEMA_signal_366, new_AGEMA_signal_365, new_AGEMA_signal_364, M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M38_U1 ( .a ({new_AGEMA_signal_357, new_AGEMA_signal_356, new_AGEMA_signal_355, M32}), .b ({new_AGEMA_signal_348, new_AGEMA_signal_347, new_AGEMA_signal_346, M33}), .c ({new_AGEMA_signal_369, new_AGEMA_signal_368, new_AGEMA_signal_367, M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M39_U1 ( .a ({new_AGEMA_signal_324, new_AGEMA_signal_323, new_AGEMA_signal_322, M23}), .b ({new_AGEMA_signal_354, new_AGEMA_signal_353, new_AGEMA_signal_352, M30}), .c ({new_AGEMA_signal_372, new_AGEMA_signal_371, new_AGEMA_signal_370, M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M40_U1 ( .a ({new_AGEMA_signal_360, new_AGEMA_signal_359, new_AGEMA_signal_358, M35}), .b ({new_AGEMA_signal_363, new_AGEMA_signal_362, new_AGEMA_signal_361, M36}), .c ({new_AGEMA_signal_375, new_AGEMA_signal_374, new_AGEMA_signal_373, M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M41_U1 ( .a ({new_AGEMA_signal_369, new_AGEMA_signal_368, new_AGEMA_signal_367, M38}), .b ({new_AGEMA_signal_375, new_AGEMA_signal_374, new_AGEMA_signal_373, M40}), .c ({new_AGEMA_signal_378, new_AGEMA_signal_377, new_AGEMA_signal_376, M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M42_U1 ( .a ({new_AGEMA_signal_366, new_AGEMA_signal_365, new_AGEMA_signal_364, M37}), .b ({new_AGEMA_signal_372, new_AGEMA_signal_371, new_AGEMA_signal_370, M39}), .c ({new_AGEMA_signal_381, new_AGEMA_signal_380, new_AGEMA_signal_379, M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M43_U1 ( .a ({new_AGEMA_signal_366, new_AGEMA_signal_365, new_AGEMA_signal_364, M37}), .b ({new_AGEMA_signal_369, new_AGEMA_signal_368, new_AGEMA_signal_367, M38}), .c ({new_AGEMA_signal_384, new_AGEMA_signal_383, new_AGEMA_signal_382, M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M44_U1 ( .a ({new_AGEMA_signal_372, new_AGEMA_signal_371, new_AGEMA_signal_370, M39}), .b ({new_AGEMA_signal_375, new_AGEMA_signal_374, new_AGEMA_signal_373, M40}), .c ({new_AGEMA_signal_387, new_AGEMA_signal_386, new_AGEMA_signal_385, M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_M45_U1 ( .a ({new_AGEMA_signal_381, new_AGEMA_signal_380, new_AGEMA_signal_379, M42}), .b ({new_AGEMA_signal_378, new_AGEMA_signal_377, new_AGEMA_signal_376, M41}), .c ({new_AGEMA_signal_414, new_AGEMA_signal_413, new_AGEMA_signal_412, M45}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M46_U1 ( .a ({new_AGEMA_signal_387, new_AGEMA_signal_386, new_AGEMA_signal_385, M44}), .b ({new_AGEMA_signal_207, new_AGEMA_signal_206, new_AGEMA_signal_205, T6}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_417, new_AGEMA_signal_416, new_AGEMA_signal_415, M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M47_U1 ( .a ({new_AGEMA_signal_375, new_AGEMA_signal_374, new_AGEMA_signal_373, M40}), .b ({new_AGEMA_signal_231, new_AGEMA_signal_230, new_AGEMA_signal_229, T8}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_390, new_AGEMA_signal_389, new_AGEMA_signal_388, M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M48_U1 ( .a ({new_AGEMA_signal_372, new_AGEMA_signal_371, new_AGEMA_signal_370, M39}), .b ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_393, new_AGEMA_signal_392, new_AGEMA_signal_391, M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M49_U1 ( .a ({new_AGEMA_signal_384, new_AGEMA_signal_383, new_AGEMA_signal_382, M43}), .b ({new_AGEMA_signal_219, new_AGEMA_signal_218, new_AGEMA_signal_217, T16}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_420, new_AGEMA_signal_419, new_AGEMA_signal_418, M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M50_U1 ( .a ({new_AGEMA_signal_369, new_AGEMA_signal_368, new_AGEMA_signal_367, M38}), .b ({new_AGEMA_signal_210, new_AGEMA_signal_209, new_AGEMA_signal_208, T9}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_396, new_AGEMA_signal_395, new_AGEMA_signal_394, M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M51_U1 ( .a ({new_AGEMA_signal_366, new_AGEMA_signal_365, new_AGEMA_signal_364, M37}), .b ({new_AGEMA_signal_240, new_AGEMA_signal_239, new_AGEMA_signal_238, T17}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_399, new_AGEMA_signal_398, new_AGEMA_signal_397, M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M52_U1 ( .a ({new_AGEMA_signal_381, new_AGEMA_signal_380, new_AGEMA_signal_379, M42}), .b ({new_AGEMA_signal_216, new_AGEMA_signal_215, new_AGEMA_signal_214, T15}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_423, new_AGEMA_signal_422, new_AGEMA_signal_421, M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M53_U1 ( .a ({new_AGEMA_signal_414, new_AGEMA_signal_413, new_AGEMA_signal_412, M45}), .b ({new_AGEMA_signal_228, new_AGEMA_signal_227, new_AGEMA_signal_226, T27}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_450, new_AGEMA_signal_449, new_AGEMA_signal_448, M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M54_U1 ( .a ({new_AGEMA_signal_378, new_AGEMA_signal_377, new_AGEMA_signal_376, M41}), .b ({new_AGEMA_signal_234, new_AGEMA_signal_233, new_AGEMA_signal_232, T10}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_426, new_AGEMA_signal_425, new_AGEMA_signal_424, M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M55_U1 ( .a ({new_AGEMA_signal_387, new_AGEMA_signal_386, new_AGEMA_signal_385, M44}), .b ({new_AGEMA_signal_213, new_AGEMA_signal_212, new_AGEMA_signal_211, T13}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_429, new_AGEMA_signal_428, new_AGEMA_signal_427, M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M56_U1 ( .a ({new_AGEMA_signal_375, new_AGEMA_signal_374, new_AGEMA_signal_373, M40}), .b ({new_AGEMA_signal_246, new_AGEMA_signal_245, new_AGEMA_signal_244, T23}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_402, new_AGEMA_signal_401, new_AGEMA_signal_400, M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M57_U1 ( .a ({new_AGEMA_signal_372, new_AGEMA_signal_371, new_AGEMA_signal_370, M39}), .b ({new_AGEMA_signal_222, new_AGEMA_signal_221, new_AGEMA_signal_220, T19}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_405, new_AGEMA_signal_404, new_AGEMA_signal_403, M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M58_U1 ( .a ({new_AGEMA_signal_384, new_AGEMA_signal_383, new_AGEMA_signal_382, M43}), .b ({new_AGEMA_signal_171, new_AGEMA_signal_170, new_AGEMA_signal_169, T3}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_432, new_AGEMA_signal_431, new_AGEMA_signal_430, M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M59_U1 ( .a ({new_AGEMA_signal_369, new_AGEMA_signal_368, new_AGEMA_signal_367, M38}), .b ({new_AGEMA_signal_225, new_AGEMA_signal_224, new_AGEMA_signal_223, T22}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_408, new_AGEMA_signal_407, new_AGEMA_signal_406, M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M60_U1 ( .a ({new_AGEMA_signal_366, new_AGEMA_signal_365, new_AGEMA_signal_364, M37}), .b ({new_AGEMA_signal_243, new_AGEMA_signal_242, new_AGEMA_signal_241, T20}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_411, new_AGEMA_signal_410, new_AGEMA_signal_409, M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M61_U1 ( .a ({new_AGEMA_signal_381, new_AGEMA_signal_380, new_AGEMA_signal_379, M42}), .b ({new_AGEMA_signal_159, new_AGEMA_signal_158, new_AGEMA_signal_157, T1}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_435, new_AGEMA_signal_434, new_AGEMA_signal_433, M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M62_U1 ( .a ({new_AGEMA_signal_414, new_AGEMA_signal_413, new_AGEMA_signal_412, M45}), .b ({new_AGEMA_signal_174, new_AGEMA_signal_173, new_AGEMA_signal_172, T4}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_453, new_AGEMA_signal_452, new_AGEMA_signal_451, M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AND_M63_U1 ( .a ({new_AGEMA_signal_378, new_AGEMA_signal_377, new_AGEMA_signal_376, M41}), .b ({new_AGEMA_signal_165, new_AGEMA_signal_164, new_AGEMA_signal_163, T2}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_438, new_AGEMA_signal_437, new_AGEMA_signal_436, M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L0_U1 ( .a ({new_AGEMA_signal_435, new_AGEMA_signal_434, new_AGEMA_signal_433, M61}), .b ({new_AGEMA_signal_453, new_AGEMA_signal_452, new_AGEMA_signal_451, M62}), .c ({new_AGEMA_signal_480, new_AGEMA_signal_479, new_AGEMA_signal_478, L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L1_U1 ( .a ({new_AGEMA_signal_396, new_AGEMA_signal_395, new_AGEMA_signal_394, M50}), .b ({new_AGEMA_signal_402, new_AGEMA_signal_401, new_AGEMA_signal_400, M56}), .c ({new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L2_U1 ( .a ({new_AGEMA_signal_417, new_AGEMA_signal_416, new_AGEMA_signal_415, M46}), .b ({new_AGEMA_signal_393, new_AGEMA_signal_392, new_AGEMA_signal_391, M48}), .c ({new_AGEMA_signal_456, new_AGEMA_signal_455, new_AGEMA_signal_454, L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L3_U1 ( .a ({new_AGEMA_signal_390, new_AGEMA_signal_389, new_AGEMA_signal_388, M47}), .b ({new_AGEMA_signal_429, new_AGEMA_signal_428, new_AGEMA_signal_427, M55}), .c ({new_AGEMA_signal_459, new_AGEMA_signal_458, new_AGEMA_signal_457, L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L4_U1 ( .a ({new_AGEMA_signal_426, new_AGEMA_signal_425, new_AGEMA_signal_424, M54}), .b ({new_AGEMA_signal_432, new_AGEMA_signal_431, new_AGEMA_signal_430, M58}), .c ({new_AGEMA_signal_462, new_AGEMA_signal_461, new_AGEMA_signal_460, L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L5_U1 ( .a ({new_AGEMA_signal_420, new_AGEMA_signal_419, new_AGEMA_signal_418, M49}), .b ({new_AGEMA_signal_435, new_AGEMA_signal_434, new_AGEMA_signal_433, M61}), .c ({new_AGEMA_signal_465, new_AGEMA_signal_464, new_AGEMA_signal_463, L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L6_U1 ( .a ({new_AGEMA_signal_453, new_AGEMA_signal_452, new_AGEMA_signal_451, M62}), .b ({new_AGEMA_signal_465, new_AGEMA_signal_464, new_AGEMA_signal_463, L5}), .c ({new_AGEMA_signal_483, new_AGEMA_signal_482, new_AGEMA_signal_481, L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L7_U1 ( .a ({new_AGEMA_signal_417, new_AGEMA_signal_416, new_AGEMA_signal_415, M46}), .b ({new_AGEMA_signal_459, new_AGEMA_signal_458, new_AGEMA_signal_457, L3}), .c ({new_AGEMA_signal_486, new_AGEMA_signal_485, new_AGEMA_signal_484, L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L8_U1 ( .a ({new_AGEMA_signal_399, new_AGEMA_signal_398, new_AGEMA_signal_397, M51}), .b ({new_AGEMA_signal_408, new_AGEMA_signal_407, new_AGEMA_signal_406, M59}), .c ({new_AGEMA_signal_444, new_AGEMA_signal_443, new_AGEMA_signal_442, L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L9_U1 ( .a ({new_AGEMA_signal_423, new_AGEMA_signal_422, new_AGEMA_signal_421, M52}), .b ({new_AGEMA_signal_450, new_AGEMA_signal_449, new_AGEMA_signal_448, M53}), .c ({new_AGEMA_signal_489, new_AGEMA_signal_488, new_AGEMA_signal_487, L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L10_U1 ( .a ({new_AGEMA_signal_450, new_AGEMA_signal_449, new_AGEMA_signal_448, M53}), .b ({new_AGEMA_signal_462, new_AGEMA_signal_461, new_AGEMA_signal_460, L4}), .c ({new_AGEMA_signal_492, new_AGEMA_signal_491, new_AGEMA_signal_490, L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L11_U1 ( .a ({new_AGEMA_signal_411, new_AGEMA_signal_410, new_AGEMA_signal_409, M60}), .b ({new_AGEMA_signal_456, new_AGEMA_signal_455, new_AGEMA_signal_454, L2}), .c ({new_AGEMA_signal_495, new_AGEMA_signal_494, new_AGEMA_signal_493, L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L12_U1 ( .a ({new_AGEMA_signal_393, new_AGEMA_signal_392, new_AGEMA_signal_391, M48}), .b ({new_AGEMA_signal_399, new_AGEMA_signal_398, new_AGEMA_signal_397, M51}), .c ({new_AGEMA_signal_447, new_AGEMA_signal_446, new_AGEMA_signal_445, L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L13_U1 ( .a ({new_AGEMA_signal_396, new_AGEMA_signal_395, new_AGEMA_signal_394, M50}), .b ({new_AGEMA_signal_480, new_AGEMA_signal_479, new_AGEMA_signal_478, L0}), .c ({new_AGEMA_signal_507, new_AGEMA_signal_506, new_AGEMA_signal_505, L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L14_U1 ( .a ({new_AGEMA_signal_423, new_AGEMA_signal_422, new_AGEMA_signal_421, M52}), .b ({new_AGEMA_signal_435, new_AGEMA_signal_434, new_AGEMA_signal_433, M61}), .c ({new_AGEMA_signal_468, new_AGEMA_signal_467, new_AGEMA_signal_466, L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L15_U1 ( .a ({new_AGEMA_signal_429, new_AGEMA_signal_428, new_AGEMA_signal_427, M55}), .b ({new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, L1}), .c ({new_AGEMA_signal_471, new_AGEMA_signal_470, new_AGEMA_signal_469, L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L16_U1 ( .a ({new_AGEMA_signal_402, new_AGEMA_signal_401, new_AGEMA_signal_400, M56}), .b ({new_AGEMA_signal_480, new_AGEMA_signal_479, new_AGEMA_signal_478, L0}), .c ({new_AGEMA_signal_510, new_AGEMA_signal_509, new_AGEMA_signal_508, L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L17_U1 ( .a ({new_AGEMA_signal_405, new_AGEMA_signal_404, new_AGEMA_signal_403, M57}), .b ({new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, L1}), .c ({new_AGEMA_signal_474, new_AGEMA_signal_473, new_AGEMA_signal_472, L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L18_U1 ( .a ({new_AGEMA_signal_432, new_AGEMA_signal_431, new_AGEMA_signal_430, M58}), .b ({new_AGEMA_signal_444, new_AGEMA_signal_443, new_AGEMA_signal_442, L8}), .c ({new_AGEMA_signal_477, new_AGEMA_signal_476, new_AGEMA_signal_475, L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L19_U1 ( .a ({new_AGEMA_signal_438, new_AGEMA_signal_437, new_AGEMA_signal_436, M63}), .b ({new_AGEMA_signal_462, new_AGEMA_signal_461, new_AGEMA_signal_460, L4}), .c ({new_AGEMA_signal_498, new_AGEMA_signal_497, new_AGEMA_signal_496, L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L20_U1 ( .a ({new_AGEMA_signal_480, new_AGEMA_signal_479, new_AGEMA_signal_478, L0}), .b ({new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, L1}), .c ({new_AGEMA_signal_513, new_AGEMA_signal_512, new_AGEMA_signal_511, L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L21_U1 ( .a ({new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, L1}), .b ({new_AGEMA_signal_486, new_AGEMA_signal_485, new_AGEMA_signal_484, L7}), .c ({new_AGEMA_signal_516, new_AGEMA_signal_515, new_AGEMA_signal_514, L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L22_U1 ( .a ({new_AGEMA_signal_459, new_AGEMA_signal_458, new_AGEMA_signal_457, L3}), .b ({new_AGEMA_signal_447, new_AGEMA_signal_446, new_AGEMA_signal_445, L12}), .c ({new_AGEMA_signal_501, new_AGEMA_signal_500, new_AGEMA_signal_499, L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L23_U1 ( .a ({new_AGEMA_signal_477, new_AGEMA_signal_476, new_AGEMA_signal_475, L18}), .b ({new_AGEMA_signal_456, new_AGEMA_signal_455, new_AGEMA_signal_454, L2}), .c ({new_AGEMA_signal_504, new_AGEMA_signal_503, new_AGEMA_signal_502, L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L24_U1 ( .a ({new_AGEMA_signal_471, new_AGEMA_signal_470, new_AGEMA_signal_469, L15}), .b ({new_AGEMA_signal_489, new_AGEMA_signal_488, new_AGEMA_signal_487, L9}), .c ({new_AGEMA_signal_519, new_AGEMA_signal_518, new_AGEMA_signal_517, L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L25_U1 ( .a ({new_AGEMA_signal_483, new_AGEMA_signal_482, new_AGEMA_signal_481, L6}), .b ({new_AGEMA_signal_492, new_AGEMA_signal_491, new_AGEMA_signal_490, L10}), .c ({new_AGEMA_signal_522, new_AGEMA_signal_521, new_AGEMA_signal_520, L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L26_U1 ( .a ({new_AGEMA_signal_486, new_AGEMA_signal_485, new_AGEMA_signal_484, L7}), .b ({new_AGEMA_signal_489, new_AGEMA_signal_488, new_AGEMA_signal_487, L9}), .c ({new_AGEMA_signal_525, new_AGEMA_signal_524, new_AGEMA_signal_523, L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L27_U1 ( .a ({new_AGEMA_signal_444, new_AGEMA_signal_443, new_AGEMA_signal_442, L8}), .b ({new_AGEMA_signal_492, new_AGEMA_signal_491, new_AGEMA_signal_490, L10}), .c ({new_AGEMA_signal_528, new_AGEMA_signal_527, new_AGEMA_signal_526, L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L28_U1 ( .a ({new_AGEMA_signal_495, new_AGEMA_signal_494, new_AGEMA_signal_493, L11}), .b ({new_AGEMA_signal_468, new_AGEMA_signal_467, new_AGEMA_signal_466, L14}), .c ({new_AGEMA_signal_531, new_AGEMA_signal_530, new_AGEMA_signal_529, L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_L29_U1 ( .a ({new_AGEMA_signal_495, new_AGEMA_signal_494, new_AGEMA_signal_493, L11}), .b ({new_AGEMA_signal_474, new_AGEMA_signal_473, new_AGEMA_signal_472, L17}), .c ({new_AGEMA_signal_534, new_AGEMA_signal_533, new_AGEMA_signal_532, L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_S0_U1 ( .a ({new_AGEMA_signal_483, new_AGEMA_signal_482, new_AGEMA_signal_481, L6}), .b ({new_AGEMA_signal_519, new_AGEMA_signal_518, new_AGEMA_signal_517, L24}), .c ({new_AGEMA_signal_540, new_AGEMA_signal_539, new_AGEMA_signal_538, O[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) XOR_S1_U1 ( .a ({new_AGEMA_signal_510, new_AGEMA_signal_509, new_AGEMA_signal_508, L16}), .b ({new_AGEMA_signal_525, new_AGEMA_signal_524, new_AGEMA_signal_523, L26}), .c ({new_AGEMA_signal_543, new_AGEMA_signal_542, new_AGEMA_signal_541, O[6]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) XOR_S2_U1 ( .a ({new_AGEMA_signal_498, new_AGEMA_signal_497, new_AGEMA_signal_496, L19}), .b ({new_AGEMA_signal_531, new_AGEMA_signal_530, new_AGEMA_signal_529, L28}), .c ({new_AGEMA_signal_546, new_AGEMA_signal_545, new_AGEMA_signal_544, O[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_S3_U1 ( .a ({new_AGEMA_signal_483, new_AGEMA_signal_482, new_AGEMA_signal_481, L6}), .b ({new_AGEMA_signal_516, new_AGEMA_signal_515, new_AGEMA_signal_514, L21}), .c ({new_AGEMA_signal_549, new_AGEMA_signal_548, new_AGEMA_signal_547, O[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_S4_U1 ( .a ({new_AGEMA_signal_513, new_AGEMA_signal_512, new_AGEMA_signal_511, L20}), .b ({new_AGEMA_signal_501, new_AGEMA_signal_500, new_AGEMA_signal_499, L22}), .c ({new_AGEMA_signal_552, new_AGEMA_signal_551, new_AGEMA_signal_550, O[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) XOR_S5_U1 ( .a ({new_AGEMA_signal_522, new_AGEMA_signal_521, new_AGEMA_signal_520, L25}), .b ({new_AGEMA_signal_534, new_AGEMA_signal_533, new_AGEMA_signal_532, L29}), .c ({new_AGEMA_signal_555, new_AGEMA_signal_554, new_AGEMA_signal_553, O[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) XOR_S6_U1 ( .a ({new_AGEMA_signal_507, new_AGEMA_signal_506, new_AGEMA_signal_505, L13}), .b ({new_AGEMA_signal_528, new_AGEMA_signal_527, new_AGEMA_signal_526, L27}), .c ({new_AGEMA_signal_558, new_AGEMA_signal_557, new_AGEMA_signal_556, O[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) XOR_S7_U1 ( .a ({new_AGEMA_signal_483, new_AGEMA_signal_482, new_AGEMA_signal_481, L6}), .b ({new_AGEMA_signal_504, new_AGEMA_signal_503, new_AGEMA_signal_502, L23}), .c ({new_AGEMA_signal_537, new_AGEMA_signal_536, new_AGEMA_signal_535, O[0]}) ) ;

    /* register cells */
    assign {Y_s3[7], Y_s2[7], Y_s1[7], Y_s0[7]} = {new_AGEMA_signal_540, new_AGEMA_signal_539, new_AGEMA_signal_538, O[7]};
    assign {Y_s3[6], Y_s2[6], Y_s1[6], Y_s0[6]} = {new_AGEMA_signal_543, new_AGEMA_signal_542, new_AGEMA_signal_541, O[6]};
    assign {Y_s3[5], Y_s2[5], Y_s1[5], Y_s0[5]} = {new_AGEMA_signal_546, new_AGEMA_signal_545, new_AGEMA_signal_544, O[5]};
    assign {Y_s3[4], Y_s2[4], Y_s1[4], Y_s0[4]} = {new_AGEMA_signal_549, new_AGEMA_signal_548, new_AGEMA_signal_547, O[4]};
    assign {Y_s3[3], Y_s2[3], Y_s1[3], Y_s0[3]} = {new_AGEMA_signal_552, new_AGEMA_signal_551, new_AGEMA_signal_550, O[3]};
    assign {Y_s3[2], Y_s2[2], Y_s1[2], Y_s0[2]} = {new_AGEMA_signal_555, new_AGEMA_signal_554, new_AGEMA_signal_553, O[2]};
    assign {Y_s3[1], Y_s2[1], Y_s1[1], Y_s0[1]} = {new_AGEMA_signal_558, new_AGEMA_signal_557, new_AGEMA_signal_556, O[1]};
    assign {Y_s3[0], Y_s2[0], Y_s1[0], Y_s0[0]} = {new_AGEMA_signal_537, new_AGEMA_signal_536, new_AGEMA_signal_535, O[0]};
endmodule
