////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module PRESENT in file /AGEMA/Designs/PRESENT_nibble-serial/AGEMA/PRESENT.v */
/* clock gating is added to the circuit, the latency increased 4 time(s)  */

module PRESENT_HPC2_ClockGating_d3 (data_in_s0, key_s0, clk, reset, data_in_s1, data_in_s2, data_in_s3, key_s1, key_s2, key_s3, Fresh, data_out_s0, done, data_out_s1, data_out_s2, data_out_s3, Synch);
    input [63:0] data_in_s0 ;
    input [79:0] key_s0 ;
    input clk ;
    input reset ;
    input [63:0] data_in_s1 ;
    input [63:0] data_in_s2 ;
    input [63:0] data_in_s3 ;
    input [79:0] key_s1 ;
    input [79:0] key_s2 ;
    input [79:0] key_s3 ;
    input [23:0] Fresh ;
    output [63:0] data_out_s0 ;
    output done ;
    output [63:0] data_out_s1 ;
    output [63:0] data_out_s2 ;
    output [63:0] data_out_s3 ;
    output Synch ;
    wire selSbox ;
    wire ctrlData_0_ ;
    wire intDone ;
    wire fsm_n15 ;
    wire fsm_n14 ;
    wire fsm_n13 ;
    wire fsm_n12 ;
    wire fsm_n11 ;
    wire fsm_n10 ;
    wire fsm_n9 ;
    wire fsm_n8 ;
    wire fsm_n7 ;
    wire fsm_n6 ;
    wire fsm_n4 ;
    wire fsm_n2 ;
    wire fsm_n5 ;
    wire fsm_n20 ;
    wire fsm_ps_state_0_ ;
    wire fsm_ps_state_1_ ;
    wire fsm_n21 ;
    wire fsm_n3 ;
    wire fsm_rst_countSerial ;
    wire fsm_en_countRound ;
    wire fsm_cnt_rnd_n33 ;
    wire fsm_cnt_rnd_n32 ;
    wire fsm_cnt_rnd_n31 ;
    wire fsm_cnt_rnd_n30 ;
    wire fsm_cnt_rnd_n29 ;
    wire fsm_cnt_rnd_n28 ;
    wire fsm_cnt_rnd_n27 ;
    wire fsm_cnt_rnd_n26 ;
    wire fsm_cnt_rnd_n23 ;
    wire fsm_cnt_rnd_n22 ;
    wire fsm_cnt_rnd_n21 ;
    wire fsm_cnt_rnd_n20 ;
    wire fsm_cnt_rnd_n19 ;
    wire fsm_cnt_rnd_n17 ;
    wire fsm_cnt_rnd_n15 ;
    wire fsm_cnt_rnd_n13 ;
    wire fsm_cnt_rnd_n12 ;
    wire fsm_cnt_rnd_n11 ;
    wire fsm_cnt_rnd_n10 ;
    wire fsm_cnt_rnd_n9 ;
    wire fsm_cnt_rnd_n8 ;
    wire fsm_cnt_rnd_n7 ;
    wire fsm_cnt_rnd_n6 ;
    wire fsm_cnt_rnd_n5 ;
    wire fsm_cnt_rnd_n3 ;
    wire fsm_cnt_rnd_n24 ;
    wire fsm_cnt_rnd_n41 ;
    wire fsm_cnt_rnd_n25 ;
    wire fsm_cnt_rnd_n1 ;
    wire fsm_cnt_rnd_n18 ;
    wire fsm_cnt_rnd_n16 ;
    wire fsm_cnt_rnd_n14 ;
    wire fsm_cnt_ser_n10 ;
    wire fsm_cnt_ser_n9 ;
    wire fsm_cnt_ser_n8 ;
    wire fsm_cnt_ser_n7 ;
    wire fsm_cnt_ser_n6 ;
    wire fsm_cnt_ser_n5 ;
    wire fsm_cnt_ser_n4 ;
    wire fsm_cnt_ser_n2 ;
    wire fsm_cnt_ser_n20 ;
    wire fsm_cnt_ser_n28 ;
    wire fsm_cnt_ser_n26 ;
    wire fsm_cnt_ser_n3 ;
    wire fsm_cnt_ser_n1 ;
    wire stateFF_state_n7 ;
    wire stateFF_state_n6 ;
    wire stateFF_state_n5 ;
    wire keyFF_keystate_n8 ;
    wire keyFF_keystate_n7 ;
    wire keyFF_keystate_n6 ;
    wire sboxInst_n3 ;
    wire sboxInst_n2 ;
    wire sboxInst_n1 ;
    wire sboxInst_L8 ;
    wire sboxInst_L7 ;
    wire sboxInst_T3 ;
    wire sboxInst_T1 ;
    wire sboxInst_Q7 ;
    wire sboxInst_Q6 ;
    wire sboxInst_L5 ;
    wire sboxInst_T2 ;
    wire sboxInst_L4 ;
    wire sboxInst_Q3 ;
    wire sboxInst_L3 ;
    wire sboxInst_Q2 ;
    wire sboxInst_T0 ;
    wire sboxInst_L2 ;
    wire sboxInst_L1 ;
    wire sboxInst_L0 ;
    wire [4:0] counter ;
    wire [3:0] serialIn ;
    wire [3:0] sboxOut ;
    wire [3:0] roundkey ;
    wire [3:1] keyRegKS ;
    wire [3:0] sboxIn ;
    wire [3:0] stateXORroundkey ;
    wire [3:0] fsm_countSerial ;
    wire [63:0] stateFF_inputPar ;
    wire [3:0] stateFF_state_gff_1_s_next_state ;
    wire [3:0] stateFF_state_gff_2_s_next_state ;
    wire [3:0] stateFF_state_gff_3_s_next_state ;
    wire [3:0] stateFF_state_gff_4_s_next_state ;
    wire [3:0] stateFF_state_gff_5_s_next_state ;
    wire [3:0] stateFF_state_gff_6_s_next_state ;
    wire [3:0] stateFF_state_gff_7_s_next_state ;
    wire [3:0] stateFF_state_gff_8_s_next_state ;
    wire [3:0] stateFF_state_gff_9_s_next_state ;
    wire [3:0] stateFF_state_gff_10_s_next_state ;
    wire [3:0] stateFF_state_gff_11_s_next_state ;
    wire [3:0] stateFF_state_gff_12_s_next_state ;
    wire [3:0] stateFF_state_gff_13_s_next_state ;
    wire [3:0] stateFF_state_gff_14_s_next_state ;
    wire [3:0] stateFF_state_gff_15_s_next_state ;
    wire [3:0] stateFF_state_gff_16_s_next_state ;
    wire [4:0] keyFF_counterAdd ;
    wire [75:3] keyFF_outputPar ;
    wire [79:0] keyFF_inputPar ;
    wire [3:0] keyFF_keystate_gff_1_s_next_state ;
    wire [3:0] keyFF_keystate_gff_2_s_next_state ;
    wire [3:0] keyFF_keystate_gff_3_s_next_state ;
    wire [3:0] keyFF_keystate_gff_4_s_next_state ;
    wire [3:0] keyFF_keystate_gff_5_s_next_state ;
    wire [3:0] keyFF_keystate_gff_6_s_next_state ;
    wire [3:0] keyFF_keystate_gff_7_s_next_state ;
    wire [3:0] keyFF_keystate_gff_8_s_next_state ;
    wire [3:0] keyFF_keystate_gff_9_s_next_state ;
    wire [3:0] keyFF_keystate_gff_10_s_next_state ;
    wire [3:0] keyFF_keystate_gff_11_s_next_state ;
    wire [3:0] keyFF_keystate_gff_12_s_next_state ;
    wire [3:0] keyFF_keystate_gff_13_s_next_state ;
    wire [3:0] keyFF_keystate_gff_14_s_next_state ;
    wire [3:0] keyFF_keystate_gff_15_s_next_state ;
    wire [3:0] keyFF_keystate_gff_16_s_next_state ;
    wire [3:0] keyFF_keystate_gff_17_s_next_state ;
    wire [3:0] keyFF_keystate_gff_18_s_next_state ;
    wire [3:0] keyFF_keystate_gff_19_s_next_state ;
    wire [3:0] keyFF_keystate_gff_20_s_next_state ;
    wire new_AGEMA_signal_856 ;
    wire new_AGEMA_signal_857 ;
    wire new_AGEMA_signal_858 ;
    wire new_AGEMA_signal_862 ;
    wire new_AGEMA_signal_863 ;
    wire new_AGEMA_signal_864 ;
    wire new_AGEMA_signal_865 ;
    wire new_AGEMA_signal_866 ;
    wire new_AGEMA_signal_867 ;
    wire new_AGEMA_signal_871 ;
    wire new_AGEMA_signal_872 ;
    wire new_AGEMA_signal_873 ;
    wire new_AGEMA_signal_874 ;
    wire new_AGEMA_signal_875 ;
    wire new_AGEMA_signal_876 ;
    wire new_AGEMA_signal_880 ;
    wire new_AGEMA_signal_881 ;
    wire new_AGEMA_signal_882 ;
    wire new_AGEMA_signal_883 ;
    wire new_AGEMA_signal_884 ;
    wire new_AGEMA_signal_885 ;
    wire new_AGEMA_signal_889 ;
    wire new_AGEMA_signal_890 ;
    wire new_AGEMA_signal_891 ;
    wire new_AGEMA_signal_898 ;
    wire new_AGEMA_signal_899 ;
    wire new_AGEMA_signal_900 ;
    wire new_AGEMA_signal_907 ;
    wire new_AGEMA_signal_908 ;
    wire new_AGEMA_signal_909 ;
    wire new_AGEMA_signal_916 ;
    wire new_AGEMA_signal_917 ;
    wire new_AGEMA_signal_918 ;
    wire new_AGEMA_signal_925 ;
    wire new_AGEMA_signal_926 ;
    wire new_AGEMA_signal_927 ;
    wire new_AGEMA_signal_934 ;
    wire new_AGEMA_signal_935 ;
    wire new_AGEMA_signal_936 ;
    wire new_AGEMA_signal_943 ;
    wire new_AGEMA_signal_944 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_952 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_954 ;
    wire new_AGEMA_signal_961 ;
    wire new_AGEMA_signal_962 ;
    wire new_AGEMA_signal_963 ;
    wire new_AGEMA_signal_970 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_972 ;
    wire new_AGEMA_signal_979 ;
    wire new_AGEMA_signal_980 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_990 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1007 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1015 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(3), .pipeline(0)) U9 ( .a ({new_AGEMA_signal_858, new_AGEMA_signal_857, new_AGEMA_signal_856, roundkey[0]}), .b ({data_out_s3[60], data_out_s2[60], data_out_s1[60], data_out_s0[60]}), .c ({new_AGEMA_signal_864, new_AGEMA_signal_863, new_AGEMA_signal_862, stateXORroundkey[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U10 ( .a ({new_AGEMA_signal_867, new_AGEMA_signal_866, new_AGEMA_signal_865, roundkey[1]}), .b ({data_out_s3[61], data_out_s2[61], data_out_s1[61], data_out_s0[61]}), .c ({new_AGEMA_signal_873, new_AGEMA_signal_872, new_AGEMA_signal_871, stateXORroundkey[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U11 ( .a ({new_AGEMA_signal_876, new_AGEMA_signal_875, new_AGEMA_signal_874, roundkey[2]}), .b ({data_out_s3[62], data_out_s2[62], data_out_s1[62], data_out_s0[62]}), .c ({new_AGEMA_signal_882, new_AGEMA_signal_881, new_AGEMA_signal_880, stateXORroundkey[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U12 ( .a ({new_AGEMA_signal_885, new_AGEMA_signal_884, new_AGEMA_signal_883, roundkey[3]}), .b ({data_out_s3[63], data_out_s2[63], data_out_s1[63], data_out_s0[63]}), .c ({new_AGEMA_signal_891, new_AGEMA_signal_890, new_AGEMA_signal_889, stateXORroundkey[3]}) ) ;
    NOR2_X1 fsm_U20 ( .A1 (reset), .A2 (fsm_n15), .ZN (fsm_n21) ) ;
    NOR2_X1 fsm_U19 ( .A1 (fsm_n14), .A2 (done), .ZN (fsm_n15) ) ;
    NOR2_X1 fsm_U18 ( .A1 (reset), .A2 (fsm_n13), .ZN (fsm_n20) ) ;
    NOR2_X1 fsm_U17 ( .A1 (fsm_ps_state_1_), .A2 (fsm_n12), .ZN (fsm_n13) ) ;
    NOR2_X1 fsm_U16 ( .A1 (fsm_n11), .A2 (fsm_n10), .ZN (fsm_n12) ) ;
    NAND2_X1 fsm_U15 ( .A1 (counter[3]), .A2 (counter[1]), .ZN (fsm_n10) ) ;
    OR2_X1 fsm_U14 ( .A1 (fsm_n9), .A2 (fsm_n8), .ZN (fsm_n11) ) ;
    NAND2_X1 fsm_U13 ( .A1 (counter[0]), .A2 (counter[4]), .ZN (fsm_n8) ) ;
    NAND2_X1 fsm_U12 ( .A1 (counter[2]), .A2 (fsm_ps_state_0_), .ZN (fsm_n9) ) ;
    NOR2_X1 fsm_U11 ( .A1 (fsm_n3), .A2 (fsm_n5), .ZN (done) ) ;
    AND2_X1 fsm_U10 ( .A1 (fsm_n14), .A2 (fsm_n5), .ZN (fsm_en_countRound) ) ;
    AND2_X1 fsm_U9 ( .A1 (fsm_countSerial[2]), .A2 (fsm_n7), .ZN (fsm_n14) ) ;
    NOR2_X1 fsm_U8 ( .A1 (fsm_n6), .A2 (fsm_n4), .ZN (fsm_n7) ) ;
    NAND2_X1 fsm_U7 ( .A1 (fsm_countSerial[1]), .A2 (fsm_countSerial[0]), .ZN (fsm_n4) ) ;
    NAND2_X1 fsm_U6 ( .A1 (fsm_n3), .A2 (fsm_countSerial[3]), .ZN (fsm_n6) ) ;
    NOR2_X1 fsm_U5 ( .A1 (fsm_ps_state_0_), .A2 (fsm_n5), .ZN (intDone) ) ;
    NOR2_X1 fsm_U4 ( .A1 (fsm_ps_state_1_), .A2 (fsm_n3), .ZN (selSbox) ) ;
    NOR2_X1 fsm_U3 ( .A1 (reset), .A2 (selSbox), .ZN (fsm_rst_countSerial) ) ;
    INV_X1 fsm_U2 ( .A (reset), .ZN (fsm_n2) ) ;
    INV_X1 fsm_U1 ( .A (fsm_rst_countSerial), .ZN (ctrlData_0_) ) ;
    NAND2_X1 fsm_cnt_rnd_U28 ( .A1 (fsm_cnt_rnd_n33), .A2 (fsm_cnt_rnd_n32), .ZN (fsm_cnt_rnd_n41) ) ;
    NAND2_X1 fsm_cnt_rnd_U27 ( .A1 (fsm_cnt_rnd_n31), .A2 (counter[1]), .ZN (fsm_cnt_rnd_n32) ) ;
    NAND2_X1 fsm_cnt_rnd_U26 ( .A1 (fsm_cnt_rnd_n30), .A2 (fsm_cnt_rnd_n24), .ZN (fsm_cnt_rnd_n33) ) ;
    NAND2_X1 fsm_cnt_rnd_U25 ( .A1 (fsm_cnt_rnd_n29), .A2 (counter[0]), .ZN (fsm_cnt_rnd_n30) ) ;
    NAND2_X1 fsm_cnt_rnd_U24 ( .A1 (fsm_cnt_rnd_n28), .A2 (fsm_cnt_rnd_n27), .ZN (fsm_cnt_rnd_n18) ) ;
    NAND2_X1 fsm_cnt_rnd_U23 ( .A1 (fsm_cnt_rnd_n26), .A2 (counter[0]), .ZN (fsm_cnt_rnd_n27) ) ;
    MUX2_X1 fsm_cnt_rnd_U22 ( .S (fsm_cnt_rnd_n5), .A (fsm_cnt_rnd_n23), .B (fsm_cnt_rnd_n22), .Z (fsm_cnt_rnd_n16) ) ;
    NAND2_X1 fsm_cnt_rnd_U21 ( .A1 (fsm_cnt_rnd_n31), .A2 (fsm_cnt_rnd_n21), .ZN (fsm_cnt_rnd_n23) ) ;
    NAND2_X1 fsm_cnt_rnd_U20 ( .A1 (fsm_cnt_rnd_n29), .A2 (fsm_cnt_rnd_n24), .ZN (fsm_cnt_rnd_n21) ) ;
    NOR2_X1 fsm_cnt_rnd_U19 ( .A1 (fsm_cnt_rnd_n20), .A2 (fsm_cnt_rnd_n26), .ZN (fsm_cnt_rnd_n31) ) ;
    NOR2_X1 fsm_cnt_rnd_U18 ( .A1 (fsm_en_countRound), .A2 (fsm_cnt_rnd_n6), .ZN (fsm_cnt_rnd_n26) ) ;
    INV_X1 fsm_cnt_rnd_U17 ( .A (fsm_cnt_rnd_n28), .ZN (fsm_cnt_rnd_n20) ) ;
    NAND2_X1 fsm_cnt_rnd_U16 ( .A1 (fsm_cnt_rnd_n29), .A2 (fsm_cnt_rnd_n3), .ZN (fsm_cnt_rnd_n28) ) ;
    MUX2_X1 fsm_cnt_rnd_U15 ( .S (counter[4]), .A (fsm_cnt_rnd_n19), .B (fsm_cnt_rnd_n17), .Z (fsm_cnt_rnd_n14) ) ;
    NAND2_X1 fsm_cnt_rnd_U14 ( .A1 (fsm_cnt_rnd_n15), .A2 (fsm_cnt_rnd_n13), .ZN (fsm_cnt_rnd_n17) ) ;
    NAND2_X1 fsm_cnt_rnd_U13 ( .A1 (fsm_cnt_rnd_n29), .A2 (fsm_cnt_rnd_n25), .ZN (fsm_cnt_rnd_n15) ) ;
    INV_X1 fsm_cnt_rnd_U12 ( .A (fsm_cnt_rnd_n12), .ZN (fsm_cnt_rnd_n29) ) ;
    NOR2_X1 fsm_cnt_rnd_U11 ( .A1 (fsm_cnt_rnd_n25), .A2 (fsm_cnt_rnd_n11), .ZN (fsm_cnt_rnd_n19) ) ;
    INV_X1 fsm_cnt_rnd_U10 ( .A (fsm_cnt_rnd_n10), .ZN (fsm_cnt_rnd_n1) ) ;
    MUX2_X1 fsm_cnt_rnd_U9 ( .S (fsm_cnt_rnd_n25), .A (fsm_cnt_rnd_n13), .B (fsm_cnt_rnd_n11), .Z (fsm_cnt_rnd_n10) ) ;
    NAND2_X1 fsm_cnt_rnd_U8 ( .A1 (counter[2]), .A2 (fsm_cnt_rnd_n22), .ZN (fsm_cnt_rnd_n11) ) ;
    NOR2_X1 fsm_cnt_rnd_U7 ( .A1 (fsm_cnt_rnd_n12), .A2 (fsm_cnt_rnd_n9), .ZN (fsm_cnt_rnd_n22) ) ;
    NAND2_X1 fsm_cnt_rnd_U6 ( .A1 (fsm_en_countRound), .A2 (fsm_n2), .ZN (fsm_cnt_rnd_n12) ) ;
    NAND2_X1 fsm_cnt_rnd_U5 ( .A1 (fsm_n2), .A2 (fsm_cnt_rnd_n8), .ZN (fsm_cnt_rnd_n13) ) ;
    NAND2_X1 fsm_cnt_rnd_U4 ( .A1 (fsm_en_countRound), .A2 (fsm_cnt_rnd_n7), .ZN (fsm_cnt_rnd_n8) ) ;
    NOR2_X1 fsm_cnt_rnd_U3 ( .A1 (fsm_cnt_rnd_n5), .A2 (fsm_cnt_rnd_n9), .ZN (fsm_cnt_rnd_n7) ) ;
    OR2_X1 fsm_cnt_rnd_U2 ( .A1 (fsm_cnt_rnd_n24), .A2 (fsm_cnt_rnd_n3), .ZN (fsm_cnt_rnd_n9) ) ;
    INV_X1 fsm_cnt_rnd_U1 ( .A (fsm_n2), .ZN (fsm_cnt_rnd_n6) ) ;
    INV_X1 fsm_cnt_rnd_count_reg_reg_2__U1 ( .A (counter[2]), .ZN (fsm_cnt_rnd_n5) ) ;
    INV_X1 fsm_cnt_rnd_count_reg_reg_0__U1 ( .A (counter[0]), .ZN (fsm_cnt_rnd_n3) ) ;
    INV_X1 fsm_cnt_rnd_count_reg_reg_3__U1 ( .A (counter[3]), .ZN (fsm_cnt_rnd_n25) ) ;
    INV_X1 fsm_cnt_rnd_count_reg_reg_1__U1 ( .A (fsm_cnt_rnd_n24), .ZN (counter[1]) ) ;
    NOR2_X1 fsm_cnt_ser_U12 ( .A1 (fsm_cnt_ser_n10), .A2 (fsm_cnt_ser_n9), .ZN (fsm_cnt_ser_n3) ) ;
    XNOR2_X1 fsm_cnt_ser_U11 ( .A (fsm_n3), .B (fsm_countSerial[0]), .ZN (fsm_cnt_ser_n10) ) ;
    NOR2_X1 fsm_cnt_ser_U10 ( .A1 (fsm_cnt_ser_n9), .A2 (fsm_cnt_ser_n8), .ZN (fsm_cnt_ser_n28) ) ;
    XOR2_X1 fsm_cnt_ser_U9 ( .A (fsm_countSerial[1]), .B (fsm_cnt_ser_n7), .Z (fsm_cnt_ser_n8) ) ;
    NOR2_X1 fsm_cnt_ser_U8 ( .A1 (fsm_cnt_ser_n9), .A2 (fsm_cnt_ser_n6), .ZN (fsm_cnt_ser_n26) ) ;
    XOR2_X1 fsm_cnt_ser_U7 ( .A (fsm_countSerial[3]), .B (fsm_cnt_ser_n5), .Z (fsm_cnt_ser_n6) ) ;
    NAND2_X1 fsm_cnt_ser_U6 ( .A1 (fsm_cnt_ser_n4), .A2 (fsm_countSerial[2]), .ZN (fsm_cnt_ser_n5) ) ;
    NOR2_X1 fsm_cnt_ser_U5 ( .A1 (fsm_cnt_ser_n2), .A2 (fsm_cnt_ser_n9), .ZN (fsm_cnt_ser_n1) ) ;
    INV_X1 fsm_cnt_ser_U4 ( .A (fsm_rst_countSerial), .ZN (fsm_cnt_ser_n9) ) ;
    XNOR2_X1 fsm_cnt_ser_U3 ( .A (fsm_cnt_ser_n4), .B (fsm_countSerial[2]), .ZN (fsm_cnt_ser_n2) ) ;
    NOR2_X1 fsm_cnt_ser_U2 ( .A1 (fsm_cnt_ser_n20), .A2 (fsm_cnt_ser_n7), .ZN (fsm_cnt_ser_n4) ) ;
    NAND2_X1 fsm_cnt_ser_U1 ( .A1 (fsm_n3), .A2 (fsm_countSerial[0]), .ZN (fsm_cnt_ser_n7) ) ;
    INV_X1 fsm_cnt_ser_count_reg_reg_1__U1 ( .A (fsm_countSerial[1]), .ZN (fsm_cnt_ser_n20) ) ;
    INV_X1 fsm_ps_state_reg_0__U1 ( .A (fsm_ps_state_0_), .ZN (fsm_n3) ) ;
    INV_X1 fsm_ps_state_reg_1__U1 ( .A (fsm_ps_state_1_), .ZN (fsm_n5) ) ;
    INV_X1 stateFF_state_U3 ( .A (stateFF_state_n7), .ZN (stateFF_state_n6) ) ;
    INV_X1 stateFF_state_U2 ( .A (stateFF_state_n7), .ZN (stateFF_state_n5) ) ;
    INV_X1 stateFF_state_U1 ( .A (ctrlData_0_), .ZN (stateFF_state_n7) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1 ( .s (ctrlData_0_), .b ({data_out_s3[0], data_out_s2[0], data_out_s1[0], data_out_s0[0]}), .a ({new_AGEMA_signal_936, new_AGEMA_signal_935, new_AGEMA_signal_934, stateFF_inputPar[4]}), .c ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, new_AGEMA_signal_2185, stateFF_state_gff_2_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1 ( .s (ctrlData_0_), .b ({data_out_s3[1], data_out_s2[1], data_out_s1[1], data_out_s0[1]}), .a ({new_AGEMA_signal_945, new_AGEMA_signal_944, new_AGEMA_signal_943, stateFF_inputPar[5]}), .c ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, new_AGEMA_signal_2188, stateFF_state_gff_2_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1 ( .s (ctrlData_0_), .b ({data_out_s3[2], data_out_s2[2], data_out_s1[2], data_out_s0[2]}), .a ({new_AGEMA_signal_954, new_AGEMA_signal_953, new_AGEMA_signal_952, stateFF_inputPar[6]}), .c ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, new_AGEMA_signal_2191, stateFF_state_gff_2_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1 ( .s (ctrlData_0_), .b ({data_out_s3[3], data_out_s2[3], data_out_s1[3], data_out_s0[3]}), .a ({new_AGEMA_signal_963, new_AGEMA_signal_962, new_AGEMA_signal_961, stateFF_inputPar[7]}), .c ({new_AGEMA_signal_2196, new_AGEMA_signal_2195, new_AGEMA_signal_2194, stateFF_state_gff_2_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[4], data_out_s2[4], data_out_s1[4], data_out_s0[4]}), .a ({new_AGEMA_signal_972, new_AGEMA_signal_971, new_AGEMA_signal_970, stateFF_inputPar[8]}), .c ({new_AGEMA_signal_2244, new_AGEMA_signal_2243, new_AGEMA_signal_2242, stateFF_state_gff_3_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[5], data_out_s2[5], data_out_s1[5], data_out_s0[5]}), .a ({new_AGEMA_signal_981, new_AGEMA_signal_980, new_AGEMA_signal_979, stateFF_inputPar[9]}), .c ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, new_AGEMA_signal_2245, stateFF_state_gff_3_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[6], data_out_s2[6], data_out_s1[6], data_out_s0[6]}), .a ({new_AGEMA_signal_990, new_AGEMA_signal_989, new_AGEMA_signal_988, stateFF_inputPar[10]}), .c ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, new_AGEMA_signal_2248, stateFF_state_gff_3_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[7], data_out_s2[7], data_out_s1[7], data_out_s0[7]}), .a ({new_AGEMA_signal_999, new_AGEMA_signal_998, new_AGEMA_signal_997, stateFF_inputPar[11]}), .c ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, new_AGEMA_signal_2251, stateFF_state_gff_3_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[8], data_out_s2[8], data_out_s1[8], data_out_s0[8]}), .a ({new_AGEMA_signal_1008, new_AGEMA_signal_1007, new_AGEMA_signal_1006, stateFF_inputPar[12]}), .c ({new_AGEMA_signal_2256, new_AGEMA_signal_2255, new_AGEMA_signal_2254, stateFF_state_gff_4_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[9], data_out_s2[9], data_out_s1[9], data_out_s0[9]}), .a ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, new_AGEMA_signal_1015, stateFF_inputPar[13]}), .c ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, new_AGEMA_signal_2257, stateFF_state_gff_4_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[10], data_out_s2[10], data_out_s1[10], data_out_s0[10]}), .a ({new_AGEMA_signal_1026, new_AGEMA_signal_1025, new_AGEMA_signal_1024, stateFF_inputPar[14]}), .c ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, new_AGEMA_signal_2260, stateFF_state_gff_4_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[11], data_out_s2[11], data_out_s1[11], data_out_s0[11]}), .a ({new_AGEMA_signal_1032, new_AGEMA_signal_1031, new_AGEMA_signal_1030, stateFF_inputPar[15]}), .c ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, new_AGEMA_signal_2263, stateFF_state_gff_4_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[12], data_out_s2[12], data_out_s1[12], data_out_s0[12]}), .a ({new_AGEMA_signal_1041, new_AGEMA_signal_1040, new_AGEMA_signal_1039, stateFF_inputPar[16]}), .c ({new_AGEMA_signal_2268, new_AGEMA_signal_2267, new_AGEMA_signal_2266, stateFF_state_gff_5_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[13], data_out_s2[13], data_out_s1[13], data_out_s0[13]}), .a ({new_AGEMA_signal_1050, new_AGEMA_signal_1049, new_AGEMA_signal_1048, stateFF_inputPar[17]}), .c ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, new_AGEMA_signal_2269, stateFF_state_gff_5_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[14], data_out_s2[14], data_out_s1[14], data_out_s0[14]}), .a ({new_AGEMA_signal_1059, new_AGEMA_signal_1058, new_AGEMA_signal_1057, stateFF_inputPar[18]}), .c ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, new_AGEMA_signal_2272, stateFF_state_gff_5_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[15], data_out_s2[15], data_out_s1[15], data_out_s0[15]}), .a ({new_AGEMA_signal_1068, new_AGEMA_signal_1067, new_AGEMA_signal_1066, stateFF_inputPar[19]}), .c ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, new_AGEMA_signal_2275, stateFF_state_gff_5_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[16], data_out_s2[16], data_out_s1[16], data_out_s0[16]}), .a ({new_AGEMA_signal_1077, new_AGEMA_signal_1076, new_AGEMA_signal_1075, stateFF_inputPar[20]}), .c ({new_AGEMA_signal_2280, new_AGEMA_signal_2279, new_AGEMA_signal_2278, stateFF_state_gff_6_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[17], data_out_s2[17], data_out_s1[17], data_out_s0[17]}), .a ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, new_AGEMA_signal_1084, stateFF_inputPar[21]}), .c ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, new_AGEMA_signal_2281, stateFF_state_gff_6_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[18], data_out_s2[18], data_out_s1[18], data_out_s0[18]}), .a ({new_AGEMA_signal_1095, new_AGEMA_signal_1094, new_AGEMA_signal_1093, stateFF_inputPar[22]}), .c ({new_AGEMA_signal_2286, new_AGEMA_signal_2285, new_AGEMA_signal_2284, stateFF_state_gff_6_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[19], data_out_s2[19], data_out_s1[19], data_out_s0[19]}), .a ({new_AGEMA_signal_1104, new_AGEMA_signal_1103, new_AGEMA_signal_1102, stateFF_inputPar[23]}), .c ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, new_AGEMA_signal_2287, stateFF_state_gff_6_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[20], data_out_s2[20], data_out_s1[20], data_out_s0[20]}), .a ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, new_AGEMA_signal_1111, stateFF_inputPar[24]}), .c ({new_AGEMA_signal_2292, new_AGEMA_signal_2291, new_AGEMA_signal_2290, stateFF_state_gff_7_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[21], data_out_s2[21], data_out_s1[21], data_out_s0[21]}), .a ({new_AGEMA_signal_1122, new_AGEMA_signal_1121, new_AGEMA_signal_1120, stateFF_inputPar[25]}), .c ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, new_AGEMA_signal_2293, stateFF_state_gff_7_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[22], data_out_s2[22], data_out_s1[22], data_out_s0[22]}), .a ({new_AGEMA_signal_1131, new_AGEMA_signal_1130, new_AGEMA_signal_1129, stateFF_inputPar[26]}), .c ({new_AGEMA_signal_2298, new_AGEMA_signal_2297, new_AGEMA_signal_2296, stateFF_state_gff_7_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[23], data_out_s2[23], data_out_s1[23], data_out_s0[23]}), .a ({new_AGEMA_signal_1140, new_AGEMA_signal_1139, new_AGEMA_signal_1138, stateFF_inputPar[27]}), .c ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, new_AGEMA_signal_2299, stateFF_state_gff_7_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[24], data_out_s2[24], data_out_s1[24], data_out_s0[24]}), .a ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, new_AGEMA_signal_1147, stateFF_inputPar[28]}), .c ({new_AGEMA_signal_2304, new_AGEMA_signal_2303, new_AGEMA_signal_2302, stateFF_state_gff_8_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[25], data_out_s2[25], data_out_s1[25], data_out_s0[25]}), .a ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, new_AGEMA_signal_1156, stateFF_inputPar[29]}), .c ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, new_AGEMA_signal_2305, stateFF_state_gff_8_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[26], data_out_s2[26], data_out_s1[26], data_out_s0[26]}), .a ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, new_AGEMA_signal_1165, stateFF_inputPar[30]}), .c ({new_AGEMA_signal_2310, new_AGEMA_signal_2309, new_AGEMA_signal_2308, stateFF_state_gff_8_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[27], data_out_s2[27], data_out_s1[27], data_out_s0[27]}), .a ({new_AGEMA_signal_1173, new_AGEMA_signal_1172, new_AGEMA_signal_1171, stateFF_inputPar[31]}), .c ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, new_AGEMA_signal_2311, stateFF_state_gff_8_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[28], data_out_s2[28], data_out_s1[28], data_out_s0[28]}), .a ({new_AGEMA_signal_1182, new_AGEMA_signal_1181, new_AGEMA_signal_1180, stateFF_inputPar[32]}), .c ({new_AGEMA_signal_2316, new_AGEMA_signal_2315, new_AGEMA_signal_2314, stateFF_state_gff_9_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[29], data_out_s2[29], data_out_s1[29], data_out_s0[29]}), .a ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, new_AGEMA_signal_1189, stateFF_inputPar[33]}), .c ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, new_AGEMA_signal_2317, stateFF_state_gff_9_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[30], data_out_s2[30], data_out_s1[30], data_out_s0[30]}), .a ({new_AGEMA_signal_1200, new_AGEMA_signal_1199, new_AGEMA_signal_1198, stateFF_inputPar[34]}), .c ({new_AGEMA_signal_2322, new_AGEMA_signal_2321, new_AGEMA_signal_2320, stateFF_state_gff_9_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s3[31], data_out_s2[31], data_out_s1[31], data_out_s0[31]}), .a ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, new_AGEMA_signal_1207, stateFF_inputPar[35]}), .c ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, new_AGEMA_signal_2323, stateFF_state_gff_9_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[32], data_out_s2[32], data_out_s1[32], data_out_s0[32]}), .a ({new_AGEMA_signal_1218, new_AGEMA_signal_1217, new_AGEMA_signal_1216, stateFF_inputPar[36]}), .c ({new_AGEMA_signal_2328, new_AGEMA_signal_2327, new_AGEMA_signal_2326, stateFF_state_gff_10_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[33], data_out_s2[33], data_out_s1[33], data_out_s0[33]}), .a ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, new_AGEMA_signal_1225, stateFF_inputPar[37]}), .c ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, new_AGEMA_signal_2329, stateFF_state_gff_10_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[34], data_out_s2[34], data_out_s1[34], data_out_s0[34]}), .a ({new_AGEMA_signal_1236, new_AGEMA_signal_1235, new_AGEMA_signal_1234, stateFF_inputPar[38]}), .c ({new_AGEMA_signal_2334, new_AGEMA_signal_2333, new_AGEMA_signal_2332, stateFF_state_gff_10_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[35], data_out_s2[35], data_out_s1[35], data_out_s0[35]}), .a ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, new_AGEMA_signal_1243, stateFF_inputPar[39]}), .c ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, new_AGEMA_signal_2335, stateFF_state_gff_10_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[36], data_out_s2[36], data_out_s1[36], data_out_s0[36]}), .a ({new_AGEMA_signal_1254, new_AGEMA_signal_1253, new_AGEMA_signal_1252, stateFF_inputPar[40]}), .c ({new_AGEMA_signal_2340, new_AGEMA_signal_2339, new_AGEMA_signal_2338, stateFF_state_gff_11_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[37], data_out_s2[37], data_out_s1[37], data_out_s0[37]}), .a ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, new_AGEMA_signal_1261, stateFF_inputPar[41]}), .c ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, new_AGEMA_signal_2341, stateFF_state_gff_11_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[38], data_out_s2[38], data_out_s1[38], data_out_s0[38]}), .a ({new_AGEMA_signal_1272, new_AGEMA_signal_1271, new_AGEMA_signal_1270, stateFF_inputPar[42]}), .c ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, new_AGEMA_signal_2344, stateFF_state_gff_11_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[39], data_out_s2[39], data_out_s1[39], data_out_s0[39]}), .a ({new_AGEMA_signal_1281, new_AGEMA_signal_1280, new_AGEMA_signal_1279, stateFF_inputPar[43]}), .c ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, new_AGEMA_signal_2347, stateFF_state_gff_11_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[40], data_out_s2[40], data_out_s1[40], data_out_s0[40]}), .a ({new_AGEMA_signal_1290, new_AGEMA_signal_1289, new_AGEMA_signal_1288, stateFF_inputPar[44]}), .c ({new_AGEMA_signal_2352, new_AGEMA_signal_2351, new_AGEMA_signal_2350, stateFF_state_gff_12_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[41], data_out_s2[41], data_out_s1[41], data_out_s0[41]}), .a ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, new_AGEMA_signal_1297, stateFF_inputPar[45]}), .c ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, new_AGEMA_signal_2353, stateFF_state_gff_12_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[42], data_out_s2[42], data_out_s1[42], data_out_s0[42]}), .a ({new_AGEMA_signal_1308, new_AGEMA_signal_1307, new_AGEMA_signal_1306, stateFF_inputPar[46]}), .c ({new_AGEMA_signal_2358, new_AGEMA_signal_2357, new_AGEMA_signal_2356, stateFF_state_gff_12_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[43], data_out_s2[43], data_out_s1[43], data_out_s0[43]}), .a ({new_AGEMA_signal_1314, new_AGEMA_signal_1313, new_AGEMA_signal_1312, stateFF_inputPar[47]}), .c ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, new_AGEMA_signal_2359, stateFF_state_gff_12_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[44], data_out_s2[44], data_out_s1[44], data_out_s0[44]}), .a ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, new_AGEMA_signal_1321, stateFF_inputPar[48]}), .c ({new_AGEMA_signal_2364, new_AGEMA_signal_2363, new_AGEMA_signal_2362, stateFF_state_gff_13_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[45], data_out_s2[45], data_out_s1[45], data_out_s0[45]}), .a ({new_AGEMA_signal_1332, new_AGEMA_signal_1331, new_AGEMA_signal_1330, stateFF_inputPar[49]}), .c ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, new_AGEMA_signal_2365, stateFF_state_gff_13_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[46], data_out_s2[46], data_out_s1[46], data_out_s0[46]}), .a ({new_AGEMA_signal_1341, new_AGEMA_signal_1340, new_AGEMA_signal_1339, stateFF_inputPar[50]}), .c ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, new_AGEMA_signal_2368, stateFF_state_gff_13_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[47], data_out_s2[47], data_out_s1[47], data_out_s0[47]}), .a ({new_AGEMA_signal_1350, new_AGEMA_signal_1349, new_AGEMA_signal_1348, stateFF_inputPar[51]}), .c ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, new_AGEMA_signal_2371, stateFF_state_gff_13_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[48], data_out_s2[48], data_out_s1[48], data_out_s0[48]}), .a ({new_AGEMA_signal_1359, new_AGEMA_signal_1358, new_AGEMA_signal_1357, stateFF_inputPar[52]}), .c ({new_AGEMA_signal_2376, new_AGEMA_signal_2375, new_AGEMA_signal_2374, stateFF_state_gff_14_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[49], data_out_s2[49], data_out_s1[49], data_out_s0[49]}), .a ({new_AGEMA_signal_1368, new_AGEMA_signal_1367, new_AGEMA_signal_1366, stateFF_inputPar[53]}), .c ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, new_AGEMA_signal_2377, stateFF_state_gff_14_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[50], data_out_s2[50], data_out_s1[50], data_out_s0[50]}), .a ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, new_AGEMA_signal_1375, stateFF_inputPar[54]}), .c ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, new_AGEMA_signal_2380, stateFF_state_gff_14_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[51], data_out_s2[51], data_out_s1[51], data_out_s0[51]}), .a ({new_AGEMA_signal_1386, new_AGEMA_signal_1385, new_AGEMA_signal_1384, stateFF_inputPar[55]}), .c ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, new_AGEMA_signal_2383, stateFF_state_gff_14_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[52], data_out_s2[52], data_out_s1[52], data_out_s0[52]}), .a ({new_AGEMA_signal_1395, new_AGEMA_signal_1394, new_AGEMA_signal_1393, stateFF_inputPar[56]}), .c ({new_AGEMA_signal_2388, new_AGEMA_signal_2387, new_AGEMA_signal_2386, stateFF_state_gff_15_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[53], data_out_s2[53], data_out_s1[53], data_out_s0[53]}), .a ({new_AGEMA_signal_1404, new_AGEMA_signal_1403, new_AGEMA_signal_1402, stateFF_inputPar[57]}), .c ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, new_AGEMA_signal_2389, stateFF_state_gff_15_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[54], data_out_s2[54], data_out_s1[54], data_out_s0[54]}), .a ({new_AGEMA_signal_1413, new_AGEMA_signal_1412, new_AGEMA_signal_1411, stateFF_inputPar[58]}), .c ({new_AGEMA_signal_2394, new_AGEMA_signal_2393, new_AGEMA_signal_2392, stateFF_state_gff_15_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[55], data_out_s2[55], data_out_s1[55], data_out_s0[55]}), .a ({new_AGEMA_signal_1422, new_AGEMA_signal_1421, new_AGEMA_signal_1420, stateFF_inputPar[59]}), .c ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, new_AGEMA_signal_2395, stateFF_state_gff_15_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[56], data_out_s2[56], data_out_s1[56], data_out_s0[56]}), .a ({new_AGEMA_signal_1431, new_AGEMA_signal_1430, new_AGEMA_signal_1429, stateFF_inputPar[60]}), .c ({new_AGEMA_signal_2400, new_AGEMA_signal_2399, new_AGEMA_signal_2398, stateFF_state_gff_16_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[57], data_out_s2[57], data_out_s1[57], data_out_s0[57]}), .a ({new_AGEMA_signal_1440, new_AGEMA_signal_1439, new_AGEMA_signal_1438, stateFF_inputPar[61]}), .c ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, new_AGEMA_signal_2401, stateFF_state_gff_16_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[58], data_out_s2[58], data_out_s1[58], data_out_s0[58]}), .a ({new_AGEMA_signal_1449, new_AGEMA_signal_1448, new_AGEMA_signal_1447, stateFF_inputPar[62]}), .c ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, new_AGEMA_signal_2404, stateFF_state_gff_16_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s3[59], data_out_s2[59], data_out_s1[59], data_out_s0[59]}), .a ({new_AGEMA_signal_1455, new_AGEMA_signal_1454, new_AGEMA_signal_1453, stateFF_inputPar[63]}), .c ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, new_AGEMA_signal_2407, stateFF_state_gff_16_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_0_U1 ( .s (reset), .b ({data_out_s3[0], data_out_s2[0], data_out_s1[0], data_out_s0[0]}), .a ({data_in_s3[0], data_in_s2[0], data_in_s1[0], data_in_s0[0]}), .c ({new_AGEMA_signal_900, new_AGEMA_signal_899, new_AGEMA_signal_898, stateFF_inputPar[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_1_U1 ( .s (reset), .b ({data_out_s3[4], data_out_s2[4], data_out_s1[4], data_out_s0[4]}), .a ({data_in_s3[1], data_in_s2[1], data_in_s1[1], data_in_s0[1]}), .c ({new_AGEMA_signal_909, new_AGEMA_signal_908, new_AGEMA_signal_907, stateFF_inputPar[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_2_U1 ( .s (reset), .b ({data_out_s3[8], data_out_s2[8], data_out_s1[8], data_out_s0[8]}), .a ({data_in_s3[2], data_in_s2[2], data_in_s1[2], data_in_s0[2]}), .c ({new_AGEMA_signal_918, new_AGEMA_signal_917, new_AGEMA_signal_916, stateFF_inputPar[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_3_U1 ( .s (reset), .b ({data_out_s3[12], data_out_s2[12], data_out_s1[12], data_out_s0[12]}), .a ({data_in_s3[3], data_in_s2[3], data_in_s1[3], data_in_s0[3]}), .c ({new_AGEMA_signal_927, new_AGEMA_signal_926, new_AGEMA_signal_925, stateFF_inputPar[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_4_U1 ( .s (reset), .b ({data_out_s3[16], data_out_s2[16], data_out_s1[16], data_out_s0[16]}), .a ({data_in_s3[4], data_in_s2[4], data_in_s1[4], data_in_s0[4]}), .c ({new_AGEMA_signal_936, new_AGEMA_signal_935, new_AGEMA_signal_934, stateFF_inputPar[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_5_U1 ( .s (reset), .b ({data_out_s3[20], data_out_s2[20], data_out_s1[20], data_out_s0[20]}), .a ({data_in_s3[5], data_in_s2[5], data_in_s1[5], data_in_s0[5]}), .c ({new_AGEMA_signal_945, new_AGEMA_signal_944, new_AGEMA_signal_943, stateFF_inputPar[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_6_U1 ( .s (reset), .b ({data_out_s3[24], data_out_s2[24], data_out_s1[24], data_out_s0[24]}), .a ({data_in_s3[6], data_in_s2[6], data_in_s1[6], data_in_s0[6]}), .c ({new_AGEMA_signal_954, new_AGEMA_signal_953, new_AGEMA_signal_952, stateFF_inputPar[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_7_U1 ( .s (reset), .b ({data_out_s3[28], data_out_s2[28], data_out_s1[28], data_out_s0[28]}), .a ({data_in_s3[7], data_in_s2[7], data_in_s1[7], data_in_s0[7]}), .c ({new_AGEMA_signal_963, new_AGEMA_signal_962, new_AGEMA_signal_961, stateFF_inputPar[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_8_U1 ( .s (reset), .b ({data_out_s3[32], data_out_s2[32], data_out_s1[32], data_out_s0[32]}), .a ({data_in_s3[8], data_in_s2[8], data_in_s1[8], data_in_s0[8]}), .c ({new_AGEMA_signal_972, new_AGEMA_signal_971, new_AGEMA_signal_970, stateFF_inputPar[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_9_U1 ( .s (reset), .b ({data_out_s3[36], data_out_s2[36], data_out_s1[36], data_out_s0[36]}), .a ({data_in_s3[9], data_in_s2[9], data_in_s1[9], data_in_s0[9]}), .c ({new_AGEMA_signal_981, new_AGEMA_signal_980, new_AGEMA_signal_979, stateFF_inputPar[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_10_U1 ( .s (reset), .b ({data_out_s3[40], data_out_s2[40], data_out_s1[40], data_out_s0[40]}), .a ({data_in_s3[10], data_in_s2[10], data_in_s1[10], data_in_s0[10]}), .c ({new_AGEMA_signal_990, new_AGEMA_signal_989, new_AGEMA_signal_988, stateFF_inputPar[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_11_U1 ( .s (reset), .b ({data_out_s3[44], data_out_s2[44], data_out_s1[44], data_out_s0[44]}), .a ({data_in_s3[11], data_in_s2[11], data_in_s1[11], data_in_s0[11]}), .c ({new_AGEMA_signal_999, new_AGEMA_signal_998, new_AGEMA_signal_997, stateFF_inputPar[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_12_U1 ( .s (reset), .b ({data_out_s3[48], data_out_s2[48], data_out_s1[48], data_out_s0[48]}), .a ({data_in_s3[12], data_in_s2[12], data_in_s1[12], data_in_s0[12]}), .c ({new_AGEMA_signal_1008, new_AGEMA_signal_1007, new_AGEMA_signal_1006, stateFF_inputPar[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_13_U1 ( .s (reset), .b ({data_out_s3[52], data_out_s2[52], data_out_s1[52], data_out_s0[52]}), .a ({data_in_s3[13], data_in_s2[13], data_in_s1[13], data_in_s0[13]}), .c ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, new_AGEMA_signal_1015, stateFF_inputPar[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_14_U1 ( .s (reset), .b ({data_out_s3[56], data_out_s2[56], data_out_s1[56], data_out_s0[56]}), .a ({data_in_s3[14], data_in_s2[14], data_in_s1[14], data_in_s0[14]}), .c ({new_AGEMA_signal_1026, new_AGEMA_signal_1025, new_AGEMA_signal_1024, stateFF_inputPar[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_15_U1 ( .s (reset), .b ({data_out_s3[60], data_out_s2[60], data_out_s1[60], data_out_s0[60]}), .a ({data_in_s3[15], data_in_s2[15], data_in_s1[15], data_in_s0[15]}), .c ({new_AGEMA_signal_1032, new_AGEMA_signal_1031, new_AGEMA_signal_1030, stateFF_inputPar[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_16_U1 ( .s (reset), .b ({data_out_s3[1], data_out_s2[1], data_out_s1[1], data_out_s0[1]}), .a ({data_in_s3[16], data_in_s2[16], data_in_s1[16], data_in_s0[16]}), .c ({new_AGEMA_signal_1041, new_AGEMA_signal_1040, new_AGEMA_signal_1039, stateFF_inputPar[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_17_U1 ( .s (reset), .b ({data_out_s3[5], data_out_s2[5], data_out_s1[5], data_out_s0[5]}), .a ({data_in_s3[17], data_in_s2[17], data_in_s1[17], data_in_s0[17]}), .c ({new_AGEMA_signal_1050, new_AGEMA_signal_1049, new_AGEMA_signal_1048, stateFF_inputPar[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_18_U1 ( .s (reset), .b ({data_out_s3[9], data_out_s2[9], data_out_s1[9], data_out_s0[9]}), .a ({data_in_s3[18], data_in_s2[18], data_in_s1[18], data_in_s0[18]}), .c ({new_AGEMA_signal_1059, new_AGEMA_signal_1058, new_AGEMA_signal_1057, stateFF_inputPar[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_19_U1 ( .s (reset), .b ({data_out_s3[13], data_out_s2[13], data_out_s1[13], data_out_s0[13]}), .a ({data_in_s3[19], data_in_s2[19], data_in_s1[19], data_in_s0[19]}), .c ({new_AGEMA_signal_1068, new_AGEMA_signal_1067, new_AGEMA_signal_1066, stateFF_inputPar[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_20_U1 ( .s (reset), .b ({data_out_s3[17], data_out_s2[17], data_out_s1[17], data_out_s0[17]}), .a ({data_in_s3[20], data_in_s2[20], data_in_s1[20], data_in_s0[20]}), .c ({new_AGEMA_signal_1077, new_AGEMA_signal_1076, new_AGEMA_signal_1075, stateFF_inputPar[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_21_U1 ( .s (reset), .b ({data_out_s3[21], data_out_s2[21], data_out_s1[21], data_out_s0[21]}), .a ({data_in_s3[21], data_in_s2[21], data_in_s1[21], data_in_s0[21]}), .c ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, new_AGEMA_signal_1084, stateFF_inputPar[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_22_U1 ( .s (reset), .b ({data_out_s3[25], data_out_s2[25], data_out_s1[25], data_out_s0[25]}), .a ({data_in_s3[22], data_in_s2[22], data_in_s1[22], data_in_s0[22]}), .c ({new_AGEMA_signal_1095, new_AGEMA_signal_1094, new_AGEMA_signal_1093, stateFF_inputPar[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_23_U1 ( .s (reset), .b ({data_out_s3[29], data_out_s2[29], data_out_s1[29], data_out_s0[29]}), .a ({data_in_s3[23], data_in_s2[23], data_in_s1[23], data_in_s0[23]}), .c ({new_AGEMA_signal_1104, new_AGEMA_signal_1103, new_AGEMA_signal_1102, stateFF_inputPar[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_24_U1 ( .s (reset), .b ({data_out_s3[33], data_out_s2[33], data_out_s1[33], data_out_s0[33]}), .a ({data_in_s3[24], data_in_s2[24], data_in_s1[24], data_in_s0[24]}), .c ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, new_AGEMA_signal_1111, stateFF_inputPar[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_25_U1 ( .s (reset), .b ({data_out_s3[37], data_out_s2[37], data_out_s1[37], data_out_s0[37]}), .a ({data_in_s3[25], data_in_s2[25], data_in_s1[25], data_in_s0[25]}), .c ({new_AGEMA_signal_1122, new_AGEMA_signal_1121, new_AGEMA_signal_1120, stateFF_inputPar[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_26_U1 ( .s (reset), .b ({data_out_s3[41], data_out_s2[41], data_out_s1[41], data_out_s0[41]}), .a ({data_in_s3[26], data_in_s2[26], data_in_s1[26], data_in_s0[26]}), .c ({new_AGEMA_signal_1131, new_AGEMA_signal_1130, new_AGEMA_signal_1129, stateFF_inputPar[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_27_U1 ( .s (reset), .b ({data_out_s3[45], data_out_s2[45], data_out_s1[45], data_out_s0[45]}), .a ({data_in_s3[27], data_in_s2[27], data_in_s1[27], data_in_s0[27]}), .c ({new_AGEMA_signal_1140, new_AGEMA_signal_1139, new_AGEMA_signal_1138, stateFF_inputPar[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_28_U1 ( .s (reset), .b ({data_out_s3[49], data_out_s2[49], data_out_s1[49], data_out_s0[49]}), .a ({data_in_s3[28], data_in_s2[28], data_in_s1[28], data_in_s0[28]}), .c ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, new_AGEMA_signal_1147, stateFF_inputPar[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_29_U1 ( .s (reset), .b ({data_out_s3[53], data_out_s2[53], data_out_s1[53], data_out_s0[53]}), .a ({data_in_s3[29], data_in_s2[29], data_in_s1[29], data_in_s0[29]}), .c ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, new_AGEMA_signal_1156, stateFF_inputPar[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_30_U1 ( .s (reset), .b ({data_out_s3[57], data_out_s2[57], data_out_s1[57], data_out_s0[57]}), .a ({data_in_s3[30], data_in_s2[30], data_in_s1[30], data_in_s0[30]}), .c ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, new_AGEMA_signal_1165, stateFF_inputPar[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_31_U1 ( .s (reset), .b ({data_out_s3[61], data_out_s2[61], data_out_s1[61], data_out_s0[61]}), .a ({data_in_s3[31], data_in_s2[31], data_in_s1[31], data_in_s0[31]}), .c ({new_AGEMA_signal_1173, new_AGEMA_signal_1172, new_AGEMA_signal_1171, stateFF_inputPar[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_32_U1 ( .s (reset), .b ({data_out_s3[2], data_out_s2[2], data_out_s1[2], data_out_s0[2]}), .a ({data_in_s3[32], data_in_s2[32], data_in_s1[32], data_in_s0[32]}), .c ({new_AGEMA_signal_1182, new_AGEMA_signal_1181, new_AGEMA_signal_1180, stateFF_inputPar[32]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_33_U1 ( .s (reset), .b ({data_out_s3[6], data_out_s2[6], data_out_s1[6], data_out_s0[6]}), .a ({data_in_s3[33], data_in_s2[33], data_in_s1[33], data_in_s0[33]}), .c ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, new_AGEMA_signal_1189, stateFF_inputPar[33]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_34_U1 ( .s (reset), .b ({data_out_s3[10], data_out_s2[10], data_out_s1[10], data_out_s0[10]}), .a ({data_in_s3[34], data_in_s2[34], data_in_s1[34], data_in_s0[34]}), .c ({new_AGEMA_signal_1200, new_AGEMA_signal_1199, new_AGEMA_signal_1198, stateFF_inputPar[34]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_35_U1 ( .s (reset), .b ({data_out_s3[14], data_out_s2[14], data_out_s1[14], data_out_s0[14]}), .a ({data_in_s3[35], data_in_s2[35], data_in_s1[35], data_in_s0[35]}), .c ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, new_AGEMA_signal_1207, stateFF_inputPar[35]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_36_U1 ( .s (reset), .b ({data_out_s3[18], data_out_s2[18], data_out_s1[18], data_out_s0[18]}), .a ({data_in_s3[36], data_in_s2[36], data_in_s1[36], data_in_s0[36]}), .c ({new_AGEMA_signal_1218, new_AGEMA_signal_1217, new_AGEMA_signal_1216, stateFF_inputPar[36]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_37_U1 ( .s (reset), .b ({data_out_s3[22], data_out_s2[22], data_out_s1[22], data_out_s0[22]}), .a ({data_in_s3[37], data_in_s2[37], data_in_s1[37], data_in_s0[37]}), .c ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, new_AGEMA_signal_1225, stateFF_inputPar[37]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_38_U1 ( .s (reset), .b ({data_out_s3[26], data_out_s2[26], data_out_s1[26], data_out_s0[26]}), .a ({data_in_s3[38], data_in_s2[38], data_in_s1[38], data_in_s0[38]}), .c ({new_AGEMA_signal_1236, new_AGEMA_signal_1235, new_AGEMA_signal_1234, stateFF_inputPar[38]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_39_U1 ( .s (reset), .b ({data_out_s3[30], data_out_s2[30], data_out_s1[30], data_out_s0[30]}), .a ({data_in_s3[39], data_in_s2[39], data_in_s1[39], data_in_s0[39]}), .c ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, new_AGEMA_signal_1243, stateFF_inputPar[39]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_40_U1 ( .s (reset), .b ({data_out_s3[34], data_out_s2[34], data_out_s1[34], data_out_s0[34]}), .a ({data_in_s3[40], data_in_s2[40], data_in_s1[40], data_in_s0[40]}), .c ({new_AGEMA_signal_1254, new_AGEMA_signal_1253, new_AGEMA_signal_1252, stateFF_inputPar[40]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_41_U1 ( .s (reset), .b ({data_out_s3[38], data_out_s2[38], data_out_s1[38], data_out_s0[38]}), .a ({data_in_s3[41], data_in_s2[41], data_in_s1[41], data_in_s0[41]}), .c ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, new_AGEMA_signal_1261, stateFF_inputPar[41]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_42_U1 ( .s (reset), .b ({data_out_s3[42], data_out_s2[42], data_out_s1[42], data_out_s0[42]}), .a ({data_in_s3[42], data_in_s2[42], data_in_s1[42], data_in_s0[42]}), .c ({new_AGEMA_signal_1272, new_AGEMA_signal_1271, new_AGEMA_signal_1270, stateFF_inputPar[42]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_43_U1 ( .s (reset), .b ({data_out_s3[46], data_out_s2[46], data_out_s1[46], data_out_s0[46]}), .a ({data_in_s3[43], data_in_s2[43], data_in_s1[43], data_in_s0[43]}), .c ({new_AGEMA_signal_1281, new_AGEMA_signal_1280, new_AGEMA_signal_1279, stateFF_inputPar[43]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_44_U1 ( .s (reset), .b ({data_out_s3[50], data_out_s2[50], data_out_s1[50], data_out_s0[50]}), .a ({data_in_s3[44], data_in_s2[44], data_in_s1[44], data_in_s0[44]}), .c ({new_AGEMA_signal_1290, new_AGEMA_signal_1289, new_AGEMA_signal_1288, stateFF_inputPar[44]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_45_U1 ( .s (reset), .b ({data_out_s3[54], data_out_s2[54], data_out_s1[54], data_out_s0[54]}), .a ({data_in_s3[45], data_in_s2[45], data_in_s1[45], data_in_s0[45]}), .c ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, new_AGEMA_signal_1297, stateFF_inputPar[45]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_46_U1 ( .s (reset), .b ({data_out_s3[58], data_out_s2[58], data_out_s1[58], data_out_s0[58]}), .a ({data_in_s3[46], data_in_s2[46], data_in_s1[46], data_in_s0[46]}), .c ({new_AGEMA_signal_1308, new_AGEMA_signal_1307, new_AGEMA_signal_1306, stateFF_inputPar[46]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_47_U1 ( .s (reset), .b ({data_out_s3[62], data_out_s2[62], data_out_s1[62], data_out_s0[62]}), .a ({data_in_s3[47], data_in_s2[47], data_in_s1[47], data_in_s0[47]}), .c ({new_AGEMA_signal_1314, new_AGEMA_signal_1313, new_AGEMA_signal_1312, stateFF_inputPar[47]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_48_U1 ( .s (reset), .b ({data_out_s3[3], data_out_s2[3], data_out_s1[3], data_out_s0[3]}), .a ({data_in_s3[48], data_in_s2[48], data_in_s1[48], data_in_s0[48]}), .c ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, new_AGEMA_signal_1321, stateFF_inputPar[48]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_49_U1 ( .s (reset), .b ({data_out_s3[7], data_out_s2[7], data_out_s1[7], data_out_s0[7]}), .a ({data_in_s3[49], data_in_s2[49], data_in_s1[49], data_in_s0[49]}), .c ({new_AGEMA_signal_1332, new_AGEMA_signal_1331, new_AGEMA_signal_1330, stateFF_inputPar[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_50_U1 ( .s (reset), .b ({data_out_s3[11], data_out_s2[11], data_out_s1[11], data_out_s0[11]}), .a ({data_in_s3[50], data_in_s2[50], data_in_s1[50], data_in_s0[50]}), .c ({new_AGEMA_signal_1341, new_AGEMA_signal_1340, new_AGEMA_signal_1339, stateFF_inputPar[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_51_U1 ( .s (reset), .b ({data_out_s3[15], data_out_s2[15], data_out_s1[15], data_out_s0[15]}), .a ({data_in_s3[51], data_in_s2[51], data_in_s1[51], data_in_s0[51]}), .c ({new_AGEMA_signal_1350, new_AGEMA_signal_1349, new_AGEMA_signal_1348, stateFF_inputPar[51]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_52_U1 ( .s (reset), .b ({data_out_s3[19], data_out_s2[19], data_out_s1[19], data_out_s0[19]}), .a ({data_in_s3[52], data_in_s2[52], data_in_s1[52], data_in_s0[52]}), .c ({new_AGEMA_signal_1359, new_AGEMA_signal_1358, new_AGEMA_signal_1357, stateFF_inputPar[52]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_53_U1 ( .s (reset), .b ({data_out_s3[23], data_out_s2[23], data_out_s1[23], data_out_s0[23]}), .a ({data_in_s3[53], data_in_s2[53], data_in_s1[53], data_in_s0[53]}), .c ({new_AGEMA_signal_1368, new_AGEMA_signal_1367, new_AGEMA_signal_1366, stateFF_inputPar[53]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_54_U1 ( .s (reset), .b ({data_out_s3[27], data_out_s2[27], data_out_s1[27], data_out_s0[27]}), .a ({data_in_s3[54], data_in_s2[54], data_in_s1[54], data_in_s0[54]}), .c ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, new_AGEMA_signal_1375, stateFF_inputPar[54]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_55_U1 ( .s (reset), .b ({data_out_s3[31], data_out_s2[31], data_out_s1[31], data_out_s0[31]}), .a ({data_in_s3[55], data_in_s2[55], data_in_s1[55], data_in_s0[55]}), .c ({new_AGEMA_signal_1386, new_AGEMA_signal_1385, new_AGEMA_signal_1384, stateFF_inputPar[55]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_56_U1 ( .s (reset), .b ({data_out_s3[35], data_out_s2[35], data_out_s1[35], data_out_s0[35]}), .a ({data_in_s3[56], data_in_s2[56], data_in_s1[56], data_in_s0[56]}), .c ({new_AGEMA_signal_1395, new_AGEMA_signal_1394, new_AGEMA_signal_1393, stateFF_inputPar[56]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_57_U1 ( .s (reset), .b ({data_out_s3[39], data_out_s2[39], data_out_s1[39], data_out_s0[39]}), .a ({data_in_s3[57], data_in_s2[57], data_in_s1[57], data_in_s0[57]}), .c ({new_AGEMA_signal_1404, new_AGEMA_signal_1403, new_AGEMA_signal_1402, stateFF_inputPar[57]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_58_U1 ( .s (reset), .b ({data_out_s3[43], data_out_s2[43], data_out_s1[43], data_out_s0[43]}), .a ({data_in_s3[58], data_in_s2[58], data_in_s1[58], data_in_s0[58]}), .c ({new_AGEMA_signal_1413, new_AGEMA_signal_1412, new_AGEMA_signal_1411, stateFF_inputPar[58]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_59_U1 ( .s (reset), .b ({data_out_s3[47], data_out_s2[47], data_out_s1[47], data_out_s0[47]}), .a ({data_in_s3[59], data_in_s2[59], data_in_s1[59], data_in_s0[59]}), .c ({new_AGEMA_signal_1422, new_AGEMA_signal_1421, new_AGEMA_signal_1420, stateFF_inputPar[59]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_60_U1 ( .s (reset), .b ({data_out_s3[51], data_out_s2[51], data_out_s1[51], data_out_s0[51]}), .a ({data_in_s3[60], data_in_s2[60], data_in_s1[60], data_in_s0[60]}), .c ({new_AGEMA_signal_1431, new_AGEMA_signal_1430, new_AGEMA_signal_1429, stateFF_inputPar[60]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_61_U1 ( .s (reset), .b ({data_out_s3[55], data_out_s2[55], data_out_s1[55], data_out_s0[55]}), .a ({data_in_s3[61], data_in_s2[61], data_in_s1[61], data_in_s0[61]}), .c ({new_AGEMA_signal_1440, new_AGEMA_signal_1439, new_AGEMA_signal_1438, stateFF_inputPar[61]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_62_U1 ( .s (reset), .b ({data_out_s3[59], data_out_s2[59], data_out_s1[59], data_out_s0[59]}), .a ({data_in_s3[62], data_in_s2[62], data_in_s1[62], data_in_s0[62]}), .c ({new_AGEMA_signal_1449, new_AGEMA_signal_1448, new_AGEMA_signal_1447, stateFF_inputPar[62]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_63_U1 ( .s (reset), .b ({data_out_s3[63], data_out_s2[63], data_out_s1[63], data_out_s0[63]}), .a ({data_in_s3[63], data_in_s2[63], data_in_s1[63], data_in_s0[63]}), .c ({new_AGEMA_signal_1455, new_AGEMA_signal_1454, new_AGEMA_signal_1453, stateFF_inputPar[63]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keyFF_U5 ( .a ({1'b0, 1'b0, 1'b0, counter[4]}), .b ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, new_AGEMA_signal_1456, keyFF_outputPar[22]}), .c ({new_AGEMA_signal_1461, new_AGEMA_signal_1460, new_AGEMA_signal_1459, keyFF_counterAdd[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keyFF_U4 ( .a ({1'b0, 1'b0, 1'b0, counter[3]}), .b ({new_AGEMA_signal_1464, new_AGEMA_signal_1463, new_AGEMA_signal_1462, keyFF_outputPar[21]}), .c ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, new_AGEMA_signal_1465, keyFF_counterAdd[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keyFF_U3 ( .a ({1'b0, 1'b0, 1'b0, counter[2]}), .b ({new_AGEMA_signal_1470, new_AGEMA_signal_1469, new_AGEMA_signal_1468, keyFF_outputPar[20]}), .c ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, new_AGEMA_signal_1471, keyFF_counterAdd[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keyFF_U2 ( .a ({1'b0, 1'b0, 1'b0, counter[1]}), .b ({new_AGEMA_signal_2112, new_AGEMA_signal_2111, new_AGEMA_signal_2110, keyFF_outputPar[19]}), .c ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, new_AGEMA_signal_2113, keyFF_counterAdd[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keyFF_U1 ( .a ({1'b0, 1'b0, 1'b0, counter[0]}), .b ({new_AGEMA_signal_1476, new_AGEMA_signal_1475, new_AGEMA_signal_1474, keyFF_outputPar[18]}), .c ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, new_AGEMA_signal_1477, keyFF_counterAdd[0]}) ) ;
    INV_X1 keyFF_keystate_U3 ( .A (keyFF_keystate_n8), .ZN (keyFF_keystate_n6) ) ;
    INV_X1 keyFF_keystate_U2 ( .A (keyFF_keystate_n8), .ZN (keyFF_keystate_n7) ) ;
    INV_X1 keyFF_keystate_U1 ( .A (ctrlData_0_), .ZN (keyFF_keystate_n8) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_858, new_AGEMA_signal_857, new_AGEMA_signal_856, roundkey[0]}), .a ({new_AGEMA_signal_1488, new_AGEMA_signal_1487, new_AGEMA_signal_1486, keyFF_inputPar[0]}), .c ({new_AGEMA_signal_2412, new_AGEMA_signal_2411, new_AGEMA_signal_2410, keyFF_keystate_gff_1_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_867, new_AGEMA_signal_866, new_AGEMA_signal_865, roundkey[1]}), .a ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, new_AGEMA_signal_1495, keyFF_inputPar[1]}), .c ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, new_AGEMA_signal_2413, keyFF_keystate_gff_1_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_876, new_AGEMA_signal_875, new_AGEMA_signal_874, roundkey[2]}), .a ({new_AGEMA_signal_1506, new_AGEMA_signal_1505, new_AGEMA_signal_1504, keyFF_inputPar[2]}), .c ({new_AGEMA_signal_2418, new_AGEMA_signal_2417, new_AGEMA_signal_2416, keyFF_keystate_gff_1_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_885, new_AGEMA_signal_884, new_AGEMA_signal_883, roundkey[3]}), .a ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, new_AGEMA_signal_1513, keyFF_inputPar[3]}), .c ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, new_AGEMA_signal_2419, keyFF_keystate_gff_1_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, new_AGEMA_signal_2149, keyRegKS[1]}), .a ({new_AGEMA_signal_1524, new_AGEMA_signal_1523, new_AGEMA_signal_1522, keyFF_inputPar[4]}), .c ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, new_AGEMA_signal_2422, keyFF_keystate_gff_2_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, new_AGEMA_signal_2155, keyRegKS[2]}), .a ({new_AGEMA_signal_1533, new_AGEMA_signal_1532, new_AGEMA_signal_1531, keyFF_inputPar[5]}), .c ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, new_AGEMA_signal_2425, keyFF_keystate_gff_2_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, new_AGEMA_signal_2161, keyRegKS[3]}), .a ({new_AGEMA_signal_1542, new_AGEMA_signal_1541, new_AGEMA_signal_1540, keyFF_inputPar[6]}), .c ({new_AGEMA_signal_2430, new_AGEMA_signal_2429, new_AGEMA_signal_2428, keyFF_keystate_gff_2_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1482, new_AGEMA_signal_1481, new_AGEMA_signal_1480, keyFF_outputPar[3]}), .a ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, new_AGEMA_signal_1549, keyFF_inputPar[7]}), .c ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, new_AGEMA_signal_2431, keyFF_keystate_gff_2_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, new_AGEMA_signal_1489, keyFF_outputPar[4]}), .a ({new_AGEMA_signal_1560, new_AGEMA_signal_1559, new_AGEMA_signal_1558, keyFF_inputPar[8]}), .c ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, new_AGEMA_signal_2434, keyFF_keystate_gff_3_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1500, new_AGEMA_signal_1499, new_AGEMA_signal_1498, keyFF_outputPar[5]}), .a ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, new_AGEMA_signal_1567, keyFF_inputPar[9]}), .c ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, new_AGEMA_signal_2437, keyFF_keystate_gff_3_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, new_AGEMA_signal_1507, keyFF_outputPar[6]}), .a ({new_AGEMA_signal_1578, new_AGEMA_signal_1577, new_AGEMA_signal_1576, keyFF_inputPar[10]}), .c ({new_AGEMA_signal_2442, new_AGEMA_signal_2441, new_AGEMA_signal_2440, keyFF_keystate_gff_3_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1518, new_AGEMA_signal_1517, new_AGEMA_signal_1516, keyFF_outputPar[7]}), .a ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, new_AGEMA_signal_1585, keyFF_inputPar[11]}), .c ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, new_AGEMA_signal_2443, keyFF_keystate_gff_3_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, new_AGEMA_signal_1525, keyFF_outputPar[8]}), .a ({new_AGEMA_signal_1596, new_AGEMA_signal_1595, new_AGEMA_signal_1594, keyFF_inputPar[12]}), .c ({new_AGEMA_signal_2448, new_AGEMA_signal_2447, new_AGEMA_signal_2446, keyFF_keystate_gff_4_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1536, new_AGEMA_signal_1535, new_AGEMA_signal_1534, keyFF_outputPar[9]}), .a ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, new_AGEMA_signal_1603, keyFF_inputPar[13]}), .c ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, new_AGEMA_signal_2449, keyFF_keystate_gff_4_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, new_AGEMA_signal_1543, keyFF_outputPar[10]}), .a ({new_AGEMA_signal_1614, new_AGEMA_signal_1613, new_AGEMA_signal_1612, keyFF_inputPar[14]}), .c ({new_AGEMA_signal_2454, new_AGEMA_signal_2453, new_AGEMA_signal_2452, keyFF_keystate_gff_4_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1554, new_AGEMA_signal_1553, new_AGEMA_signal_1552, keyFF_outputPar[11]}), .a ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, new_AGEMA_signal_2119, keyFF_inputPar[15]}), .c ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, new_AGEMA_signal_2455, keyFF_keystate_gff_4_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1563, new_AGEMA_signal_1562, new_AGEMA_signal_1561, keyFF_outputPar[12]}), .a ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, new_AGEMA_signal_2143, keyFF_inputPar[16]}), .c ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, new_AGEMA_signal_2197, keyFF_keystate_gff_5_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, new_AGEMA_signal_1570, keyFF_outputPar[13]}), .a ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, new_AGEMA_signal_2125, keyFF_inputPar[17]}), .c ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, new_AGEMA_signal_2200, keyFF_keystate_gff_5_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, new_AGEMA_signal_1579, keyFF_outputPar[14]}), .a ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, new_AGEMA_signal_2131, keyFF_inputPar[18]}), .c ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, new_AGEMA_signal_2203, keyFF_keystate_gff_5_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1590, new_AGEMA_signal_1589, new_AGEMA_signal_1588, keyFF_outputPar[15]}), .a ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, new_AGEMA_signal_2137, keyFF_inputPar[19]}), .c ({new_AGEMA_signal_2208, new_AGEMA_signal_2207, new_AGEMA_signal_2206, keyFF_keystate_gff_5_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, new_AGEMA_signal_1597, keyFF_outputPar[16]}), .a ({new_AGEMA_signal_1623, new_AGEMA_signal_1622, new_AGEMA_signal_1621, keyFF_inputPar[20]}), .c ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, new_AGEMA_signal_2209, keyFF_keystate_gff_6_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, new_AGEMA_signal_1606, keyFF_outputPar[17]}), .a ({new_AGEMA_signal_1632, new_AGEMA_signal_1631, new_AGEMA_signal_1630, keyFF_inputPar[21]}), .c ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, new_AGEMA_signal_2212, keyFF_keystate_gff_6_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1476, new_AGEMA_signal_1475, new_AGEMA_signal_1474, keyFF_outputPar[18]}), .a ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, new_AGEMA_signal_1639, keyFF_inputPar[22]}), .c ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, new_AGEMA_signal_2215, keyFF_keystate_gff_6_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_2112, new_AGEMA_signal_2111, new_AGEMA_signal_2110, keyFF_outputPar[19]}), .a ({new_AGEMA_signal_1650, new_AGEMA_signal_1649, new_AGEMA_signal_1648, keyFF_inputPar[23]}), .c ({new_AGEMA_signal_2220, new_AGEMA_signal_2219, new_AGEMA_signal_2218, keyFF_keystate_gff_6_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1470, new_AGEMA_signal_1469, new_AGEMA_signal_1468, keyFF_outputPar[20]}), .a ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, new_AGEMA_signal_1657, keyFF_inputPar[24]}), .c ({new_AGEMA_signal_2460, new_AGEMA_signal_2459, new_AGEMA_signal_2458, keyFF_keystate_gff_7_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1464, new_AGEMA_signal_1463, new_AGEMA_signal_1462, keyFF_outputPar[21]}), .a ({new_AGEMA_signal_1668, new_AGEMA_signal_1667, new_AGEMA_signal_1666, keyFF_inputPar[25]}), .c ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, new_AGEMA_signal_2461, keyFF_keystate_gff_7_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, new_AGEMA_signal_1456, keyFF_outputPar[22]}), .a ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, new_AGEMA_signal_1675, keyFF_inputPar[26]}), .c ({new_AGEMA_signal_2466, new_AGEMA_signal_2465, new_AGEMA_signal_2464, keyFF_keystate_gff_7_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, new_AGEMA_signal_1615, keyFF_outputPar[23]}), .a ({new_AGEMA_signal_1686, new_AGEMA_signal_1685, new_AGEMA_signal_1684, keyFF_inputPar[27]}), .c ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, new_AGEMA_signal_2467, keyFF_keystate_gff_7_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1626, new_AGEMA_signal_1625, new_AGEMA_signal_1624, keyFF_outputPar[24]}), .a ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, new_AGEMA_signal_1693, keyFF_inputPar[28]}), .c ({new_AGEMA_signal_2472, new_AGEMA_signal_2471, new_AGEMA_signal_2470, keyFF_keystate_gff_8_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, new_AGEMA_signal_1633, keyFF_outputPar[25]}), .a ({new_AGEMA_signal_1704, new_AGEMA_signal_1703, new_AGEMA_signal_1702, keyFF_inputPar[29]}), .c ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, new_AGEMA_signal_2473, keyFF_keystate_gff_8_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1644, new_AGEMA_signal_1643, new_AGEMA_signal_1642, keyFF_outputPar[26]}), .a ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, new_AGEMA_signal_1711, keyFF_inputPar[30]}), .c ({new_AGEMA_signal_2478, new_AGEMA_signal_2477, new_AGEMA_signal_2476, keyFF_keystate_gff_8_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, new_AGEMA_signal_1651, keyFF_outputPar[27]}), .a ({new_AGEMA_signal_1722, new_AGEMA_signal_1721, new_AGEMA_signal_1720, keyFF_inputPar[31]}), .c ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, new_AGEMA_signal_2479, keyFF_keystate_gff_8_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1662, new_AGEMA_signal_1661, new_AGEMA_signal_1660, keyFF_outputPar[28]}), .a ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, new_AGEMA_signal_1729, keyFF_inputPar[32]}), .c ({new_AGEMA_signal_2484, new_AGEMA_signal_2483, new_AGEMA_signal_2482, keyFF_keystate_gff_9_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, new_AGEMA_signal_1669, keyFF_outputPar[29]}), .a ({new_AGEMA_signal_1740, new_AGEMA_signal_1739, new_AGEMA_signal_1738, keyFF_inputPar[33]}), .c ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, new_AGEMA_signal_2485, keyFF_keystate_gff_9_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1680, new_AGEMA_signal_1679, new_AGEMA_signal_1678, keyFF_outputPar[30]}), .a ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, new_AGEMA_signal_1747, keyFF_inputPar[34]}), .c ({new_AGEMA_signal_2490, new_AGEMA_signal_2489, new_AGEMA_signal_2488, keyFF_keystate_gff_9_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, new_AGEMA_signal_1687, keyFF_outputPar[31]}), .a ({new_AGEMA_signal_1758, new_AGEMA_signal_1757, new_AGEMA_signal_1756, keyFF_inputPar[35]}), .c ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, new_AGEMA_signal_2491, keyFF_keystate_gff_9_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, new_AGEMA_signal_1696, keyFF_outputPar[32]}), .a ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, new_AGEMA_signal_1765, keyFF_inputPar[36]}), .c ({new_AGEMA_signal_2496, new_AGEMA_signal_2495, new_AGEMA_signal_2494, keyFF_keystate_gff_10_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, new_AGEMA_signal_1705, keyFF_outputPar[33]}), .a ({new_AGEMA_signal_1776, new_AGEMA_signal_1775, new_AGEMA_signal_1774, keyFF_inputPar[37]}), .c ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, new_AGEMA_signal_2497, keyFF_keystate_gff_10_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1716, new_AGEMA_signal_1715, new_AGEMA_signal_1714, keyFF_outputPar[34]}), .a ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, new_AGEMA_signal_1783, keyFF_inputPar[38]}), .c ({new_AGEMA_signal_2502, new_AGEMA_signal_2501, new_AGEMA_signal_2500, keyFF_keystate_gff_10_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, new_AGEMA_signal_1723, keyFF_outputPar[35]}), .a ({new_AGEMA_signal_1794, new_AGEMA_signal_1793, new_AGEMA_signal_1792, keyFF_inputPar[39]}), .c ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, new_AGEMA_signal_2503, keyFF_keystate_gff_10_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1734, new_AGEMA_signal_1733, new_AGEMA_signal_1732, keyFF_outputPar[36]}), .a ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, new_AGEMA_signal_1801, keyFF_inputPar[40]}), .c ({new_AGEMA_signal_2508, new_AGEMA_signal_2507, new_AGEMA_signal_2506, keyFF_keystate_gff_11_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, new_AGEMA_signal_1741, keyFF_outputPar[37]}), .a ({new_AGEMA_signal_1812, new_AGEMA_signal_1811, new_AGEMA_signal_1810, keyFF_inputPar[41]}), .c ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, new_AGEMA_signal_2509, keyFF_keystate_gff_11_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1752, new_AGEMA_signal_1751, new_AGEMA_signal_1750, keyFF_outputPar[38]}), .a ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, new_AGEMA_signal_1819, keyFF_inputPar[42]}), .c ({new_AGEMA_signal_2514, new_AGEMA_signal_2513, new_AGEMA_signal_2512, keyFF_keystate_gff_11_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, new_AGEMA_signal_1759, keyFF_outputPar[39]}), .a ({new_AGEMA_signal_1830, new_AGEMA_signal_1829, new_AGEMA_signal_1828, keyFF_inputPar[43]}), .c ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, new_AGEMA_signal_2515, keyFF_keystate_gff_11_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, new_AGEMA_signal_1768, keyFF_outputPar[40]}), .a ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, new_AGEMA_signal_1837, keyFF_inputPar[44]}), .c ({new_AGEMA_signal_2520, new_AGEMA_signal_2519, new_AGEMA_signal_2518, keyFF_keystate_gff_12_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, new_AGEMA_signal_1777, keyFF_outputPar[41]}), .a ({new_AGEMA_signal_1848, new_AGEMA_signal_1847, new_AGEMA_signal_1846, keyFF_inputPar[45]}), .c ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, new_AGEMA_signal_2521, keyFF_keystate_gff_12_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, new_AGEMA_signal_1786, keyFF_outputPar[42]}), .a ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, new_AGEMA_signal_1855, keyFF_inputPar[46]}), .c ({new_AGEMA_signal_2526, new_AGEMA_signal_2525, new_AGEMA_signal_2524, keyFF_keystate_gff_12_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, new_AGEMA_signal_1795, keyFF_outputPar[43]}), .a ({new_AGEMA_signal_1866, new_AGEMA_signal_1865, new_AGEMA_signal_1864, keyFF_inputPar[47]}), .c ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, new_AGEMA_signal_2527, keyFF_keystate_gff_12_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1806, new_AGEMA_signal_1805, new_AGEMA_signal_1804, keyFF_outputPar[44]}), .a ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, new_AGEMA_signal_1873, keyFF_inputPar[48]}), .c ({new_AGEMA_signal_2532, new_AGEMA_signal_2531, new_AGEMA_signal_2530, keyFF_keystate_gff_13_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, new_AGEMA_signal_1813, keyFF_outputPar[45]}), .a ({new_AGEMA_signal_1884, new_AGEMA_signal_1883, new_AGEMA_signal_1882, keyFF_inputPar[49]}), .c ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, new_AGEMA_signal_2533, keyFF_keystate_gff_13_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1824, new_AGEMA_signal_1823, new_AGEMA_signal_1822, keyFF_outputPar[46]}), .a ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, new_AGEMA_signal_1891, keyFF_inputPar[50]}), .c ({new_AGEMA_signal_2538, new_AGEMA_signal_2537, new_AGEMA_signal_2536, keyFF_keystate_gff_13_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, new_AGEMA_signal_1831, keyFF_outputPar[47]}), .a ({new_AGEMA_signal_1902, new_AGEMA_signal_1901, new_AGEMA_signal_1900, keyFF_inputPar[51]}), .c ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, new_AGEMA_signal_2539, keyFF_keystate_gff_13_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1842, new_AGEMA_signal_1841, new_AGEMA_signal_1840, keyFF_outputPar[48]}), .a ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, new_AGEMA_signal_1909, keyFF_inputPar[52]}), .c ({new_AGEMA_signal_2544, new_AGEMA_signal_2543, new_AGEMA_signal_2542, keyFF_keystate_gff_14_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, new_AGEMA_signal_1849, keyFF_outputPar[49]}), .a ({new_AGEMA_signal_1920, new_AGEMA_signal_1919, new_AGEMA_signal_1918, keyFF_inputPar[53]}), .c ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, new_AGEMA_signal_2545, keyFF_keystate_gff_14_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1860, new_AGEMA_signal_1859, new_AGEMA_signal_1858, keyFF_outputPar[50]}), .a ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, new_AGEMA_signal_1927, keyFF_inputPar[54]}), .c ({new_AGEMA_signal_2550, new_AGEMA_signal_2549, new_AGEMA_signal_2548, keyFF_keystate_gff_14_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, new_AGEMA_signal_1867, keyFF_outputPar[51]}), .a ({new_AGEMA_signal_1938, new_AGEMA_signal_1937, new_AGEMA_signal_1936, keyFF_inputPar[55]}), .c ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, new_AGEMA_signal_2551, keyFF_keystate_gff_14_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1878, new_AGEMA_signal_1877, new_AGEMA_signal_1876, keyFF_outputPar[52]}), .a ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, new_AGEMA_signal_1945, keyFF_inputPar[56]}), .c ({new_AGEMA_signal_2556, new_AGEMA_signal_2555, new_AGEMA_signal_2554, keyFF_keystate_gff_15_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, new_AGEMA_signal_1885, keyFF_outputPar[53]}), .a ({new_AGEMA_signal_1956, new_AGEMA_signal_1955, new_AGEMA_signal_1954, keyFF_inputPar[57]}), .c ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, new_AGEMA_signal_2557, keyFF_keystate_gff_15_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1896, new_AGEMA_signal_1895, new_AGEMA_signal_1894, keyFF_outputPar[54]}), .a ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, new_AGEMA_signal_1963, keyFF_inputPar[58]}), .c ({new_AGEMA_signal_2562, new_AGEMA_signal_2561, new_AGEMA_signal_2560, keyFF_keystate_gff_15_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, new_AGEMA_signal_1903, keyFF_outputPar[55]}), .a ({new_AGEMA_signal_1974, new_AGEMA_signal_1973, new_AGEMA_signal_1972, keyFF_inputPar[59]}), .c ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, new_AGEMA_signal_2563, keyFF_keystate_gff_15_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1914, new_AGEMA_signal_1913, new_AGEMA_signal_1912, keyFF_outputPar[56]}), .a ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, new_AGEMA_signal_1981, keyFF_inputPar[60]}), .c ({new_AGEMA_signal_2568, new_AGEMA_signal_2567, new_AGEMA_signal_2566, keyFF_keystate_gff_16_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, new_AGEMA_signal_1921, keyFF_outputPar[57]}), .a ({new_AGEMA_signal_1992, new_AGEMA_signal_1991, new_AGEMA_signal_1990, keyFF_inputPar[61]}), .c ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, new_AGEMA_signal_2569, keyFF_keystate_gff_16_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1932, new_AGEMA_signal_1931, new_AGEMA_signal_1930, keyFF_outputPar[58]}), .a ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, new_AGEMA_signal_1999, keyFF_inputPar[62]}), .c ({new_AGEMA_signal_2574, new_AGEMA_signal_2573, new_AGEMA_signal_2572, keyFF_keystate_gff_16_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, new_AGEMA_signal_1939, keyFF_outputPar[59]}), .a ({new_AGEMA_signal_2010, new_AGEMA_signal_2009, new_AGEMA_signal_2008, keyFF_inputPar[63]}), .c ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, new_AGEMA_signal_2575, keyFF_keystate_gff_16_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1950, new_AGEMA_signal_1949, new_AGEMA_signal_1948, keyFF_outputPar[60]}), .a ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, new_AGEMA_signal_2017, keyFF_inputPar[64]}), .c ({new_AGEMA_signal_2580, new_AGEMA_signal_2579, new_AGEMA_signal_2578, keyFF_keystate_gff_17_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, new_AGEMA_signal_1957, keyFF_outputPar[61]}), .a ({new_AGEMA_signal_2028, new_AGEMA_signal_2027, new_AGEMA_signal_2026, keyFF_inputPar[65]}), .c ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, new_AGEMA_signal_2581, keyFF_keystate_gff_17_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1968, new_AGEMA_signal_1967, new_AGEMA_signal_1966, keyFF_outputPar[62]}), .a ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, new_AGEMA_signal_2035, keyFF_inputPar[66]}), .c ({new_AGEMA_signal_2586, new_AGEMA_signal_2585, new_AGEMA_signal_2584, keyFF_keystate_gff_17_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, new_AGEMA_signal_1975, keyFF_outputPar[63]}), .a ({new_AGEMA_signal_2046, new_AGEMA_signal_2045, new_AGEMA_signal_2044, keyFF_inputPar[67]}), .c ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, new_AGEMA_signal_2587, keyFF_keystate_gff_17_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1986, new_AGEMA_signal_1985, new_AGEMA_signal_1984, keyFF_outputPar[64]}), .a ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, new_AGEMA_signal_2053, keyFF_inputPar[68]}), .c ({new_AGEMA_signal_2592, new_AGEMA_signal_2591, new_AGEMA_signal_2590, keyFF_keystate_gff_18_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, new_AGEMA_signal_1993, keyFF_outputPar[65]}), .a ({new_AGEMA_signal_2064, new_AGEMA_signal_2063, new_AGEMA_signal_2062, keyFF_inputPar[69]}), .c ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, new_AGEMA_signal_2593, keyFF_keystate_gff_18_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_2004, new_AGEMA_signal_2003, new_AGEMA_signal_2002, keyFF_outputPar[66]}), .a ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, new_AGEMA_signal_2071, keyFF_inputPar[70]}), .c ({new_AGEMA_signal_2598, new_AGEMA_signal_2597, new_AGEMA_signal_2596, keyFF_keystate_gff_18_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, new_AGEMA_signal_2011, keyFF_outputPar[67]}), .a ({new_AGEMA_signal_2082, new_AGEMA_signal_2081, new_AGEMA_signal_2080, keyFF_inputPar[71]}), .c ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, new_AGEMA_signal_2599, keyFF_keystate_gff_18_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_2022, new_AGEMA_signal_2021, new_AGEMA_signal_2020, keyFF_outputPar[68]}), .a ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, new_AGEMA_signal_2089, keyFF_inputPar[72]}), .c ({new_AGEMA_signal_2604, new_AGEMA_signal_2603, new_AGEMA_signal_2602, keyFF_keystate_gff_19_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, new_AGEMA_signal_2029, keyFF_outputPar[69]}), .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, new_AGEMA_signal_2095, keyFF_inputPar[73]}), .c ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, new_AGEMA_signal_2605, keyFF_keystate_gff_19_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_2040, new_AGEMA_signal_2039, new_AGEMA_signal_2038, keyFF_outputPar[70]}), .a ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, new_AGEMA_signal_2101, keyFF_inputPar[74]}), .c ({new_AGEMA_signal_2610, new_AGEMA_signal_2609, new_AGEMA_signal_2608, keyFF_keystate_gff_19_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, new_AGEMA_signal_2047, keyFF_outputPar[71]}), .a ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, new_AGEMA_signal_2107, keyFF_inputPar[75]}), .c ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, new_AGEMA_signal_2611, keyFF_keystate_gff_19_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_0_U1 ( .s (reset), .b ({new_AGEMA_signal_1482, new_AGEMA_signal_1481, new_AGEMA_signal_1480, keyFF_outputPar[3]}), .a ({key_s3[0], key_s2[0], key_s1[0], key_s0[0]}), .c ({new_AGEMA_signal_1488, new_AGEMA_signal_1487, new_AGEMA_signal_1486, keyFF_inputPar[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_1_U1 ( .s (reset), .b ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, new_AGEMA_signal_1489, keyFF_outputPar[4]}), .a ({key_s3[1], key_s2[1], key_s1[1], key_s0[1]}), .c ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, new_AGEMA_signal_1495, keyFF_inputPar[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_2_U1 ( .s (reset), .b ({new_AGEMA_signal_1500, new_AGEMA_signal_1499, new_AGEMA_signal_1498, keyFF_outputPar[5]}), .a ({key_s3[2], key_s2[2], key_s1[2], key_s0[2]}), .c ({new_AGEMA_signal_1506, new_AGEMA_signal_1505, new_AGEMA_signal_1504, keyFF_inputPar[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_3_U1 ( .s (reset), .b ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, new_AGEMA_signal_1507, keyFF_outputPar[6]}), .a ({key_s3[3], key_s2[3], key_s1[3], key_s0[3]}), .c ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, new_AGEMA_signal_1513, keyFF_inputPar[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_4_U1 ( .s (reset), .b ({new_AGEMA_signal_1518, new_AGEMA_signal_1517, new_AGEMA_signal_1516, keyFF_outputPar[7]}), .a ({key_s3[4], key_s2[4], key_s1[4], key_s0[4]}), .c ({new_AGEMA_signal_1524, new_AGEMA_signal_1523, new_AGEMA_signal_1522, keyFF_inputPar[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_5_U1 ( .s (reset), .b ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, new_AGEMA_signal_1525, keyFF_outputPar[8]}), .a ({key_s3[5], key_s2[5], key_s1[5], key_s0[5]}), .c ({new_AGEMA_signal_1533, new_AGEMA_signal_1532, new_AGEMA_signal_1531, keyFF_inputPar[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_6_U1 ( .s (reset), .b ({new_AGEMA_signal_1536, new_AGEMA_signal_1535, new_AGEMA_signal_1534, keyFF_outputPar[9]}), .a ({key_s3[6], key_s2[6], key_s1[6], key_s0[6]}), .c ({new_AGEMA_signal_1542, new_AGEMA_signal_1541, new_AGEMA_signal_1540, keyFF_inputPar[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_7_U1 ( .s (reset), .b ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, new_AGEMA_signal_1543, keyFF_outputPar[10]}), .a ({key_s3[7], key_s2[7], key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, new_AGEMA_signal_1549, keyFF_inputPar[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_8_U1 ( .s (reset), .b ({new_AGEMA_signal_1554, new_AGEMA_signal_1553, new_AGEMA_signal_1552, keyFF_outputPar[11]}), .a ({key_s3[8], key_s2[8], key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_1560, new_AGEMA_signal_1559, new_AGEMA_signal_1558, keyFF_inputPar[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_9_U1 ( .s (reset), .b ({new_AGEMA_signal_1563, new_AGEMA_signal_1562, new_AGEMA_signal_1561, keyFF_outputPar[12]}), .a ({key_s3[9], key_s2[9], key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, new_AGEMA_signal_1567, keyFF_inputPar[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_10_U1 ( .s (reset), .b ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, new_AGEMA_signal_1570, keyFF_outputPar[13]}), .a ({key_s3[10], key_s2[10], key_s1[10], key_s0[10]}), .c ({new_AGEMA_signal_1578, new_AGEMA_signal_1577, new_AGEMA_signal_1576, keyFF_inputPar[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_11_U1 ( .s (reset), .b ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, new_AGEMA_signal_1579, keyFF_outputPar[14]}), .a ({key_s3[11], key_s2[11], key_s1[11], key_s0[11]}), .c ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, new_AGEMA_signal_1585, keyFF_inputPar[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_12_U1 ( .s (reset), .b ({new_AGEMA_signal_1590, new_AGEMA_signal_1589, new_AGEMA_signal_1588, keyFF_outputPar[15]}), .a ({key_s3[12], key_s2[12], key_s1[12], key_s0[12]}), .c ({new_AGEMA_signal_1596, new_AGEMA_signal_1595, new_AGEMA_signal_1594, keyFF_inputPar[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_13_U1 ( .s (reset), .b ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, new_AGEMA_signal_1597, keyFF_outputPar[16]}), .a ({key_s3[13], key_s2[13], key_s1[13], key_s0[13]}), .c ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, new_AGEMA_signal_1603, keyFF_inputPar[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_14_U1 ( .s (reset), .b ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, new_AGEMA_signal_1606, keyFF_outputPar[17]}), .a ({key_s3[14], key_s2[14], key_s1[14], key_s0[14]}), .c ({new_AGEMA_signal_1614, new_AGEMA_signal_1613, new_AGEMA_signal_1612, keyFF_inputPar[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_15_U1 ( .s (reset), .b ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, new_AGEMA_signal_1477, keyFF_counterAdd[0]}), .a ({key_s3[15], key_s2[15], key_s1[15], key_s0[15]}), .c ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, new_AGEMA_signal_2119, keyFF_inputPar[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_16_U1 ( .s (reset), .b ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, new_AGEMA_signal_2113, keyFF_counterAdd[1]}), .a ({key_s3[16], key_s2[16], key_s1[16], key_s0[16]}), .c ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, new_AGEMA_signal_2143, keyFF_inputPar[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_17_U1 ( .s (reset), .b ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, new_AGEMA_signal_1471, keyFF_counterAdd[2]}), .a ({key_s3[17], key_s2[17], key_s1[17], key_s0[17]}), .c ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, new_AGEMA_signal_2125, keyFF_inputPar[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_18_U1 ( .s (reset), .b ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, new_AGEMA_signal_1465, keyFF_counterAdd[3]}), .a ({key_s3[18], key_s2[18], key_s1[18], key_s0[18]}), .c ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, new_AGEMA_signal_2131, keyFF_inputPar[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_19_U1 ( .s (reset), .b ({new_AGEMA_signal_1461, new_AGEMA_signal_1460, new_AGEMA_signal_1459, keyFF_counterAdd[4]}), .a ({key_s3[19], key_s2[19], key_s1[19], key_s0[19]}), .c ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, new_AGEMA_signal_2137, keyFF_inputPar[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_20_U1 ( .s (reset), .b ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, new_AGEMA_signal_1615, keyFF_outputPar[23]}), .a ({key_s3[20], key_s2[20], key_s1[20], key_s0[20]}), .c ({new_AGEMA_signal_1623, new_AGEMA_signal_1622, new_AGEMA_signal_1621, keyFF_inputPar[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_21_U1 ( .s (reset), .b ({new_AGEMA_signal_1626, new_AGEMA_signal_1625, new_AGEMA_signal_1624, keyFF_outputPar[24]}), .a ({key_s3[21], key_s2[21], key_s1[21], key_s0[21]}), .c ({new_AGEMA_signal_1632, new_AGEMA_signal_1631, new_AGEMA_signal_1630, keyFF_inputPar[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_22_U1 ( .s (reset), .b ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, new_AGEMA_signal_1633, keyFF_outputPar[25]}), .a ({key_s3[22], key_s2[22], key_s1[22], key_s0[22]}), .c ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, new_AGEMA_signal_1639, keyFF_inputPar[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_23_U1 ( .s (reset), .b ({new_AGEMA_signal_1644, new_AGEMA_signal_1643, new_AGEMA_signal_1642, keyFF_outputPar[26]}), .a ({key_s3[23], key_s2[23], key_s1[23], key_s0[23]}), .c ({new_AGEMA_signal_1650, new_AGEMA_signal_1649, new_AGEMA_signal_1648, keyFF_inputPar[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_24_U1 ( .s (reset), .b ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, new_AGEMA_signal_1651, keyFF_outputPar[27]}), .a ({key_s3[24], key_s2[24], key_s1[24], key_s0[24]}), .c ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, new_AGEMA_signal_1657, keyFF_inputPar[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_25_U1 ( .s (reset), .b ({new_AGEMA_signal_1662, new_AGEMA_signal_1661, new_AGEMA_signal_1660, keyFF_outputPar[28]}), .a ({key_s3[25], key_s2[25], key_s1[25], key_s0[25]}), .c ({new_AGEMA_signal_1668, new_AGEMA_signal_1667, new_AGEMA_signal_1666, keyFF_inputPar[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_26_U1 ( .s (reset), .b ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, new_AGEMA_signal_1669, keyFF_outputPar[29]}), .a ({key_s3[26], key_s2[26], key_s1[26], key_s0[26]}), .c ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, new_AGEMA_signal_1675, keyFF_inputPar[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_27_U1 ( .s (reset), .b ({new_AGEMA_signal_1680, new_AGEMA_signal_1679, new_AGEMA_signal_1678, keyFF_outputPar[30]}), .a ({key_s3[27], key_s2[27], key_s1[27], key_s0[27]}), .c ({new_AGEMA_signal_1686, new_AGEMA_signal_1685, new_AGEMA_signal_1684, keyFF_inputPar[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_28_U1 ( .s (reset), .b ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, new_AGEMA_signal_1687, keyFF_outputPar[31]}), .a ({key_s3[28], key_s2[28], key_s1[28], key_s0[28]}), .c ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, new_AGEMA_signal_1693, keyFF_inputPar[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_29_U1 ( .s (reset), .b ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, new_AGEMA_signal_1696, keyFF_outputPar[32]}), .a ({key_s3[29], key_s2[29], key_s1[29], key_s0[29]}), .c ({new_AGEMA_signal_1704, new_AGEMA_signal_1703, new_AGEMA_signal_1702, keyFF_inputPar[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_30_U1 ( .s (reset), .b ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, new_AGEMA_signal_1705, keyFF_outputPar[33]}), .a ({key_s3[30], key_s2[30], key_s1[30], key_s0[30]}), .c ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, new_AGEMA_signal_1711, keyFF_inputPar[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_31_U1 ( .s (reset), .b ({new_AGEMA_signal_1716, new_AGEMA_signal_1715, new_AGEMA_signal_1714, keyFF_outputPar[34]}), .a ({key_s3[31], key_s2[31], key_s1[31], key_s0[31]}), .c ({new_AGEMA_signal_1722, new_AGEMA_signal_1721, new_AGEMA_signal_1720, keyFF_inputPar[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_32_U1 ( .s (reset), .b ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, new_AGEMA_signal_1723, keyFF_outputPar[35]}), .a ({key_s3[32], key_s2[32], key_s1[32], key_s0[32]}), .c ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, new_AGEMA_signal_1729, keyFF_inputPar[32]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_33_U1 ( .s (reset), .b ({new_AGEMA_signal_1734, new_AGEMA_signal_1733, new_AGEMA_signal_1732, keyFF_outputPar[36]}), .a ({key_s3[33], key_s2[33], key_s1[33], key_s0[33]}), .c ({new_AGEMA_signal_1740, new_AGEMA_signal_1739, new_AGEMA_signal_1738, keyFF_inputPar[33]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_34_U1 ( .s (reset), .b ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, new_AGEMA_signal_1741, keyFF_outputPar[37]}), .a ({key_s3[34], key_s2[34], key_s1[34], key_s0[34]}), .c ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, new_AGEMA_signal_1747, keyFF_inputPar[34]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_35_U1 ( .s (reset), .b ({new_AGEMA_signal_1752, new_AGEMA_signal_1751, new_AGEMA_signal_1750, keyFF_outputPar[38]}), .a ({key_s3[35], key_s2[35], key_s1[35], key_s0[35]}), .c ({new_AGEMA_signal_1758, new_AGEMA_signal_1757, new_AGEMA_signal_1756, keyFF_inputPar[35]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_36_U1 ( .s (reset), .b ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, new_AGEMA_signal_1759, keyFF_outputPar[39]}), .a ({key_s3[36], key_s2[36], key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, new_AGEMA_signal_1765, keyFF_inputPar[36]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_37_U1 ( .s (reset), .b ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, new_AGEMA_signal_1768, keyFF_outputPar[40]}), .a ({key_s3[37], key_s2[37], key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_1776, new_AGEMA_signal_1775, new_AGEMA_signal_1774, keyFF_inputPar[37]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_38_U1 ( .s (reset), .b ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, new_AGEMA_signal_1777, keyFF_outputPar[41]}), .a ({key_s3[38], key_s2[38], key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, new_AGEMA_signal_1783, keyFF_inputPar[38]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_39_U1 ( .s (reset), .b ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, new_AGEMA_signal_1786, keyFF_outputPar[42]}), .a ({key_s3[39], key_s2[39], key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_1794, new_AGEMA_signal_1793, new_AGEMA_signal_1792, keyFF_inputPar[39]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_40_U1 ( .s (reset), .b ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, new_AGEMA_signal_1795, keyFF_outputPar[43]}), .a ({key_s3[40], key_s2[40], key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, new_AGEMA_signal_1801, keyFF_inputPar[40]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_41_U1 ( .s (reset), .b ({new_AGEMA_signal_1806, new_AGEMA_signal_1805, new_AGEMA_signal_1804, keyFF_outputPar[44]}), .a ({key_s3[41], key_s2[41], key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_1812, new_AGEMA_signal_1811, new_AGEMA_signal_1810, keyFF_inputPar[41]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_42_U1 ( .s (reset), .b ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, new_AGEMA_signal_1813, keyFF_outputPar[45]}), .a ({key_s3[42], key_s2[42], key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, new_AGEMA_signal_1819, keyFF_inputPar[42]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_43_U1 ( .s (reset), .b ({new_AGEMA_signal_1824, new_AGEMA_signal_1823, new_AGEMA_signal_1822, keyFF_outputPar[46]}), .a ({key_s3[43], key_s2[43], key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_1830, new_AGEMA_signal_1829, new_AGEMA_signal_1828, keyFF_inputPar[43]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_44_U1 ( .s (reset), .b ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, new_AGEMA_signal_1831, keyFF_outputPar[47]}), .a ({key_s3[44], key_s2[44], key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, new_AGEMA_signal_1837, keyFF_inputPar[44]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_45_U1 ( .s (reset), .b ({new_AGEMA_signal_1842, new_AGEMA_signal_1841, new_AGEMA_signal_1840, keyFF_outputPar[48]}), .a ({key_s3[45], key_s2[45], key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_1848, new_AGEMA_signal_1847, new_AGEMA_signal_1846, keyFF_inputPar[45]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_46_U1 ( .s (reset), .b ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, new_AGEMA_signal_1849, keyFF_outputPar[49]}), .a ({key_s3[46], key_s2[46], key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, new_AGEMA_signal_1855, keyFF_inputPar[46]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_47_U1 ( .s (reset), .b ({new_AGEMA_signal_1860, new_AGEMA_signal_1859, new_AGEMA_signal_1858, keyFF_outputPar[50]}), .a ({key_s3[47], key_s2[47], key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_1866, new_AGEMA_signal_1865, new_AGEMA_signal_1864, keyFF_inputPar[47]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_48_U1 ( .s (reset), .b ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, new_AGEMA_signal_1867, keyFF_outputPar[51]}), .a ({key_s3[48], key_s2[48], key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, new_AGEMA_signal_1873, keyFF_inputPar[48]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_49_U1 ( .s (reset), .b ({new_AGEMA_signal_1878, new_AGEMA_signal_1877, new_AGEMA_signal_1876, keyFF_outputPar[52]}), .a ({key_s3[49], key_s2[49], key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_1884, new_AGEMA_signal_1883, new_AGEMA_signal_1882, keyFF_inputPar[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_50_U1 ( .s (reset), .b ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, new_AGEMA_signal_1885, keyFF_outputPar[53]}), .a ({key_s3[50], key_s2[50], key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, new_AGEMA_signal_1891, keyFF_inputPar[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_51_U1 ( .s (reset), .b ({new_AGEMA_signal_1896, new_AGEMA_signal_1895, new_AGEMA_signal_1894, keyFF_outputPar[54]}), .a ({key_s3[51], key_s2[51], key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_1902, new_AGEMA_signal_1901, new_AGEMA_signal_1900, keyFF_inputPar[51]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_52_U1 ( .s (reset), .b ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, new_AGEMA_signal_1903, keyFF_outputPar[55]}), .a ({key_s3[52], key_s2[52], key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, new_AGEMA_signal_1909, keyFF_inputPar[52]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_53_U1 ( .s (reset), .b ({new_AGEMA_signal_1914, new_AGEMA_signal_1913, new_AGEMA_signal_1912, keyFF_outputPar[56]}), .a ({key_s3[53], key_s2[53], key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_1920, new_AGEMA_signal_1919, new_AGEMA_signal_1918, keyFF_inputPar[53]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_54_U1 ( .s (reset), .b ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, new_AGEMA_signal_1921, keyFF_outputPar[57]}), .a ({key_s3[54], key_s2[54], key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, new_AGEMA_signal_1927, keyFF_inputPar[54]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_55_U1 ( .s (reset), .b ({new_AGEMA_signal_1932, new_AGEMA_signal_1931, new_AGEMA_signal_1930, keyFF_outputPar[58]}), .a ({key_s3[55], key_s2[55], key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_1938, new_AGEMA_signal_1937, new_AGEMA_signal_1936, keyFF_inputPar[55]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_56_U1 ( .s (reset), .b ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, new_AGEMA_signal_1939, keyFF_outputPar[59]}), .a ({key_s3[56], key_s2[56], key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, new_AGEMA_signal_1945, keyFF_inputPar[56]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_57_U1 ( .s (reset), .b ({new_AGEMA_signal_1950, new_AGEMA_signal_1949, new_AGEMA_signal_1948, keyFF_outputPar[60]}), .a ({key_s3[57], key_s2[57], key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_1956, new_AGEMA_signal_1955, new_AGEMA_signal_1954, keyFF_inputPar[57]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_58_U1 ( .s (reset), .b ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, new_AGEMA_signal_1957, keyFF_outputPar[61]}), .a ({key_s3[58], key_s2[58], key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, new_AGEMA_signal_1963, keyFF_inputPar[58]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_59_U1 ( .s (reset), .b ({new_AGEMA_signal_1968, new_AGEMA_signal_1967, new_AGEMA_signal_1966, keyFF_outputPar[62]}), .a ({key_s3[59], key_s2[59], key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_1974, new_AGEMA_signal_1973, new_AGEMA_signal_1972, keyFF_inputPar[59]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_60_U1 ( .s (reset), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, new_AGEMA_signal_1975, keyFF_outputPar[63]}), .a ({key_s3[60], key_s2[60], key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, new_AGEMA_signal_1981, keyFF_inputPar[60]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_61_U1 ( .s (reset), .b ({new_AGEMA_signal_1986, new_AGEMA_signal_1985, new_AGEMA_signal_1984, keyFF_outputPar[64]}), .a ({key_s3[61], key_s2[61], key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_1992, new_AGEMA_signal_1991, new_AGEMA_signal_1990, keyFF_inputPar[61]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_62_U1 ( .s (reset), .b ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, new_AGEMA_signal_1993, keyFF_outputPar[65]}), .a ({key_s3[62], key_s2[62], key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, new_AGEMA_signal_1999, keyFF_inputPar[62]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_63_U1 ( .s (reset), .b ({new_AGEMA_signal_2004, new_AGEMA_signal_2003, new_AGEMA_signal_2002, keyFF_outputPar[66]}), .a ({key_s3[63], key_s2[63], key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_2010, new_AGEMA_signal_2009, new_AGEMA_signal_2008, keyFF_inputPar[63]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_64_U1 ( .s (reset), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, new_AGEMA_signal_2011, keyFF_outputPar[67]}), .a ({key_s3[64], key_s2[64], key_s1[64], key_s0[64]}), .c ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, new_AGEMA_signal_2017, keyFF_inputPar[64]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_65_U1 ( .s (reset), .b ({new_AGEMA_signal_2022, new_AGEMA_signal_2021, new_AGEMA_signal_2020, keyFF_outputPar[68]}), .a ({key_s3[65], key_s2[65], key_s1[65], key_s0[65]}), .c ({new_AGEMA_signal_2028, new_AGEMA_signal_2027, new_AGEMA_signal_2026, keyFF_inputPar[65]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_66_U1 ( .s (reset), .b ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, new_AGEMA_signal_2029, keyFF_outputPar[69]}), .a ({key_s3[66], key_s2[66], key_s1[66], key_s0[66]}), .c ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, new_AGEMA_signal_2035, keyFF_inputPar[66]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_67_U1 ( .s (reset), .b ({new_AGEMA_signal_2040, new_AGEMA_signal_2039, new_AGEMA_signal_2038, keyFF_outputPar[70]}), .a ({key_s3[67], key_s2[67], key_s1[67], key_s0[67]}), .c ({new_AGEMA_signal_2046, new_AGEMA_signal_2045, new_AGEMA_signal_2044, keyFF_inputPar[67]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_68_U1 ( .s (reset), .b ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, new_AGEMA_signal_2047, keyFF_outputPar[71]}), .a ({key_s3[68], key_s2[68], key_s1[68], key_s0[68]}), .c ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, new_AGEMA_signal_2053, keyFF_inputPar[68]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_69_U1 ( .s (reset), .b ({new_AGEMA_signal_2058, new_AGEMA_signal_2057, new_AGEMA_signal_2056, keyFF_outputPar[72]}), .a ({key_s3[69], key_s2[69], key_s1[69], key_s0[69]}), .c ({new_AGEMA_signal_2064, new_AGEMA_signal_2063, new_AGEMA_signal_2062, keyFF_inputPar[69]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_70_U1 ( .s (reset), .b ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, new_AGEMA_signal_2065, keyFF_outputPar[73]}), .a ({key_s3[70], key_s2[70], key_s1[70], key_s0[70]}), .c ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, new_AGEMA_signal_2071, keyFF_inputPar[70]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_71_U1 ( .s (reset), .b ({new_AGEMA_signal_2076, new_AGEMA_signal_2075, new_AGEMA_signal_2074, keyFF_outputPar[74]}), .a ({key_s3[71], key_s2[71], key_s1[71], key_s0[71]}), .c ({new_AGEMA_signal_2082, new_AGEMA_signal_2081, new_AGEMA_signal_2080, keyFF_inputPar[71]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_72_U1 ( .s (reset), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, new_AGEMA_signal_2083, keyFF_outputPar[75]}), .a ({key_s3[72], key_s2[72], key_s1[72], key_s0[72]}), .c ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, new_AGEMA_signal_2089, keyFF_inputPar[72]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_73_U1 ( .s (reset), .b ({new_AGEMA_signal_858, new_AGEMA_signal_857, new_AGEMA_signal_856, roundkey[0]}), .a ({key_s3[73], key_s2[73], key_s1[73], key_s0[73]}), .c ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, new_AGEMA_signal_2095, keyFF_inputPar[73]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_74_U1 ( .s (reset), .b ({new_AGEMA_signal_867, new_AGEMA_signal_866, new_AGEMA_signal_865, roundkey[1]}), .a ({key_s3[74], key_s2[74], key_s1[74], key_s0[74]}), .c ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, new_AGEMA_signal_2101, keyFF_inputPar[74]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_75_U1 ( .s (reset), .b ({new_AGEMA_signal_876, new_AGEMA_signal_875, new_AGEMA_signal_874, roundkey[2]}), .a ({key_s3[75], key_s2[75], key_s1[75], key_s0[75]}), .c ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, new_AGEMA_signal_2107, keyFF_inputPar[75]}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sboxInst_U3 ( .a ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, new_AGEMA_signal_2173, sboxInst_L0}), .b ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, new_AGEMA_signal_2221, sboxInst_n1}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sboxInst_U2 ( .a ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, new_AGEMA_signal_2164, sboxIn[3]}), .b ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, new_AGEMA_signal_2167, sboxInst_n2}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sboxInst_U1 ( .a ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, new_AGEMA_signal_2152, sboxIn[1]}), .b ({new_AGEMA_signal_2172, new_AGEMA_signal_2171, new_AGEMA_signal_2170, sboxInst_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_XOR1_U1 ( .a ({new_AGEMA_signal_2160, new_AGEMA_signal_2159, new_AGEMA_signal_2158, sboxIn[2]}), .b ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, new_AGEMA_signal_2152, sboxIn[1]}), .c ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, new_AGEMA_signal_2173, sboxInst_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_XOR2_U1 ( .a ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, new_AGEMA_signal_2152, sboxIn[1]}), .b ({new_AGEMA_signal_2148, new_AGEMA_signal_2147, new_AGEMA_signal_2146, sboxIn[0]}), .c ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, new_AGEMA_signal_2176, sboxInst_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_XOR3_U1 ( .a ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, new_AGEMA_signal_2176, sboxInst_L1}), .b ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, new_AGEMA_signal_2164, sboxIn[3]}), .c ({new_AGEMA_signal_2226, new_AGEMA_signal_2225, new_AGEMA_signal_2224, sboxInst_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_XOR4_U1 ( .a ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, new_AGEMA_signal_2164, sboxIn[3]}), .b ({new_AGEMA_signal_2148, new_AGEMA_signal_2147, new_AGEMA_signal_2146, sboxIn[0]}), .c ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, new_AGEMA_signal_2179, sboxInst_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_XOR5_U1 ( .a ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, new_AGEMA_signal_2179, sboxInst_L3}), .b ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, new_AGEMA_signal_2173, sboxInst_L0}), .c ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, new_AGEMA_signal_2227, sboxInst_Q3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_XOR6_U1 ( .a ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, new_AGEMA_signal_2164, sboxIn[3]}), .b ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, new_AGEMA_signal_2152, sboxIn[1]}), .c ({new_AGEMA_signal_2184, new_AGEMA_signal_2183, new_AGEMA_signal_2182, sboxInst_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_XOR9_U1 ( .a ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, new_AGEMA_signal_2176, sboxInst_L1}), .b ({new_AGEMA_signal_2160, new_AGEMA_signal_2159, new_AGEMA_signal_2158, sboxIn[2]}), .c ({new_AGEMA_signal_2232, new_AGEMA_signal_2231, new_AGEMA_signal_2230, sboxInst_Q7}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_sboxin_mux_inst_0_U1 ( .s (selSbox), .b ({new_AGEMA_signal_864, new_AGEMA_signal_863, new_AGEMA_signal_862, stateXORroundkey[0]}), .a ({new_AGEMA_signal_885, new_AGEMA_signal_884, new_AGEMA_signal_883, roundkey[3]}), .c ({new_AGEMA_signal_2148, new_AGEMA_signal_2147, new_AGEMA_signal_2146, sboxIn[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_sboxin_mux_inst_1_U1 ( .s (selSbox), .b ({new_AGEMA_signal_873, new_AGEMA_signal_872, new_AGEMA_signal_871, stateXORroundkey[1]}), .a ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, new_AGEMA_signal_2149, keyRegKS[1]}), .c ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, new_AGEMA_signal_2152, sboxIn[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_sboxin_mux_inst_2_U1 ( .s (selSbox), .b ({new_AGEMA_signal_882, new_AGEMA_signal_881, new_AGEMA_signal_880, stateXORroundkey[2]}), .a ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, new_AGEMA_signal_2155, keyRegKS[2]}), .c ({new_AGEMA_signal_2160, new_AGEMA_signal_2159, new_AGEMA_signal_2158, sboxIn[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_sboxin_mux_inst_3_U1 ( .s (selSbox), .b ({new_AGEMA_signal_891, new_AGEMA_signal_890, new_AGEMA_signal_889, stateXORroundkey[3]}), .a ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, new_AGEMA_signal_2161, keyRegKS[3]}), .c ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, new_AGEMA_signal_2164, sboxIn[3]}) ) ;
    ClockGatingController #(5) ClockGatingInst ( .clk (clk), .rst (reset), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_2628, new_AGEMA_signal_2627, new_AGEMA_signal_2626, serialIn[0]}), .a ({new_AGEMA_signal_900, new_AGEMA_signal_899, new_AGEMA_signal_898, stateFF_inputPar[0]}), .c ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, new_AGEMA_signal_2629, stateFF_state_gff_1_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_2058, new_AGEMA_signal_2057, new_AGEMA_signal_2056, keyFF_outputPar[72]}), .a ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, new_AGEMA_signal_2617, keyFF_inputPar[76]}), .c ({new_AGEMA_signal_2634, new_AGEMA_signal_2633, new_AGEMA_signal_2632, keyFF_keystate_gff_20_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_76_U1 ( .s (reset), .b ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, new_AGEMA_signal_2239, sboxOut[0]}), .a ({key_s3[76], key_s2[76], key_s1[76], key_s0[76]}), .c ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, new_AGEMA_signal_2617, keyFF_inputPar[76]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_XOR16_U1 ( .a ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, new_AGEMA_signal_2236, sboxInst_T0}), .b ({new_AGEMA_signal_2226, new_AGEMA_signal_2225, new_AGEMA_signal_2224, sboxInst_L2}), .c ({new_AGEMA_signal_2622, new_AGEMA_signal_2621, new_AGEMA_signal_2620, sboxInst_Q2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_XOR7_U1 ( .a ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, new_AGEMA_signal_2236, sboxInst_T0}), .b ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, new_AGEMA_signal_2233, sboxInst_T2}), .c ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, new_AGEMA_signal_2623, sboxInst_L5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_XOR8_U1 ( .a ({new_AGEMA_signal_2184, new_AGEMA_signal_2183, new_AGEMA_signal_2182, sboxInst_L4}), .b ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, new_AGEMA_signal_2623, sboxInst_L5}), .c ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, new_AGEMA_signal_2635, sboxInst_Q6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_AND1_U1 ( .a ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, new_AGEMA_signal_2221, sboxInst_n1}), .b ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, new_AGEMA_signal_2167, sboxInst_n2}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, new_AGEMA_signal_2236, sboxInst_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_AND3_U1 ( .a ({new_AGEMA_signal_2172, new_AGEMA_signal_2171, new_AGEMA_signal_2170, sboxInst_n3}), .b ({new_AGEMA_signal_2160, new_AGEMA_signal_2159, new_AGEMA_signal_2158, sboxIn[2]}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, new_AGEMA_signal_2233, sboxInst_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_XOR15_U1 ( .a ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, new_AGEMA_signal_2179, sboxInst_L3}), .b ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, new_AGEMA_signal_2233, sboxInst_T2}), .c ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, new_AGEMA_signal_2239, sboxOut[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_serialIn_mux_inst_0_U1 ( .s (intDone), .b ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, new_AGEMA_signal_2239, sboxOut[0]}), .a ({new_AGEMA_signal_864, new_AGEMA_signal_863, new_AGEMA_signal_862, stateXORroundkey[0]}), .c ({new_AGEMA_signal_2628, new_AGEMA_signal_2627, new_AGEMA_signal_2626, serialIn[0]}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, new_AGEMA_signal_2671, serialIn[1]}), .a ({new_AGEMA_signal_909, new_AGEMA_signal_908, new_AGEMA_signal_907, stateFF_inputPar[1]}), .c ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, new_AGEMA_signal_2677, stateFF_state_gff_1_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, new_AGEMA_signal_2674, serialIn[2]}), .a ({new_AGEMA_signal_918, new_AGEMA_signal_917, new_AGEMA_signal_916, stateFF_inputPar[2]}), .c ({new_AGEMA_signal_2682, new_AGEMA_signal_2681, new_AGEMA_signal_2680, stateFF_state_gff_1_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, new_AGEMA_signal_2695, serialIn[3]}), .a ({new_AGEMA_signal_927, new_AGEMA_signal_926, new_AGEMA_signal_925, stateFF_inputPar[3]}), .c ({new_AGEMA_signal_2700, new_AGEMA_signal_2699, new_AGEMA_signal_2698, stateFF_state_gff_1_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, new_AGEMA_signal_2065, keyFF_outputPar[73]}), .a ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, new_AGEMA_signal_2659, keyFF_inputPar[77]}), .c ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, new_AGEMA_signal_2683, keyFF_keystate_gff_20_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_2076, new_AGEMA_signal_2075, new_AGEMA_signal_2074, keyFF_outputPar[74]}), .a ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, new_AGEMA_signal_2665, keyFF_inputPar[78]}), .c ({new_AGEMA_signal_2688, new_AGEMA_signal_2687, new_AGEMA_signal_2686, keyFF_keystate_gff_20_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, new_AGEMA_signal_2083, keyFF_outputPar[75]}), .a ({new_AGEMA_signal_2694, new_AGEMA_signal_2693, new_AGEMA_signal_2692, keyFF_inputPar[79]}), .c ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, new_AGEMA_signal_2701, keyFF_keystate_gff_20_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_77_U1 ( .s (reset), .b ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, new_AGEMA_signal_2653, sboxOut[1]}), .a ({key_s3[77], key_s2[77], key_s1[77], key_s0[77]}), .c ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, new_AGEMA_signal_2659, keyFF_inputPar[77]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_78_U1 ( .s (reset), .b ({new_AGEMA_signal_2652, new_AGEMA_signal_2651, new_AGEMA_signal_2650, sboxOut[2]}), .a ({key_s3[78], key_s2[78], key_s1[78], key_s0[78]}), .c ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, new_AGEMA_signal_2665, keyFF_inputPar[78]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_79_U1 ( .s (reset), .b ({new_AGEMA_signal_2670, new_AGEMA_signal_2669, new_AGEMA_signal_2668, sboxOut[3]}), .a ({key_s3[79], key_s2[79], key_s1[79], key_s0[79]}), .c ({new_AGEMA_signal_2694, new_AGEMA_signal_2693, new_AGEMA_signal_2692, keyFF_inputPar[79]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_AND2_U1 ( .a ({new_AGEMA_signal_2622, new_AGEMA_signal_2621, new_AGEMA_signal_2620, sboxInst_Q2}), .b ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, new_AGEMA_signal_2227, sboxInst_Q3}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_2640, new_AGEMA_signal_2639, new_AGEMA_signal_2638, sboxInst_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_AND4_U1 ( .a ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, new_AGEMA_signal_2635, sboxInst_Q6}), .b ({new_AGEMA_signal_2232, new_AGEMA_signal_2231, new_AGEMA_signal_2230, sboxInst_Q7}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, new_AGEMA_signal_2641, sboxInst_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_XOR10_U1 ( .a ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, new_AGEMA_signal_2623, sboxInst_L5}), .b ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, new_AGEMA_signal_2641, sboxInst_T3}), .c ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, new_AGEMA_signal_2647, sboxInst_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_XOR11_U1 ( .a ({new_AGEMA_signal_2148, new_AGEMA_signal_2147, new_AGEMA_signal_2146, sboxIn[0]}), .b ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, new_AGEMA_signal_2647, sboxInst_L7}), .c ({new_AGEMA_signal_2670, new_AGEMA_signal_2669, new_AGEMA_signal_2668, sboxOut[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_XOR12_U1 ( .a ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, new_AGEMA_signal_2623, sboxInst_L5}), .b ({new_AGEMA_signal_2640, new_AGEMA_signal_2639, new_AGEMA_signal_2638, sboxInst_T1}), .c ({new_AGEMA_signal_2646, new_AGEMA_signal_2645, new_AGEMA_signal_2644, sboxInst_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_XOR13_U1 ( .a ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, new_AGEMA_signal_2176, sboxInst_L1}), .b ({new_AGEMA_signal_2646, new_AGEMA_signal_2645, new_AGEMA_signal_2644, sboxInst_L8}), .c ({new_AGEMA_signal_2652, new_AGEMA_signal_2651, new_AGEMA_signal_2650, sboxOut[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sboxInst_XOR14_U1 ( .a ({new_AGEMA_signal_2184, new_AGEMA_signal_2183, new_AGEMA_signal_2182, sboxInst_L4}), .b ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, new_AGEMA_signal_2641, sboxInst_T3}), .c ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, new_AGEMA_signal_2653, sboxOut[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_serialIn_mux_inst_1_U1 ( .s (intDone), .b ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, new_AGEMA_signal_2653, sboxOut[1]}), .a ({new_AGEMA_signal_873, new_AGEMA_signal_872, new_AGEMA_signal_871, stateXORroundkey[1]}), .c ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, new_AGEMA_signal_2671, serialIn[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_serialIn_mux_inst_2_U1 ( .s (intDone), .b ({new_AGEMA_signal_2652, new_AGEMA_signal_2651, new_AGEMA_signal_2650, sboxOut[2]}), .a ({new_AGEMA_signal_882, new_AGEMA_signal_881, new_AGEMA_signal_880, stateXORroundkey[2]}), .c ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, new_AGEMA_signal_2674, serialIn[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_serialIn_mux_inst_3_U1 ( .s (intDone), .b ({new_AGEMA_signal_2670, new_AGEMA_signal_2669, new_AGEMA_signal_2668, sboxOut[3]}), .a ({new_AGEMA_signal_891, new_AGEMA_signal_890, new_AGEMA_signal_889, stateXORroundkey[3]}), .c ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, new_AGEMA_signal_2695, serialIn[3]}) ) ;

    /* register cells */
    DFF_X1 fsm_cnt_rnd_count_reg_reg_4__FF_FF ( .CK (clk_gated), .D (fsm_cnt_rnd_n14), .Q (counter[4]), .QN () ) ;
    DFF_X1 fsm_cnt_rnd_count_reg_reg_2__FF_FF ( .CK (clk_gated), .D (fsm_cnt_rnd_n16), .Q (counter[2]), .QN () ) ;
    DFF_X1 fsm_cnt_rnd_count_reg_reg_0__FF_FF ( .CK (clk_gated), .D (fsm_cnt_rnd_n18), .Q (counter[0]), .QN () ) ;
    DFF_X1 fsm_cnt_rnd_count_reg_reg_3__FF_FF ( .CK (clk_gated), .D (fsm_cnt_rnd_n1), .Q (counter[3]), .QN () ) ;
    DFF_X1 fsm_cnt_rnd_count_reg_reg_1__FF_FF ( .CK (clk_gated), .D (fsm_cnt_rnd_n41), .Q (fsm_cnt_rnd_n24), .QN () ) ;
    DFF_X1 fsm_cnt_ser_count_reg_reg_2__FF_FF ( .CK (clk_gated), .D (fsm_cnt_ser_n1), .Q (fsm_countSerial[2]), .QN () ) ;
    DFF_X1 fsm_cnt_ser_count_reg_reg_0__FF_FF ( .CK (clk_gated), .D (fsm_cnt_ser_n3), .Q (fsm_countSerial[0]), .QN () ) ;
    DFF_X1 fsm_cnt_ser_count_reg_reg_3__FF_FF ( .CK (clk_gated), .D (fsm_cnt_ser_n26), .Q (fsm_countSerial[3]), .QN () ) ;
    DFF_X1 fsm_cnt_ser_count_reg_reg_1__FF_FF ( .CK (clk_gated), .D (fsm_cnt_ser_n28), .Q (fsm_countSerial[1]), .QN () ) ;
    DFF_X1 fsm_ps_state_reg_0__FF_FF ( .CK (clk_gated), .D (fsm_n21), .Q (fsm_ps_state_0_), .QN () ) ;
    DFF_X1 fsm_ps_state_reg_1__FF_FF ( .CK (clk_gated), .D (fsm_n20), .Q (fsm_ps_state_1_), .QN () ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_1_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, new_AGEMA_signal_2629, stateFF_state_gff_1_s_next_state[0]}), .Q ({data_out_s3[0], data_out_s2[0], data_out_s1[0], data_out_s0[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_1_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2682, new_AGEMA_signal_2681, new_AGEMA_signal_2680, stateFF_state_gff_1_s_next_state[2]}), .Q ({data_out_s3[2], data_out_s2[2], data_out_s1[2], data_out_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_1_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, new_AGEMA_signal_2677, stateFF_state_gff_1_s_next_state[1]}), .Q ({data_out_s3[1], data_out_s2[1], data_out_s1[1], data_out_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_1_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2700, new_AGEMA_signal_2699, new_AGEMA_signal_2698, stateFF_state_gff_1_s_next_state[3]}), .Q ({data_out_s3[3], data_out_s2[3], data_out_s1[3], data_out_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_2_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2196, new_AGEMA_signal_2195, new_AGEMA_signal_2194, stateFF_state_gff_2_s_next_state[3]}), .Q ({data_out_s3[7], data_out_s2[7], data_out_s1[7], data_out_s0[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_2_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, new_AGEMA_signal_2191, stateFF_state_gff_2_s_next_state[2]}), .Q ({data_out_s3[6], data_out_s2[6], data_out_s1[6], data_out_s0[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_2_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, new_AGEMA_signal_2188, stateFF_state_gff_2_s_next_state[1]}), .Q ({data_out_s3[5], data_out_s2[5], data_out_s1[5], data_out_s0[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_2_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, new_AGEMA_signal_2185, stateFF_state_gff_2_s_next_state[0]}), .Q ({data_out_s3[4], data_out_s2[4], data_out_s1[4], data_out_s0[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_3_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, new_AGEMA_signal_2251, stateFF_state_gff_3_s_next_state[3]}), .Q ({data_out_s3[11], data_out_s2[11], data_out_s1[11], data_out_s0[11]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_3_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, new_AGEMA_signal_2248, stateFF_state_gff_3_s_next_state[2]}), .Q ({data_out_s3[10], data_out_s2[10], data_out_s1[10], data_out_s0[10]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_3_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, new_AGEMA_signal_2245, stateFF_state_gff_3_s_next_state[1]}), .Q ({data_out_s3[9], data_out_s2[9], data_out_s1[9], data_out_s0[9]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_3_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2244, new_AGEMA_signal_2243, new_AGEMA_signal_2242, stateFF_state_gff_3_s_next_state[0]}), .Q ({data_out_s3[8], data_out_s2[8], data_out_s1[8], data_out_s0[8]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_4_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, new_AGEMA_signal_2263, stateFF_state_gff_4_s_next_state[3]}), .Q ({data_out_s3[15], data_out_s2[15], data_out_s1[15], data_out_s0[15]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_4_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, new_AGEMA_signal_2260, stateFF_state_gff_4_s_next_state[2]}), .Q ({data_out_s3[14], data_out_s2[14], data_out_s1[14], data_out_s0[14]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_4_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, new_AGEMA_signal_2257, stateFF_state_gff_4_s_next_state[1]}), .Q ({data_out_s3[13], data_out_s2[13], data_out_s1[13], data_out_s0[13]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_4_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2256, new_AGEMA_signal_2255, new_AGEMA_signal_2254, stateFF_state_gff_4_s_next_state[0]}), .Q ({data_out_s3[12], data_out_s2[12], data_out_s1[12], data_out_s0[12]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_5_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, new_AGEMA_signal_2275, stateFF_state_gff_5_s_next_state[3]}), .Q ({data_out_s3[19], data_out_s2[19], data_out_s1[19], data_out_s0[19]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_5_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, new_AGEMA_signal_2272, stateFF_state_gff_5_s_next_state[2]}), .Q ({data_out_s3[18], data_out_s2[18], data_out_s1[18], data_out_s0[18]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_5_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, new_AGEMA_signal_2269, stateFF_state_gff_5_s_next_state[1]}), .Q ({data_out_s3[17], data_out_s2[17], data_out_s1[17], data_out_s0[17]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_5_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2268, new_AGEMA_signal_2267, new_AGEMA_signal_2266, stateFF_state_gff_5_s_next_state[0]}), .Q ({data_out_s3[16], data_out_s2[16], data_out_s1[16], data_out_s0[16]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_6_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, new_AGEMA_signal_2287, stateFF_state_gff_6_s_next_state[3]}), .Q ({data_out_s3[23], data_out_s2[23], data_out_s1[23], data_out_s0[23]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_6_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2286, new_AGEMA_signal_2285, new_AGEMA_signal_2284, stateFF_state_gff_6_s_next_state[2]}), .Q ({data_out_s3[22], data_out_s2[22], data_out_s1[22], data_out_s0[22]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_6_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, new_AGEMA_signal_2281, stateFF_state_gff_6_s_next_state[1]}), .Q ({data_out_s3[21], data_out_s2[21], data_out_s1[21], data_out_s0[21]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_6_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2280, new_AGEMA_signal_2279, new_AGEMA_signal_2278, stateFF_state_gff_6_s_next_state[0]}), .Q ({data_out_s3[20], data_out_s2[20], data_out_s1[20], data_out_s0[20]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_7_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, new_AGEMA_signal_2299, stateFF_state_gff_7_s_next_state[3]}), .Q ({data_out_s3[27], data_out_s2[27], data_out_s1[27], data_out_s0[27]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_7_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2298, new_AGEMA_signal_2297, new_AGEMA_signal_2296, stateFF_state_gff_7_s_next_state[2]}), .Q ({data_out_s3[26], data_out_s2[26], data_out_s1[26], data_out_s0[26]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_7_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, new_AGEMA_signal_2293, stateFF_state_gff_7_s_next_state[1]}), .Q ({data_out_s3[25], data_out_s2[25], data_out_s1[25], data_out_s0[25]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_7_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2292, new_AGEMA_signal_2291, new_AGEMA_signal_2290, stateFF_state_gff_7_s_next_state[0]}), .Q ({data_out_s3[24], data_out_s2[24], data_out_s1[24], data_out_s0[24]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_8_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, new_AGEMA_signal_2311, stateFF_state_gff_8_s_next_state[3]}), .Q ({data_out_s3[31], data_out_s2[31], data_out_s1[31], data_out_s0[31]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_8_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2310, new_AGEMA_signal_2309, new_AGEMA_signal_2308, stateFF_state_gff_8_s_next_state[2]}), .Q ({data_out_s3[30], data_out_s2[30], data_out_s1[30], data_out_s0[30]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_8_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, new_AGEMA_signal_2305, stateFF_state_gff_8_s_next_state[1]}), .Q ({data_out_s3[29], data_out_s2[29], data_out_s1[29], data_out_s0[29]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_8_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2304, new_AGEMA_signal_2303, new_AGEMA_signal_2302, stateFF_state_gff_8_s_next_state[0]}), .Q ({data_out_s3[28], data_out_s2[28], data_out_s1[28], data_out_s0[28]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_9_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, new_AGEMA_signal_2323, stateFF_state_gff_9_s_next_state[3]}), .Q ({data_out_s3[35], data_out_s2[35], data_out_s1[35], data_out_s0[35]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_9_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2322, new_AGEMA_signal_2321, new_AGEMA_signal_2320, stateFF_state_gff_9_s_next_state[2]}), .Q ({data_out_s3[34], data_out_s2[34], data_out_s1[34], data_out_s0[34]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_9_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, new_AGEMA_signal_2317, stateFF_state_gff_9_s_next_state[1]}), .Q ({data_out_s3[33], data_out_s2[33], data_out_s1[33], data_out_s0[33]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_9_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2316, new_AGEMA_signal_2315, new_AGEMA_signal_2314, stateFF_state_gff_9_s_next_state[0]}), .Q ({data_out_s3[32], data_out_s2[32], data_out_s1[32], data_out_s0[32]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_10_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, new_AGEMA_signal_2335, stateFF_state_gff_10_s_next_state[3]}), .Q ({data_out_s3[39], data_out_s2[39], data_out_s1[39], data_out_s0[39]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_10_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2334, new_AGEMA_signal_2333, new_AGEMA_signal_2332, stateFF_state_gff_10_s_next_state[2]}), .Q ({data_out_s3[38], data_out_s2[38], data_out_s1[38], data_out_s0[38]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_10_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, new_AGEMA_signal_2329, stateFF_state_gff_10_s_next_state[1]}), .Q ({data_out_s3[37], data_out_s2[37], data_out_s1[37], data_out_s0[37]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_10_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2328, new_AGEMA_signal_2327, new_AGEMA_signal_2326, stateFF_state_gff_10_s_next_state[0]}), .Q ({data_out_s3[36], data_out_s2[36], data_out_s1[36], data_out_s0[36]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_11_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, new_AGEMA_signal_2347, stateFF_state_gff_11_s_next_state[3]}), .Q ({data_out_s3[43], data_out_s2[43], data_out_s1[43], data_out_s0[43]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_11_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, new_AGEMA_signal_2344, stateFF_state_gff_11_s_next_state[2]}), .Q ({data_out_s3[42], data_out_s2[42], data_out_s1[42], data_out_s0[42]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_11_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, new_AGEMA_signal_2341, stateFF_state_gff_11_s_next_state[1]}), .Q ({data_out_s3[41], data_out_s2[41], data_out_s1[41], data_out_s0[41]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_11_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2340, new_AGEMA_signal_2339, new_AGEMA_signal_2338, stateFF_state_gff_11_s_next_state[0]}), .Q ({data_out_s3[40], data_out_s2[40], data_out_s1[40], data_out_s0[40]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_12_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, new_AGEMA_signal_2359, stateFF_state_gff_12_s_next_state[3]}), .Q ({data_out_s3[47], data_out_s2[47], data_out_s1[47], data_out_s0[47]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_12_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2358, new_AGEMA_signal_2357, new_AGEMA_signal_2356, stateFF_state_gff_12_s_next_state[2]}), .Q ({data_out_s3[46], data_out_s2[46], data_out_s1[46], data_out_s0[46]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_12_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, new_AGEMA_signal_2353, stateFF_state_gff_12_s_next_state[1]}), .Q ({data_out_s3[45], data_out_s2[45], data_out_s1[45], data_out_s0[45]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_12_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2352, new_AGEMA_signal_2351, new_AGEMA_signal_2350, stateFF_state_gff_12_s_next_state[0]}), .Q ({data_out_s3[44], data_out_s2[44], data_out_s1[44], data_out_s0[44]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_13_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, new_AGEMA_signal_2371, stateFF_state_gff_13_s_next_state[3]}), .Q ({data_out_s3[51], data_out_s2[51], data_out_s1[51], data_out_s0[51]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_13_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, new_AGEMA_signal_2368, stateFF_state_gff_13_s_next_state[2]}), .Q ({data_out_s3[50], data_out_s2[50], data_out_s1[50], data_out_s0[50]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_13_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, new_AGEMA_signal_2365, stateFF_state_gff_13_s_next_state[1]}), .Q ({data_out_s3[49], data_out_s2[49], data_out_s1[49], data_out_s0[49]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_13_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2364, new_AGEMA_signal_2363, new_AGEMA_signal_2362, stateFF_state_gff_13_s_next_state[0]}), .Q ({data_out_s3[48], data_out_s2[48], data_out_s1[48], data_out_s0[48]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_14_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, new_AGEMA_signal_2383, stateFF_state_gff_14_s_next_state[3]}), .Q ({data_out_s3[55], data_out_s2[55], data_out_s1[55], data_out_s0[55]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_14_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, new_AGEMA_signal_2380, stateFF_state_gff_14_s_next_state[2]}), .Q ({data_out_s3[54], data_out_s2[54], data_out_s1[54], data_out_s0[54]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_14_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, new_AGEMA_signal_2377, stateFF_state_gff_14_s_next_state[1]}), .Q ({data_out_s3[53], data_out_s2[53], data_out_s1[53], data_out_s0[53]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_14_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2376, new_AGEMA_signal_2375, new_AGEMA_signal_2374, stateFF_state_gff_14_s_next_state[0]}), .Q ({data_out_s3[52], data_out_s2[52], data_out_s1[52], data_out_s0[52]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_15_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, new_AGEMA_signal_2395, stateFF_state_gff_15_s_next_state[3]}), .Q ({data_out_s3[59], data_out_s2[59], data_out_s1[59], data_out_s0[59]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_15_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2394, new_AGEMA_signal_2393, new_AGEMA_signal_2392, stateFF_state_gff_15_s_next_state[2]}), .Q ({data_out_s3[58], data_out_s2[58], data_out_s1[58], data_out_s0[58]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_15_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, new_AGEMA_signal_2389, stateFF_state_gff_15_s_next_state[1]}), .Q ({data_out_s3[57], data_out_s2[57], data_out_s1[57], data_out_s0[57]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_15_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2388, new_AGEMA_signal_2387, new_AGEMA_signal_2386, stateFF_state_gff_15_s_next_state[0]}), .Q ({data_out_s3[56], data_out_s2[56], data_out_s1[56], data_out_s0[56]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_16_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, new_AGEMA_signal_2407, stateFF_state_gff_16_s_next_state[3]}), .Q ({data_out_s3[63], data_out_s2[63], data_out_s1[63], data_out_s0[63]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_16_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, new_AGEMA_signal_2404, stateFF_state_gff_16_s_next_state[2]}), .Q ({data_out_s3[62], data_out_s2[62], data_out_s1[62], data_out_s0[62]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_16_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, new_AGEMA_signal_2401, stateFF_state_gff_16_s_next_state[1]}), .Q ({data_out_s3[61], data_out_s2[61], data_out_s1[61], data_out_s0[61]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) stateFF_state_gff_16_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2400, new_AGEMA_signal_2399, new_AGEMA_signal_2398, stateFF_state_gff_16_s_next_state[0]}), .Q ({data_out_s3[60], data_out_s2[60], data_out_s1[60], data_out_s0[60]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_1_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, new_AGEMA_signal_2419, keyFF_keystate_gff_1_s_next_state[3]}), .Q ({new_AGEMA_signal_1482, new_AGEMA_signal_1481, new_AGEMA_signal_1480, keyFF_outputPar[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_1_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2418, new_AGEMA_signal_2417, new_AGEMA_signal_2416, keyFF_keystate_gff_1_s_next_state[2]}), .Q ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, new_AGEMA_signal_2161, keyRegKS[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_1_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, new_AGEMA_signal_2413, keyFF_keystate_gff_1_s_next_state[1]}), .Q ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, new_AGEMA_signal_2155, keyRegKS[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_1_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2412, new_AGEMA_signal_2411, new_AGEMA_signal_2410, keyFF_keystate_gff_1_s_next_state[0]}), .Q ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, new_AGEMA_signal_2149, keyRegKS[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_2_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, new_AGEMA_signal_2431, keyFF_keystate_gff_2_s_next_state[3]}), .Q ({new_AGEMA_signal_1518, new_AGEMA_signal_1517, new_AGEMA_signal_1516, keyFF_outputPar[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_2_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2430, new_AGEMA_signal_2429, new_AGEMA_signal_2428, keyFF_keystate_gff_2_s_next_state[2]}), .Q ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, new_AGEMA_signal_1507, keyFF_outputPar[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_2_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, new_AGEMA_signal_2425, keyFF_keystate_gff_2_s_next_state[1]}), .Q ({new_AGEMA_signal_1500, new_AGEMA_signal_1499, new_AGEMA_signal_1498, keyFF_outputPar[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_2_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, new_AGEMA_signal_2422, keyFF_keystate_gff_2_s_next_state[0]}), .Q ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, new_AGEMA_signal_1489, keyFF_outputPar[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_3_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, new_AGEMA_signal_2443, keyFF_keystate_gff_3_s_next_state[3]}), .Q ({new_AGEMA_signal_1554, new_AGEMA_signal_1553, new_AGEMA_signal_1552, keyFF_outputPar[11]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_3_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2442, new_AGEMA_signal_2441, new_AGEMA_signal_2440, keyFF_keystate_gff_3_s_next_state[2]}), .Q ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, new_AGEMA_signal_1543, keyFF_outputPar[10]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_3_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, new_AGEMA_signal_2437, keyFF_keystate_gff_3_s_next_state[1]}), .Q ({new_AGEMA_signal_1536, new_AGEMA_signal_1535, new_AGEMA_signal_1534, keyFF_outputPar[9]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_3_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, new_AGEMA_signal_2434, keyFF_keystate_gff_3_s_next_state[0]}), .Q ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, new_AGEMA_signal_1525, keyFF_outputPar[8]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_4_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, new_AGEMA_signal_2455, keyFF_keystate_gff_4_s_next_state[3]}), .Q ({new_AGEMA_signal_1590, new_AGEMA_signal_1589, new_AGEMA_signal_1588, keyFF_outputPar[15]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_4_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2454, new_AGEMA_signal_2453, new_AGEMA_signal_2452, keyFF_keystate_gff_4_s_next_state[2]}), .Q ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, new_AGEMA_signal_1579, keyFF_outputPar[14]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_4_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, new_AGEMA_signal_2449, keyFF_keystate_gff_4_s_next_state[1]}), .Q ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, new_AGEMA_signal_1570, keyFF_outputPar[13]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_4_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2448, new_AGEMA_signal_2447, new_AGEMA_signal_2446, keyFF_keystate_gff_4_s_next_state[0]}), .Q ({new_AGEMA_signal_1563, new_AGEMA_signal_1562, new_AGEMA_signal_1561, keyFF_outputPar[12]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_5_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2208, new_AGEMA_signal_2207, new_AGEMA_signal_2206, keyFF_keystate_gff_5_s_next_state[3]}), .Q ({new_AGEMA_signal_2112, new_AGEMA_signal_2111, new_AGEMA_signal_2110, keyFF_outputPar[19]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_5_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, new_AGEMA_signal_2203, keyFF_keystate_gff_5_s_next_state[2]}), .Q ({new_AGEMA_signal_1476, new_AGEMA_signal_1475, new_AGEMA_signal_1474, keyFF_outputPar[18]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_5_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, new_AGEMA_signal_2200, keyFF_keystate_gff_5_s_next_state[1]}), .Q ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, new_AGEMA_signal_1606, keyFF_outputPar[17]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_5_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, new_AGEMA_signal_2197, keyFF_keystate_gff_5_s_next_state[0]}), .Q ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, new_AGEMA_signal_1597, keyFF_outputPar[16]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_6_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2220, new_AGEMA_signal_2219, new_AGEMA_signal_2218, keyFF_keystate_gff_6_s_next_state[3]}), .Q ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, new_AGEMA_signal_1615, keyFF_outputPar[23]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_6_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, new_AGEMA_signal_2215, keyFF_keystate_gff_6_s_next_state[2]}), .Q ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, new_AGEMA_signal_1456, keyFF_outputPar[22]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_6_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, new_AGEMA_signal_2212, keyFF_keystate_gff_6_s_next_state[1]}), .Q ({new_AGEMA_signal_1464, new_AGEMA_signal_1463, new_AGEMA_signal_1462, keyFF_outputPar[21]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_6_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, new_AGEMA_signal_2209, keyFF_keystate_gff_6_s_next_state[0]}), .Q ({new_AGEMA_signal_1470, new_AGEMA_signal_1469, new_AGEMA_signal_1468, keyFF_outputPar[20]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_7_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, new_AGEMA_signal_2467, keyFF_keystate_gff_7_s_next_state[3]}), .Q ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, new_AGEMA_signal_1651, keyFF_outputPar[27]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_7_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2466, new_AGEMA_signal_2465, new_AGEMA_signal_2464, keyFF_keystate_gff_7_s_next_state[2]}), .Q ({new_AGEMA_signal_1644, new_AGEMA_signal_1643, new_AGEMA_signal_1642, keyFF_outputPar[26]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_7_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, new_AGEMA_signal_2461, keyFF_keystate_gff_7_s_next_state[1]}), .Q ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, new_AGEMA_signal_1633, keyFF_outputPar[25]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_7_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2460, new_AGEMA_signal_2459, new_AGEMA_signal_2458, keyFF_keystate_gff_7_s_next_state[0]}), .Q ({new_AGEMA_signal_1626, new_AGEMA_signal_1625, new_AGEMA_signal_1624, keyFF_outputPar[24]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_8_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, new_AGEMA_signal_2479, keyFF_keystate_gff_8_s_next_state[3]}), .Q ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, new_AGEMA_signal_1687, keyFF_outputPar[31]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_8_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2478, new_AGEMA_signal_2477, new_AGEMA_signal_2476, keyFF_keystate_gff_8_s_next_state[2]}), .Q ({new_AGEMA_signal_1680, new_AGEMA_signal_1679, new_AGEMA_signal_1678, keyFF_outputPar[30]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_8_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, new_AGEMA_signal_2473, keyFF_keystate_gff_8_s_next_state[1]}), .Q ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, new_AGEMA_signal_1669, keyFF_outputPar[29]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_8_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2472, new_AGEMA_signal_2471, new_AGEMA_signal_2470, keyFF_keystate_gff_8_s_next_state[0]}), .Q ({new_AGEMA_signal_1662, new_AGEMA_signal_1661, new_AGEMA_signal_1660, keyFF_outputPar[28]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_9_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, new_AGEMA_signal_2491, keyFF_keystate_gff_9_s_next_state[3]}), .Q ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, new_AGEMA_signal_1723, keyFF_outputPar[35]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_9_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2490, new_AGEMA_signal_2489, new_AGEMA_signal_2488, keyFF_keystate_gff_9_s_next_state[2]}), .Q ({new_AGEMA_signal_1716, new_AGEMA_signal_1715, new_AGEMA_signal_1714, keyFF_outputPar[34]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_9_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, new_AGEMA_signal_2485, keyFF_keystate_gff_9_s_next_state[1]}), .Q ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, new_AGEMA_signal_1705, keyFF_outputPar[33]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_9_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2484, new_AGEMA_signal_2483, new_AGEMA_signal_2482, keyFF_keystate_gff_9_s_next_state[0]}), .Q ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, new_AGEMA_signal_1696, keyFF_outputPar[32]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_10_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, new_AGEMA_signal_2503, keyFF_keystate_gff_10_s_next_state[3]}), .Q ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, new_AGEMA_signal_1759, keyFF_outputPar[39]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_10_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2502, new_AGEMA_signal_2501, new_AGEMA_signal_2500, keyFF_keystate_gff_10_s_next_state[2]}), .Q ({new_AGEMA_signal_1752, new_AGEMA_signal_1751, new_AGEMA_signal_1750, keyFF_outputPar[38]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_10_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, new_AGEMA_signal_2497, keyFF_keystate_gff_10_s_next_state[1]}), .Q ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, new_AGEMA_signal_1741, keyFF_outputPar[37]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_10_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2496, new_AGEMA_signal_2495, new_AGEMA_signal_2494, keyFF_keystate_gff_10_s_next_state[0]}), .Q ({new_AGEMA_signal_1734, new_AGEMA_signal_1733, new_AGEMA_signal_1732, keyFF_outputPar[36]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_11_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, new_AGEMA_signal_2515, keyFF_keystate_gff_11_s_next_state[3]}), .Q ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, new_AGEMA_signal_1795, keyFF_outputPar[43]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_11_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2514, new_AGEMA_signal_2513, new_AGEMA_signal_2512, keyFF_keystate_gff_11_s_next_state[2]}), .Q ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, new_AGEMA_signal_1786, keyFF_outputPar[42]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_11_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, new_AGEMA_signal_2509, keyFF_keystate_gff_11_s_next_state[1]}), .Q ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, new_AGEMA_signal_1777, keyFF_outputPar[41]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_11_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2508, new_AGEMA_signal_2507, new_AGEMA_signal_2506, keyFF_keystate_gff_11_s_next_state[0]}), .Q ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, new_AGEMA_signal_1768, keyFF_outputPar[40]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_12_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, new_AGEMA_signal_2527, keyFF_keystate_gff_12_s_next_state[3]}), .Q ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, new_AGEMA_signal_1831, keyFF_outputPar[47]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_12_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2526, new_AGEMA_signal_2525, new_AGEMA_signal_2524, keyFF_keystate_gff_12_s_next_state[2]}), .Q ({new_AGEMA_signal_1824, new_AGEMA_signal_1823, new_AGEMA_signal_1822, keyFF_outputPar[46]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_12_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, new_AGEMA_signal_2521, keyFF_keystate_gff_12_s_next_state[1]}), .Q ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, new_AGEMA_signal_1813, keyFF_outputPar[45]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_12_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2520, new_AGEMA_signal_2519, new_AGEMA_signal_2518, keyFF_keystate_gff_12_s_next_state[0]}), .Q ({new_AGEMA_signal_1806, new_AGEMA_signal_1805, new_AGEMA_signal_1804, keyFF_outputPar[44]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_13_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, new_AGEMA_signal_2539, keyFF_keystate_gff_13_s_next_state[3]}), .Q ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, new_AGEMA_signal_1867, keyFF_outputPar[51]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_13_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2538, new_AGEMA_signal_2537, new_AGEMA_signal_2536, keyFF_keystate_gff_13_s_next_state[2]}), .Q ({new_AGEMA_signal_1860, new_AGEMA_signal_1859, new_AGEMA_signal_1858, keyFF_outputPar[50]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_13_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, new_AGEMA_signal_2533, keyFF_keystate_gff_13_s_next_state[1]}), .Q ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, new_AGEMA_signal_1849, keyFF_outputPar[49]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_13_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2532, new_AGEMA_signal_2531, new_AGEMA_signal_2530, keyFF_keystate_gff_13_s_next_state[0]}), .Q ({new_AGEMA_signal_1842, new_AGEMA_signal_1841, new_AGEMA_signal_1840, keyFF_outputPar[48]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_14_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, new_AGEMA_signal_2551, keyFF_keystate_gff_14_s_next_state[3]}), .Q ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, new_AGEMA_signal_1903, keyFF_outputPar[55]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_14_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2550, new_AGEMA_signal_2549, new_AGEMA_signal_2548, keyFF_keystate_gff_14_s_next_state[2]}), .Q ({new_AGEMA_signal_1896, new_AGEMA_signal_1895, new_AGEMA_signal_1894, keyFF_outputPar[54]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_14_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, new_AGEMA_signal_2545, keyFF_keystate_gff_14_s_next_state[1]}), .Q ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, new_AGEMA_signal_1885, keyFF_outputPar[53]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_14_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2544, new_AGEMA_signal_2543, new_AGEMA_signal_2542, keyFF_keystate_gff_14_s_next_state[0]}), .Q ({new_AGEMA_signal_1878, new_AGEMA_signal_1877, new_AGEMA_signal_1876, keyFF_outputPar[52]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_15_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, new_AGEMA_signal_2563, keyFF_keystate_gff_15_s_next_state[3]}), .Q ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, new_AGEMA_signal_1939, keyFF_outputPar[59]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_15_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2562, new_AGEMA_signal_2561, new_AGEMA_signal_2560, keyFF_keystate_gff_15_s_next_state[2]}), .Q ({new_AGEMA_signal_1932, new_AGEMA_signal_1931, new_AGEMA_signal_1930, keyFF_outputPar[58]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_15_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, new_AGEMA_signal_2557, keyFF_keystate_gff_15_s_next_state[1]}), .Q ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, new_AGEMA_signal_1921, keyFF_outputPar[57]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_15_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2556, new_AGEMA_signal_2555, new_AGEMA_signal_2554, keyFF_keystate_gff_15_s_next_state[0]}), .Q ({new_AGEMA_signal_1914, new_AGEMA_signal_1913, new_AGEMA_signal_1912, keyFF_outputPar[56]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_16_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, new_AGEMA_signal_2575, keyFF_keystate_gff_16_s_next_state[3]}), .Q ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, new_AGEMA_signal_1975, keyFF_outputPar[63]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_16_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2574, new_AGEMA_signal_2573, new_AGEMA_signal_2572, keyFF_keystate_gff_16_s_next_state[2]}), .Q ({new_AGEMA_signal_1968, new_AGEMA_signal_1967, new_AGEMA_signal_1966, keyFF_outputPar[62]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_16_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, new_AGEMA_signal_2569, keyFF_keystate_gff_16_s_next_state[1]}), .Q ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, new_AGEMA_signal_1957, keyFF_outputPar[61]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_16_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2568, new_AGEMA_signal_2567, new_AGEMA_signal_2566, keyFF_keystate_gff_16_s_next_state[0]}), .Q ({new_AGEMA_signal_1950, new_AGEMA_signal_1949, new_AGEMA_signal_1948, keyFF_outputPar[60]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_17_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, new_AGEMA_signal_2587, keyFF_keystate_gff_17_s_next_state[3]}), .Q ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, new_AGEMA_signal_2011, keyFF_outputPar[67]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_17_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2586, new_AGEMA_signal_2585, new_AGEMA_signal_2584, keyFF_keystate_gff_17_s_next_state[2]}), .Q ({new_AGEMA_signal_2004, new_AGEMA_signal_2003, new_AGEMA_signal_2002, keyFF_outputPar[66]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_17_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, new_AGEMA_signal_2581, keyFF_keystate_gff_17_s_next_state[1]}), .Q ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, new_AGEMA_signal_1993, keyFF_outputPar[65]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_17_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2580, new_AGEMA_signal_2579, new_AGEMA_signal_2578, keyFF_keystate_gff_17_s_next_state[0]}), .Q ({new_AGEMA_signal_1986, new_AGEMA_signal_1985, new_AGEMA_signal_1984, keyFF_outputPar[64]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_18_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, new_AGEMA_signal_2599, keyFF_keystate_gff_18_s_next_state[3]}), .Q ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, new_AGEMA_signal_2047, keyFF_outputPar[71]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_18_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2598, new_AGEMA_signal_2597, new_AGEMA_signal_2596, keyFF_keystate_gff_18_s_next_state[2]}), .Q ({new_AGEMA_signal_2040, new_AGEMA_signal_2039, new_AGEMA_signal_2038, keyFF_outputPar[70]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_18_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, new_AGEMA_signal_2593, keyFF_keystate_gff_18_s_next_state[1]}), .Q ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, new_AGEMA_signal_2029, keyFF_outputPar[69]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_18_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2592, new_AGEMA_signal_2591, new_AGEMA_signal_2590, keyFF_keystate_gff_18_s_next_state[0]}), .Q ({new_AGEMA_signal_2022, new_AGEMA_signal_2021, new_AGEMA_signal_2020, keyFF_outputPar[68]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_19_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, new_AGEMA_signal_2611, keyFF_keystate_gff_19_s_next_state[3]}), .Q ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, new_AGEMA_signal_2083, keyFF_outputPar[75]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_19_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2610, new_AGEMA_signal_2609, new_AGEMA_signal_2608, keyFF_keystate_gff_19_s_next_state[2]}), .Q ({new_AGEMA_signal_2076, new_AGEMA_signal_2075, new_AGEMA_signal_2074, keyFF_outputPar[74]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_19_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, new_AGEMA_signal_2605, keyFF_keystate_gff_19_s_next_state[1]}), .Q ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, new_AGEMA_signal_2065, keyFF_outputPar[73]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_19_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2604, new_AGEMA_signal_2603, new_AGEMA_signal_2602, keyFF_keystate_gff_19_s_next_state[0]}), .Q ({new_AGEMA_signal_2058, new_AGEMA_signal_2057, new_AGEMA_signal_2056, keyFF_outputPar[72]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_20_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, new_AGEMA_signal_2701, keyFF_keystate_gff_20_s_next_state[3]}), .Q ({new_AGEMA_signal_885, new_AGEMA_signal_884, new_AGEMA_signal_883, roundkey[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_20_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2688, new_AGEMA_signal_2687, new_AGEMA_signal_2686, keyFF_keystate_gff_20_s_next_state[2]}), .Q ({new_AGEMA_signal_876, new_AGEMA_signal_875, new_AGEMA_signal_874, roundkey[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_20_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, new_AGEMA_signal_2683, keyFF_keystate_gff_20_s_next_state[1]}), .Q ({new_AGEMA_signal_867, new_AGEMA_signal_866, new_AGEMA_signal_865, roundkey[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) keyFF_keystate_gff_20_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2634, new_AGEMA_signal_2633, new_AGEMA_signal_2632, keyFF_keystate_gff_20_s_next_state[0]}), .Q ({new_AGEMA_signal_858, new_AGEMA_signal_857, new_AGEMA_signal_856, roundkey[0]}) ) ;
endmodule
