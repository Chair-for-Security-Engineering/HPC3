////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module LED in file /AGEMA/Designs/LED_round-based/AGEMA/LED.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module LED_HPC2_Pipeline_d2 (IN_plaintext_s0, IN_key_s0, IN_reset, CLK, IN_key_s1, IN_key_s2, IN_plaintext_s1, IN_plaintext_s2, Fresh, OUT_ciphertext_s0, OUT_done, OUT_ciphertext_s1, OUT_ciphertext_s2);
    input [63:0] IN_plaintext_s0 ;
    input [127:0] IN_key_s0 ;
    input IN_reset ;
    input CLK ;
    input [127:0] IN_key_s1 ;
    input [127:0] IN_key_s2 ;
    input [63:0] IN_plaintext_s1 ;
    input [63:0] IN_plaintext_s2 ;
    input [191:0] Fresh ;
    output [63:0] OUT_ciphertext_s0 ;
    output OUT_done ;
    output [63:0] OUT_ciphertext_s1 ;
    output [63:0] OUT_ciphertext_s2 ;
    wire n15 ;
    wire n14 ;
    wire n16 ;
    wire n17 ;
    wire n18 ;
    wire n19 ;
    wire n20 ;
    wire LED_128_Instance_n34 ;
    wire LED_128_Instance_n33 ;
    wire LED_128_Instance_n32 ;
    wire LED_128_Instance_n23 ;
    wire LED_128_Instance_n21 ;
    wire LED_128_Instance_n20 ;
    wire LED_128_Instance_n19 ;
    wire LED_128_Instance_n18 ;
    wire LED_128_Instance_n17 ;
    wire LED_128_Instance_n16 ;
    wire LED_128_Instance_n15 ;
    wire LED_128_Instance_n14 ;
    wire LED_128_Instance_n13 ;
    wire LED_128_Instance_n12 ;
    wire LED_128_Instance_n11 ;
    wire LED_128_Instance_n10 ;
    wire LED_128_Instance_n2 ;
    wire LED_128_Instance_n1 ;
    wire LED_128_Instance_n27 ;
    wire LED_128_Instance_N9 ;
    wire LED_128_Instance_n28 ;
    wire LED_128_Instance_N8 ;
    wire LED_128_Instance_n30 ;
    wire LED_128_Instance_N7 ;
    wire LED_128_Instance_n5 ;
    wire LED_128_Instance_N6 ;
    wire LED_128_Instance_n29 ;
    wire LED_128_Instance_N5 ;
    wire LED_128_Instance_n6 ;
    wire LED_128_Instance_N4 ;
    wire LED_128_Instance_n24 ;
    wire LED_128_Instance_N13 ;
    wire LED_128_Instance_n25 ;
    wire LED_128_Instance_N12 ;
    wire LED_128_Instance_n8 ;
    wire LED_128_Instance_n26 ;
    wire LED_128_Instance_N11 ;
    wire LED_128_Instance_n4 ;
    wire LED_128_Instance_N10 ;
    wire LED_128_Instance_n31 ;
    wire LED_128_Instance_addroundkey_out_0_ ;
    wire LED_128_Instance_addroundkey_out_1_ ;
    wire LED_128_Instance_addroundkey_out_2_ ;
    wire LED_128_Instance_addroundkey_out_3_ ;
    wire LED_128_Instance_addroundkey_out_4_ ;
    wire LED_128_Instance_addroundkey_out_5_ ;
    wire LED_128_Instance_addroundkey_out_6_ ;
    wire LED_128_Instance_addroundkey_out_16_ ;
    wire LED_128_Instance_addroundkey_out_17_ ;
    wire LED_128_Instance_addroundkey_out_18_ ;
    wire LED_128_Instance_addroundkey_out_19_ ;
    wire LED_128_Instance_addroundkey_out_20_ ;
    wire LED_128_Instance_addroundkey_out_21_ ;
    wire LED_128_Instance_addroundkey_out_22_ ;
    wire LED_128_Instance_addroundkey_out_32_ ;
    wire LED_128_Instance_addroundkey_out_33_ ;
    wire LED_128_Instance_addroundkey_out_34_ ;
    wire LED_128_Instance_addroundkey_out_35_ ;
    wire LED_128_Instance_addroundkey_out_36_ ;
    wire LED_128_Instance_addroundkey_out_37_ ;
    wire LED_128_Instance_addroundkey_out_38_ ;
    wire LED_128_Instance_addroundkey_out_48_ ;
    wire LED_128_Instance_addroundkey_out_49_ ;
    wire LED_128_Instance_addroundkey_out_50_ ;
    wire LED_128_Instance_addroundkey_out_51_ ;
    wire LED_128_Instance_addroundkey_out_52_ ;
    wire LED_128_Instance_addroundkey_out_53_ ;
    wire LED_128_Instance_addroundkey_out_54_ ;
    wire LED_128_Instance_n22 ;
    wire LED_128_Instance_MUX_state0_n11 ;
    wire LED_128_Instance_MUX_state0_n10 ;
    wire LED_128_Instance_MUX_state0_n9 ;
    wire LED_128_Instance_MUX_state0_n8 ;
    wire LED_128_Instance_MUX_current_roundkey_n10 ;
    wire LED_128_Instance_MUX_current_roundkey_n9 ;
    wire LED_128_Instance_MUX_current_roundkey_n8 ;
    wire LED_128_Instance_MUX_current_roundkey_n7 ;
    wire LED_128_Instance_MUX_addroundkey_out_n9 ;
    wire LED_128_Instance_MUX_addroundkey_out_n8 ;
    wire LED_128_Instance_MUX_addroundkey_out_n7 ;
    wire LED_128_Instance_SBox_Instance_0_n3 ;
    wire LED_128_Instance_SBox_Instance_0_n2 ;
    wire LED_128_Instance_SBox_Instance_0_n1 ;
    wire LED_128_Instance_SBox_Instance_0_L8 ;
    wire LED_128_Instance_SBox_Instance_0_L7 ;
    wire LED_128_Instance_SBox_Instance_0_T3 ;
    wire LED_128_Instance_SBox_Instance_0_T1 ;
    wire LED_128_Instance_SBox_Instance_0_Q7 ;
    wire LED_128_Instance_SBox_Instance_0_Q6 ;
    wire LED_128_Instance_SBox_Instance_0_L5 ;
    wire LED_128_Instance_SBox_Instance_0_T2 ;
    wire LED_128_Instance_SBox_Instance_0_L4 ;
    wire LED_128_Instance_SBox_Instance_0_Q3 ;
    wire LED_128_Instance_SBox_Instance_0_L3 ;
    wire LED_128_Instance_SBox_Instance_0_Q2 ;
    wire LED_128_Instance_SBox_Instance_0_T0 ;
    wire LED_128_Instance_SBox_Instance_0_L2 ;
    wire LED_128_Instance_SBox_Instance_0_L1 ;
    wire LED_128_Instance_SBox_Instance_0_L0 ;
    wire LED_128_Instance_SBox_Instance_1_n3 ;
    wire LED_128_Instance_SBox_Instance_1_n2 ;
    wire LED_128_Instance_SBox_Instance_1_n1 ;
    wire LED_128_Instance_SBox_Instance_1_L8 ;
    wire LED_128_Instance_SBox_Instance_1_L7 ;
    wire LED_128_Instance_SBox_Instance_1_T3 ;
    wire LED_128_Instance_SBox_Instance_1_T1 ;
    wire LED_128_Instance_SBox_Instance_1_Q7 ;
    wire LED_128_Instance_SBox_Instance_1_Q6 ;
    wire LED_128_Instance_SBox_Instance_1_L5 ;
    wire LED_128_Instance_SBox_Instance_1_T2 ;
    wire LED_128_Instance_SBox_Instance_1_L4 ;
    wire LED_128_Instance_SBox_Instance_1_Q3 ;
    wire LED_128_Instance_SBox_Instance_1_L3 ;
    wire LED_128_Instance_SBox_Instance_1_Q2 ;
    wire LED_128_Instance_SBox_Instance_1_T0 ;
    wire LED_128_Instance_SBox_Instance_1_L2 ;
    wire LED_128_Instance_SBox_Instance_1_L1 ;
    wire LED_128_Instance_SBox_Instance_1_L0 ;
    wire LED_128_Instance_SBox_Instance_2_n3 ;
    wire LED_128_Instance_SBox_Instance_2_n2 ;
    wire LED_128_Instance_SBox_Instance_2_n1 ;
    wire LED_128_Instance_SBox_Instance_2_L8 ;
    wire LED_128_Instance_SBox_Instance_2_L7 ;
    wire LED_128_Instance_SBox_Instance_2_T3 ;
    wire LED_128_Instance_SBox_Instance_2_T1 ;
    wire LED_128_Instance_SBox_Instance_2_Q7 ;
    wire LED_128_Instance_SBox_Instance_2_Q6 ;
    wire LED_128_Instance_SBox_Instance_2_L5 ;
    wire LED_128_Instance_SBox_Instance_2_T2 ;
    wire LED_128_Instance_SBox_Instance_2_L4 ;
    wire LED_128_Instance_SBox_Instance_2_Q3 ;
    wire LED_128_Instance_SBox_Instance_2_L3 ;
    wire LED_128_Instance_SBox_Instance_2_Q2 ;
    wire LED_128_Instance_SBox_Instance_2_T0 ;
    wire LED_128_Instance_SBox_Instance_2_L2 ;
    wire LED_128_Instance_SBox_Instance_2_L1 ;
    wire LED_128_Instance_SBox_Instance_2_L0 ;
    wire LED_128_Instance_SBox_Instance_3_n3 ;
    wire LED_128_Instance_SBox_Instance_3_n2 ;
    wire LED_128_Instance_SBox_Instance_3_n1 ;
    wire LED_128_Instance_SBox_Instance_3_L8 ;
    wire LED_128_Instance_SBox_Instance_3_L7 ;
    wire LED_128_Instance_SBox_Instance_3_T3 ;
    wire LED_128_Instance_SBox_Instance_3_T1 ;
    wire LED_128_Instance_SBox_Instance_3_Q7 ;
    wire LED_128_Instance_SBox_Instance_3_Q6 ;
    wire LED_128_Instance_SBox_Instance_3_L5 ;
    wire LED_128_Instance_SBox_Instance_3_T2 ;
    wire LED_128_Instance_SBox_Instance_3_L4 ;
    wire LED_128_Instance_SBox_Instance_3_Q3 ;
    wire LED_128_Instance_SBox_Instance_3_L3 ;
    wire LED_128_Instance_SBox_Instance_3_Q2 ;
    wire LED_128_Instance_SBox_Instance_3_T0 ;
    wire LED_128_Instance_SBox_Instance_3_L2 ;
    wire LED_128_Instance_SBox_Instance_3_L1 ;
    wire LED_128_Instance_SBox_Instance_3_L0 ;
    wire LED_128_Instance_SBox_Instance_4_n3 ;
    wire LED_128_Instance_SBox_Instance_4_n2 ;
    wire LED_128_Instance_SBox_Instance_4_n1 ;
    wire LED_128_Instance_SBox_Instance_4_L8 ;
    wire LED_128_Instance_SBox_Instance_4_L7 ;
    wire LED_128_Instance_SBox_Instance_4_T3 ;
    wire LED_128_Instance_SBox_Instance_4_T1 ;
    wire LED_128_Instance_SBox_Instance_4_Q7 ;
    wire LED_128_Instance_SBox_Instance_4_Q6 ;
    wire LED_128_Instance_SBox_Instance_4_L5 ;
    wire LED_128_Instance_SBox_Instance_4_T2 ;
    wire LED_128_Instance_SBox_Instance_4_L4 ;
    wire LED_128_Instance_SBox_Instance_4_Q3 ;
    wire LED_128_Instance_SBox_Instance_4_L3 ;
    wire LED_128_Instance_SBox_Instance_4_Q2 ;
    wire LED_128_Instance_SBox_Instance_4_T0 ;
    wire LED_128_Instance_SBox_Instance_4_L2 ;
    wire LED_128_Instance_SBox_Instance_4_L1 ;
    wire LED_128_Instance_SBox_Instance_4_L0 ;
    wire LED_128_Instance_SBox_Instance_5_n3 ;
    wire LED_128_Instance_SBox_Instance_5_n2 ;
    wire LED_128_Instance_SBox_Instance_5_n1 ;
    wire LED_128_Instance_SBox_Instance_5_L8 ;
    wire LED_128_Instance_SBox_Instance_5_L7 ;
    wire LED_128_Instance_SBox_Instance_5_T3 ;
    wire LED_128_Instance_SBox_Instance_5_T1 ;
    wire LED_128_Instance_SBox_Instance_5_Q7 ;
    wire LED_128_Instance_SBox_Instance_5_Q6 ;
    wire LED_128_Instance_SBox_Instance_5_L5 ;
    wire LED_128_Instance_SBox_Instance_5_T2 ;
    wire LED_128_Instance_SBox_Instance_5_L4 ;
    wire LED_128_Instance_SBox_Instance_5_Q3 ;
    wire LED_128_Instance_SBox_Instance_5_L3 ;
    wire LED_128_Instance_SBox_Instance_5_Q2 ;
    wire LED_128_Instance_SBox_Instance_5_T0 ;
    wire LED_128_Instance_SBox_Instance_5_L2 ;
    wire LED_128_Instance_SBox_Instance_5_L1 ;
    wire LED_128_Instance_SBox_Instance_5_L0 ;
    wire LED_128_Instance_SBox_Instance_6_n3 ;
    wire LED_128_Instance_SBox_Instance_6_n2 ;
    wire LED_128_Instance_SBox_Instance_6_n1 ;
    wire LED_128_Instance_SBox_Instance_6_L8 ;
    wire LED_128_Instance_SBox_Instance_6_L7 ;
    wire LED_128_Instance_SBox_Instance_6_T3 ;
    wire LED_128_Instance_SBox_Instance_6_T1 ;
    wire LED_128_Instance_SBox_Instance_6_Q7 ;
    wire LED_128_Instance_SBox_Instance_6_Q6 ;
    wire LED_128_Instance_SBox_Instance_6_L5 ;
    wire LED_128_Instance_SBox_Instance_6_T2 ;
    wire LED_128_Instance_SBox_Instance_6_L4 ;
    wire LED_128_Instance_SBox_Instance_6_Q3 ;
    wire LED_128_Instance_SBox_Instance_6_L3 ;
    wire LED_128_Instance_SBox_Instance_6_Q2 ;
    wire LED_128_Instance_SBox_Instance_6_T0 ;
    wire LED_128_Instance_SBox_Instance_6_L2 ;
    wire LED_128_Instance_SBox_Instance_6_L1 ;
    wire LED_128_Instance_SBox_Instance_6_L0 ;
    wire LED_128_Instance_SBox_Instance_7_n3 ;
    wire LED_128_Instance_SBox_Instance_7_n2 ;
    wire LED_128_Instance_SBox_Instance_7_n1 ;
    wire LED_128_Instance_SBox_Instance_7_L8 ;
    wire LED_128_Instance_SBox_Instance_7_L7 ;
    wire LED_128_Instance_SBox_Instance_7_T3 ;
    wire LED_128_Instance_SBox_Instance_7_T1 ;
    wire LED_128_Instance_SBox_Instance_7_Q7 ;
    wire LED_128_Instance_SBox_Instance_7_Q6 ;
    wire LED_128_Instance_SBox_Instance_7_L5 ;
    wire LED_128_Instance_SBox_Instance_7_T2 ;
    wire LED_128_Instance_SBox_Instance_7_L4 ;
    wire LED_128_Instance_SBox_Instance_7_Q3 ;
    wire LED_128_Instance_SBox_Instance_7_L3 ;
    wire LED_128_Instance_SBox_Instance_7_Q2 ;
    wire LED_128_Instance_SBox_Instance_7_T0 ;
    wire LED_128_Instance_SBox_Instance_7_L2 ;
    wire LED_128_Instance_SBox_Instance_7_L1 ;
    wire LED_128_Instance_SBox_Instance_7_L0 ;
    wire LED_128_Instance_SBox_Instance_8_n3 ;
    wire LED_128_Instance_SBox_Instance_8_n2 ;
    wire LED_128_Instance_SBox_Instance_8_n1 ;
    wire LED_128_Instance_SBox_Instance_8_L8 ;
    wire LED_128_Instance_SBox_Instance_8_L7 ;
    wire LED_128_Instance_SBox_Instance_8_T3 ;
    wire LED_128_Instance_SBox_Instance_8_T1 ;
    wire LED_128_Instance_SBox_Instance_8_Q7 ;
    wire LED_128_Instance_SBox_Instance_8_Q6 ;
    wire LED_128_Instance_SBox_Instance_8_L5 ;
    wire LED_128_Instance_SBox_Instance_8_T2 ;
    wire LED_128_Instance_SBox_Instance_8_L4 ;
    wire LED_128_Instance_SBox_Instance_8_Q3 ;
    wire LED_128_Instance_SBox_Instance_8_L3 ;
    wire LED_128_Instance_SBox_Instance_8_Q2 ;
    wire LED_128_Instance_SBox_Instance_8_T0 ;
    wire LED_128_Instance_SBox_Instance_8_L2 ;
    wire LED_128_Instance_SBox_Instance_8_L1 ;
    wire LED_128_Instance_SBox_Instance_8_L0 ;
    wire LED_128_Instance_SBox_Instance_9_n3 ;
    wire LED_128_Instance_SBox_Instance_9_n2 ;
    wire LED_128_Instance_SBox_Instance_9_n1 ;
    wire LED_128_Instance_SBox_Instance_9_L8 ;
    wire LED_128_Instance_SBox_Instance_9_L7 ;
    wire LED_128_Instance_SBox_Instance_9_T3 ;
    wire LED_128_Instance_SBox_Instance_9_T1 ;
    wire LED_128_Instance_SBox_Instance_9_Q7 ;
    wire LED_128_Instance_SBox_Instance_9_Q6 ;
    wire LED_128_Instance_SBox_Instance_9_L5 ;
    wire LED_128_Instance_SBox_Instance_9_T2 ;
    wire LED_128_Instance_SBox_Instance_9_L4 ;
    wire LED_128_Instance_SBox_Instance_9_Q3 ;
    wire LED_128_Instance_SBox_Instance_9_L3 ;
    wire LED_128_Instance_SBox_Instance_9_Q2 ;
    wire LED_128_Instance_SBox_Instance_9_T0 ;
    wire LED_128_Instance_SBox_Instance_9_L2 ;
    wire LED_128_Instance_SBox_Instance_9_L1 ;
    wire LED_128_Instance_SBox_Instance_9_L0 ;
    wire LED_128_Instance_SBox_Instance_10_n3 ;
    wire LED_128_Instance_SBox_Instance_10_n2 ;
    wire LED_128_Instance_SBox_Instance_10_n1 ;
    wire LED_128_Instance_SBox_Instance_10_L8 ;
    wire LED_128_Instance_SBox_Instance_10_L7 ;
    wire LED_128_Instance_SBox_Instance_10_T3 ;
    wire LED_128_Instance_SBox_Instance_10_T1 ;
    wire LED_128_Instance_SBox_Instance_10_Q7 ;
    wire LED_128_Instance_SBox_Instance_10_Q6 ;
    wire LED_128_Instance_SBox_Instance_10_L5 ;
    wire LED_128_Instance_SBox_Instance_10_T2 ;
    wire LED_128_Instance_SBox_Instance_10_L4 ;
    wire LED_128_Instance_SBox_Instance_10_Q3 ;
    wire LED_128_Instance_SBox_Instance_10_L3 ;
    wire LED_128_Instance_SBox_Instance_10_Q2 ;
    wire LED_128_Instance_SBox_Instance_10_T0 ;
    wire LED_128_Instance_SBox_Instance_10_L2 ;
    wire LED_128_Instance_SBox_Instance_10_L1 ;
    wire LED_128_Instance_SBox_Instance_10_L0 ;
    wire LED_128_Instance_SBox_Instance_11_n3 ;
    wire LED_128_Instance_SBox_Instance_11_n2 ;
    wire LED_128_Instance_SBox_Instance_11_n1 ;
    wire LED_128_Instance_SBox_Instance_11_L8 ;
    wire LED_128_Instance_SBox_Instance_11_L7 ;
    wire LED_128_Instance_SBox_Instance_11_T3 ;
    wire LED_128_Instance_SBox_Instance_11_T1 ;
    wire LED_128_Instance_SBox_Instance_11_Q7 ;
    wire LED_128_Instance_SBox_Instance_11_Q6 ;
    wire LED_128_Instance_SBox_Instance_11_L5 ;
    wire LED_128_Instance_SBox_Instance_11_T2 ;
    wire LED_128_Instance_SBox_Instance_11_L4 ;
    wire LED_128_Instance_SBox_Instance_11_Q3 ;
    wire LED_128_Instance_SBox_Instance_11_L3 ;
    wire LED_128_Instance_SBox_Instance_11_Q2 ;
    wire LED_128_Instance_SBox_Instance_11_T0 ;
    wire LED_128_Instance_SBox_Instance_11_L2 ;
    wire LED_128_Instance_SBox_Instance_11_L1 ;
    wire LED_128_Instance_SBox_Instance_11_L0 ;
    wire LED_128_Instance_SBox_Instance_12_n3 ;
    wire LED_128_Instance_SBox_Instance_12_n2 ;
    wire LED_128_Instance_SBox_Instance_12_n1 ;
    wire LED_128_Instance_SBox_Instance_12_L8 ;
    wire LED_128_Instance_SBox_Instance_12_L7 ;
    wire LED_128_Instance_SBox_Instance_12_T3 ;
    wire LED_128_Instance_SBox_Instance_12_T1 ;
    wire LED_128_Instance_SBox_Instance_12_Q7 ;
    wire LED_128_Instance_SBox_Instance_12_Q6 ;
    wire LED_128_Instance_SBox_Instance_12_L5 ;
    wire LED_128_Instance_SBox_Instance_12_T2 ;
    wire LED_128_Instance_SBox_Instance_12_L4 ;
    wire LED_128_Instance_SBox_Instance_12_Q3 ;
    wire LED_128_Instance_SBox_Instance_12_L3 ;
    wire LED_128_Instance_SBox_Instance_12_Q2 ;
    wire LED_128_Instance_SBox_Instance_12_T0 ;
    wire LED_128_Instance_SBox_Instance_12_L2 ;
    wire LED_128_Instance_SBox_Instance_12_L1 ;
    wire LED_128_Instance_SBox_Instance_12_L0 ;
    wire LED_128_Instance_SBox_Instance_13_n3 ;
    wire LED_128_Instance_SBox_Instance_13_n2 ;
    wire LED_128_Instance_SBox_Instance_13_n1 ;
    wire LED_128_Instance_SBox_Instance_13_L8 ;
    wire LED_128_Instance_SBox_Instance_13_L7 ;
    wire LED_128_Instance_SBox_Instance_13_T3 ;
    wire LED_128_Instance_SBox_Instance_13_T1 ;
    wire LED_128_Instance_SBox_Instance_13_Q7 ;
    wire LED_128_Instance_SBox_Instance_13_Q6 ;
    wire LED_128_Instance_SBox_Instance_13_L5 ;
    wire LED_128_Instance_SBox_Instance_13_T2 ;
    wire LED_128_Instance_SBox_Instance_13_L4 ;
    wire LED_128_Instance_SBox_Instance_13_Q3 ;
    wire LED_128_Instance_SBox_Instance_13_L3 ;
    wire LED_128_Instance_SBox_Instance_13_Q2 ;
    wire LED_128_Instance_SBox_Instance_13_T0 ;
    wire LED_128_Instance_SBox_Instance_13_L2 ;
    wire LED_128_Instance_SBox_Instance_13_L1 ;
    wire LED_128_Instance_SBox_Instance_13_L0 ;
    wire LED_128_Instance_SBox_Instance_14_n3 ;
    wire LED_128_Instance_SBox_Instance_14_n2 ;
    wire LED_128_Instance_SBox_Instance_14_n1 ;
    wire LED_128_Instance_SBox_Instance_14_L8 ;
    wire LED_128_Instance_SBox_Instance_14_L7 ;
    wire LED_128_Instance_SBox_Instance_14_T3 ;
    wire LED_128_Instance_SBox_Instance_14_T1 ;
    wire LED_128_Instance_SBox_Instance_14_Q7 ;
    wire LED_128_Instance_SBox_Instance_14_Q6 ;
    wire LED_128_Instance_SBox_Instance_14_L5 ;
    wire LED_128_Instance_SBox_Instance_14_T2 ;
    wire LED_128_Instance_SBox_Instance_14_L4 ;
    wire LED_128_Instance_SBox_Instance_14_Q3 ;
    wire LED_128_Instance_SBox_Instance_14_L3 ;
    wire LED_128_Instance_SBox_Instance_14_Q2 ;
    wire LED_128_Instance_SBox_Instance_14_T0 ;
    wire LED_128_Instance_SBox_Instance_14_L2 ;
    wire LED_128_Instance_SBox_Instance_14_L1 ;
    wire LED_128_Instance_SBox_Instance_14_L0 ;
    wire LED_128_Instance_SBox_Instance_15_n3 ;
    wire LED_128_Instance_SBox_Instance_15_n2 ;
    wire LED_128_Instance_SBox_Instance_15_n1 ;
    wire LED_128_Instance_SBox_Instance_15_L8 ;
    wire LED_128_Instance_SBox_Instance_15_L7 ;
    wire LED_128_Instance_SBox_Instance_15_T3 ;
    wire LED_128_Instance_SBox_Instance_15_T1 ;
    wire LED_128_Instance_SBox_Instance_15_Q7 ;
    wire LED_128_Instance_SBox_Instance_15_Q6 ;
    wire LED_128_Instance_SBox_Instance_15_L5 ;
    wire LED_128_Instance_SBox_Instance_15_T2 ;
    wire LED_128_Instance_SBox_Instance_15_L4 ;
    wire LED_128_Instance_SBox_Instance_15_Q3 ;
    wire LED_128_Instance_SBox_Instance_15_L3 ;
    wire LED_128_Instance_SBox_Instance_15_Q2 ;
    wire LED_128_Instance_SBox_Instance_15_T0 ;
    wire LED_128_Instance_SBox_Instance_15_L2 ;
    wire LED_128_Instance_SBox_Instance_15_L1 ;
    wire LED_128_Instance_SBox_Instance_15_L0 ;
    wire LED_128_Instance_MCS_Instance_0_n38 ;
    wire LED_128_Instance_MCS_Instance_0_n37 ;
    wire LED_128_Instance_MCS_Instance_0_n36 ;
    wire LED_128_Instance_MCS_Instance_0_n35 ;
    wire LED_128_Instance_MCS_Instance_0_n34 ;
    wire LED_128_Instance_MCS_Instance_0_n33 ;
    wire LED_128_Instance_MCS_Instance_0_n32 ;
    wire LED_128_Instance_MCS_Instance_0_n31 ;
    wire LED_128_Instance_MCS_Instance_0_n30 ;
    wire LED_128_Instance_MCS_Instance_0_n29 ;
    wire LED_128_Instance_MCS_Instance_0_n28 ;
    wire LED_128_Instance_MCS_Instance_0_n27 ;
    wire LED_128_Instance_MCS_Instance_0_n26 ;
    wire LED_128_Instance_MCS_Instance_0_n25 ;
    wire LED_128_Instance_MCS_Instance_0_n24 ;
    wire LED_128_Instance_MCS_Instance_0_n23 ;
    wire LED_128_Instance_MCS_Instance_0_n22 ;
    wire LED_128_Instance_MCS_Instance_0_n21 ;
    wire LED_128_Instance_MCS_Instance_0_n20 ;
    wire LED_128_Instance_MCS_Instance_0_n19 ;
    wire LED_128_Instance_MCS_Instance_0_n18 ;
    wire LED_128_Instance_MCS_Instance_0_n17 ;
    wire LED_128_Instance_MCS_Instance_0_n16 ;
    wire LED_128_Instance_MCS_Instance_0_n15 ;
    wire LED_128_Instance_MCS_Instance_0_n14 ;
    wire LED_128_Instance_MCS_Instance_0_n13 ;
    wire LED_128_Instance_MCS_Instance_0_n12 ;
    wire LED_128_Instance_MCS_Instance_0_n11 ;
    wire LED_128_Instance_MCS_Instance_0_n10 ;
    wire LED_128_Instance_MCS_Instance_0_n9 ;
    wire LED_128_Instance_MCS_Instance_0_n8 ;
    wire LED_128_Instance_MCS_Instance_0_n7 ;
    wire LED_128_Instance_MCS_Instance_0_n6 ;
    wire LED_128_Instance_MCS_Instance_0_n5 ;
    wire LED_128_Instance_MCS_Instance_0_n4 ;
    wire LED_128_Instance_MCS_Instance_0_n3 ;
    wire LED_128_Instance_MCS_Instance_0_n2 ;
    wire LED_128_Instance_MCS_Instance_0_n1 ;
    wire LED_128_Instance_MCS_Instance_1_n38 ;
    wire LED_128_Instance_MCS_Instance_1_n37 ;
    wire LED_128_Instance_MCS_Instance_1_n36 ;
    wire LED_128_Instance_MCS_Instance_1_n35 ;
    wire LED_128_Instance_MCS_Instance_1_n34 ;
    wire LED_128_Instance_MCS_Instance_1_n33 ;
    wire LED_128_Instance_MCS_Instance_1_n32 ;
    wire LED_128_Instance_MCS_Instance_1_n31 ;
    wire LED_128_Instance_MCS_Instance_1_n30 ;
    wire LED_128_Instance_MCS_Instance_1_n29 ;
    wire LED_128_Instance_MCS_Instance_1_n28 ;
    wire LED_128_Instance_MCS_Instance_1_n27 ;
    wire LED_128_Instance_MCS_Instance_1_n26 ;
    wire LED_128_Instance_MCS_Instance_1_n25 ;
    wire LED_128_Instance_MCS_Instance_1_n24 ;
    wire LED_128_Instance_MCS_Instance_1_n23 ;
    wire LED_128_Instance_MCS_Instance_1_n22 ;
    wire LED_128_Instance_MCS_Instance_1_n21 ;
    wire LED_128_Instance_MCS_Instance_1_n20 ;
    wire LED_128_Instance_MCS_Instance_1_n19 ;
    wire LED_128_Instance_MCS_Instance_1_n18 ;
    wire LED_128_Instance_MCS_Instance_1_n17 ;
    wire LED_128_Instance_MCS_Instance_1_n16 ;
    wire LED_128_Instance_MCS_Instance_1_n15 ;
    wire LED_128_Instance_MCS_Instance_1_n14 ;
    wire LED_128_Instance_MCS_Instance_1_n13 ;
    wire LED_128_Instance_MCS_Instance_1_n12 ;
    wire LED_128_Instance_MCS_Instance_1_n11 ;
    wire LED_128_Instance_MCS_Instance_1_n10 ;
    wire LED_128_Instance_MCS_Instance_1_n9 ;
    wire LED_128_Instance_MCS_Instance_1_n8 ;
    wire LED_128_Instance_MCS_Instance_1_n7 ;
    wire LED_128_Instance_MCS_Instance_1_n6 ;
    wire LED_128_Instance_MCS_Instance_1_n5 ;
    wire LED_128_Instance_MCS_Instance_1_n4 ;
    wire LED_128_Instance_MCS_Instance_1_n3 ;
    wire LED_128_Instance_MCS_Instance_1_n2 ;
    wire LED_128_Instance_MCS_Instance_1_n1 ;
    wire LED_128_Instance_MCS_Instance_2_n38 ;
    wire LED_128_Instance_MCS_Instance_2_n37 ;
    wire LED_128_Instance_MCS_Instance_2_n36 ;
    wire LED_128_Instance_MCS_Instance_2_n35 ;
    wire LED_128_Instance_MCS_Instance_2_n34 ;
    wire LED_128_Instance_MCS_Instance_2_n33 ;
    wire LED_128_Instance_MCS_Instance_2_n32 ;
    wire LED_128_Instance_MCS_Instance_2_n31 ;
    wire LED_128_Instance_MCS_Instance_2_n30 ;
    wire LED_128_Instance_MCS_Instance_2_n29 ;
    wire LED_128_Instance_MCS_Instance_2_n28 ;
    wire LED_128_Instance_MCS_Instance_2_n27 ;
    wire LED_128_Instance_MCS_Instance_2_n26 ;
    wire LED_128_Instance_MCS_Instance_2_n25 ;
    wire LED_128_Instance_MCS_Instance_2_n24 ;
    wire LED_128_Instance_MCS_Instance_2_n23 ;
    wire LED_128_Instance_MCS_Instance_2_n22 ;
    wire LED_128_Instance_MCS_Instance_2_n21 ;
    wire LED_128_Instance_MCS_Instance_2_n20 ;
    wire LED_128_Instance_MCS_Instance_2_n19 ;
    wire LED_128_Instance_MCS_Instance_2_n18 ;
    wire LED_128_Instance_MCS_Instance_2_n17 ;
    wire LED_128_Instance_MCS_Instance_2_n16 ;
    wire LED_128_Instance_MCS_Instance_2_n15 ;
    wire LED_128_Instance_MCS_Instance_2_n14 ;
    wire LED_128_Instance_MCS_Instance_2_n13 ;
    wire LED_128_Instance_MCS_Instance_2_n12 ;
    wire LED_128_Instance_MCS_Instance_2_n11 ;
    wire LED_128_Instance_MCS_Instance_2_n10 ;
    wire LED_128_Instance_MCS_Instance_2_n9 ;
    wire LED_128_Instance_MCS_Instance_2_n8 ;
    wire LED_128_Instance_MCS_Instance_2_n7 ;
    wire LED_128_Instance_MCS_Instance_2_n6 ;
    wire LED_128_Instance_MCS_Instance_2_n5 ;
    wire LED_128_Instance_MCS_Instance_2_n4 ;
    wire LED_128_Instance_MCS_Instance_2_n3 ;
    wire LED_128_Instance_MCS_Instance_2_n2 ;
    wire LED_128_Instance_MCS_Instance_2_n1 ;
    wire LED_128_Instance_MCS_Instance_3_n38 ;
    wire LED_128_Instance_MCS_Instance_3_n37 ;
    wire LED_128_Instance_MCS_Instance_3_n36 ;
    wire LED_128_Instance_MCS_Instance_3_n35 ;
    wire LED_128_Instance_MCS_Instance_3_n34 ;
    wire LED_128_Instance_MCS_Instance_3_n33 ;
    wire LED_128_Instance_MCS_Instance_3_n32 ;
    wire LED_128_Instance_MCS_Instance_3_n31 ;
    wire LED_128_Instance_MCS_Instance_3_n30 ;
    wire LED_128_Instance_MCS_Instance_3_n29 ;
    wire LED_128_Instance_MCS_Instance_3_n28 ;
    wire LED_128_Instance_MCS_Instance_3_n27 ;
    wire LED_128_Instance_MCS_Instance_3_n26 ;
    wire LED_128_Instance_MCS_Instance_3_n25 ;
    wire LED_128_Instance_MCS_Instance_3_n24 ;
    wire LED_128_Instance_MCS_Instance_3_n23 ;
    wire LED_128_Instance_MCS_Instance_3_n22 ;
    wire LED_128_Instance_MCS_Instance_3_n21 ;
    wire LED_128_Instance_MCS_Instance_3_n20 ;
    wire LED_128_Instance_MCS_Instance_3_n19 ;
    wire LED_128_Instance_MCS_Instance_3_n18 ;
    wire LED_128_Instance_MCS_Instance_3_n17 ;
    wire LED_128_Instance_MCS_Instance_3_n16 ;
    wire LED_128_Instance_MCS_Instance_3_n15 ;
    wire LED_128_Instance_MCS_Instance_3_n14 ;
    wire LED_128_Instance_MCS_Instance_3_n13 ;
    wire LED_128_Instance_MCS_Instance_3_n12 ;
    wire LED_128_Instance_MCS_Instance_3_n11 ;
    wire LED_128_Instance_MCS_Instance_3_n10 ;
    wire LED_128_Instance_MCS_Instance_3_n9 ;
    wire LED_128_Instance_MCS_Instance_3_n8 ;
    wire LED_128_Instance_MCS_Instance_3_n7 ;
    wire LED_128_Instance_MCS_Instance_3_n6 ;
    wire LED_128_Instance_MCS_Instance_3_n5 ;
    wire LED_128_Instance_MCS_Instance_3_n4 ;
    wire LED_128_Instance_MCS_Instance_3_n3 ;
    wire LED_128_Instance_MCS_Instance_3_n2 ;
    wire LED_128_Instance_MCS_Instance_3_n1 ;
    wire LED_128_Instance_ks_reg_0__Q ;
    wire [5:0] roundconstant ;
    wire [63:0] LED_128_Instance_subcells_out ;
    wire [63:0] LED_128_Instance_addconst_out ;
    wire [63:0] LED_128_Instance_addroundkey_tmp ;
    wire [63:0] LED_128_Instance_current_roundkey ;
    wire [63:0] LED_128_Instance_state1 ;
    wire [63:0] LED_128_Instance_state0 ;
    wire [63:0] LED_128_Instance_mixcolumns_out ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4235 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4282 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4290 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4308 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4318 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4325 ;
    wire new_AGEMA_signal_4326 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4336 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4354 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4361 ;
    wire new_AGEMA_signal_4362 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4372 ;
    wire new_AGEMA_signal_4373 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4378 ;
    wire new_AGEMA_signal_4379 ;
    wire new_AGEMA_signal_4380 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4382 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4497 ;
    wire new_AGEMA_signal_4498 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5195 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5202 ;
    wire new_AGEMA_signal_5203 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5207 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5213 ;
    wire new_AGEMA_signal_5214 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5219 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5226 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5231 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5238 ;
    wire new_AGEMA_signal_5239 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5249 ;
    wire new_AGEMA_signal_5250 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5255 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5262 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5273 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5291 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5303 ;
    wire new_AGEMA_signal_5304 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5309 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;

    /* cells in depth 0 */
    NOR2_X1 U16 ( .A1 (roundconstant[4]), .A2 (roundconstant[1]), .ZN (n14) ) ;
    NAND2_X1 U17 ( .A1 (roundconstant[0]), .A2 (n14), .ZN (n16) ) ;
    NOR2_X1 U18 ( .A1 (roundconstant[5]), .A2 (n16), .ZN (n17) ) ;
    NAND2_X1 U19 ( .A1 (roundconstant[3]), .A2 (n17), .ZN (n18) ) ;
    NOR2_X1 U20 ( .A1 (roundconstant[2]), .A2 (n18), .ZN (n19) ) ;
    NOR2_X1 U21 ( .A1 (OUT_done), .A2 (n19), .ZN (n20) ) ;
    NOR2_X1 U22 ( .A1 (IN_reset), .A2 (n20), .ZN (n15) ) ;
    NAND2_X1 LED_128_Instance_U30 ( .A1 (LED_128_Instance_n33), .A2 (LED_128_Instance_n32), .ZN (LED_128_Instance_n34) ) ;
    XNOR2_X1 LED_128_Instance_U29 ( .A (LED_128_Instance_n25), .B (LED_128_Instance_n23), .ZN (LED_128_Instance_n32) ) ;
    XOR2_X1 LED_128_Instance_U28 ( .A (LED_128_Instance_n4), .B (LED_128_Instance_n26), .Z (LED_128_Instance_n23) ) ;
    NAND2_X1 LED_128_Instance_U27 ( .A1 (LED_128_Instance_n21), .A2 (LED_128_Instance_n20), .ZN (LED_128_Instance_n33) ) ;
    NAND2_X1 LED_128_Instance_U26 ( .A1 (LED_128_Instance_n19), .A2 (LED_128_Instance_n18), .ZN (LED_128_Instance_n20) ) ;
    NOR2_X1 LED_128_Instance_U25 ( .A1 (LED_128_Instance_n24), .A2 (LED_128_Instance_n1), .ZN (LED_128_Instance_n18) ) ;
    NOR2_X1 LED_128_Instance_U24 ( .A1 (LED_128_Instance_n8), .A2 (LED_128_Instance_n4), .ZN (LED_128_Instance_n19) ) ;
    NAND2_X1 LED_128_Instance_U23 ( .A1 (LED_128_Instance_n1), .A2 (LED_128_Instance_n17), .ZN (LED_128_Instance_n21) ) ;
    AND2_X1 LED_128_Instance_U22 ( .A1 (LED_128_Instance_n8), .A2 (LED_128_Instance_n4), .ZN (LED_128_Instance_n17) ) ;
    NAND2_X1 LED_128_Instance_U21 ( .A1 (LED_128_Instance_n29), .A2 (LED_128_Instance_n14), .ZN (LED_128_Instance_n15) ) ;
    NOR2_X1 LED_128_Instance_U20 ( .A1 (LED_128_Instance_n6), .A2 (LED_128_Instance_n13), .ZN (LED_128_Instance_n14) ) ;
    NAND2_X1 LED_128_Instance_U19 ( .A1 (LED_128_Instance_n5), .A2 (roundconstant[3]), .ZN (LED_128_Instance_n13) ) ;
    NAND2_X1 LED_128_Instance_U18 ( .A1 (LED_128_Instance_n28), .A2 (LED_128_Instance_n27), .ZN (LED_128_Instance_n16) ) ;
    NOR2_X1 LED_128_Instance_U17 ( .A1 (LED_128_Instance_n28), .A2 (IN_reset), .ZN (LED_128_Instance_N9) ) ;
    NOR2_X1 LED_128_Instance_U16 ( .A1 (IN_reset), .A2 (LED_128_Instance_n30), .ZN (LED_128_Instance_N8) ) ;
    NOR2_X1 LED_128_Instance_U15 ( .A1 (IN_reset), .A2 (LED_128_Instance_n5), .ZN (LED_128_Instance_N7) ) ;
    NOR2_X1 LED_128_Instance_U14 ( .A1 (IN_reset), .A2 (LED_128_Instance_n29), .ZN (LED_128_Instance_N6) ) ;
    NOR2_X1 LED_128_Instance_U13 ( .A1 (IN_reset), .A2 (LED_128_Instance_n6), .ZN (LED_128_Instance_N5) ) ;
    NOR2_X1 LED_128_Instance_U12 ( .A1 (LED_128_Instance_n1), .A2 (IN_reset), .ZN (LED_128_Instance_N13) ) ;
    NOR2_X1 LED_128_Instance_U11 ( .A1 (LED_128_Instance_n8), .A2 (IN_reset), .ZN (LED_128_Instance_N12) ) ;
    NOR2_X1 LED_128_Instance_U10 ( .A1 (LED_128_Instance_n4), .A2 (IN_reset), .ZN (LED_128_Instance_N11) ) ;
    NOR2_X1 LED_128_Instance_U9 ( .A1 (LED_128_Instance_n2), .A2 (IN_reset), .ZN (LED_128_Instance_N10) ) ;
    OR2_X1 LED_128_Instance_U8 ( .A1 (LED_128_Instance_n2), .A2 (LED_128_Instance_n21), .ZN (LED_128_Instance_n11) ) ;
    NAND2_X1 LED_128_Instance_U7 ( .A1 (LED_128_Instance_n34), .A2 (LED_128_Instance_n11), .ZN (LED_128_Instance_n31) ) ;
    NOR2_X1 LED_128_Instance_U6 ( .A1 (LED_128_Instance_n16), .A2 (LED_128_Instance_n15), .ZN (LED_128_Instance_n22) ) ;
    INV_X1 LED_128_Instance_U5 ( .A (LED_128_Instance_n11), .ZN (LED_128_Instance_n12) ) ;
    OR2_X1 LED_128_Instance_U4 ( .A1 (IN_reset), .A2 (LED_128_Instance_n10), .ZN (LED_128_Instance_N4) ) ;
    XNOR2_X1 LED_128_Instance_U3 ( .A (LED_128_Instance_n28), .B (LED_128_Instance_n27), .ZN (LED_128_Instance_n10) ) ;
    INV_X1 LED_128_Instance_MUX_state0_U4 ( .A (LED_128_Instance_n22), .ZN (LED_128_Instance_MUX_state0_n11) ) ;
    INV_X1 LED_128_Instance_MUX_state0_U3 ( .A (LED_128_Instance_MUX_state0_n11), .ZN (LED_128_Instance_MUX_state0_n8) ) ;
    INV_X1 LED_128_Instance_MUX_state0_U2 ( .A (LED_128_Instance_MUX_state0_n11), .ZN (LED_128_Instance_MUX_state0_n10) ) ;
    INV_X1 LED_128_Instance_MUX_state0_U1 ( .A (LED_128_Instance_MUX_state0_n11), .ZN (LED_128_Instance_MUX_state0_n9) ) ;
    INV_X1 LED_128_Instance_MUX_current_roundkey_U4 ( .A (LED_128_Instance_MUX_current_roundkey_n10), .ZN (LED_128_Instance_MUX_current_roundkey_n9) ) ;
    INV_X1 LED_128_Instance_MUX_current_roundkey_U3 ( .A (LED_128_Instance_n12), .ZN (LED_128_Instance_MUX_current_roundkey_n10) ) ;
    INV_X1 LED_128_Instance_MUX_current_roundkey_U2 ( .A (LED_128_Instance_MUX_current_roundkey_n10), .ZN (LED_128_Instance_MUX_current_roundkey_n7) ) ;
    INV_X1 LED_128_Instance_MUX_current_roundkey_U1 ( .A (LED_128_Instance_MUX_current_roundkey_n10), .ZN (LED_128_Instance_MUX_current_roundkey_n8) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s2[64], IN_key_s1[64], IN_key_s0[64]}), .a ({IN_key_s2[0], IN_key_s1[0], IN_key_s0[0]}), .c ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, LED_128_Instance_current_roundkey[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s2[65], IN_key_s1[65], IN_key_s0[65]}), .a ({IN_key_s2[1], IN_key_s1[1], IN_key_s0[1]}), .c ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, LED_128_Instance_current_roundkey[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s2[66], IN_key_s1[66], IN_key_s0[66]}), .a ({IN_key_s2[2], IN_key_s1[2], IN_key_s0[2]}), .c ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, LED_128_Instance_current_roundkey[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s2[67], IN_key_s1[67], IN_key_s0[67]}), .a ({IN_key_s2[3], IN_key_s1[3], IN_key_s0[3]}), .c ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, LED_128_Instance_current_roundkey[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s2[68], IN_key_s1[68], IN_key_s0[68]}), .a ({IN_key_s2[4], IN_key_s1[4], IN_key_s0[4]}), .c ({new_AGEMA_signal_1475, new_AGEMA_signal_1474, LED_128_Instance_current_roundkey[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s2[69], IN_key_s1[69], IN_key_s0[69]}), .a ({IN_key_s2[5], IN_key_s1[5], IN_key_s0[5]}), .c ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, LED_128_Instance_current_roundkey[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s2[70], IN_key_s1[70], IN_key_s0[70]}), .a ({IN_key_s2[6], IN_key_s1[6], IN_key_s0[6]}), .c ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, LED_128_Instance_current_roundkey[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s2[71], IN_key_s1[71], IN_key_s0[71]}), .a ({IN_key_s2[7], IN_key_s1[7], IN_key_s0[7]}), .c ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, LED_128_Instance_current_roundkey[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s2[72], IN_key_s1[72], IN_key_s0[72]}), .a ({IN_key_s2[8], IN_key_s1[8], IN_key_s0[8]}), .c ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, LED_128_Instance_current_roundkey[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s2[73], IN_key_s1[73], IN_key_s0[73]}), .a ({IN_key_s2[9], IN_key_s1[9], IN_key_s0[9]}), .c ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, LED_128_Instance_current_roundkey[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s2[74], IN_key_s1[74], IN_key_s0[74]}), .a ({IN_key_s2[10], IN_key_s1[10], IN_key_s0[10]}), .c ({new_AGEMA_signal_1511, new_AGEMA_signal_1510, LED_128_Instance_current_roundkey[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s2[75], IN_key_s1[75], IN_key_s0[75]}), .a ({IN_key_s2[11], IN_key_s1[11], IN_key_s0[11]}), .c ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, LED_128_Instance_current_roundkey[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s2[76], IN_key_s1[76], IN_key_s0[76]}), .a ({IN_key_s2[12], IN_key_s1[12], IN_key_s0[12]}), .c ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, LED_128_Instance_current_roundkey[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s2[77], IN_key_s1[77], IN_key_s0[77]}), .a ({IN_key_s2[13], IN_key_s1[13], IN_key_s0[13]}), .c ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, LED_128_Instance_current_roundkey[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s2[78], IN_key_s1[78], IN_key_s0[78]}), .a ({IN_key_s2[14], IN_key_s1[14], IN_key_s0[14]}), .c ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, LED_128_Instance_current_roundkey[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s2[79], IN_key_s1[79], IN_key_s0[79]}), .a ({IN_key_s2[15], IN_key_s1[15], IN_key_s0[15]}), .c ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, LED_128_Instance_current_roundkey[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s2[80], IN_key_s1[80], IN_key_s0[80]}), .a ({IN_key_s2[16], IN_key_s1[16], IN_key_s0[16]}), .c ({new_AGEMA_signal_1345, new_AGEMA_signal_1344, LED_128_Instance_current_roundkey[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s2[81], IN_key_s1[81], IN_key_s0[81]}), .a ({IN_key_s2[17], IN_key_s1[17], IN_key_s0[17]}), .c ({new_AGEMA_signal_1547, new_AGEMA_signal_1546, LED_128_Instance_current_roundkey[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s2[82], IN_key_s1[82], IN_key_s0[82]}), .a ({IN_key_s2[18], IN_key_s1[18], IN_key_s0[18]}), .c ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, LED_128_Instance_current_roundkey[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s2[83], IN_key_s1[83], IN_key_s0[83]}), .a ({IN_key_s2[19], IN_key_s1[19], IN_key_s0[19]}), .c ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, LED_128_Instance_current_roundkey[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s2[84], IN_key_s1[84], IN_key_s0[84]}), .a ({IN_key_s2[20], IN_key_s1[20], IN_key_s0[20]}), .c ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_current_roundkey[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s2[85], IN_key_s1[85], IN_key_s0[85]}), .a ({IN_key_s2[21], IN_key_s1[21], IN_key_s0[21]}), .c ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, LED_128_Instance_current_roundkey[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s2[86], IN_key_s1[86], IN_key_s0[86]}), .a ({IN_key_s2[22], IN_key_s1[22], IN_key_s0[22]}), .c ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, LED_128_Instance_current_roundkey[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s2[87], IN_key_s1[87], IN_key_s0[87]}), .a ({IN_key_s2[23], IN_key_s1[23], IN_key_s0[23]}), .c ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, LED_128_Instance_current_roundkey[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s2[88], IN_key_s1[88], IN_key_s0[88]}), .a ({IN_key_s2[24], IN_key_s1[24], IN_key_s0[24]}), .c ({new_AGEMA_signal_1363, new_AGEMA_signal_1362, LED_128_Instance_current_roundkey[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s2[89], IN_key_s1[89], IN_key_s0[89]}), .a ({IN_key_s2[25], IN_key_s1[25], IN_key_s0[25]}), .c ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, LED_128_Instance_current_roundkey[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s2[90], IN_key_s1[90], IN_key_s0[90]}), .a ({IN_key_s2[26], IN_key_s1[26], IN_key_s0[26]}), .c ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, LED_128_Instance_current_roundkey[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s2[91], IN_key_s1[91], IN_key_s0[91]}), .a ({IN_key_s2[27], IN_key_s1[27], IN_key_s0[27]}), .c ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, LED_128_Instance_current_roundkey[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s2[92], IN_key_s1[92], IN_key_s0[92]}), .a ({IN_key_s2[28], IN_key_s1[28], IN_key_s0[28]}), .c ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, LED_128_Instance_current_roundkey[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s2[93], IN_key_s1[93], IN_key_s0[93]}), .a ({IN_key_s2[29], IN_key_s1[29], IN_key_s0[29]}), .c ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, LED_128_Instance_current_roundkey[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s2[94], IN_key_s1[94], IN_key_s0[94]}), .a ({IN_key_s2[30], IN_key_s1[30], IN_key_s0[30]}), .c ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, LED_128_Instance_current_roundkey[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s2[95], IN_key_s1[95], IN_key_s0[95]}), .a ({IN_key_s2[31], IN_key_s1[31], IN_key_s0[31]}), .c ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, LED_128_Instance_current_roundkey[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s2[96], IN_key_s1[96], IN_key_s0[96]}), .a ({IN_key_s2[32], IN_key_s1[32], IN_key_s0[32]}), .c ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, LED_128_Instance_current_roundkey[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s2[97], IN_key_s1[97], IN_key_s0[97]}), .a ({IN_key_s2[33], IN_key_s1[33], IN_key_s0[33]}), .c ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, LED_128_Instance_current_roundkey[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s2[98], IN_key_s1[98], IN_key_s0[98]}), .a ({IN_key_s2[34], IN_key_s1[34], IN_key_s0[34]}), .c ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, LED_128_Instance_current_roundkey[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s2[99], IN_key_s1[99], IN_key_s0[99]}), .a ({IN_key_s2[35], IN_key_s1[35], IN_key_s0[35]}), .c ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, LED_128_Instance_current_roundkey[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s2[100], IN_key_s1[100], IN_key_s0[100]}), .a ({IN_key_s2[36], IN_key_s1[36], IN_key_s0[36]}), .c ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, LED_128_Instance_current_roundkey[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s2[101], IN_key_s1[101], IN_key_s0[101]}), .a ({IN_key_s2[37], IN_key_s1[37], IN_key_s0[37]}), .c ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, LED_128_Instance_current_roundkey[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s2[102], IN_key_s1[102], IN_key_s0[102]}), .a ({IN_key_s2[38], IN_key_s1[38], IN_key_s0[38]}), .c ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, LED_128_Instance_current_roundkey[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s2[103], IN_key_s1[103], IN_key_s0[103]}), .a ({IN_key_s2[39], IN_key_s1[39], IN_key_s0[39]}), .c ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, LED_128_Instance_current_roundkey[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s2[104], IN_key_s1[104], IN_key_s0[104]}), .a ({IN_key_s2[40], IN_key_s1[40], IN_key_s0[40]}), .c ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, LED_128_Instance_current_roundkey[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s2[105], IN_key_s1[105], IN_key_s0[105]}), .a ({IN_key_s2[41], IN_key_s1[41], IN_key_s0[41]}), .c ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, LED_128_Instance_current_roundkey[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s2[106], IN_key_s1[106], IN_key_s0[106]}), .a ({IN_key_s2[42], IN_key_s1[42], IN_key_s0[42]}), .c ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, LED_128_Instance_current_roundkey[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s2[107], IN_key_s1[107], IN_key_s0[107]}), .a ({IN_key_s2[43], IN_key_s1[43], IN_key_s0[43]}), .c ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, LED_128_Instance_current_roundkey[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s2[108], IN_key_s1[108], IN_key_s0[108]}), .a ({IN_key_s2[44], IN_key_s1[44], IN_key_s0[44]}), .c ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, LED_128_Instance_current_roundkey[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s2[109], IN_key_s1[109], IN_key_s0[109]}), .a ({IN_key_s2[45], IN_key_s1[45], IN_key_s0[45]}), .c ({new_AGEMA_signal_1655, new_AGEMA_signal_1654, LED_128_Instance_current_roundkey[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s2[110], IN_key_s1[110], IN_key_s0[110]}), .a ({IN_key_s2[46], IN_key_s1[46], IN_key_s0[46]}), .c ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, LED_128_Instance_current_roundkey[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s2[111], IN_key_s1[111], IN_key_s0[111]}), .a ({IN_key_s2[47], IN_key_s1[47], IN_key_s0[47]}), .c ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, LED_128_Instance_current_roundkey[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s2[112], IN_key_s1[112], IN_key_s0[112]}), .a ({IN_key_s2[48], IN_key_s1[48], IN_key_s0[48]}), .c ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, LED_128_Instance_current_roundkey[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s2[113], IN_key_s1[113], IN_key_s0[113]}), .a ({IN_key_s2[49], IN_key_s1[49], IN_key_s0[49]}), .c ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, LED_128_Instance_current_roundkey[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s2[114], IN_key_s1[114], IN_key_s0[114]}), .a ({IN_key_s2[50], IN_key_s1[50], IN_key_s0[50]}), .c ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, LED_128_Instance_current_roundkey[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s2[115], IN_key_s1[115], IN_key_s0[115]}), .a ({IN_key_s2[51], IN_key_s1[51], IN_key_s0[51]}), .c ({new_AGEMA_signal_1691, new_AGEMA_signal_1690, LED_128_Instance_current_roundkey[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s2[116], IN_key_s1[116], IN_key_s0[116]}), .a ({IN_key_s2[52], IN_key_s1[52], IN_key_s0[52]}), .c ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, LED_128_Instance_current_roundkey[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s2[117], IN_key_s1[117], IN_key_s0[117]}), .a ({IN_key_s2[53], IN_key_s1[53], IN_key_s0[53]}), .c ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, LED_128_Instance_current_roundkey[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s2[118], IN_key_s1[118], IN_key_s0[118]}), .a ({IN_key_s2[54], IN_key_s1[54], IN_key_s0[54]}), .c ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, LED_128_Instance_current_roundkey[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s2[119], IN_key_s1[119], IN_key_s0[119]}), .a ({IN_key_s2[55], IN_key_s1[55], IN_key_s0[55]}), .c ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, LED_128_Instance_current_roundkey[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s2[120], IN_key_s1[120], IN_key_s0[120]}), .a ({IN_key_s2[56], IN_key_s1[56], IN_key_s0[56]}), .c ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, LED_128_Instance_current_roundkey[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s2[121], IN_key_s1[121], IN_key_s0[121]}), .a ({IN_key_s2[57], IN_key_s1[57], IN_key_s0[57]}), .c ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, LED_128_Instance_current_roundkey[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s2[122], IN_key_s1[122], IN_key_s0[122]}), .a ({IN_key_s2[58], IN_key_s1[58], IN_key_s0[58]}), .c ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, LED_128_Instance_current_roundkey[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s2[123], IN_key_s1[123], IN_key_s0[123]}), .a ({IN_key_s2[59], IN_key_s1[59], IN_key_s0[59]}), .c ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, LED_128_Instance_current_roundkey[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s2[124], IN_key_s1[124], IN_key_s0[124]}), .a ({IN_key_s2[60], IN_key_s1[60], IN_key_s0[60]}), .c ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, LED_128_Instance_current_roundkey[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s2[125], IN_key_s1[125], IN_key_s0[125]}), .a ({IN_key_s2[61], IN_key_s1[61], IN_key_s0[61]}), .c ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, LED_128_Instance_current_roundkey[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s2[126], IN_key_s1[126], IN_key_s0[126]}), .a ({IN_key_s2[62], IN_key_s1[62], IN_key_s0[62]}), .c ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, LED_128_Instance_current_roundkey[62]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s2[127], IN_key_s1[127], IN_key_s0[127]}), .a ({IN_key_s2[63], IN_key_s1[63], IN_key_s0[63]}), .c ({new_AGEMA_signal_1763, new_AGEMA_signal_1762, LED_128_Instance_current_roundkey[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U64 ( .a ({OUT_ciphertext_s2[9], OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .b ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, LED_128_Instance_current_roundkey[9]}), .c ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, LED_128_Instance_addroundkey_tmp[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U63 ( .a ({OUT_ciphertext_s2[8], OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .b ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, LED_128_Instance_current_roundkey[8]}), .c ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, LED_128_Instance_addroundkey_tmp[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U62 ( .a ({OUT_ciphertext_s2[7], OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .b ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, LED_128_Instance_current_roundkey[7]}), .c ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, LED_128_Instance_addroundkey_tmp[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U61 ( .a ({OUT_ciphertext_s2[6], OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .b ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, LED_128_Instance_current_roundkey[6]}), .c ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, LED_128_Instance_addroundkey_tmp[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U60 ( .a ({OUT_ciphertext_s2[63], OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .b ({new_AGEMA_signal_1763, new_AGEMA_signal_1762, LED_128_Instance_current_roundkey[63]}), .c ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, LED_128_Instance_addroundkey_tmp[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U59 ( .a ({OUT_ciphertext_s2[62], OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .b ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, LED_128_Instance_current_roundkey[62]}), .c ({new_AGEMA_signal_1801, new_AGEMA_signal_1800, LED_128_Instance_addroundkey_tmp[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U58 ( .a ({OUT_ciphertext_s2[61], OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .b ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, LED_128_Instance_current_roundkey[61]}), .c ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, LED_128_Instance_addroundkey_tmp[61]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U57 ( .a ({OUT_ciphertext_s2[60], OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .b ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, LED_128_Instance_current_roundkey[60]}), .c ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, LED_128_Instance_addroundkey_tmp[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U56 ( .a ({OUT_ciphertext_s2[5], OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .b ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, LED_128_Instance_current_roundkey[5]}), .c ({new_AGEMA_signal_1813, new_AGEMA_signal_1812, LED_128_Instance_addroundkey_tmp[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U55 ( .a ({OUT_ciphertext_s2[59], OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .b ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, LED_128_Instance_current_roundkey[59]}), .c ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, LED_128_Instance_addroundkey_tmp[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U54 ( .a ({OUT_ciphertext_s2[58], OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .b ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, LED_128_Instance_current_roundkey[58]}), .c ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, LED_128_Instance_addroundkey_tmp[58]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U53 ( .a ({OUT_ciphertext_s2[57], OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .b ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, LED_128_Instance_current_roundkey[57]}), .c ({new_AGEMA_signal_1825, new_AGEMA_signal_1824, LED_128_Instance_addroundkey_tmp[57]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U52 ( .a ({OUT_ciphertext_s2[56], OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .b ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, LED_128_Instance_current_roundkey[56]}), .c ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, LED_128_Instance_addroundkey_tmp[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U51 ( .a ({OUT_ciphertext_s2[55], OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .b ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, LED_128_Instance_current_roundkey[55]}), .c ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, LED_128_Instance_addroundkey_tmp[55]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U50 ( .a ({OUT_ciphertext_s2[54], OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .b ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, LED_128_Instance_current_roundkey[54]}), .c ({new_AGEMA_signal_1837, new_AGEMA_signal_1836, LED_128_Instance_addroundkey_tmp[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U49 ( .a ({OUT_ciphertext_s2[53], OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .b ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, LED_128_Instance_current_roundkey[53]}), .c ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, LED_128_Instance_addroundkey_tmp[53]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U48 ( .a ({OUT_ciphertext_s2[52], OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .b ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, LED_128_Instance_current_roundkey[52]}), .c ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, LED_128_Instance_addroundkey_tmp[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U47 ( .a ({OUT_ciphertext_s2[51], OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .b ({new_AGEMA_signal_1691, new_AGEMA_signal_1690, LED_128_Instance_current_roundkey[51]}), .c ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, LED_128_Instance_addroundkey_tmp[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U46 ( .a ({OUT_ciphertext_s2[50], OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .b ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, LED_128_Instance_current_roundkey[50]}), .c ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, LED_128_Instance_addroundkey_tmp[50]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U45 ( .a ({OUT_ciphertext_s2[4], OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .b ({new_AGEMA_signal_1475, new_AGEMA_signal_1474, LED_128_Instance_current_roundkey[4]}), .c ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, LED_128_Instance_addroundkey_tmp[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U44 ( .a ({OUT_ciphertext_s2[49], OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .b ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, LED_128_Instance_current_roundkey[49]}), .c ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, LED_128_Instance_addroundkey_tmp[49]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U43 ( .a ({OUT_ciphertext_s2[48], OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .b ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, LED_128_Instance_current_roundkey[48]}), .c ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, LED_128_Instance_addroundkey_tmp[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U42 ( .a ({OUT_ciphertext_s2[47], OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .b ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, LED_128_Instance_current_roundkey[47]}), .c ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, LED_128_Instance_addroundkey_tmp[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U41 ( .a ({OUT_ciphertext_s2[46], OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .b ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, LED_128_Instance_current_roundkey[46]}), .c ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, LED_128_Instance_addroundkey_tmp[46]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U40 ( .a ({OUT_ciphertext_s2[45], OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .b ({new_AGEMA_signal_1655, new_AGEMA_signal_1654, LED_128_Instance_current_roundkey[45]}), .c ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, LED_128_Instance_addroundkey_tmp[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U39 ( .a ({OUT_ciphertext_s2[44], OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .b ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, LED_128_Instance_current_roundkey[44]}), .c ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, LED_128_Instance_addroundkey_tmp[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U38 ( .a ({OUT_ciphertext_s2[43], OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .b ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, LED_128_Instance_current_roundkey[43]}), .c ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, LED_128_Instance_addroundkey_tmp[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U37 ( .a ({OUT_ciphertext_s2[42], OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .b ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, LED_128_Instance_current_roundkey[42]}), .c ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, LED_128_Instance_addroundkey_tmp[42]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U36 ( .a ({OUT_ciphertext_s2[41], OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .b ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, LED_128_Instance_current_roundkey[41]}), .c ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, LED_128_Instance_addroundkey_tmp[41]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U35 ( .a ({OUT_ciphertext_s2[40], OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .b ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, LED_128_Instance_current_roundkey[40]}), .c ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, LED_128_Instance_addroundkey_tmp[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U34 ( .a ({OUT_ciphertext_s2[3], OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .b ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, LED_128_Instance_current_roundkey[3]}), .c ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, LED_128_Instance_addroundkey_tmp[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U33 ( .a ({OUT_ciphertext_s2[39], OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .b ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, LED_128_Instance_current_roundkey[39]}), .c ({new_AGEMA_signal_1413, new_AGEMA_signal_1412, LED_128_Instance_addroundkey_tmp[39]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U32 ( .a ({OUT_ciphertext_s2[38], OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .b ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, LED_128_Instance_current_roundkey[38]}), .c ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, LED_128_Instance_addroundkey_tmp[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U31 ( .a ({OUT_ciphertext_s2[37], OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .b ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, LED_128_Instance_current_roundkey[37]}), .c ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, LED_128_Instance_addroundkey_tmp[37]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U30 ( .a ({OUT_ciphertext_s2[36], OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .b ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, LED_128_Instance_current_roundkey[36]}), .c ({new_AGEMA_signal_1417, new_AGEMA_signal_1416, LED_128_Instance_addroundkey_tmp[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U29 ( .a ({OUT_ciphertext_s2[35], OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .b ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, LED_128_Instance_current_roundkey[35]}), .c ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, LED_128_Instance_addroundkey_tmp[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U28 ( .a ({OUT_ciphertext_s2[34], OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .b ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, LED_128_Instance_current_roundkey[34]}), .c ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, LED_128_Instance_addroundkey_tmp[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U27 ( .a ({OUT_ciphertext_s2[33], OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .b ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, LED_128_Instance_current_roundkey[33]}), .c ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, LED_128_Instance_addroundkey_tmp[33]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U26 ( .a ({OUT_ciphertext_s2[32], OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .b ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, LED_128_Instance_current_roundkey[32]}), .c ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, LED_128_Instance_addroundkey_tmp[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U25 ( .a ({OUT_ciphertext_s2[31], OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .b ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, LED_128_Instance_current_roundkey[31]}), .c ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, LED_128_Instance_addroundkey_tmp[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U24 ( .a ({OUT_ciphertext_s2[30], OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .b ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, LED_128_Instance_current_roundkey[30]}), .c ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, LED_128_Instance_addroundkey_tmp[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U23 ( .a ({OUT_ciphertext_s2[2], OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .b ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, LED_128_Instance_current_roundkey[2]}), .c ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, LED_128_Instance_addroundkey_tmp[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U22 ( .a ({OUT_ciphertext_s2[29], OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .b ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, LED_128_Instance_current_roundkey[29]}), .c ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, LED_128_Instance_addroundkey_tmp[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U21 ( .a ({OUT_ciphertext_s2[28], OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .b ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, LED_128_Instance_current_roundkey[28]}), .c ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, LED_128_Instance_addroundkey_tmp[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U20 ( .a ({OUT_ciphertext_s2[27], OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .b ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, LED_128_Instance_current_roundkey[27]}), .c ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, LED_128_Instance_addroundkey_tmp[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U19 ( .a ({OUT_ciphertext_s2[26], OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .b ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, LED_128_Instance_current_roundkey[26]}), .c ({new_AGEMA_signal_1437, new_AGEMA_signal_1436, LED_128_Instance_addroundkey_tmp[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U18 ( .a ({OUT_ciphertext_s2[25], OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .b ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, LED_128_Instance_current_roundkey[25]}), .c ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, LED_128_Instance_addroundkey_tmp[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U17 ( .a ({OUT_ciphertext_s2[24], OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .b ({new_AGEMA_signal_1363, new_AGEMA_signal_1362, LED_128_Instance_current_roundkey[24]}), .c ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, LED_128_Instance_addroundkey_tmp[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U16 ( .a ({OUT_ciphertext_s2[23], OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .b ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, LED_128_Instance_current_roundkey[23]}), .c ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, LED_128_Instance_addroundkey_tmp[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U15 ( .a ({OUT_ciphertext_s2[22], OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .b ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, LED_128_Instance_current_roundkey[22]}), .c ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, LED_128_Instance_addroundkey_tmp[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U14 ( .a ({OUT_ciphertext_s2[21], OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .b ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, LED_128_Instance_current_roundkey[21]}), .c ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, LED_128_Instance_addroundkey_tmp[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U13 ( .a ({OUT_ciphertext_s2[20], OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .b ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_current_roundkey[20]}), .c ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, LED_128_Instance_addroundkey_tmp[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U12 ( .a ({OUT_ciphertext_s2[1], OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .b ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, LED_128_Instance_current_roundkey[1]}), .c ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, LED_128_Instance_addroundkey_tmp[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U11 ( .a ({OUT_ciphertext_s2[19], OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .b ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, LED_128_Instance_current_roundkey[19]}), .c ({new_AGEMA_signal_1449, new_AGEMA_signal_1448, LED_128_Instance_addroundkey_tmp[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U10 ( .a ({OUT_ciphertext_s2[18], OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .b ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, LED_128_Instance_current_roundkey[18]}), .c ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, LED_128_Instance_addroundkey_tmp[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U9 ( .a ({OUT_ciphertext_s2[17], OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .b ({new_AGEMA_signal_1547, new_AGEMA_signal_1546, LED_128_Instance_current_roundkey[17]}), .c ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, LED_128_Instance_addroundkey_tmp[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U8 ( .a ({OUT_ciphertext_s2[16], OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .b ({new_AGEMA_signal_1345, new_AGEMA_signal_1344, LED_128_Instance_current_roundkey[16]}), .c ({new_AGEMA_signal_1453, new_AGEMA_signal_1452, LED_128_Instance_addroundkey_tmp[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U7 ( .a ({OUT_ciphertext_s2[15], OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .b ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, LED_128_Instance_current_roundkey[15]}), .c ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, LED_128_Instance_addroundkey_tmp[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U6 ( .a ({OUT_ciphertext_s2[14], OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .b ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, LED_128_Instance_current_roundkey[14]}), .c ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, LED_128_Instance_addroundkey_tmp[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U5 ( .a ({OUT_ciphertext_s2[13], OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .b ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, LED_128_Instance_current_roundkey[13]}), .c ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, LED_128_Instance_addroundkey_tmp[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U4 ( .a ({OUT_ciphertext_s2[12], OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .b ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, LED_128_Instance_current_roundkey[12]}), .c ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, LED_128_Instance_addroundkey_tmp[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U3 ( .a ({OUT_ciphertext_s2[11], OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .b ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, LED_128_Instance_current_roundkey[11]}), .c ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, LED_128_Instance_addroundkey_tmp[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U2 ( .a ({OUT_ciphertext_s2[10], OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .b ({new_AGEMA_signal_1511, new_AGEMA_signal_1510, LED_128_Instance_current_roundkey[10]}), .c ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, LED_128_Instance_addroundkey_tmp[10]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U1 ( .a ({OUT_ciphertext_s2[0], OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .b ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, LED_128_Instance_current_roundkey[0]}), .c ({new_AGEMA_signal_1457, new_AGEMA_signal_1456, LED_128_Instance_addroundkey_tmp[0]}) ) ;
    INV_X1 LED_128_Instance_MUX_addroundkey_out_U3 ( .A (LED_128_Instance_MUX_addroundkey_out_n9), .ZN (LED_128_Instance_MUX_addroundkey_out_n7) ) ;
    INV_X1 LED_128_Instance_MUX_addroundkey_out_U2 ( .A (LED_128_Instance_n31), .ZN (LED_128_Instance_MUX_addroundkey_out_n9) ) ;
    INV_X1 LED_128_Instance_MUX_addroundkey_out_U1 ( .A (LED_128_Instance_MUX_addroundkey_out_n9), .ZN (LED_128_Instance_MUX_addroundkey_out_n8) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s2[0], OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .a ({new_AGEMA_signal_1457, new_AGEMA_signal_1456, LED_128_Instance_addroundkey_tmp[0]}), .c ({new_AGEMA_signal_1765, new_AGEMA_signal_1764, LED_128_Instance_addroundkey_out_0_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s2[1], OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .a ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, LED_128_Instance_addroundkey_tmp[1]}), .c ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, LED_128_Instance_addroundkey_out_1_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s2[2], OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .a ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, LED_128_Instance_addroundkey_tmp[2]}), .c ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, LED_128_Instance_addroundkey_out_2_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s2[3], OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .a ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, LED_128_Instance_addroundkey_tmp[3]}), .c ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, LED_128_Instance_addroundkey_out_3_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s2[4], OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .a ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, LED_128_Instance_addroundkey_tmp[4]}), .c ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, LED_128_Instance_addroundkey_out_4_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s2[5], OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .a ({new_AGEMA_signal_1813, new_AGEMA_signal_1812, LED_128_Instance_addroundkey_tmp[5]}), .c ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, LED_128_Instance_addroundkey_out_5_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s2[6], OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .a ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, LED_128_Instance_addroundkey_tmp[6]}), .c ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, LED_128_Instance_addroundkey_out_6_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s2[7], OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .a ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, LED_128_Instance_addroundkey_tmp[7]}), .c ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, LED_128_Instance_addconst_out[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s2[8], OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .a ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, LED_128_Instance_addroundkey_tmp[8]}), .c ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, LED_128_Instance_addconst_out[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s2[9], OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .a ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, LED_128_Instance_addroundkey_tmp[9]}), .c ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, LED_128_Instance_addconst_out[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s2[10], OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .a ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, LED_128_Instance_addroundkey_tmp[10]}), .c ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, LED_128_Instance_addconst_out[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s2[11], OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .a ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, LED_128_Instance_addroundkey_tmp[11]}), .c ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, LED_128_Instance_addconst_out[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s2[12], OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .a ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, LED_128_Instance_addroundkey_tmp[12]}), .c ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, LED_128_Instance_addconst_out[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s2[13], OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .a ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, LED_128_Instance_addroundkey_tmp[13]}), .c ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, LED_128_Instance_addconst_out[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s2[14], OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .a ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, LED_128_Instance_addroundkey_tmp[14]}), .c ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, LED_128_Instance_addconst_out[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s2[15], OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .a ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, LED_128_Instance_addroundkey_tmp[15]}), .c ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, LED_128_Instance_addconst_out[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s2[16], OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .a ({new_AGEMA_signal_1453, new_AGEMA_signal_1452, LED_128_Instance_addroundkey_tmp[16]}), .c ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, LED_128_Instance_addroundkey_out_16_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s2[17], OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .a ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, LED_128_Instance_addroundkey_tmp[17]}), .c ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, LED_128_Instance_addroundkey_out_17_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s2[18], OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .a ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, LED_128_Instance_addroundkey_tmp[18]}), .c ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, LED_128_Instance_addroundkey_out_18_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s2[19], OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .a ({new_AGEMA_signal_1449, new_AGEMA_signal_1448, LED_128_Instance_addroundkey_tmp[19]}), .c ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, LED_128_Instance_addroundkey_out_19_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s2[20], OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .a ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, LED_128_Instance_addroundkey_tmp[20]}), .c ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, LED_128_Instance_addroundkey_out_20_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s2[21], OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .a ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, LED_128_Instance_addroundkey_tmp[21]}), .c ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, LED_128_Instance_addroundkey_out_21_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s2[22], OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .a ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, LED_128_Instance_addroundkey_tmp[22]}), .c ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, LED_128_Instance_addroundkey_out_22_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s2[23], OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .a ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, LED_128_Instance_addroundkey_tmp[23]}), .c ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, LED_128_Instance_addconst_out[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s2[24], OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .a ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, LED_128_Instance_addroundkey_tmp[24]}), .c ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, LED_128_Instance_addconst_out[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s2[25], OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .a ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, LED_128_Instance_addroundkey_tmp[25]}), .c ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, LED_128_Instance_addconst_out[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s2[26], OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .a ({new_AGEMA_signal_1437, new_AGEMA_signal_1436, LED_128_Instance_addroundkey_tmp[26]}), .c ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_addconst_out[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s2[27], OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .a ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, LED_128_Instance_addroundkey_tmp[27]}), .c ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, LED_128_Instance_addconst_out[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[28], OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .a ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, LED_128_Instance_addroundkey_tmp[28]}), .c ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, LED_128_Instance_addconst_out[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[29], OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .a ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, LED_128_Instance_addroundkey_tmp[29]}), .c ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, LED_128_Instance_addconst_out[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[30], OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .a ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, LED_128_Instance_addroundkey_tmp[30]}), .c ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, LED_128_Instance_addconst_out[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[31], OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .a ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, LED_128_Instance_addroundkey_tmp[31]}), .c ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, LED_128_Instance_addconst_out[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[32], OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .a ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, LED_128_Instance_addroundkey_tmp[32]}), .c ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, LED_128_Instance_addroundkey_out_32_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[33], OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .a ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, LED_128_Instance_addroundkey_tmp[33]}), .c ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, LED_128_Instance_addroundkey_out_33_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[34], OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .a ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, LED_128_Instance_addroundkey_tmp[34]}), .c ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, LED_128_Instance_addroundkey_out_34_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[35], OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .a ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, LED_128_Instance_addroundkey_tmp[35]}), .c ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, LED_128_Instance_addroundkey_out_35_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[36], OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .a ({new_AGEMA_signal_1417, new_AGEMA_signal_1416, LED_128_Instance_addroundkey_tmp[36]}), .c ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, LED_128_Instance_addroundkey_out_36_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s2[37], OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .a ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, LED_128_Instance_addroundkey_tmp[37]}), .c ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, LED_128_Instance_addroundkey_out_37_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[38], OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .a ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, LED_128_Instance_addroundkey_tmp[38]}), .c ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, LED_128_Instance_addroundkey_out_38_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[39], OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .a ({new_AGEMA_signal_1413, new_AGEMA_signal_1412, LED_128_Instance_addroundkey_tmp[39]}), .c ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, LED_128_Instance_addconst_out[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[40], OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .a ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, LED_128_Instance_addroundkey_tmp[40]}), .c ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, LED_128_Instance_addconst_out[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[41], OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .a ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, LED_128_Instance_addroundkey_tmp[41]}), .c ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, LED_128_Instance_addconst_out[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[42], OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .a ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, LED_128_Instance_addroundkey_tmp[42]}), .c ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, LED_128_Instance_addconst_out[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[43], OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .a ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, LED_128_Instance_addroundkey_tmp[43]}), .c ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, LED_128_Instance_addconst_out[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[44], OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .a ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, LED_128_Instance_addroundkey_tmp[44]}), .c ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, LED_128_Instance_addconst_out[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[45], OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .a ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, LED_128_Instance_addroundkey_tmp[45]}), .c ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, LED_128_Instance_addconst_out[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[46], OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .a ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, LED_128_Instance_addroundkey_tmp[46]}), .c ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, LED_128_Instance_addconst_out[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[47], OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .a ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, LED_128_Instance_addroundkey_tmp[47]}), .c ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, LED_128_Instance_addconst_out[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[48], OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .a ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, LED_128_Instance_addroundkey_tmp[48]}), .c ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, LED_128_Instance_addroundkey_out_48_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[49], OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .a ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, LED_128_Instance_addroundkey_tmp[49]}), .c ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, LED_128_Instance_addroundkey_out_49_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s2[50], OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .a ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, LED_128_Instance_addroundkey_tmp[50]}), .c ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, LED_128_Instance_addroundkey_out_50_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[51], OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .a ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, LED_128_Instance_addroundkey_tmp[51]}), .c ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, LED_128_Instance_addroundkey_out_51_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[52], OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .a ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, LED_128_Instance_addroundkey_tmp[52]}), .c ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, LED_128_Instance_addroundkey_out_52_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[53], OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .a ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, LED_128_Instance_addroundkey_tmp[53]}), .c ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, LED_128_Instance_addroundkey_out_53_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[54], OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .a ({new_AGEMA_signal_1837, new_AGEMA_signal_1836, LED_128_Instance_addroundkey_tmp[54]}), .c ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, LED_128_Instance_addroundkey_out_54_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[55], OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .a ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, LED_128_Instance_addroundkey_tmp[55]}), .c ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, LED_128_Instance_addconst_out[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[56], OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .a ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, LED_128_Instance_addroundkey_tmp[56]}), .c ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, LED_128_Instance_addconst_out[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[57], OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .a ({new_AGEMA_signal_1825, new_AGEMA_signal_1824, LED_128_Instance_addroundkey_tmp[57]}), .c ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, LED_128_Instance_addconst_out[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[58], OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .a ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, LED_128_Instance_addroundkey_tmp[58]}), .c ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, LED_128_Instance_addconst_out[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[59], OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .a ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, LED_128_Instance_addroundkey_tmp[59]}), .c ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, LED_128_Instance_addconst_out[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[60], OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .a ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, LED_128_Instance_addroundkey_tmp[60]}), .c ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, LED_128_Instance_addconst_out[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[61], OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .a ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, LED_128_Instance_addroundkey_tmp[61]}), .c ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, LED_128_Instance_addconst_out[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[62], OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .a ({new_AGEMA_signal_1801, new_AGEMA_signal_1800, LED_128_Instance_addroundkey_tmp[62]}), .c ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, LED_128_Instance_addconst_out[62]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s2[63], OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .a ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, LED_128_Instance_addroundkey_tmp[63]}), .c ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, LED_128_Instance_addconst_out[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U28 ( .a ({1'b0, 1'b0, roundconstant[5]}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, LED_128_Instance_addroundkey_out_6_}), .c ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, LED_128_Instance_addconst_out[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U27 ( .a ({1'b0, 1'b0, roundconstant[4]}), .b ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, LED_128_Instance_addroundkey_out_5_}), .c ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, LED_128_Instance_addconst_out[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U26 ( .a ({1'b0, 1'b0, roundconstant[2]}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, LED_128_Instance_addroundkey_out_54_}), .c ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, LED_128_Instance_addconst_out[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U25 ( .a ({1'b0, 1'b0, roundconstant[1]}), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, LED_128_Instance_addroundkey_out_53_}), .c ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, LED_128_Instance_addconst_out[53]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U24 ( .a ({1'b0, 1'b0, roundconstant[0]}), .b ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, LED_128_Instance_addroundkey_out_52_}), .c ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, LED_128_Instance_addconst_out[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U23 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, LED_128_Instance_addroundkey_out_51_}), .c ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, LED_128_Instance_addconst_out[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U22 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, LED_128_Instance_addroundkey_out_50_}), .c ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, LED_128_Instance_addconst_out[50]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U21 ( .a ({1'b0, 1'b0, roundconstant[3]}), .b ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, LED_128_Instance_addroundkey_out_4_}), .c ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, LED_128_Instance_addconst_out[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U20 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, LED_128_Instance_addroundkey_out_49_}), .c ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, LED_128_Instance_addconst_out[49]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U19 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, LED_128_Instance_addroundkey_out_48_}), .c ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, LED_128_Instance_addconst_out[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U18 ( .a ({1'b0, 1'b0, 1'b1}), .b ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, LED_128_Instance_addroundkey_out_3_}), .c ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, LED_128_Instance_addconst_out[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U17 ( .a ({1'b0, 1'b0, roundconstant[5]}), .b ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, LED_128_Instance_addroundkey_out_38_}), .c ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, LED_128_Instance_addconst_out[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U16 ( .a ({1'b0, 1'b0, roundconstant[4]}), .b ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, LED_128_Instance_addroundkey_out_37_}), .c ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, LED_128_Instance_addconst_out[37]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U15 ( .a ({1'b0, 1'b0, roundconstant[3]}), .b ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, LED_128_Instance_addroundkey_out_36_}), .c ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, LED_128_Instance_addconst_out[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U14 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, LED_128_Instance_addroundkey_out_35_}), .c ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, LED_128_Instance_addconst_out[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U13 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, LED_128_Instance_addroundkey_out_34_}), .c ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, LED_128_Instance_addconst_out[34]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U12 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, LED_128_Instance_addroundkey_out_33_}), .c ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, LED_128_Instance_addconst_out[33]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U11 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, LED_128_Instance_addroundkey_out_32_}), .c ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, LED_128_Instance_addconst_out[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U10 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, LED_128_Instance_addroundkey_out_2_}), .c ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, LED_128_Instance_addconst_out[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U9 ( .a ({1'b0, 1'b0, roundconstant[2]}), .b ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, LED_128_Instance_addroundkey_out_22_}), .c ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_addconst_out[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U8 ( .a ({1'b0, 1'b0, roundconstant[1]}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, LED_128_Instance_addroundkey_out_21_}), .c ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, LED_128_Instance_addconst_out[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U7 ( .a ({1'b0, 1'b0, roundconstant[0]}), .b ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, LED_128_Instance_addroundkey_out_20_}), .c ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, LED_128_Instance_addconst_out[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U6 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, LED_128_Instance_addroundkey_out_1_}), .c ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, LED_128_Instance_addconst_out[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U5 ( .a ({1'b0, 1'b0, 1'b1}), .b ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, LED_128_Instance_addroundkey_out_19_}), .c ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, LED_128_Instance_addconst_out[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U4 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, LED_128_Instance_addroundkey_out_18_}), .c ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, LED_128_Instance_addconst_out[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U3 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, LED_128_Instance_addroundkey_out_17_}), .c ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, LED_128_Instance_addconst_out[17]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U2 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, LED_128_Instance_addroundkey_out_16_}), .c ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, LED_128_Instance_addconst_out[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_AddConstants_instance_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_1765, new_AGEMA_signal_1764, LED_128_Instance_addroundkey_out_0_}), .c ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, LED_128_Instance_addconst_out[0]}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_U3 ( .a ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, LED_128_Instance_SBox_Instance_0_L0}), .b ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, LED_128_Instance_SBox_Instance_0_n1}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_U2 ( .a ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, LED_128_Instance_addconst_out[3]}), .b ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, LED_128_Instance_SBox_Instance_0_n2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_U1 ( .a ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, LED_128_Instance_addconst_out[1]}), .b ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, LED_128_Instance_SBox_Instance_0_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR1_U1 ( .a ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, LED_128_Instance_addconst_out[2]}), .b ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, LED_128_Instance_addconst_out[1]}), .c ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, LED_128_Instance_SBox_Instance_0_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR2_U1 ( .a ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, LED_128_Instance_addconst_out[1]}), .b ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, LED_128_Instance_addconst_out[0]}), .c ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, LED_128_Instance_SBox_Instance_0_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR3_U1 ( .a ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, LED_128_Instance_SBox_Instance_0_L1}), .b ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, LED_128_Instance_addconst_out[3]}), .c ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, LED_128_Instance_SBox_Instance_0_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR4_U1 ( .a ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, LED_128_Instance_addconst_out[3]}), .b ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, LED_128_Instance_addconst_out[0]}), .c ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, LED_128_Instance_SBox_Instance_0_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR5_U1 ( .a ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, LED_128_Instance_SBox_Instance_0_L3}), .b ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, LED_128_Instance_SBox_Instance_0_L0}), .c ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, LED_128_Instance_SBox_Instance_0_Q3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR6_U1 ( .a ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, LED_128_Instance_addconst_out[3]}), .b ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, LED_128_Instance_addconst_out[1]}), .c ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, LED_128_Instance_SBox_Instance_0_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR9_U1 ( .a ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, LED_128_Instance_SBox_Instance_0_L1}), .b ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, LED_128_Instance_addconst_out[2]}), .c ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, LED_128_Instance_SBox_Instance_0_Q7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_U3 ( .a ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, LED_128_Instance_SBox_Instance_1_L0}), .b ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, LED_128_Instance_SBox_Instance_1_n1}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_U2 ( .a ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, LED_128_Instance_addconst_out[7]}), .b ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, LED_128_Instance_SBox_Instance_1_n2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_U1 ( .a ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, LED_128_Instance_addconst_out[5]}), .b ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, LED_128_Instance_SBox_Instance_1_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR1_U1 ( .a ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, LED_128_Instance_addconst_out[6]}), .b ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, LED_128_Instance_addconst_out[5]}), .c ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, LED_128_Instance_SBox_Instance_1_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR2_U1 ( .a ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, LED_128_Instance_addconst_out[5]}), .b ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, LED_128_Instance_addconst_out[4]}), .c ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, LED_128_Instance_SBox_Instance_1_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR3_U1 ( .a ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, LED_128_Instance_SBox_Instance_1_L1}), .b ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, LED_128_Instance_addconst_out[7]}), .c ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, LED_128_Instance_SBox_Instance_1_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR4_U1 ( .a ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, LED_128_Instance_addconst_out[7]}), .b ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, LED_128_Instance_addconst_out[4]}), .c ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, LED_128_Instance_SBox_Instance_1_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR5_U1 ( .a ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, LED_128_Instance_SBox_Instance_1_L3}), .b ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, LED_128_Instance_SBox_Instance_1_L0}), .c ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, LED_128_Instance_SBox_Instance_1_Q3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR6_U1 ( .a ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, LED_128_Instance_addconst_out[7]}), .b ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, LED_128_Instance_addconst_out[5]}), .c ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, LED_128_Instance_SBox_Instance_1_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR9_U1 ( .a ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, LED_128_Instance_SBox_Instance_1_L1}), .b ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, LED_128_Instance_addconst_out[6]}), .c ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, LED_128_Instance_SBox_Instance_1_Q7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_U3 ( .a ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, LED_128_Instance_SBox_Instance_2_L0}), .b ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, LED_128_Instance_SBox_Instance_2_n1}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_U2 ( .a ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, LED_128_Instance_addconst_out[11]}), .b ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, LED_128_Instance_SBox_Instance_2_n2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_U1 ( .a ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, LED_128_Instance_addconst_out[9]}), .b ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, LED_128_Instance_SBox_Instance_2_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR1_U1 ( .a ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, LED_128_Instance_addconst_out[10]}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, LED_128_Instance_addconst_out[9]}), .c ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, LED_128_Instance_SBox_Instance_2_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR2_U1 ( .a ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, LED_128_Instance_addconst_out[9]}), .b ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, LED_128_Instance_addconst_out[8]}), .c ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, LED_128_Instance_SBox_Instance_2_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR3_U1 ( .a ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, LED_128_Instance_SBox_Instance_2_L1}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, LED_128_Instance_addconst_out[11]}), .c ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, LED_128_Instance_SBox_Instance_2_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR4_U1 ( .a ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, LED_128_Instance_addconst_out[11]}), .b ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, LED_128_Instance_addconst_out[8]}), .c ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, LED_128_Instance_SBox_Instance_2_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR5_U1 ( .a ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, LED_128_Instance_SBox_Instance_2_L3}), .b ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, LED_128_Instance_SBox_Instance_2_L0}), .c ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, LED_128_Instance_SBox_Instance_2_Q3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR6_U1 ( .a ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, LED_128_Instance_addconst_out[11]}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, LED_128_Instance_addconst_out[9]}), .c ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, LED_128_Instance_SBox_Instance_2_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR9_U1 ( .a ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, LED_128_Instance_SBox_Instance_2_L1}), .b ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, LED_128_Instance_addconst_out[10]}), .c ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, LED_128_Instance_SBox_Instance_2_Q7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_U3 ( .a ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, LED_128_Instance_SBox_Instance_3_L0}), .b ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, LED_128_Instance_SBox_Instance_3_n1}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_U2 ( .a ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, LED_128_Instance_addconst_out[15]}), .b ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, LED_128_Instance_SBox_Instance_3_n2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_U1 ( .a ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, LED_128_Instance_addconst_out[13]}), .b ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, LED_128_Instance_SBox_Instance_3_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR1_U1 ( .a ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, LED_128_Instance_addconst_out[14]}), .b ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, LED_128_Instance_addconst_out[13]}), .c ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, LED_128_Instance_SBox_Instance_3_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR2_U1 ( .a ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, LED_128_Instance_addconst_out[13]}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, LED_128_Instance_addconst_out[12]}), .c ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, LED_128_Instance_SBox_Instance_3_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR3_U1 ( .a ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, LED_128_Instance_SBox_Instance_3_L1}), .b ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, LED_128_Instance_addconst_out[15]}), .c ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, LED_128_Instance_SBox_Instance_3_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR4_U1 ( .a ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, LED_128_Instance_addconst_out[15]}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, LED_128_Instance_addconst_out[12]}), .c ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, LED_128_Instance_SBox_Instance_3_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR5_U1 ( .a ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, LED_128_Instance_SBox_Instance_3_L3}), .b ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, LED_128_Instance_SBox_Instance_3_L0}), .c ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, LED_128_Instance_SBox_Instance_3_Q3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR6_U1 ( .a ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, LED_128_Instance_addconst_out[15]}), .b ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, LED_128_Instance_addconst_out[13]}), .c ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, LED_128_Instance_SBox_Instance_3_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR9_U1 ( .a ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, LED_128_Instance_SBox_Instance_3_L1}), .b ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, LED_128_Instance_addconst_out[14]}), .c ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, LED_128_Instance_SBox_Instance_3_Q7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_U3 ( .a ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, LED_128_Instance_SBox_Instance_4_L0}), .b ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, LED_128_Instance_SBox_Instance_4_n1}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_U2 ( .a ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, LED_128_Instance_addconst_out[19]}), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, LED_128_Instance_SBox_Instance_4_n2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_U1 ( .a ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, LED_128_Instance_addconst_out[17]}), .b ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, LED_128_Instance_SBox_Instance_4_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR1_U1 ( .a ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, LED_128_Instance_addconst_out[18]}), .b ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, LED_128_Instance_addconst_out[17]}), .c ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, LED_128_Instance_SBox_Instance_4_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR2_U1 ( .a ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, LED_128_Instance_addconst_out[17]}), .b ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, LED_128_Instance_addconst_out[16]}), .c ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, LED_128_Instance_SBox_Instance_4_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR3_U1 ( .a ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, LED_128_Instance_SBox_Instance_4_L1}), .b ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, LED_128_Instance_addconst_out[19]}), .c ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, LED_128_Instance_SBox_Instance_4_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR4_U1 ( .a ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, LED_128_Instance_addconst_out[19]}), .b ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, LED_128_Instance_addconst_out[16]}), .c ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, LED_128_Instance_SBox_Instance_4_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR5_U1 ( .a ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, LED_128_Instance_SBox_Instance_4_L3}), .b ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, LED_128_Instance_SBox_Instance_4_L0}), .c ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, LED_128_Instance_SBox_Instance_4_Q3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR6_U1 ( .a ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, LED_128_Instance_addconst_out[19]}), .b ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, LED_128_Instance_addconst_out[17]}), .c ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, LED_128_Instance_SBox_Instance_4_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR9_U1 ( .a ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, LED_128_Instance_SBox_Instance_4_L1}), .b ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, LED_128_Instance_addconst_out[18]}), .c ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, LED_128_Instance_SBox_Instance_4_Q7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_U3 ( .a ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, LED_128_Instance_SBox_Instance_5_L0}), .b ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, LED_128_Instance_SBox_Instance_5_n1}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_U2 ( .a ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, LED_128_Instance_addconst_out[23]}), .b ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, LED_128_Instance_SBox_Instance_5_n2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_U1 ( .a ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, LED_128_Instance_addconst_out[21]}), .b ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, LED_128_Instance_SBox_Instance_5_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR1_U1 ( .a ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_addconst_out[22]}), .b ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, LED_128_Instance_addconst_out[21]}), .c ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, LED_128_Instance_SBox_Instance_5_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR2_U1 ( .a ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, LED_128_Instance_addconst_out[21]}), .b ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, LED_128_Instance_addconst_out[20]}), .c ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, LED_128_Instance_SBox_Instance_5_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR3_U1 ( .a ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, LED_128_Instance_SBox_Instance_5_L1}), .b ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, LED_128_Instance_addconst_out[23]}), .c ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, LED_128_Instance_SBox_Instance_5_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR4_U1 ( .a ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, LED_128_Instance_addconst_out[23]}), .b ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, LED_128_Instance_addconst_out[20]}), .c ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, LED_128_Instance_SBox_Instance_5_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR5_U1 ( .a ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, LED_128_Instance_SBox_Instance_5_L3}), .b ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, LED_128_Instance_SBox_Instance_5_L0}), .c ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, LED_128_Instance_SBox_Instance_5_Q3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR6_U1 ( .a ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, LED_128_Instance_addconst_out[23]}), .b ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, LED_128_Instance_addconst_out[21]}), .c ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, LED_128_Instance_SBox_Instance_5_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR9_U1 ( .a ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, LED_128_Instance_SBox_Instance_5_L1}), .b ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_addconst_out[22]}), .c ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, LED_128_Instance_SBox_Instance_5_Q7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_U3 ( .a ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, LED_128_Instance_SBox_Instance_6_L0}), .b ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, LED_128_Instance_SBox_Instance_6_n1}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_U2 ( .a ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, LED_128_Instance_addconst_out[27]}), .b ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, LED_128_Instance_SBox_Instance_6_n2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_U1 ( .a ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, LED_128_Instance_addconst_out[25]}), .b ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, LED_128_Instance_SBox_Instance_6_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR1_U1 ( .a ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_addconst_out[26]}), .b ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, LED_128_Instance_addconst_out[25]}), .c ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, LED_128_Instance_SBox_Instance_6_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR2_U1 ( .a ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, LED_128_Instance_addconst_out[25]}), .b ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, LED_128_Instance_addconst_out[24]}), .c ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, LED_128_Instance_SBox_Instance_6_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR3_U1 ( .a ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, LED_128_Instance_SBox_Instance_6_L1}), .b ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, LED_128_Instance_addconst_out[27]}), .c ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, LED_128_Instance_SBox_Instance_6_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR4_U1 ( .a ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, LED_128_Instance_addconst_out[27]}), .b ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, LED_128_Instance_addconst_out[24]}), .c ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, LED_128_Instance_SBox_Instance_6_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR5_U1 ( .a ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, LED_128_Instance_SBox_Instance_6_L3}), .b ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, LED_128_Instance_SBox_Instance_6_L0}), .c ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, LED_128_Instance_SBox_Instance_6_Q3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR6_U1 ( .a ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, LED_128_Instance_addconst_out[27]}), .b ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, LED_128_Instance_addconst_out[25]}), .c ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, LED_128_Instance_SBox_Instance_6_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR9_U1 ( .a ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, LED_128_Instance_SBox_Instance_6_L1}), .b ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_addconst_out[26]}), .c ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, LED_128_Instance_SBox_Instance_6_Q7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_U3 ( .a ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, LED_128_Instance_SBox_Instance_7_L0}), .b ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, LED_128_Instance_SBox_Instance_7_n1}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_U2 ( .a ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, LED_128_Instance_addconst_out[31]}), .b ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, LED_128_Instance_SBox_Instance_7_n2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_U1 ( .a ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, LED_128_Instance_addconst_out[29]}), .b ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, LED_128_Instance_SBox_Instance_7_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR1_U1 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, LED_128_Instance_addconst_out[30]}), .b ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, LED_128_Instance_addconst_out[29]}), .c ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, LED_128_Instance_SBox_Instance_7_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR2_U1 ( .a ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, LED_128_Instance_addconst_out[29]}), .b ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, LED_128_Instance_addconst_out[28]}), .c ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, LED_128_Instance_SBox_Instance_7_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR3_U1 ( .a ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, LED_128_Instance_SBox_Instance_7_L1}), .b ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, LED_128_Instance_addconst_out[31]}), .c ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, LED_128_Instance_SBox_Instance_7_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR4_U1 ( .a ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, LED_128_Instance_addconst_out[31]}), .b ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, LED_128_Instance_addconst_out[28]}), .c ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, LED_128_Instance_SBox_Instance_7_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR5_U1 ( .a ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, LED_128_Instance_SBox_Instance_7_L3}), .b ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, LED_128_Instance_SBox_Instance_7_L0}), .c ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, LED_128_Instance_SBox_Instance_7_Q3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR6_U1 ( .a ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, LED_128_Instance_addconst_out[31]}), .b ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, LED_128_Instance_addconst_out[29]}), .c ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, LED_128_Instance_SBox_Instance_7_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR9_U1 ( .a ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, LED_128_Instance_SBox_Instance_7_L1}), .b ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, LED_128_Instance_addconst_out[30]}), .c ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, LED_128_Instance_SBox_Instance_7_Q7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_U3 ( .a ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, LED_128_Instance_SBox_Instance_8_L0}), .b ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, LED_128_Instance_SBox_Instance_8_n1}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_U2 ( .a ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, LED_128_Instance_addconst_out[35]}), .b ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, LED_128_Instance_SBox_Instance_8_n2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_U1 ( .a ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, LED_128_Instance_addconst_out[33]}), .b ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, LED_128_Instance_SBox_Instance_8_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR1_U1 ( .a ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, LED_128_Instance_addconst_out[34]}), .b ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, LED_128_Instance_addconst_out[33]}), .c ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, LED_128_Instance_SBox_Instance_8_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR2_U1 ( .a ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, LED_128_Instance_addconst_out[33]}), .b ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, LED_128_Instance_addconst_out[32]}), .c ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, LED_128_Instance_SBox_Instance_8_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR3_U1 ( .a ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, LED_128_Instance_SBox_Instance_8_L1}), .b ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, LED_128_Instance_addconst_out[35]}), .c ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, LED_128_Instance_SBox_Instance_8_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR4_U1 ( .a ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, LED_128_Instance_addconst_out[35]}), .b ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, LED_128_Instance_addconst_out[32]}), .c ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, LED_128_Instance_SBox_Instance_8_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR5_U1 ( .a ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, LED_128_Instance_SBox_Instance_8_L3}), .b ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, LED_128_Instance_SBox_Instance_8_L0}), .c ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, LED_128_Instance_SBox_Instance_8_Q3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR6_U1 ( .a ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, LED_128_Instance_addconst_out[35]}), .b ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, LED_128_Instance_addconst_out[33]}), .c ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, LED_128_Instance_SBox_Instance_8_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR9_U1 ( .a ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, LED_128_Instance_SBox_Instance_8_L1}), .b ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, LED_128_Instance_addconst_out[34]}), .c ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, LED_128_Instance_SBox_Instance_8_Q7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_U3 ( .a ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, LED_128_Instance_SBox_Instance_9_L0}), .b ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, LED_128_Instance_SBox_Instance_9_n1}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_U2 ( .a ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, LED_128_Instance_addconst_out[39]}), .b ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, LED_128_Instance_SBox_Instance_9_n2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_U1 ( .a ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, LED_128_Instance_addconst_out[37]}), .b ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, LED_128_Instance_SBox_Instance_9_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR1_U1 ( .a ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, LED_128_Instance_addconst_out[38]}), .b ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, LED_128_Instance_addconst_out[37]}), .c ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, LED_128_Instance_SBox_Instance_9_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR2_U1 ( .a ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, LED_128_Instance_addconst_out[37]}), .b ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, LED_128_Instance_addconst_out[36]}), .c ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, LED_128_Instance_SBox_Instance_9_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR3_U1 ( .a ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, LED_128_Instance_SBox_Instance_9_L1}), .b ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, LED_128_Instance_addconst_out[39]}), .c ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, LED_128_Instance_SBox_Instance_9_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR4_U1 ( .a ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, LED_128_Instance_addconst_out[39]}), .b ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, LED_128_Instance_addconst_out[36]}), .c ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, LED_128_Instance_SBox_Instance_9_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR5_U1 ( .a ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, LED_128_Instance_SBox_Instance_9_L3}), .b ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, LED_128_Instance_SBox_Instance_9_L0}), .c ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, LED_128_Instance_SBox_Instance_9_Q3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR6_U1 ( .a ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, LED_128_Instance_addconst_out[39]}), .b ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, LED_128_Instance_addconst_out[37]}), .c ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, LED_128_Instance_SBox_Instance_9_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR9_U1 ( .a ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, LED_128_Instance_SBox_Instance_9_L1}), .b ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, LED_128_Instance_addconst_out[38]}), .c ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, LED_128_Instance_SBox_Instance_9_Q7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_U3 ( .a ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, LED_128_Instance_SBox_Instance_10_L0}), .b ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, LED_128_Instance_SBox_Instance_10_n1}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_U2 ( .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, LED_128_Instance_addconst_out[43]}), .b ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, LED_128_Instance_SBox_Instance_10_n2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_U1 ( .a ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, LED_128_Instance_addconst_out[41]}), .b ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, LED_128_Instance_SBox_Instance_10_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR1_U1 ( .a ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, LED_128_Instance_addconst_out[42]}), .b ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, LED_128_Instance_addconst_out[41]}), .c ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, LED_128_Instance_SBox_Instance_10_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR2_U1 ( .a ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, LED_128_Instance_addconst_out[41]}), .b ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, LED_128_Instance_addconst_out[40]}), .c ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, LED_128_Instance_SBox_Instance_10_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR3_U1 ( .a ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, LED_128_Instance_SBox_Instance_10_L1}), .b ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, LED_128_Instance_addconst_out[43]}), .c ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, LED_128_Instance_SBox_Instance_10_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR4_U1 ( .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, LED_128_Instance_addconst_out[43]}), .b ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, LED_128_Instance_addconst_out[40]}), .c ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, LED_128_Instance_SBox_Instance_10_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR5_U1 ( .a ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, LED_128_Instance_SBox_Instance_10_L3}), .b ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, LED_128_Instance_SBox_Instance_10_L0}), .c ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, LED_128_Instance_SBox_Instance_10_Q3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR6_U1 ( .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, LED_128_Instance_addconst_out[43]}), .b ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, LED_128_Instance_addconst_out[41]}), .c ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, LED_128_Instance_SBox_Instance_10_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR9_U1 ( .a ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, LED_128_Instance_SBox_Instance_10_L1}), .b ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, LED_128_Instance_addconst_out[42]}), .c ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, LED_128_Instance_SBox_Instance_10_Q7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_U3 ( .a ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, LED_128_Instance_SBox_Instance_11_L0}), .b ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, LED_128_Instance_SBox_Instance_11_n1}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_U2 ( .a ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, LED_128_Instance_addconst_out[47]}), .b ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, LED_128_Instance_SBox_Instance_11_n2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_U1 ( .a ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, LED_128_Instance_addconst_out[45]}), .b ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, LED_128_Instance_SBox_Instance_11_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR1_U1 ( .a ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, LED_128_Instance_addconst_out[46]}), .b ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, LED_128_Instance_addconst_out[45]}), .c ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, LED_128_Instance_SBox_Instance_11_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR2_U1 ( .a ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, LED_128_Instance_addconst_out[45]}), .b ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, LED_128_Instance_addconst_out[44]}), .c ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, LED_128_Instance_SBox_Instance_11_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR3_U1 ( .a ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, LED_128_Instance_SBox_Instance_11_L1}), .b ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, LED_128_Instance_addconst_out[47]}), .c ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, LED_128_Instance_SBox_Instance_11_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR4_U1 ( .a ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, LED_128_Instance_addconst_out[47]}), .b ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, LED_128_Instance_addconst_out[44]}), .c ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, LED_128_Instance_SBox_Instance_11_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR5_U1 ( .a ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, LED_128_Instance_SBox_Instance_11_L3}), .b ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, LED_128_Instance_SBox_Instance_11_L0}), .c ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, LED_128_Instance_SBox_Instance_11_Q3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR6_U1 ( .a ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, LED_128_Instance_addconst_out[47]}), .b ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, LED_128_Instance_addconst_out[45]}), .c ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, LED_128_Instance_SBox_Instance_11_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR9_U1 ( .a ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, LED_128_Instance_SBox_Instance_11_L1}), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, LED_128_Instance_addconst_out[46]}), .c ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, LED_128_Instance_SBox_Instance_11_Q7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_U3 ( .a ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, LED_128_Instance_SBox_Instance_12_L0}), .b ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, LED_128_Instance_SBox_Instance_12_n1}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_U2 ( .a ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, LED_128_Instance_addconst_out[51]}), .b ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, LED_128_Instance_SBox_Instance_12_n2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_U1 ( .a ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, LED_128_Instance_addconst_out[49]}), .b ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, LED_128_Instance_SBox_Instance_12_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR1_U1 ( .a ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, LED_128_Instance_addconst_out[50]}), .b ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, LED_128_Instance_addconst_out[49]}), .c ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, LED_128_Instance_SBox_Instance_12_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR2_U1 ( .a ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, LED_128_Instance_addconst_out[49]}), .b ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, LED_128_Instance_addconst_out[48]}), .c ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, LED_128_Instance_SBox_Instance_12_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR3_U1 ( .a ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, LED_128_Instance_SBox_Instance_12_L1}), .b ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, LED_128_Instance_addconst_out[51]}), .c ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, LED_128_Instance_SBox_Instance_12_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR4_U1 ( .a ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, LED_128_Instance_addconst_out[51]}), .b ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, LED_128_Instance_addconst_out[48]}), .c ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, LED_128_Instance_SBox_Instance_12_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR5_U1 ( .a ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, LED_128_Instance_SBox_Instance_12_L3}), .b ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, LED_128_Instance_SBox_Instance_12_L0}), .c ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, LED_128_Instance_SBox_Instance_12_Q3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR6_U1 ( .a ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, LED_128_Instance_addconst_out[51]}), .b ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, LED_128_Instance_addconst_out[49]}), .c ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, LED_128_Instance_SBox_Instance_12_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR9_U1 ( .a ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, LED_128_Instance_SBox_Instance_12_L1}), .b ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, LED_128_Instance_addconst_out[50]}), .c ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, LED_128_Instance_SBox_Instance_12_Q7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_U3 ( .a ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, LED_128_Instance_SBox_Instance_13_L0}), .b ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, LED_128_Instance_SBox_Instance_13_n1}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_U2 ( .a ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, LED_128_Instance_addconst_out[55]}), .b ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, LED_128_Instance_SBox_Instance_13_n2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_U1 ( .a ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, LED_128_Instance_addconst_out[53]}), .b ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, LED_128_Instance_SBox_Instance_13_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR1_U1 ( .a ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, LED_128_Instance_addconst_out[54]}), .b ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, LED_128_Instance_addconst_out[53]}), .c ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, LED_128_Instance_SBox_Instance_13_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR2_U1 ( .a ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, LED_128_Instance_addconst_out[53]}), .b ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, LED_128_Instance_addconst_out[52]}), .c ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, LED_128_Instance_SBox_Instance_13_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR3_U1 ( .a ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, LED_128_Instance_SBox_Instance_13_L1}), .b ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, LED_128_Instance_addconst_out[55]}), .c ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, LED_128_Instance_SBox_Instance_13_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR4_U1 ( .a ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, LED_128_Instance_addconst_out[55]}), .b ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, LED_128_Instance_addconst_out[52]}), .c ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, LED_128_Instance_SBox_Instance_13_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR5_U1 ( .a ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, LED_128_Instance_SBox_Instance_13_L3}), .b ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, LED_128_Instance_SBox_Instance_13_L0}), .c ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, LED_128_Instance_SBox_Instance_13_Q3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR6_U1 ( .a ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, LED_128_Instance_addconst_out[55]}), .b ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, LED_128_Instance_addconst_out[53]}), .c ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, LED_128_Instance_SBox_Instance_13_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR9_U1 ( .a ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, LED_128_Instance_SBox_Instance_13_L1}), .b ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, LED_128_Instance_addconst_out[54]}), .c ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, LED_128_Instance_SBox_Instance_13_Q7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_U3 ( .a ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, LED_128_Instance_SBox_Instance_14_L0}), .b ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, LED_128_Instance_SBox_Instance_14_n1}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_U2 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, LED_128_Instance_addconst_out[59]}), .b ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, LED_128_Instance_SBox_Instance_14_n2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_U1 ( .a ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, LED_128_Instance_addconst_out[57]}), .b ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, LED_128_Instance_SBox_Instance_14_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR1_U1 ( .a ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, LED_128_Instance_addconst_out[58]}), .b ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, LED_128_Instance_addconst_out[57]}), .c ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, LED_128_Instance_SBox_Instance_14_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR2_U1 ( .a ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, LED_128_Instance_addconst_out[57]}), .b ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, LED_128_Instance_addconst_out[56]}), .c ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, LED_128_Instance_SBox_Instance_14_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR3_U1 ( .a ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, LED_128_Instance_SBox_Instance_14_L1}), .b ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, LED_128_Instance_addconst_out[59]}), .c ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, LED_128_Instance_SBox_Instance_14_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR4_U1 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, LED_128_Instance_addconst_out[59]}), .b ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, LED_128_Instance_addconst_out[56]}), .c ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, LED_128_Instance_SBox_Instance_14_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR5_U1 ( .a ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, LED_128_Instance_SBox_Instance_14_L3}), .b ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, LED_128_Instance_SBox_Instance_14_L0}), .c ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, LED_128_Instance_SBox_Instance_14_Q3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR6_U1 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, LED_128_Instance_addconst_out[59]}), .b ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, LED_128_Instance_addconst_out[57]}), .c ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, LED_128_Instance_SBox_Instance_14_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR9_U1 ( .a ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, LED_128_Instance_SBox_Instance_14_L1}), .b ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, LED_128_Instance_addconst_out[58]}), .c ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, LED_128_Instance_SBox_Instance_14_Q7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_U3 ( .a ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, LED_128_Instance_SBox_Instance_15_L0}), .b ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, LED_128_Instance_SBox_Instance_15_n1}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_U2 ( .a ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, LED_128_Instance_addconst_out[63]}), .b ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, LED_128_Instance_SBox_Instance_15_n2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_U1 ( .a ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, LED_128_Instance_addconst_out[61]}), .b ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, LED_128_Instance_SBox_Instance_15_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR1_U1 ( .a ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, LED_128_Instance_addconst_out[62]}), .b ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, LED_128_Instance_addconst_out[61]}), .c ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, LED_128_Instance_SBox_Instance_15_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR2_U1 ( .a ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, LED_128_Instance_addconst_out[61]}), .b ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, LED_128_Instance_addconst_out[60]}), .c ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, LED_128_Instance_SBox_Instance_15_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR3_U1 ( .a ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, LED_128_Instance_SBox_Instance_15_L1}), .b ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, LED_128_Instance_addconst_out[63]}), .c ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, LED_128_Instance_SBox_Instance_15_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR4_U1 ( .a ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, LED_128_Instance_addconst_out[63]}), .b ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, LED_128_Instance_addconst_out[60]}), .c ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, LED_128_Instance_SBox_Instance_15_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR5_U1 ( .a ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, LED_128_Instance_SBox_Instance_15_L3}), .b ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, LED_128_Instance_SBox_Instance_15_L0}), .c ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, LED_128_Instance_SBox_Instance_15_Q3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR6_U1 ( .a ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, LED_128_Instance_addconst_out[63]}), .b ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, LED_128_Instance_addconst_out[61]}), .c ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, LED_128_Instance_SBox_Instance_15_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR9_U1 ( .a ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, LED_128_Instance_SBox_Instance_15_L1}), .b ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, LED_128_Instance_addconst_out[62]}), .c ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, LED_128_Instance_SBox_Instance_15_Q7}) ) ;
    INV_X1 LED_128_Instance_ks_reg_0__U1 ( .A (LED_128_Instance_ks_reg_0__Q), .ZN (LED_128_Instance_n4) ) ;
    INV_X1 LED_128_Instance_ks_reg_1__U1 ( .A (LED_128_Instance_n26), .ZN (LED_128_Instance_n8) ) ;
    INV_X1 LED_128_Instance_ks_reg_2__U1 ( .A (LED_128_Instance_n25), .ZN (LED_128_Instance_n1) ) ;
    INV_X1 LED_128_Instance_ks_reg_3__U1 ( .A (LED_128_Instance_n2), .ZN (LED_128_Instance_n24) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_0__U1 ( .A (roundconstant[0]), .ZN (LED_128_Instance_n6) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_1__U1 ( .A (roundconstant[1]), .ZN (LED_128_Instance_n29) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_2__U1 ( .A (roundconstant[2]), .ZN (LED_128_Instance_n5) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_3__U1 ( .A (roundconstant[3]), .ZN (LED_128_Instance_n30) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_4__U1 ( .A (roundconstant[4]), .ZN (LED_128_Instance_n28) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_5__U1 ( .A (roundconstant[5]), .ZN (LED_128_Instance_n27) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_1128 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_0_L2), .Q (new_AGEMA_signal_3896) ) ;
    buf_clk new_AGEMA_reg_buffer_1130 ( .C (CLK), .D (new_AGEMA_signal_2426), .Q (new_AGEMA_signal_3898) ) ;
    buf_clk new_AGEMA_reg_buffer_1132 ( .C (CLK), .D (new_AGEMA_signal_2427), .Q (new_AGEMA_signal_3900) ) ;
    buf_clk new_AGEMA_reg_buffer_1134 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_0_L4), .Q (new_AGEMA_signal_3902) ) ;
    buf_clk new_AGEMA_reg_buffer_1136 ( .C (CLK), .D (new_AGEMA_signal_2276), .Q (new_AGEMA_signal_3904) ) ;
    buf_clk new_AGEMA_reg_buffer_1138 ( .C (CLK), .D (new_AGEMA_signal_2277), .Q (new_AGEMA_signal_3906) ) ;
    buf_clk new_AGEMA_reg_buffer_1140 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_0_L3), .Q (new_AGEMA_signal_3908) ) ;
    buf_clk new_AGEMA_reg_buffer_1142 ( .C (CLK), .D (new_AGEMA_signal_2116), .Q (new_AGEMA_signal_3910) ) ;
    buf_clk new_AGEMA_reg_buffer_1144 ( .C (CLK), .D (new_AGEMA_signal_2117), .Q (new_AGEMA_signal_3912) ) ;
    buf_clk new_AGEMA_reg_buffer_1146 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_1_L2), .Q (new_AGEMA_signal_3914) ) ;
    buf_clk new_AGEMA_reg_buffer_1148 ( .C (CLK), .D (new_AGEMA_signal_2436), .Q (new_AGEMA_signal_3916) ) ;
    buf_clk new_AGEMA_reg_buffer_1150 ( .C (CLK), .D (new_AGEMA_signal_2437), .Q (new_AGEMA_signal_3918) ) ;
    buf_clk new_AGEMA_reg_buffer_1152 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_1_L4), .Q (new_AGEMA_signal_3920) ) ;
    buf_clk new_AGEMA_reg_buffer_1154 ( .C (CLK), .D (new_AGEMA_signal_2286), .Q (new_AGEMA_signal_3922) ) ;
    buf_clk new_AGEMA_reg_buffer_1156 ( .C (CLK), .D (new_AGEMA_signal_2287), .Q (new_AGEMA_signal_3924) ) ;
    buf_clk new_AGEMA_reg_buffer_1158 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_1_L3), .Q (new_AGEMA_signal_3926) ) ;
    buf_clk new_AGEMA_reg_buffer_1160 ( .C (CLK), .D (new_AGEMA_signal_2284), .Q (new_AGEMA_signal_3928) ) ;
    buf_clk new_AGEMA_reg_buffer_1162 ( .C (CLK), .D (new_AGEMA_signal_2285), .Q (new_AGEMA_signal_3930) ) ;
    buf_clk new_AGEMA_reg_buffer_1164 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_2_L2), .Q (new_AGEMA_signal_3932) ) ;
    buf_clk new_AGEMA_reg_buffer_1166 ( .C (CLK), .D (new_AGEMA_signal_2290), .Q (new_AGEMA_signal_3934) ) ;
    buf_clk new_AGEMA_reg_buffer_1168 ( .C (CLK), .D (new_AGEMA_signal_2291), .Q (new_AGEMA_signal_3936) ) ;
    buf_clk new_AGEMA_reg_buffer_1170 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_2_L4), .Q (new_AGEMA_signal_3938) ) ;
    buf_clk new_AGEMA_reg_buffer_1172 ( .C (CLK), .D (new_AGEMA_signal_2174), .Q (new_AGEMA_signal_3940) ) ;
    buf_clk new_AGEMA_reg_buffer_1174 ( .C (CLK), .D (new_AGEMA_signal_2175), .Q (new_AGEMA_signal_3942) ) ;
    buf_clk new_AGEMA_reg_buffer_1176 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_2_L3), .Q (new_AGEMA_signal_3944) ) ;
    buf_clk new_AGEMA_reg_buffer_1178 ( .C (CLK), .D (new_AGEMA_signal_2172), .Q (new_AGEMA_signal_3946) ) ;
    buf_clk new_AGEMA_reg_buffer_1180 ( .C (CLK), .D (new_AGEMA_signal_2173), .Q (new_AGEMA_signal_3948) ) ;
    buf_clk new_AGEMA_reg_buffer_1182 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_3_L2), .Q (new_AGEMA_signal_3950) ) ;
    buf_clk new_AGEMA_reg_buffer_1184 ( .C (CLK), .D (new_AGEMA_signal_2300), .Q (new_AGEMA_signal_3952) ) ;
    buf_clk new_AGEMA_reg_buffer_1186 ( .C (CLK), .D (new_AGEMA_signal_2301), .Q (new_AGEMA_signal_3954) ) ;
    buf_clk new_AGEMA_reg_buffer_1188 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_3_L4), .Q (new_AGEMA_signal_3956) ) ;
    buf_clk new_AGEMA_reg_buffer_1190 ( .C (CLK), .D (new_AGEMA_signal_2186), .Q (new_AGEMA_signal_3958) ) ;
    buf_clk new_AGEMA_reg_buffer_1192 ( .C (CLK), .D (new_AGEMA_signal_2187), .Q (new_AGEMA_signal_3960) ) ;
    buf_clk new_AGEMA_reg_buffer_1194 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_3_L3), .Q (new_AGEMA_signal_3962) ) ;
    buf_clk new_AGEMA_reg_buffer_1196 ( .C (CLK), .D (new_AGEMA_signal_2184), .Q (new_AGEMA_signal_3964) ) ;
    buf_clk new_AGEMA_reg_buffer_1198 ( .C (CLK), .D (new_AGEMA_signal_2185), .Q (new_AGEMA_signal_3966) ) ;
    buf_clk new_AGEMA_reg_buffer_1200 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_4_L2), .Q (new_AGEMA_signal_3968) ) ;
    buf_clk new_AGEMA_reg_buffer_1202 ( .C (CLK), .D (new_AGEMA_signal_2454), .Q (new_AGEMA_signal_3970) ) ;
    buf_clk new_AGEMA_reg_buffer_1204 ( .C (CLK), .D (new_AGEMA_signal_2455), .Q (new_AGEMA_signal_3972) ) ;
    buf_clk new_AGEMA_reg_buffer_1206 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_4_L4), .Q (new_AGEMA_signal_3974) ) ;
    buf_clk new_AGEMA_reg_buffer_1208 ( .C (CLK), .D (new_AGEMA_signal_2314), .Q (new_AGEMA_signal_3976) ) ;
    buf_clk new_AGEMA_reg_buffer_1210 ( .C (CLK), .D (new_AGEMA_signal_2315), .Q (new_AGEMA_signal_3978) ) ;
    buf_clk new_AGEMA_reg_buffer_1212 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_4_L3), .Q (new_AGEMA_signal_3980) ) ;
    buf_clk new_AGEMA_reg_buffer_1214 ( .C (CLK), .D (new_AGEMA_signal_2120), .Q (new_AGEMA_signal_3982) ) ;
    buf_clk new_AGEMA_reg_buffer_1216 ( .C (CLK), .D (new_AGEMA_signal_2121), .Q (new_AGEMA_signal_3984) ) ;
    buf_clk new_AGEMA_reg_buffer_1218 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_5_L2), .Q (new_AGEMA_signal_3986) ) ;
    buf_clk new_AGEMA_reg_buffer_1220 ( .C (CLK), .D (new_AGEMA_signal_2464), .Q (new_AGEMA_signal_3988) ) ;
    buf_clk new_AGEMA_reg_buffer_1222 ( .C (CLK), .D (new_AGEMA_signal_2465), .Q (new_AGEMA_signal_3990) ) ;
    buf_clk new_AGEMA_reg_buffer_1224 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_5_L4), .Q (new_AGEMA_signal_3992) ) ;
    buf_clk new_AGEMA_reg_buffer_1226 ( .C (CLK), .D (new_AGEMA_signal_2324), .Q (new_AGEMA_signal_3994) ) ;
    buf_clk new_AGEMA_reg_buffer_1228 ( .C (CLK), .D (new_AGEMA_signal_2325), .Q (new_AGEMA_signal_3996) ) ;
    buf_clk new_AGEMA_reg_buffer_1230 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_5_L3), .Q (new_AGEMA_signal_3998) ) ;
    buf_clk new_AGEMA_reg_buffer_1232 ( .C (CLK), .D (new_AGEMA_signal_2322), .Q (new_AGEMA_signal_4000) ) ;
    buf_clk new_AGEMA_reg_buffer_1234 ( .C (CLK), .D (new_AGEMA_signal_2323), .Q (new_AGEMA_signal_4002) ) ;
    buf_clk new_AGEMA_reg_buffer_1236 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_6_L2), .Q (new_AGEMA_signal_4004) ) ;
    buf_clk new_AGEMA_reg_buffer_1238 ( .C (CLK), .D (new_AGEMA_signal_2328), .Q (new_AGEMA_signal_4006) ) ;
    buf_clk new_AGEMA_reg_buffer_1240 ( .C (CLK), .D (new_AGEMA_signal_2329), .Q (new_AGEMA_signal_4008) ) ;
    buf_clk new_AGEMA_reg_buffer_1242 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_6_L4), .Q (new_AGEMA_signal_4010) ) ;
    buf_clk new_AGEMA_reg_buffer_1244 ( .C (CLK), .D (new_AGEMA_signal_2200), .Q (new_AGEMA_signal_4012) ) ;
    buf_clk new_AGEMA_reg_buffer_1246 ( .C (CLK), .D (new_AGEMA_signal_2201), .Q (new_AGEMA_signal_4014) ) ;
    buf_clk new_AGEMA_reg_buffer_1248 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_6_L3), .Q (new_AGEMA_signal_4016) ) ;
    buf_clk new_AGEMA_reg_buffer_1250 ( .C (CLK), .D (new_AGEMA_signal_2198), .Q (new_AGEMA_signal_4018) ) ;
    buf_clk new_AGEMA_reg_buffer_1252 ( .C (CLK), .D (new_AGEMA_signal_2199), .Q (new_AGEMA_signal_4020) ) ;
    buf_clk new_AGEMA_reg_buffer_1254 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_7_L2), .Q (new_AGEMA_signal_4022) ) ;
    buf_clk new_AGEMA_reg_buffer_1256 ( .C (CLK), .D (new_AGEMA_signal_2338), .Q (new_AGEMA_signal_4024) ) ;
    buf_clk new_AGEMA_reg_buffer_1258 ( .C (CLK), .D (new_AGEMA_signal_2339), .Q (new_AGEMA_signal_4026) ) ;
    buf_clk new_AGEMA_reg_buffer_1260 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_7_L4), .Q (new_AGEMA_signal_4028) ) ;
    buf_clk new_AGEMA_reg_buffer_1262 ( .C (CLK), .D (new_AGEMA_signal_2212), .Q (new_AGEMA_signal_4030) ) ;
    buf_clk new_AGEMA_reg_buffer_1264 ( .C (CLK), .D (new_AGEMA_signal_2213), .Q (new_AGEMA_signal_4032) ) ;
    buf_clk new_AGEMA_reg_buffer_1266 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_7_L3), .Q (new_AGEMA_signal_4034) ) ;
    buf_clk new_AGEMA_reg_buffer_1268 ( .C (CLK), .D (new_AGEMA_signal_2210), .Q (new_AGEMA_signal_4036) ) ;
    buf_clk new_AGEMA_reg_buffer_1270 ( .C (CLK), .D (new_AGEMA_signal_2211), .Q (new_AGEMA_signal_4038) ) ;
    buf_clk new_AGEMA_reg_buffer_1272 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_8_L2), .Q (new_AGEMA_signal_4040) ) ;
    buf_clk new_AGEMA_reg_buffer_1274 ( .C (CLK), .D (new_AGEMA_signal_2482), .Q (new_AGEMA_signal_4042) ) ;
    buf_clk new_AGEMA_reg_buffer_1276 ( .C (CLK), .D (new_AGEMA_signal_2483), .Q (new_AGEMA_signal_4044) ) ;
    buf_clk new_AGEMA_reg_buffer_1278 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_8_L4), .Q (new_AGEMA_signal_4046) ) ;
    buf_clk new_AGEMA_reg_buffer_1280 ( .C (CLK), .D (new_AGEMA_signal_2352), .Q (new_AGEMA_signal_4048) ) ;
    buf_clk new_AGEMA_reg_buffer_1282 ( .C (CLK), .D (new_AGEMA_signal_2353), .Q (new_AGEMA_signal_4050) ) ;
    buf_clk new_AGEMA_reg_buffer_1284 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_8_L3), .Q (new_AGEMA_signal_4052) ) ;
    buf_clk new_AGEMA_reg_buffer_1286 ( .C (CLK), .D (new_AGEMA_signal_2216), .Q (new_AGEMA_signal_4054) ) ;
    buf_clk new_AGEMA_reg_buffer_1288 ( .C (CLK), .D (new_AGEMA_signal_2217), .Q (new_AGEMA_signal_4056) ) ;
    buf_clk new_AGEMA_reg_buffer_1290 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_9_L2), .Q (new_AGEMA_signal_4058) ) ;
    buf_clk new_AGEMA_reg_buffer_1292 ( .C (CLK), .D (new_AGEMA_signal_2492), .Q (new_AGEMA_signal_4060) ) ;
    buf_clk new_AGEMA_reg_buffer_1294 ( .C (CLK), .D (new_AGEMA_signal_2493), .Q (new_AGEMA_signal_4062) ) ;
    buf_clk new_AGEMA_reg_buffer_1296 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_9_L4), .Q (new_AGEMA_signal_4064) ) ;
    buf_clk new_AGEMA_reg_buffer_1298 ( .C (CLK), .D (new_AGEMA_signal_2360), .Q (new_AGEMA_signal_4066) ) ;
    buf_clk new_AGEMA_reg_buffer_1300 ( .C (CLK), .D (new_AGEMA_signal_2361), .Q (new_AGEMA_signal_4068) ) ;
    buf_clk new_AGEMA_reg_buffer_1302 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_9_L3), .Q (new_AGEMA_signal_4070) ) ;
    buf_clk new_AGEMA_reg_buffer_1304 ( .C (CLK), .D (new_AGEMA_signal_2218), .Q (new_AGEMA_signal_4072) ) ;
    buf_clk new_AGEMA_reg_buffer_1306 ( .C (CLK), .D (new_AGEMA_signal_2219), .Q (new_AGEMA_signal_4074) ) ;
    buf_clk new_AGEMA_reg_buffer_1308 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_10_L2), .Q (new_AGEMA_signal_4076) ) ;
    buf_clk new_AGEMA_reg_buffer_1310 ( .C (CLK), .D (new_AGEMA_signal_2364), .Q (new_AGEMA_signal_4078) ) ;
    buf_clk new_AGEMA_reg_buffer_1312 ( .C (CLK), .D (new_AGEMA_signal_2365), .Q (new_AGEMA_signal_4080) ) ;
    buf_clk new_AGEMA_reg_buffer_1314 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_10_L4), .Q (new_AGEMA_signal_4082) ) ;
    buf_clk new_AGEMA_reg_buffer_1316 ( .C (CLK), .D (new_AGEMA_signal_2230), .Q (new_AGEMA_signal_4084) ) ;
    buf_clk new_AGEMA_reg_buffer_1318 ( .C (CLK), .D (new_AGEMA_signal_2231), .Q (new_AGEMA_signal_4086) ) ;
    buf_clk new_AGEMA_reg_buffer_1320 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_10_L3), .Q (new_AGEMA_signal_4088) ) ;
    buf_clk new_AGEMA_reg_buffer_1322 ( .C (CLK), .D (new_AGEMA_signal_2228), .Q (new_AGEMA_signal_4090) ) ;
    buf_clk new_AGEMA_reg_buffer_1324 ( .C (CLK), .D (new_AGEMA_signal_2229), .Q (new_AGEMA_signal_4092) ) ;
    buf_clk new_AGEMA_reg_buffer_1326 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_11_L2), .Q (new_AGEMA_signal_4094) ) ;
    buf_clk new_AGEMA_reg_buffer_1328 ( .C (CLK), .D (new_AGEMA_signal_2374), .Q (new_AGEMA_signal_4096) ) ;
    buf_clk new_AGEMA_reg_buffer_1330 ( .C (CLK), .D (new_AGEMA_signal_2375), .Q (new_AGEMA_signal_4098) ) ;
    buf_clk new_AGEMA_reg_buffer_1332 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_11_L4), .Q (new_AGEMA_signal_4100) ) ;
    buf_clk new_AGEMA_reg_buffer_1334 ( .C (CLK), .D (new_AGEMA_signal_2242), .Q (new_AGEMA_signal_4102) ) ;
    buf_clk new_AGEMA_reg_buffer_1336 ( .C (CLK), .D (new_AGEMA_signal_2243), .Q (new_AGEMA_signal_4104) ) ;
    buf_clk new_AGEMA_reg_buffer_1338 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_11_L3), .Q (new_AGEMA_signal_4106) ) ;
    buf_clk new_AGEMA_reg_buffer_1340 ( .C (CLK), .D (new_AGEMA_signal_2240), .Q (new_AGEMA_signal_4108) ) ;
    buf_clk new_AGEMA_reg_buffer_1342 ( .C (CLK), .D (new_AGEMA_signal_2241), .Q (new_AGEMA_signal_4110) ) ;
    buf_clk new_AGEMA_reg_buffer_1344 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_12_L2), .Q (new_AGEMA_signal_4112) ) ;
    buf_clk new_AGEMA_reg_buffer_1346 ( .C (CLK), .D (new_AGEMA_signal_2510), .Q (new_AGEMA_signal_4114) ) ;
    buf_clk new_AGEMA_reg_buffer_1348 ( .C (CLK), .D (new_AGEMA_signal_2511), .Q (new_AGEMA_signal_4116) ) ;
    buf_clk new_AGEMA_reg_buffer_1350 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_12_L4), .Q (new_AGEMA_signal_4118) ) ;
    buf_clk new_AGEMA_reg_buffer_1352 ( .C (CLK), .D (new_AGEMA_signal_2392), .Q (new_AGEMA_signal_4120) ) ;
    buf_clk new_AGEMA_reg_buffer_1354 ( .C (CLK), .D (new_AGEMA_signal_2393), .Q (new_AGEMA_signal_4122) ) ;
    buf_clk new_AGEMA_reg_buffer_1356 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_12_L3), .Q (new_AGEMA_signal_4124) ) ;
    buf_clk new_AGEMA_reg_buffer_1358 ( .C (CLK), .D (new_AGEMA_signal_2390), .Q (new_AGEMA_signal_4126) ) ;
    buf_clk new_AGEMA_reg_buffer_1360 ( .C (CLK), .D (new_AGEMA_signal_2391), .Q (new_AGEMA_signal_4128) ) ;
    buf_clk new_AGEMA_reg_buffer_1362 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_13_L2), .Q (new_AGEMA_signal_4130) ) ;
    buf_clk new_AGEMA_reg_buffer_1364 ( .C (CLK), .D (new_AGEMA_signal_2520), .Q (new_AGEMA_signal_4132) ) ;
    buf_clk new_AGEMA_reg_buffer_1366 ( .C (CLK), .D (new_AGEMA_signal_2521), .Q (new_AGEMA_signal_4134) ) ;
    buf_clk new_AGEMA_reg_buffer_1368 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_13_L4), .Q (new_AGEMA_signal_4136) ) ;
    buf_clk new_AGEMA_reg_buffer_1370 ( .C (CLK), .D (new_AGEMA_signal_2402), .Q (new_AGEMA_signal_4138) ) ;
    buf_clk new_AGEMA_reg_buffer_1372 ( .C (CLK), .D (new_AGEMA_signal_2403), .Q (new_AGEMA_signal_4140) ) ;
    buf_clk new_AGEMA_reg_buffer_1374 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_13_L3), .Q (new_AGEMA_signal_4142) ) ;
    buf_clk new_AGEMA_reg_buffer_1376 ( .C (CLK), .D (new_AGEMA_signal_2400), .Q (new_AGEMA_signal_4144) ) ;
    buf_clk new_AGEMA_reg_buffer_1378 ( .C (CLK), .D (new_AGEMA_signal_2401), .Q (new_AGEMA_signal_4146) ) ;
    buf_clk new_AGEMA_reg_buffer_1380 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_14_L2), .Q (new_AGEMA_signal_4148) ) ;
    buf_clk new_AGEMA_reg_buffer_1382 ( .C (CLK), .D (new_AGEMA_signal_2406), .Q (new_AGEMA_signal_4150) ) ;
    buf_clk new_AGEMA_reg_buffer_1384 ( .C (CLK), .D (new_AGEMA_signal_2407), .Q (new_AGEMA_signal_4152) ) ;
    buf_clk new_AGEMA_reg_buffer_1386 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_14_L4), .Q (new_AGEMA_signal_4154) ) ;
    buf_clk new_AGEMA_reg_buffer_1388 ( .C (CLK), .D (new_AGEMA_signal_2256), .Q (new_AGEMA_signal_4156) ) ;
    buf_clk new_AGEMA_reg_buffer_1390 ( .C (CLK), .D (new_AGEMA_signal_2257), .Q (new_AGEMA_signal_4158) ) ;
    buf_clk new_AGEMA_reg_buffer_1392 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_14_L3), .Q (new_AGEMA_signal_4160) ) ;
    buf_clk new_AGEMA_reg_buffer_1394 ( .C (CLK), .D (new_AGEMA_signal_2254), .Q (new_AGEMA_signal_4162) ) ;
    buf_clk new_AGEMA_reg_buffer_1396 ( .C (CLK), .D (new_AGEMA_signal_2255), .Q (new_AGEMA_signal_4164) ) ;
    buf_clk new_AGEMA_reg_buffer_1398 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_15_L2), .Q (new_AGEMA_signal_4166) ) ;
    buf_clk new_AGEMA_reg_buffer_1400 ( .C (CLK), .D (new_AGEMA_signal_2416), .Q (new_AGEMA_signal_4168) ) ;
    buf_clk new_AGEMA_reg_buffer_1402 ( .C (CLK), .D (new_AGEMA_signal_2417), .Q (new_AGEMA_signal_4170) ) ;
    buf_clk new_AGEMA_reg_buffer_1404 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_15_L4), .Q (new_AGEMA_signal_4172) ) ;
    buf_clk new_AGEMA_reg_buffer_1406 ( .C (CLK), .D (new_AGEMA_signal_2268), .Q (new_AGEMA_signal_4174) ) ;
    buf_clk new_AGEMA_reg_buffer_1408 ( .C (CLK), .D (new_AGEMA_signal_2269), .Q (new_AGEMA_signal_4176) ) ;
    buf_clk new_AGEMA_reg_buffer_1410 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_15_L3), .Q (new_AGEMA_signal_4178) ) ;
    buf_clk new_AGEMA_reg_buffer_1412 ( .C (CLK), .D (new_AGEMA_signal_2266), .Q (new_AGEMA_signal_4180) ) ;
    buf_clk new_AGEMA_reg_buffer_1414 ( .C (CLK), .D (new_AGEMA_signal_2267), .Q (new_AGEMA_signal_4182) ) ;
    buf_clk new_AGEMA_reg_buffer_1416 ( .C (CLK), .D (LED_128_Instance_MUX_state0_n9), .Q (new_AGEMA_signal_4184) ) ;
    buf_clk new_AGEMA_reg_buffer_1420 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_0_), .Q (new_AGEMA_signal_4188) ) ;
    buf_clk new_AGEMA_reg_buffer_1424 ( .C (CLK), .D (new_AGEMA_signal_1764), .Q (new_AGEMA_signal_4192) ) ;
    buf_clk new_AGEMA_reg_buffer_1428 ( .C (CLK), .D (new_AGEMA_signal_1765), .Q (new_AGEMA_signal_4196) ) ;
    buf_clk new_AGEMA_reg_buffer_1432 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_1_), .Q (new_AGEMA_signal_4200) ) ;
    buf_clk new_AGEMA_reg_buffer_1436 ( .C (CLK), .D (new_AGEMA_signal_2004), .Q (new_AGEMA_signal_4204) ) ;
    buf_clk new_AGEMA_reg_buffer_1440 ( .C (CLK), .D (new_AGEMA_signal_2005), .Q (new_AGEMA_signal_4208) ) ;
    buf_clk new_AGEMA_reg_buffer_1444 ( .C (CLK), .D (LED_128_Instance_MUX_state0_n8), .Q (new_AGEMA_signal_4212) ) ;
    buf_clk new_AGEMA_reg_buffer_1448 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_2_), .Q (new_AGEMA_signal_4216) ) ;
    buf_clk new_AGEMA_reg_buffer_1452 ( .C (CLK), .D (new_AGEMA_signal_2006), .Q (new_AGEMA_signal_4220) ) ;
    buf_clk new_AGEMA_reg_buffer_1456 ( .C (CLK), .D (new_AGEMA_signal_2007), .Q (new_AGEMA_signal_4224) ) ;
    buf_clk new_AGEMA_reg_buffer_1460 ( .C (CLK), .D (LED_128_Instance_MUX_state0_n10), .Q (new_AGEMA_signal_4228) ) ;
    buf_clk new_AGEMA_reg_buffer_1464 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_3_), .Q (new_AGEMA_signal_4232) ) ;
    buf_clk new_AGEMA_reg_buffer_1468 ( .C (CLK), .D (new_AGEMA_signal_1766), .Q (new_AGEMA_signal_4236) ) ;
    buf_clk new_AGEMA_reg_buffer_1472 ( .C (CLK), .D (new_AGEMA_signal_1767), .Q (new_AGEMA_signal_4240) ) ;
    buf_clk new_AGEMA_reg_buffer_1476 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_4_), .Q (new_AGEMA_signal_4244) ) ;
    buf_clk new_AGEMA_reg_buffer_1480 ( .C (CLK), .D (new_AGEMA_signal_2008), .Q (new_AGEMA_signal_4248) ) ;
    buf_clk new_AGEMA_reg_buffer_1484 ( .C (CLK), .D (new_AGEMA_signal_2009), .Q (new_AGEMA_signal_4252) ) ;
    buf_clk new_AGEMA_reg_buffer_1488 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_5_), .Q (new_AGEMA_signal_4256) ) ;
    buf_clk new_AGEMA_reg_buffer_1492 ( .C (CLK), .D (new_AGEMA_signal_2010), .Q (new_AGEMA_signal_4260) ) ;
    buf_clk new_AGEMA_reg_buffer_1496 ( .C (CLK), .D (new_AGEMA_signal_2011), .Q (new_AGEMA_signal_4264) ) ;
    buf_clk new_AGEMA_reg_buffer_1500 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_6_), .Q (new_AGEMA_signal_4268) ) ;
    buf_clk new_AGEMA_reg_buffer_1504 ( .C (CLK), .D (new_AGEMA_signal_2012), .Q (new_AGEMA_signal_4272) ) ;
    buf_clk new_AGEMA_reg_buffer_1508 ( .C (CLK), .D (new_AGEMA_signal_2013), .Q (new_AGEMA_signal_4276) ) ;
    buf_clk new_AGEMA_reg_buffer_1512 ( .C (CLK), .D (LED_128_Instance_addconst_out[7]), .Q (new_AGEMA_signal_4280) ) ;
    buf_clk new_AGEMA_reg_buffer_1516 ( .C (CLK), .D (new_AGEMA_signal_2014), .Q (new_AGEMA_signal_4284) ) ;
    buf_clk new_AGEMA_reg_buffer_1520 ( .C (CLK), .D (new_AGEMA_signal_2015), .Q (new_AGEMA_signal_4288) ) ;
    buf_clk new_AGEMA_reg_buffer_1524 ( .C (CLK), .D (LED_128_Instance_addconst_out[8]), .Q (new_AGEMA_signal_4292) ) ;
    buf_clk new_AGEMA_reg_buffer_1528 ( .C (CLK), .D (new_AGEMA_signal_2016), .Q (new_AGEMA_signal_4296) ) ;
    buf_clk new_AGEMA_reg_buffer_1532 ( .C (CLK), .D (new_AGEMA_signal_2017), .Q (new_AGEMA_signal_4300) ) ;
    buf_clk new_AGEMA_reg_buffer_1536 ( .C (CLK), .D (LED_128_Instance_addconst_out[9]), .Q (new_AGEMA_signal_4304) ) ;
    buf_clk new_AGEMA_reg_buffer_1540 ( .C (CLK), .D (new_AGEMA_signal_2018), .Q (new_AGEMA_signal_4308) ) ;
    buf_clk new_AGEMA_reg_buffer_1544 ( .C (CLK), .D (new_AGEMA_signal_2019), .Q (new_AGEMA_signal_4312) ) ;
    buf_clk new_AGEMA_reg_buffer_1548 ( .C (CLK), .D (LED_128_Instance_addconst_out[10]), .Q (new_AGEMA_signal_4316) ) ;
    buf_clk new_AGEMA_reg_buffer_1552 ( .C (CLK), .D (new_AGEMA_signal_2020), .Q (new_AGEMA_signal_4320) ) ;
    buf_clk new_AGEMA_reg_buffer_1556 ( .C (CLK), .D (new_AGEMA_signal_2021), .Q (new_AGEMA_signal_4324) ) ;
    buf_clk new_AGEMA_reg_buffer_1560 ( .C (CLK), .D (LED_128_Instance_addconst_out[11]), .Q (new_AGEMA_signal_4328) ) ;
    buf_clk new_AGEMA_reg_buffer_1564 ( .C (CLK), .D (new_AGEMA_signal_2022), .Q (new_AGEMA_signal_4332) ) ;
    buf_clk new_AGEMA_reg_buffer_1568 ( .C (CLK), .D (new_AGEMA_signal_2023), .Q (new_AGEMA_signal_4336) ) ;
    buf_clk new_AGEMA_reg_buffer_1572 ( .C (CLK), .D (LED_128_Instance_addconst_out[12]), .Q (new_AGEMA_signal_4340) ) ;
    buf_clk new_AGEMA_reg_buffer_1576 ( .C (CLK), .D (new_AGEMA_signal_2024), .Q (new_AGEMA_signal_4344) ) ;
    buf_clk new_AGEMA_reg_buffer_1580 ( .C (CLK), .D (new_AGEMA_signal_2025), .Q (new_AGEMA_signal_4348) ) ;
    buf_clk new_AGEMA_reg_buffer_1584 ( .C (CLK), .D (LED_128_Instance_addconst_out[13]), .Q (new_AGEMA_signal_4352) ) ;
    buf_clk new_AGEMA_reg_buffer_1588 ( .C (CLK), .D (new_AGEMA_signal_2026), .Q (new_AGEMA_signal_4356) ) ;
    buf_clk new_AGEMA_reg_buffer_1592 ( .C (CLK), .D (new_AGEMA_signal_2027), .Q (new_AGEMA_signal_4360) ) ;
    buf_clk new_AGEMA_reg_buffer_1596 ( .C (CLK), .D (LED_128_Instance_addconst_out[14]), .Q (new_AGEMA_signal_4364) ) ;
    buf_clk new_AGEMA_reg_buffer_1600 ( .C (CLK), .D (new_AGEMA_signal_2028), .Q (new_AGEMA_signal_4368) ) ;
    buf_clk new_AGEMA_reg_buffer_1604 ( .C (CLK), .D (new_AGEMA_signal_2029), .Q (new_AGEMA_signal_4372) ) ;
    buf_clk new_AGEMA_reg_buffer_1608 ( .C (CLK), .D (LED_128_Instance_addconst_out[15]), .Q (new_AGEMA_signal_4376) ) ;
    buf_clk new_AGEMA_reg_buffer_1612 ( .C (CLK), .D (new_AGEMA_signal_2030), .Q (new_AGEMA_signal_4380) ) ;
    buf_clk new_AGEMA_reg_buffer_1616 ( .C (CLK), .D (new_AGEMA_signal_2031), .Q (new_AGEMA_signal_4384) ) ;
    buf_clk new_AGEMA_reg_buffer_1620 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_16_), .Q (new_AGEMA_signal_4388) ) ;
    buf_clk new_AGEMA_reg_buffer_1624 ( .C (CLK), .D (new_AGEMA_signal_1768), .Q (new_AGEMA_signal_4392) ) ;
    buf_clk new_AGEMA_reg_buffer_1628 ( .C (CLK), .D (new_AGEMA_signal_1769), .Q (new_AGEMA_signal_4396) ) ;
    buf_clk new_AGEMA_reg_buffer_1632 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_17_), .Q (new_AGEMA_signal_4400) ) ;
    buf_clk new_AGEMA_reg_buffer_1636 ( .C (CLK), .D (new_AGEMA_signal_2032), .Q (new_AGEMA_signal_4404) ) ;
    buf_clk new_AGEMA_reg_buffer_1640 ( .C (CLK), .D (new_AGEMA_signal_2033), .Q (new_AGEMA_signal_4408) ) ;
    buf_clk new_AGEMA_reg_buffer_1644 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_18_), .Q (new_AGEMA_signal_4412) ) ;
    buf_clk new_AGEMA_reg_buffer_1648 ( .C (CLK), .D (new_AGEMA_signal_2034), .Q (new_AGEMA_signal_4416) ) ;
    buf_clk new_AGEMA_reg_buffer_1652 ( .C (CLK), .D (new_AGEMA_signal_2035), .Q (new_AGEMA_signal_4420) ) ;
    buf_clk new_AGEMA_reg_buffer_1656 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_19_), .Q (new_AGEMA_signal_4424) ) ;
    buf_clk new_AGEMA_reg_buffer_1660 ( .C (CLK), .D (new_AGEMA_signal_1770), .Q (new_AGEMA_signal_4428) ) ;
    buf_clk new_AGEMA_reg_buffer_1664 ( .C (CLK), .D (new_AGEMA_signal_1771), .Q (new_AGEMA_signal_4432) ) ;
    buf_clk new_AGEMA_reg_buffer_1668 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_20_), .Q (new_AGEMA_signal_4436) ) ;
    buf_clk new_AGEMA_reg_buffer_1672 ( .C (CLK), .D (new_AGEMA_signal_2036), .Q (new_AGEMA_signal_4440) ) ;
    buf_clk new_AGEMA_reg_buffer_1676 ( .C (CLK), .D (new_AGEMA_signal_2037), .Q (new_AGEMA_signal_4444) ) ;
    buf_clk new_AGEMA_reg_buffer_1680 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_21_), .Q (new_AGEMA_signal_4448) ) ;
    buf_clk new_AGEMA_reg_buffer_1684 ( .C (CLK), .D (new_AGEMA_signal_2038), .Q (new_AGEMA_signal_4452) ) ;
    buf_clk new_AGEMA_reg_buffer_1688 ( .C (CLK), .D (new_AGEMA_signal_2039), .Q (new_AGEMA_signal_4456) ) ;
    buf_clk new_AGEMA_reg_buffer_1692 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_22_), .Q (new_AGEMA_signal_4460) ) ;
    buf_clk new_AGEMA_reg_buffer_1696 ( .C (CLK), .D (new_AGEMA_signal_1772), .Q (new_AGEMA_signal_4464) ) ;
    buf_clk new_AGEMA_reg_buffer_1700 ( .C (CLK), .D (new_AGEMA_signal_1773), .Q (new_AGEMA_signal_4468) ) ;
    buf_clk new_AGEMA_reg_buffer_1704 ( .C (CLK), .D (LED_128_Instance_addconst_out[23]), .Q (new_AGEMA_signal_4472) ) ;
    buf_clk new_AGEMA_reg_buffer_1708 ( .C (CLK), .D (new_AGEMA_signal_2040), .Q (new_AGEMA_signal_4476) ) ;
    buf_clk new_AGEMA_reg_buffer_1712 ( .C (CLK), .D (new_AGEMA_signal_2041), .Q (new_AGEMA_signal_4480) ) ;
    buf_clk new_AGEMA_reg_buffer_1716 ( .C (CLK), .D (LED_128_Instance_addconst_out[24]), .Q (new_AGEMA_signal_4484) ) ;
    buf_clk new_AGEMA_reg_buffer_1720 ( .C (CLK), .D (new_AGEMA_signal_1774), .Q (new_AGEMA_signal_4488) ) ;
    buf_clk new_AGEMA_reg_buffer_1724 ( .C (CLK), .D (new_AGEMA_signal_1775), .Q (new_AGEMA_signal_4492) ) ;
    buf_clk new_AGEMA_reg_buffer_1728 ( .C (CLK), .D (LED_128_Instance_addconst_out[25]), .Q (new_AGEMA_signal_4496) ) ;
    buf_clk new_AGEMA_reg_buffer_1732 ( .C (CLK), .D (new_AGEMA_signal_2042), .Q (new_AGEMA_signal_4500) ) ;
    buf_clk new_AGEMA_reg_buffer_1736 ( .C (CLK), .D (new_AGEMA_signal_2043), .Q (new_AGEMA_signal_4504) ) ;
    buf_clk new_AGEMA_reg_buffer_1740 ( .C (CLK), .D (LED_128_Instance_addconst_out[26]), .Q (new_AGEMA_signal_4508) ) ;
    buf_clk new_AGEMA_reg_buffer_1744 ( .C (CLK), .D (new_AGEMA_signal_1776), .Q (new_AGEMA_signal_4512) ) ;
    buf_clk new_AGEMA_reg_buffer_1748 ( .C (CLK), .D (new_AGEMA_signal_1777), .Q (new_AGEMA_signal_4516) ) ;
    buf_clk new_AGEMA_reg_buffer_1752 ( .C (CLK), .D (LED_128_Instance_addconst_out[27]), .Q (new_AGEMA_signal_4520) ) ;
    buf_clk new_AGEMA_reg_buffer_1756 ( .C (CLK), .D (new_AGEMA_signal_2044), .Q (new_AGEMA_signal_4524) ) ;
    buf_clk new_AGEMA_reg_buffer_1760 ( .C (CLK), .D (new_AGEMA_signal_2045), .Q (new_AGEMA_signal_4528) ) ;
    buf_clk new_AGEMA_reg_buffer_1764 ( .C (CLK), .D (LED_128_Instance_addconst_out[28]), .Q (new_AGEMA_signal_4532) ) ;
    buf_clk new_AGEMA_reg_buffer_1768 ( .C (CLK), .D (new_AGEMA_signal_1982), .Q (new_AGEMA_signal_4536) ) ;
    buf_clk new_AGEMA_reg_buffer_1772 ( .C (CLK), .D (new_AGEMA_signal_1983), .Q (new_AGEMA_signal_4540) ) ;
    buf_clk new_AGEMA_reg_buffer_1776 ( .C (CLK), .D (LED_128_Instance_addconst_out[29]), .Q (new_AGEMA_signal_4544) ) ;
    buf_clk new_AGEMA_reg_buffer_1780 ( .C (CLK), .D (new_AGEMA_signal_2046), .Q (new_AGEMA_signal_4548) ) ;
    buf_clk new_AGEMA_reg_buffer_1784 ( .C (CLK), .D (new_AGEMA_signal_2047), .Q (new_AGEMA_signal_4552) ) ;
    buf_clk new_AGEMA_reg_buffer_1788 ( .C (CLK), .D (LED_128_Instance_addconst_out[30]), .Q (new_AGEMA_signal_4556) ) ;
    buf_clk new_AGEMA_reg_buffer_1792 ( .C (CLK), .D (new_AGEMA_signal_2048), .Q (new_AGEMA_signal_4560) ) ;
    buf_clk new_AGEMA_reg_buffer_1796 ( .C (CLK), .D (new_AGEMA_signal_2049), .Q (new_AGEMA_signal_4564) ) ;
    buf_clk new_AGEMA_reg_buffer_1800 ( .C (CLK), .D (LED_128_Instance_addconst_out[31]), .Q (new_AGEMA_signal_4568) ) ;
    buf_clk new_AGEMA_reg_buffer_1804 ( .C (CLK), .D (new_AGEMA_signal_2050), .Q (new_AGEMA_signal_4572) ) ;
    buf_clk new_AGEMA_reg_buffer_1808 ( .C (CLK), .D (new_AGEMA_signal_2051), .Q (new_AGEMA_signal_4576) ) ;
    buf_clk new_AGEMA_reg_buffer_1812 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_32_), .Q (new_AGEMA_signal_4580) ) ;
    buf_clk new_AGEMA_reg_buffer_1816 ( .C (CLK), .D (new_AGEMA_signal_1984), .Q (new_AGEMA_signal_4584) ) ;
    buf_clk new_AGEMA_reg_buffer_1820 ( .C (CLK), .D (new_AGEMA_signal_1985), .Q (new_AGEMA_signal_4588) ) ;
    buf_clk new_AGEMA_reg_buffer_1824 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_33_), .Q (new_AGEMA_signal_4592) ) ;
    buf_clk new_AGEMA_reg_buffer_1828 ( .C (CLK), .D (new_AGEMA_signal_2052), .Q (new_AGEMA_signal_4596) ) ;
    buf_clk new_AGEMA_reg_buffer_1832 ( .C (CLK), .D (new_AGEMA_signal_2053), .Q (new_AGEMA_signal_4600) ) ;
    buf_clk new_AGEMA_reg_buffer_1836 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_34_), .Q (new_AGEMA_signal_4604) ) ;
    buf_clk new_AGEMA_reg_buffer_1840 ( .C (CLK), .D (new_AGEMA_signal_1986), .Q (new_AGEMA_signal_4608) ) ;
    buf_clk new_AGEMA_reg_buffer_1844 ( .C (CLK), .D (new_AGEMA_signal_1987), .Q (new_AGEMA_signal_4612) ) ;
    buf_clk new_AGEMA_reg_buffer_1848 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_35_), .Q (new_AGEMA_signal_4616) ) ;
    buf_clk new_AGEMA_reg_buffer_1852 ( .C (CLK), .D (new_AGEMA_signal_1988), .Q (new_AGEMA_signal_4620) ) ;
    buf_clk new_AGEMA_reg_buffer_1856 ( .C (CLK), .D (new_AGEMA_signal_1989), .Q (new_AGEMA_signal_4624) ) ;
    buf_clk new_AGEMA_reg_buffer_1860 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_36_), .Q (new_AGEMA_signal_4628) ) ;
    buf_clk new_AGEMA_reg_buffer_1864 ( .C (CLK), .D (new_AGEMA_signal_1990), .Q (new_AGEMA_signal_4632) ) ;
    buf_clk new_AGEMA_reg_buffer_1868 ( .C (CLK), .D (new_AGEMA_signal_1991), .Q (new_AGEMA_signal_4636) ) ;
    buf_clk new_AGEMA_reg_buffer_1872 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_37_), .Q (new_AGEMA_signal_4640) ) ;
    buf_clk new_AGEMA_reg_buffer_1876 ( .C (CLK), .D (new_AGEMA_signal_2054), .Q (new_AGEMA_signal_4644) ) ;
    buf_clk new_AGEMA_reg_buffer_1880 ( .C (CLK), .D (new_AGEMA_signal_2055), .Q (new_AGEMA_signal_4648) ) ;
    buf_clk new_AGEMA_reg_buffer_1884 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_38_), .Q (new_AGEMA_signal_4652) ) ;
    buf_clk new_AGEMA_reg_buffer_1888 ( .C (CLK), .D (new_AGEMA_signal_2056), .Q (new_AGEMA_signal_4656) ) ;
    buf_clk new_AGEMA_reg_buffer_1892 ( .C (CLK), .D (new_AGEMA_signal_2057), .Q (new_AGEMA_signal_4660) ) ;
    buf_clk new_AGEMA_reg_buffer_1896 ( .C (CLK), .D (LED_128_Instance_addconst_out[39]), .Q (new_AGEMA_signal_4664) ) ;
    buf_clk new_AGEMA_reg_buffer_1900 ( .C (CLK), .D (new_AGEMA_signal_1992), .Q (new_AGEMA_signal_4668) ) ;
    buf_clk new_AGEMA_reg_buffer_1904 ( .C (CLK), .D (new_AGEMA_signal_1993), .Q (new_AGEMA_signal_4672) ) ;
    buf_clk new_AGEMA_reg_buffer_1908 ( .C (CLK), .D (LED_128_Instance_addconst_out[40]), .Q (new_AGEMA_signal_4676) ) ;
    buf_clk new_AGEMA_reg_buffer_1912 ( .C (CLK), .D (new_AGEMA_signal_2058), .Q (new_AGEMA_signal_4680) ) ;
    buf_clk new_AGEMA_reg_buffer_1916 ( .C (CLK), .D (new_AGEMA_signal_2059), .Q (new_AGEMA_signal_4684) ) ;
    buf_clk new_AGEMA_reg_buffer_1920 ( .C (CLK), .D (LED_128_Instance_addconst_out[41]), .Q (new_AGEMA_signal_4688) ) ;
    buf_clk new_AGEMA_reg_buffer_1924 ( .C (CLK), .D (new_AGEMA_signal_2060), .Q (new_AGEMA_signal_4692) ) ;
    buf_clk new_AGEMA_reg_buffer_1928 ( .C (CLK), .D (new_AGEMA_signal_2061), .Q (new_AGEMA_signal_4696) ) ;
    buf_clk new_AGEMA_reg_buffer_1932 ( .C (CLK), .D (LED_128_Instance_addconst_out[42]), .Q (new_AGEMA_signal_4700) ) ;
    buf_clk new_AGEMA_reg_buffer_1936 ( .C (CLK), .D (new_AGEMA_signal_2062), .Q (new_AGEMA_signal_4704) ) ;
    buf_clk new_AGEMA_reg_buffer_1940 ( .C (CLK), .D (new_AGEMA_signal_2063), .Q (new_AGEMA_signal_4708) ) ;
    buf_clk new_AGEMA_reg_buffer_1944 ( .C (CLK), .D (LED_128_Instance_n22), .Q (new_AGEMA_signal_4712) ) ;
    buf_clk new_AGEMA_reg_buffer_1948 ( .C (CLK), .D (LED_128_Instance_addconst_out[43]), .Q (new_AGEMA_signal_4716) ) ;
    buf_clk new_AGEMA_reg_buffer_1952 ( .C (CLK), .D (new_AGEMA_signal_2064), .Q (new_AGEMA_signal_4720) ) ;
    buf_clk new_AGEMA_reg_buffer_1956 ( .C (CLK), .D (new_AGEMA_signal_2065), .Q (new_AGEMA_signal_4724) ) ;
    buf_clk new_AGEMA_reg_buffer_1960 ( .C (CLK), .D (LED_128_Instance_addconst_out[44]), .Q (new_AGEMA_signal_4728) ) ;
    buf_clk new_AGEMA_reg_buffer_1964 ( .C (CLK), .D (new_AGEMA_signal_2066), .Q (new_AGEMA_signal_4732) ) ;
    buf_clk new_AGEMA_reg_buffer_1968 ( .C (CLK), .D (new_AGEMA_signal_2067), .Q (new_AGEMA_signal_4736) ) ;
    buf_clk new_AGEMA_reg_buffer_1972 ( .C (CLK), .D (LED_128_Instance_addconst_out[45]), .Q (new_AGEMA_signal_4740) ) ;
    buf_clk new_AGEMA_reg_buffer_1976 ( .C (CLK), .D (new_AGEMA_signal_2068), .Q (new_AGEMA_signal_4744) ) ;
    buf_clk new_AGEMA_reg_buffer_1980 ( .C (CLK), .D (new_AGEMA_signal_2069), .Q (new_AGEMA_signal_4748) ) ;
    buf_clk new_AGEMA_reg_buffer_1984 ( .C (CLK), .D (LED_128_Instance_addconst_out[46]), .Q (new_AGEMA_signal_4752) ) ;
    buf_clk new_AGEMA_reg_buffer_1988 ( .C (CLK), .D (new_AGEMA_signal_2070), .Q (new_AGEMA_signal_4756) ) ;
    buf_clk new_AGEMA_reg_buffer_1992 ( .C (CLK), .D (new_AGEMA_signal_2071), .Q (new_AGEMA_signal_4760) ) ;
    buf_clk new_AGEMA_reg_buffer_1996 ( .C (CLK), .D (LED_128_Instance_addconst_out[47]), .Q (new_AGEMA_signal_4764) ) ;
    buf_clk new_AGEMA_reg_buffer_2000 ( .C (CLK), .D (new_AGEMA_signal_2072), .Q (new_AGEMA_signal_4768) ) ;
    buf_clk new_AGEMA_reg_buffer_2004 ( .C (CLK), .D (new_AGEMA_signal_2073), .Q (new_AGEMA_signal_4772) ) ;
    buf_clk new_AGEMA_reg_buffer_2008 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_48_), .Q (new_AGEMA_signal_4776) ) ;
    buf_clk new_AGEMA_reg_buffer_2012 ( .C (CLK), .D (new_AGEMA_signal_2074), .Q (new_AGEMA_signal_4780) ) ;
    buf_clk new_AGEMA_reg_buffer_2016 ( .C (CLK), .D (new_AGEMA_signal_2075), .Q (new_AGEMA_signal_4784) ) ;
    buf_clk new_AGEMA_reg_buffer_2020 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_49_), .Q (new_AGEMA_signal_4788) ) ;
    buf_clk new_AGEMA_reg_buffer_2024 ( .C (CLK), .D (new_AGEMA_signal_2076), .Q (new_AGEMA_signal_4792) ) ;
    buf_clk new_AGEMA_reg_buffer_2028 ( .C (CLK), .D (new_AGEMA_signal_2077), .Q (new_AGEMA_signal_4796) ) ;
    buf_clk new_AGEMA_reg_buffer_2032 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_50_), .Q (new_AGEMA_signal_4800) ) ;
    buf_clk new_AGEMA_reg_buffer_2036 ( .C (CLK), .D (new_AGEMA_signal_2078), .Q (new_AGEMA_signal_4804) ) ;
    buf_clk new_AGEMA_reg_buffer_2040 ( .C (CLK), .D (new_AGEMA_signal_2079), .Q (new_AGEMA_signal_4808) ) ;
    buf_clk new_AGEMA_reg_buffer_2044 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_51_), .Q (new_AGEMA_signal_4812) ) ;
    buf_clk new_AGEMA_reg_buffer_2048 ( .C (CLK), .D (new_AGEMA_signal_2080), .Q (new_AGEMA_signal_4816) ) ;
    buf_clk new_AGEMA_reg_buffer_2052 ( .C (CLK), .D (new_AGEMA_signal_2081), .Q (new_AGEMA_signal_4820) ) ;
    buf_clk new_AGEMA_reg_buffer_2056 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_52_), .Q (new_AGEMA_signal_4824) ) ;
    buf_clk new_AGEMA_reg_buffer_2060 ( .C (CLK), .D (new_AGEMA_signal_2082), .Q (new_AGEMA_signal_4828) ) ;
    buf_clk new_AGEMA_reg_buffer_2064 ( .C (CLK), .D (new_AGEMA_signal_2083), .Q (new_AGEMA_signal_4832) ) ;
    buf_clk new_AGEMA_reg_buffer_2068 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_53_), .Q (new_AGEMA_signal_4836) ) ;
    buf_clk new_AGEMA_reg_buffer_2072 ( .C (CLK), .D (new_AGEMA_signal_2084), .Q (new_AGEMA_signal_4840) ) ;
    buf_clk new_AGEMA_reg_buffer_2076 ( .C (CLK), .D (new_AGEMA_signal_2085), .Q (new_AGEMA_signal_4844) ) ;
    buf_clk new_AGEMA_reg_buffer_2080 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_54_), .Q (new_AGEMA_signal_4848) ) ;
    buf_clk new_AGEMA_reg_buffer_2084 ( .C (CLK), .D (new_AGEMA_signal_2086), .Q (new_AGEMA_signal_4852) ) ;
    buf_clk new_AGEMA_reg_buffer_2088 ( .C (CLK), .D (new_AGEMA_signal_2087), .Q (new_AGEMA_signal_4856) ) ;
    buf_clk new_AGEMA_reg_buffer_2092 ( .C (CLK), .D (LED_128_Instance_addconst_out[55]), .Q (new_AGEMA_signal_4860) ) ;
    buf_clk new_AGEMA_reg_buffer_2096 ( .C (CLK), .D (new_AGEMA_signal_2088), .Q (new_AGEMA_signal_4864) ) ;
    buf_clk new_AGEMA_reg_buffer_2100 ( .C (CLK), .D (new_AGEMA_signal_2089), .Q (new_AGEMA_signal_4868) ) ;
    buf_clk new_AGEMA_reg_buffer_2104 ( .C (CLK), .D (LED_128_Instance_addconst_out[56]), .Q (new_AGEMA_signal_4872) ) ;
    buf_clk new_AGEMA_reg_buffer_2108 ( .C (CLK), .D (new_AGEMA_signal_2090), .Q (new_AGEMA_signal_4876) ) ;
    buf_clk new_AGEMA_reg_buffer_2112 ( .C (CLK), .D (new_AGEMA_signal_2091), .Q (new_AGEMA_signal_4880) ) ;
    buf_clk new_AGEMA_reg_buffer_2116 ( .C (CLK), .D (LED_128_Instance_addconst_out[57]), .Q (new_AGEMA_signal_4884) ) ;
    buf_clk new_AGEMA_reg_buffer_2120 ( .C (CLK), .D (new_AGEMA_signal_2092), .Q (new_AGEMA_signal_4888) ) ;
    buf_clk new_AGEMA_reg_buffer_2124 ( .C (CLK), .D (new_AGEMA_signal_2093), .Q (new_AGEMA_signal_4892) ) ;
    buf_clk new_AGEMA_reg_buffer_2128 ( .C (CLK), .D (LED_128_Instance_addconst_out[58]), .Q (new_AGEMA_signal_4896) ) ;
    buf_clk new_AGEMA_reg_buffer_2132 ( .C (CLK), .D (new_AGEMA_signal_2094), .Q (new_AGEMA_signal_4900) ) ;
    buf_clk new_AGEMA_reg_buffer_2136 ( .C (CLK), .D (new_AGEMA_signal_2095), .Q (new_AGEMA_signal_4904) ) ;
    buf_clk new_AGEMA_reg_buffer_2140 ( .C (CLK), .D (LED_128_Instance_addconst_out[59]), .Q (new_AGEMA_signal_4908) ) ;
    buf_clk new_AGEMA_reg_buffer_2144 ( .C (CLK), .D (new_AGEMA_signal_2096), .Q (new_AGEMA_signal_4912) ) ;
    buf_clk new_AGEMA_reg_buffer_2148 ( .C (CLK), .D (new_AGEMA_signal_2097), .Q (new_AGEMA_signal_4916) ) ;
    buf_clk new_AGEMA_reg_buffer_2152 ( .C (CLK), .D (LED_128_Instance_addconst_out[60]), .Q (new_AGEMA_signal_4920) ) ;
    buf_clk new_AGEMA_reg_buffer_2156 ( .C (CLK), .D (new_AGEMA_signal_2098), .Q (new_AGEMA_signal_4924) ) ;
    buf_clk new_AGEMA_reg_buffer_2160 ( .C (CLK), .D (new_AGEMA_signal_2099), .Q (new_AGEMA_signal_4928) ) ;
    buf_clk new_AGEMA_reg_buffer_2164 ( .C (CLK), .D (LED_128_Instance_addconst_out[61]), .Q (new_AGEMA_signal_4932) ) ;
    buf_clk new_AGEMA_reg_buffer_2168 ( .C (CLK), .D (new_AGEMA_signal_2100), .Q (new_AGEMA_signal_4936) ) ;
    buf_clk new_AGEMA_reg_buffer_2172 ( .C (CLK), .D (new_AGEMA_signal_2101), .Q (new_AGEMA_signal_4940) ) ;
    buf_clk new_AGEMA_reg_buffer_2176 ( .C (CLK), .D (LED_128_Instance_addconst_out[62]), .Q (new_AGEMA_signal_4944) ) ;
    buf_clk new_AGEMA_reg_buffer_2180 ( .C (CLK), .D (new_AGEMA_signal_2102), .Q (new_AGEMA_signal_4948) ) ;
    buf_clk new_AGEMA_reg_buffer_2184 ( .C (CLK), .D (new_AGEMA_signal_2103), .Q (new_AGEMA_signal_4952) ) ;
    buf_clk new_AGEMA_reg_buffer_2188 ( .C (CLK), .D (LED_128_Instance_addconst_out[63]), .Q (new_AGEMA_signal_4956) ) ;
    buf_clk new_AGEMA_reg_buffer_2192 ( .C (CLK), .D (new_AGEMA_signal_2104), .Q (new_AGEMA_signal_4960) ) ;
    buf_clk new_AGEMA_reg_buffer_2196 ( .C (CLK), .D (new_AGEMA_signal_2105), .Q (new_AGEMA_signal_4964) ) ;
    buf_clk new_AGEMA_reg_buffer_2200 ( .C (CLK), .D (IN_reset), .Q (new_AGEMA_signal_4968) ) ;
    buf_clk new_AGEMA_reg_buffer_2204 ( .C (CLK), .D (IN_plaintext_s0[0]), .Q (new_AGEMA_signal_4972) ) ;
    buf_clk new_AGEMA_reg_buffer_2208 ( .C (CLK), .D (IN_plaintext_s1[0]), .Q (new_AGEMA_signal_4976) ) ;
    buf_clk new_AGEMA_reg_buffer_2212 ( .C (CLK), .D (IN_plaintext_s2[0]), .Q (new_AGEMA_signal_4980) ) ;
    buf_clk new_AGEMA_reg_buffer_2216 ( .C (CLK), .D (IN_plaintext_s0[1]), .Q (new_AGEMA_signal_4984) ) ;
    buf_clk new_AGEMA_reg_buffer_2220 ( .C (CLK), .D (IN_plaintext_s1[1]), .Q (new_AGEMA_signal_4988) ) ;
    buf_clk new_AGEMA_reg_buffer_2224 ( .C (CLK), .D (IN_plaintext_s2[1]), .Q (new_AGEMA_signal_4992) ) ;
    buf_clk new_AGEMA_reg_buffer_2228 ( .C (CLK), .D (IN_plaintext_s0[2]), .Q (new_AGEMA_signal_4996) ) ;
    buf_clk new_AGEMA_reg_buffer_2232 ( .C (CLK), .D (IN_plaintext_s1[2]), .Q (new_AGEMA_signal_5000) ) ;
    buf_clk new_AGEMA_reg_buffer_2236 ( .C (CLK), .D (IN_plaintext_s2[2]), .Q (new_AGEMA_signal_5004) ) ;
    buf_clk new_AGEMA_reg_buffer_2240 ( .C (CLK), .D (IN_plaintext_s0[3]), .Q (new_AGEMA_signal_5008) ) ;
    buf_clk new_AGEMA_reg_buffer_2244 ( .C (CLK), .D (IN_plaintext_s1[3]), .Q (new_AGEMA_signal_5012) ) ;
    buf_clk new_AGEMA_reg_buffer_2248 ( .C (CLK), .D (IN_plaintext_s2[3]), .Q (new_AGEMA_signal_5016) ) ;
    buf_clk new_AGEMA_reg_buffer_2252 ( .C (CLK), .D (IN_plaintext_s0[4]), .Q (new_AGEMA_signal_5020) ) ;
    buf_clk new_AGEMA_reg_buffer_2256 ( .C (CLK), .D (IN_plaintext_s1[4]), .Q (new_AGEMA_signal_5024) ) ;
    buf_clk new_AGEMA_reg_buffer_2260 ( .C (CLK), .D (IN_plaintext_s2[4]), .Q (new_AGEMA_signal_5028) ) ;
    buf_clk new_AGEMA_reg_buffer_2264 ( .C (CLK), .D (IN_plaintext_s0[5]), .Q (new_AGEMA_signal_5032) ) ;
    buf_clk new_AGEMA_reg_buffer_2268 ( .C (CLK), .D (IN_plaintext_s1[5]), .Q (new_AGEMA_signal_5036) ) ;
    buf_clk new_AGEMA_reg_buffer_2272 ( .C (CLK), .D (IN_plaintext_s2[5]), .Q (new_AGEMA_signal_5040) ) ;
    buf_clk new_AGEMA_reg_buffer_2276 ( .C (CLK), .D (IN_plaintext_s0[6]), .Q (new_AGEMA_signal_5044) ) ;
    buf_clk new_AGEMA_reg_buffer_2280 ( .C (CLK), .D (IN_plaintext_s1[6]), .Q (new_AGEMA_signal_5048) ) ;
    buf_clk new_AGEMA_reg_buffer_2284 ( .C (CLK), .D (IN_plaintext_s2[6]), .Q (new_AGEMA_signal_5052) ) ;
    buf_clk new_AGEMA_reg_buffer_2288 ( .C (CLK), .D (IN_plaintext_s0[7]), .Q (new_AGEMA_signal_5056) ) ;
    buf_clk new_AGEMA_reg_buffer_2292 ( .C (CLK), .D (IN_plaintext_s1[7]), .Q (new_AGEMA_signal_5060) ) ;
    buf_clk new_AGEMA_reg_buffer_2296 ( .C (CLK), .D (IN_plaintext_s2[7]), .Q (new_AGEMA_signal_5064) ) ;
    buf_clk new_AGEMA_reg_buffer_2300 ( .C (CLK), .D (IN_plaintext_s0[8]), .Q (new_AGEMA_signal_5068) ) ;
    buf_clk new_AGEMA_reg_buffer_2304 ( .C (CLK), .D (IN_plaintext_s1[8]), .Q (new_AGEMA_signal_5072) ) ;
    buf_clk new_AGEMA_reg_buffer_2308 ( .C (CLK), .D (IN_plaintext_s2[8]), .Q (new_AGEMA_signal_5076) ) ;
    buf_clk new_AGEMA_reg_buffer_2312 ( .C (CLK), .D (IN_plaintext_s0[9]), .Q (new_AGEMA_signal_5080) ) ;
    buf_clk new_AGEMA_reg_buffer_2316 ( .C (CLK), .D (IN_plaintext_s1[9]), .Q (new_AGEMA_signal_5084) ) ;
    buf_clk new_AGEMA_reg_buffer_2320 ( .C (CLK), .D (IN_plaintext_s2[9]), .Q (new_AGEMA_signal_5088) ) ;
    buf_clk new_AGEMA_reg_buffer_2324 ( .C (CLK), .D (IN_plaintext_s0[10]), .Q (new_AGEMA_signal_5092) ) ;
    buf_clk new_AGEMA_reg_buffer_2328 ( .C (CLK), .D (IN_plaintext_s1[10]), .Q (new_AGEMA_signal_5096) ) ;
    buf_clk new_AGEMA_reg_buffer_2332 ( .C (CLK), .D (IN_plaintext_s2[10]), .Q (new_AGEMA_signal_5100) ) ;
    buf_clk new_AGEMA_reg_buffer_2336 ( .C (CLK), .D (IN_plaintext_s0[11]), .Q (new_AGEMA_signal_5104) ) ;
    buf_clk new_AGEMA_reg_buffer_2340 ( .C (CLK), .D (IN_plaintext_s1[11]), .Q (new_AGEMA_signal_5108) ) ;
    buf_clk new_AGEMA_reg_buffer_2344 ( .C (CLK), .D (IN_plaintext_s2[11]), .Q (new_AGEMA_signal_5112) ) ;
    buf_clk new_AGEMA_reg_buffer_2348 ( .C (CLK), .D (IN_plaintext_s0[12]), .Q (new_AGEMA_signal_5116) ) ;
    buf_clk new_AGEMA_reg_buffer_2352 ( .C (CLK), .D (IN_plaintext_s1[12]), .Q (new_AGEMA_signal_5120) ) ;
    buf_clk new_AGEMA_reg_buffer_2356 ( .C (CLK), .D (IN_plaintext_s2[12]), .Q (new_AGEMA_signal_5124) ) ;
    buf_clk new_AGEMA_reg_buffer_2360 ( .C (CLK), .D (IN_plaintext_s0[13]), .Q (new_AGEMA_signal_5128) ) ;
    buf_clk new_AGEMA_reg_buffer_2364 ( .C (CLK), .D (IN_plaintext_s1[13]), .Q (new_AGEMA_signal_5132) ) ;
    buf_clk new_AGEMA_reg_buffer_2368 ( .C (CLK), .D (IN_plaintext_s2[13]), .Q (new_AGEMA_signal_5136) ) ;
    buf_clk new_AGEMA_reg_buffer_2372 ( .C (CLK), .D (IN_plaintext_s0[14]), .Q (new_AGEMA_signal_5140) ) ;
    buf_clk new_AGEMA_reg_buffer_2376 ( .C (CLK), .D (IN_plaintext_s1[14]), .Q (new_AGEMA_signal_5144) ) ;
    buf_clk new_AGEMA_reg_buffer_2380 ( .C (CLK), .D (IN_plaintext_s2[14]), .Q (new_AGEMA_signal_5148) ) ;
    buf_clk new_AGEMA_reg_buffer_2384 ( .C (CLK), .D (IN_plaintext_s0[15]), .Q (new_AGEMA_signal_5152) ) ;
    buf_clk new_AGEMA_reg_buffer_2388 ( .C (CLK), .D (IN_plaintext_s1[15]), .Q (new_AGEMA_signal_5156) ) ;
    buf_clk new_AGEMA_reg_buffer_2392 ( .C (CLK), .D (IN_plaintext_s2[15]), .Q (new_AGEMA_signal_5160) ) ;
    buf_clk new_AGEMA_reg_buffer_2396 ( .C (CLK), .D (IN_plaintext_s0[16]), .Q (new_AGEMA_signal_5164) ) ;
    buf_clk new_AGEMA_reg_buffer_2400 ( .C (CLK), .D (IN_plaintext_s1[16]), .Q (new_AGEMA_signal_5168) ) ;
    buf_clk new_AGEMA_reg_buffer_2404 ( .C (CLK), .D (IN_plaintext_s2[16]), .Q (new_AGEMA_signal_5172) ) ;
    buf_clk new_AGEMA_reg_buffer_2408 ( .C (CLK), .D (IN_plaintext_s0[17]), .Q (new_AGEMA_signal_5176) ) ;
    buf_clk new_AGEMA_reg_buffer_2412 ( .C (CLK), .D (IN_plaintext_s1[17]), .Q (new_AGEMA_signal_5180) ) ;
    buf_clk new_AGEMA_reg_buffer_2416 ( .C (CLK), .D (IN_plaintext_s2[17]), .Q (new_AGEMA_signal_5184) ) ;
    buf_clk new_AGEMA_reg_buffer_2420 ( .C (CLK), .D (IN_plaintext_s0[18]), .Q (new_AGEMA_signal_5188) ) ;
    buf_clk new_AGEMA_reg_buffer_2424 ( .C (CLK), .D (IN_plaintext_s1[18]), .Q (new_AGEMA_signal_5192) ) ;
    buf_clk new_AGEMA_reg_buffer_2428 ( .C (CLK), .D (IN_plaintext_s2[18]), .Q (new_AGEMA_signal_5196) ) ;
    buf_clk new_AGEMA_reg_buffer_2432 ( .C (CLK), .D (IN_plaintext_s0[19]), .Q (new_AGEMA_signal_5200) ) ;
    buf_clk new_AGEMA_reg_buffer_2436 ( .C (CLK), .D (IN_plaintext_s1[19]), .Q (new_AGEMA_signal_5204) ) ;
    buf_clk new_AGEMA_reg_buffer_2440 ( .C (CLK), .D (IN_plaintext_s2[19]), .Q (new_AGEMA_signal_5208) ) ;
    buf_clk new_AGEMA_reg_buffer_2444 ( .C (CLK), .D (IN_plaintext_s0[20]), .Q (new_AGEMA_signal_5212) ) ;
    buf_clk new_AGEMA_reg_buffer_2448 ( .C (CLK), .D (IN_plaintext_s1[20]), .Q (new_AGEMA_signal_5216) ) ;
    buf_clk new_AGEMA_reg_buffer_2452 ( .C (CLK), .D (IN_plaintext_s2[20]), .Q (new_AGEMA_signal_5220) ) ;
    buf_clk new_AGEMA_reg_buffer_2456 ( .C (CLK), .D (IN_plaintext_s0[21]), .Q (new_AGEMA_signal_5224) ) ;
    buf_clk new_AGEMA_reg_buffer_2460 ( .C (CLK), .D (IN_plaintext_s1[21]), .Q (new_AGEMA_signal_5228) ) ;
    buf_clk new_AGEMA_reg_buffer_2464 ( .C (CLK), .D (IN_plaintext_s2[21]), .Q (new_AGEMA_signal_5232) ) ;
    buf_clk new_AGEMA_reg_buffer_2468 ( .C (CLK), .D (IN_plaintext_s0[22]), .Q (new_AGEMA_signal_5236) ) ;
    buf_clk new_AGEMA_reg_buffer_2472 ( .C (CLK), .D (IN_plaintext_s1[22]), .Q (new_AGEMA_signal_5240) ) ;
    buf_clk new_AGEMA_reg_buffer_2476 ( .C (CLK), .D (IN_plaintext_s2[22]), .Q (new_AGEMA_signal_5244) ) ;
    buf_clk new_AGEMA_reg_buffer_2480 ( .C (CLK), .D (IN_plaintext_s0[23]), .Q (new_AGEMA_signal_5248) ) ;
    buf_clk new_AGEMA_reg_buffer_2484 ( .C (CLK), .D (IN_plaintext_s1[23]), .Q (new_AGEMA_signal_5252) ) ;
    buf_clk new_AGEMA_reg_buffer_2488 ( .C (CLK), .D (IN_plaintext_s2[23]), .Q (new_AGEMA_signal_5256) ) ;
    buf_clk new_AGEMA_reg_buffer_2492 ( .C (CLK), .D (IN_plaintext_s0[24]), .Q (new_AGEMA_signal_5260) ) ;
    buf_clk new_AGEMA_reg_buffer_2496 ( .C (CLK), .D (IN_plaintext_s1[24]), .Q (new_AGEMA_signal_5264) ) ;
    buf_clk new_AGEMA_reg_buffer_2500 ( .C (CLK), .D (IN_plaintext_s2[24]), .Q (new_AGEMA_signal_5268) ) ;
    buf_clk new_AGEMA_reg_buffer_2504 ( .C (CLK), .D (IN_plaintext_s0[25]), .Q (new_AGEMA_signal_5272) ) ;
    buf_clk new_AGEMA_reg_buffer_2508 ( .C (CLK), .D (IN_plaintext_s1[25]), .Q (new_AGEMA_signal_5276) ) ;
    buf_clk new_AGEMA_reg_buffer_2512 ( .C (CLK), .D (IN_plaintext_s2[25]), .Q (new_AGEMA_signal_5280) ) ;
    buf_clk new_AGEMA_reg_buffer_2516 ( .C (CLK), .D (IN_plaintext_s0[26]), .Q (new_AGEMA_signal_5284) ) ;
    buf_clk new_AGEMA_reg_buffer_2520 ( .C (CLK), .D (IN_plaintext_s1[26]), .Q (new_AGEMA_signal_5288) ) ;
    buf_clk new_AGEMA_reg_buffer_2524 ( .C (CLK), .D (IN_plaintext_s2[26]), .Q (new_AGEMA_signal_5292) ) ;
    buf_clk new_AGEMA_reg_buffer_2528 ( .C (CLK), .D (IN_plaintext_s0[27]), .Q (new_AGEMA_signal_5296) ) ;
    buf_clk new_AGEMA_reg_buffer_2532 ( .C (CLK), .D (IN_plaintext_s1[27]), .Q (new_AGEMA_signal_5300) ) ;
    buf_clk new_AGEMA_reg_buffer_2536 ( .C (CLK), .D (IN_plaintext_s2[27]), .Q (new_AGEMA_signal_5304) ) ;
    buf_clk new_AGEMA_reg_buffer_2540 ( .C (CLK), .D (IN_plaintext_s0[28]), .Q (new_AGEMA_signal_5308) ) ;
    buf_clk new_AGEMA_reg_buffer_2544 ( .C (CLK), .D (IN_plaintext_s1[28]), .Q (new_AGEMA_signal_5312) ) ;
    buf_clk new_AGEMA_reg_buffer_2548 ( .C (CLK), .D (IN_plaintext_s2[28]), .Q (new_AGEMA_signal_5316) ) ;
    buf_clk new_AGEMA_reg_buffer_2552 ( .C (CLK), .D (IN_plaintext_s0[29]), .Q (new_AGEMA_signal_5320) ) ;
    buf_clk new_AGEMA_reg_buffer_2556 ( .C (CLK), .D (IN_plaintext_s1[29]), .Q (new_AGEMA_signal_5324) ) ;
    buf_clk new_AGEMA_reg_buffer_2560 ( .C (CLK), .D (IN_plaintext_s2[29]), .Q (new_AGEMA_signal_5328) ) ;
    buf_clk new_AGEMA_reg_buffer_2564 ( .C (CLK), .D (IN_plaintext_s0[30]), .Q (new_AGEMA_signal_5332) ) ;
    buf_clk new_AGEMA_reg_buffer_2568 ( .C (CLK), .D (IN_plaintext_s1[30]), .Q (new_AGEMA_signal_5336) ) ;
    buf_clk new_AGEMA_reg_buffer_2572 ( .C (CLK), .D (IN_plaintext_s2[30]), .Q (new_AGEMA_signal_5340) ) ;
    buf_clk new_AGEMA_reg_buffer_2576 ( .C (CLK), .D (IN_plaintext_s0[31]), .Q (new_AGEMA_signal_5344) ) ;
    buf_clk new_AGEMA_reg_buffer_2580 ( .C (CLK), .D (IN_plaintext_s1[31]), .Q (new_AGEMA_signal_5348) ) ;
    buf_clk new_AGEMA_reg_buffer_2584 ( .C (CLK), .D (IN_plaintext_s2[31]), .Q (new_AGEMA_signal_5352) ) ;
    buf_clk new_AGEMA_reg_buffer_2588 ( .C (CLK), .D (IN_plaintext_s0[32]), .Q (new_AGEMA_signal_5356) ) ;
    buf_clk new_AGEMA_reg_buffer_2592 ( .C (CLK), .D (IN_plaintext_s1[32]), .Q (new_AGEMA_signal_5360) ) ;
    buf_clk new_AGEMA_reg_buffer_2596 ( .C (CLK), .D (IN_plaintext_s2[32]), .Q (new_AGEMA_signal_5364) ) ;
    buf_clk new_AGEMA_reg_buffer_2600 ( .C (CLK), .D (IN_plaintext_s0[33]), .Q (new_AGEMA_signal_5368) ) ;
    buf_clk new_AGEMA_reg_buffer_2604 ( .C (CLK), .D (IN_plaintext_s1[33]), .Q (new_AGEMA_signal_5372) ) ;
    buf_clk new_AGEMA_reg_buffer_2608 ( .C (CLK), .D (IN_plaintext_s2[33]), .Q (new_AGEMA_signal_5376) ) ;
    buf_clk new_AGEMA_reg_buffer_2612 ( .C (CLK), .D (IN_plaintext_s0[34]), .Q (new_AGEMA_signal_5380) ) ;
    buf_clk new_AGEMA_reg_buffer_2616 ( .C (CLK), .D (IN_plaintext_s1[34]), .Q (new_AGEMA_signal_5384) ) ;
    buf_clk new_AGEMA_reg_buffer_2620 ( .C (CLK), .D (IN_plaintext_s2[34]), .Q (new_AGEMA_signal_5388) ) ;
    buf_clk new_AGEMA_reg_buffer_2624 ( .C (CLK), .D (IN_plaintext_s0[35]), .Q (new_AGEMA_signal_5392) ) ;
    buf_clk new_AGEMA_reg_buffer_2628 ( .C (CLK), .D (IN_plaintext_s1[35]), .Q (new_AGEMA_signal_5396) ) ;
    buf_clk new_AGEMA_reg_buffer_2632 ( .C (CLK), .D (IN_plaintext_s2[35]), .Q (new_AGEMA_signal_5400) ) ;
    buf_clk new_AGEMA_reg_buffer_2636 ( .C (CLK), .D (IN_plaintext_s0[36]), .Q (new_AGEMA_signal_5404) ) ;
    buf_clk new_AGEMA_reg_buffer_2640 ( .C (CLK), .D (IN_plaintext_s1[36]), .Q (new_AGEMA_signal_5408) ) ;
    buf_clk new_AGEMA_reg_buffer_2644 ( .C (CLK), .D (IN_plaintext_s2[36]), .Q (new_AGEMA_signal_5412) ) ;
    buf_clk new_AGEMA_reg_buffer_2648 ( .C (CLK), .D (IN_plaintext_s0[37]), .Q (new_AGEMA_signal_5416) ) ;
    buf_clk new_AGEMA_reg_buffer_2652 ( .C (CLK), .D (IN_plaintext_s1[37]), .Q (new_AGEMA_signal_5420) ) ;
    buf_clk new_AGEMA_reg_buffer_2656 ( .C (CLK), .D (IN_plaintext_s2[37]), .Q (new_AGEMA_signal_5424) ) ;
    buf_clk new_AGEMA_reg_buffer_2660 ( .C (CLK), .D (IN_plaintext_s0[38]), .Q (new_AGEMA_signal_5428) ) ;
    buf_clk new_AGEMA_reg_buffer_2664 ( .C (CLK), .D (IN_plaintext_s1[38]), .Q (new_AGEMA_signal_5432) ) ;
    buf_clk new_AGEMA_reg_buffer_2668 ( .C (CLK), .D (IN_plaintext_s2[38]), .Q (new_AGEMA_signal_5436) ) ;
    buf_clk new_AGEMA_reg_buffer_2672 ( .C (CLK), .D (IN_plaintext_s0[39]), .Q (new_AGEMA_signal_5440) ) ;
    buf_clk new_AGEMA_reg_buffer_2676 ( .C (CLK), .D (IN_plaintext_s1[39]), .Q (new_AGEMA_signal_5444) ) ;
    buf_clk new_AGEMA_reg_buffer_2680 ( .C (CLK), .D (IN_plaintext_s2[39]), .Q (new_AGEMA_signal_5448) ) ;
    buf_clk new_AGEMA_reg_buffer_2684 ( .C (CLK), .D (IN_plaintext_s0[40]), .Q (new_AGEMA_signal_5452) ) ;
    buf_clk new_AGEMA_reg_buffer_2688 ( .C (CLK), .D (IN_plaintext_s1[40]), .Q (new_AGEMA_signal_5456) ) ;
    buf_clk new_AGEMA_reg_buffer_2692 ( .C (CLK), .D (IN_plaintext_s2[40]), .Q (new_AGEMA_signal_5460) ) ;
    buf_clk new_AGEMA_reg_buffer_2696 ( .C (CLK), .D (IN_plaintext_s0[41]), .Q (new_AGEMA_signal_5464) ) ;
    buf_clk new_AGEMA_reg_buffer_2700 ( .C (CLK), .D (IN_plaintext_s1[41]), .Q (new_AGEMA_signal_5468) ) ;
    buf_clk new_AGEMA_reg_buffer_2704 ( .C (CLK), .D (IN_plaintext_s2[41]), .Q (new_AGEMA_signal_5472) ) ;
    buf_clk new_AGEMA_reg_buffer_2708 ( .C (CLK), .D (IN_plaintext_s0[42]), .Q (new_AGEMA_signal_5476) ) ;
    buf_clk new_AGEMA_reg_buffer_2712 ( .C (CLK), .D (IN_plaintext_s1[42]), .Q (new_AGEMA_signal_5480) ) ;
    buf_clk new_AGEMA_reg_buffer_2716 ( .C (CLK), .D (IN_plaintext_s2[42]), .Q (new_AGEMA_signal_5484) ) ;
    buf_clk new_AGEMA_reg_buffer_2720 ( .C (CLK), .D (IN_plaintext_s0[43]), .Q (new_AGEMA_signal_5488) ) ;
    buf_clk new_AGEMA_reg_buffer_2724 ( .C (CLK), .D (IN_plaintext_s1[43]), .Q (new_AGEMA_signal_5492) ) ;
    buf_clk new_AGEMA_reg_buffer_2728 ( .C (CLK), .D (IN_plaintext_s2[43]), .Q (new_AGEMA_signal_5496) ) ;
    buf_clk new_AGEMA_reg_buffer_2732 ( .C (CLK), .D (IN_plaintext_s0[44]), .Q (new_AGEMA_signal_5500) ) ;
    buf_clk new_AGEMA_reg_buffer_2736 ( .C (CLK), .D (IN_plaintext_s1[44]), .Q (new_AGEMA_signal_5504) ) ;
    buf_clk new_AGEMA_reg_buffer_2740 ( .C (CLK), .D (IN_plaintext_s2[44]), .Q (new_AGEMA_signal_5508) ) ;
    buf_clk new_AGEMA_reg_buffer_2744 ( .C (CLK), .D (IN_plaintext_s0[45]), .Q (new_AGEMA_signal_5512) ) ;
    buf_clk new_AGEMA_reg_buffer_2748 ( .C (CLK), .D (IN_plaintext_s1[45]), .Q (new_AGEMA_signal_5516) ) ;
    buf_clk new_AGEMA_reg_buffer_2752 ( .C (CLK), .D (IN_plaintext_s2[45]), .Q (new_AGEMA_signal_5520) ) ;
    buf_clk new_AGEMA_reg_buffer_2756 ( .C (CLK), .D (IN_plaintext_s0[46]), .Q (new_AGEMA_signal_5524) ) ;
    buf_clk new_AGEMA_reg_buffer_2760 ( .C (CLK), .D (IN_plaintext_s1[46]), .Q (new_AGEMA_signal_5528) ) ;
    buf_clk new_AGEMA_reg_buffer_2764 ( .C (CLK), .D (IN_plaintext_s2[46]), .Q (new_AGEMA_signal_5532) ) ;
    buf_clk new_AGEMA_reg_buffer_2768 ( .C (CLK), .D (IN_plaintext_s0[47]), .Q (new_AGEMA_signal_5536) ) ;
    buf_clk new_AGEMA_reg_buffer_2772 ( .C (CLK), .D (IN_plaintext_s1[47]), .Q (new_AGEMA_signal_5540) ) ;
    buf_clk new_AGEMA_reg_buffer_2776 ( .C (CLK), .D (IN_plaintext_s2[47]), .Q (new_AGEMA_signal_5544) ) ;
    buf_clk new_AGEMA_reg_buffer_2780 ( .C (CLK), .D (IN_plaintext_s0[48]), .Q (new_AGEMA_signal_5548) ) ;
    buf_clk new_AGEMA_reg_buffer_2784 ( .C (CLK), .D (IN_plaintext_s1[48]), .Q (new_AGEMA_signal_5552) ) ;
    buf_clk new_AGEMA_reg_buffer_2788 ( .C (CLK), .D (IN_plaintext_s2[48]), .Q (new_AGEMA_signal_5556) ) ;
    buf_clk new_AGEMA_reg_buffer_2792 ( .C (CLK), .D (IN_plaintext_s0[49]), .Q (new_AGEMA_signal_5560) ) ;
    buf_clk new_AGEMA_reg_buffer_2796 ( .C (CLK), .D (IN_plaintext_s1[49]), .Q (new_AGEMA_signal_5564) ) ;
    buf_clk new_AGEMA_reg_buffer_2800 ( .C (CLK), .D (IN_plaintext_s2[49]), .Q (new_AGEMA_signal_5568) ) ;
    buf_clk new_AGEMA_reg_buffer_2804 ( .C (CLK), .D (IN_plaintext_s0[50]), .Q (new_AGEMA_signal_5572) ) ;
    buf_clk new_AGEMA_reg_buffer_2808 ( .C (CLK), .D (IN_plaintext_s1[50]), .Q (new_AGEMA_signal_5576) ) ;
    buf_clk new_AGEMA_reg_buffer_2812 ( .C (CLK), .D (IN_plaintext_s2[50]), .Q (new_AGEMA_signal_5580) ) ;
    buf_clk new_AGEMA_reg_buffer_2816 ( .C (CLK), .D (IN_plaintext_s0[51]), .Q (new_AGEMA_signal_5584) ) ;
    buf_clk new_AGEMA_reg_buffer_2820 ( .C (CLK), .D (IN_plaintext_s1[51]), .Q (new_AGEMA_signal_5588) ) ;
    buf_clk new_AGEMA_reg_buffer_2824 ( .C (CLK), .D (IN_plaintext_s2[51]), .Q (new_AGEMA_signal_5592) ) ;
    buf_clk new_AGEMA_reg_buffer_2828 ( .C (CLK), .D (IN_plaintext_s0[52]), .Q (new_AGEMA_signal_5596) ) ;
    buf_clk new_AGEMA_reg_buffer_2832 ( .C (CLK), .D (IN_plaintext_s1[52]), .Q (new_AGEMA_signal_5600) ) ;
    buf_clk new_AGEMA_reg_buffer_2836 ( .C (CLK), .D (IN_plaintext_s2[52]), .Q (new_AGEMA_signal_5604) ) ;
    buf_clk new_AGEMA_reg_buffer_2840 ( .C (CLK), .D (IN_plaintext_s0[53]), .Q (new_AGEMA_signal_5608) ) ;
    buf_clk new_AGEMA_reg_buffer_2844 ( .C (CLK), .D (IN_plaintext_s1[53]), .Q (new_AGEMA_signal_5612) ) ;
    buf_clk new_AGEMA_reg_buffer_2848 ( .C (CLK), .D (IN_plaintext_s2[53]), .Q (new_AGEMA_signal_5616) ) ;
    buf_clk new_AGEMA_reg_buffer_2852 ( .C (CLK), .D (IN_plaintext_s0[54]), .Q (new_AGEMA_signal_5620) ) ;
    buf_clk new_AGEMA_reg_buffer_2856 ( .C (CLK), .D (IN_plaintext_s1[54]), .Q (new_AGEMA_signal_5624) ) ;
    buf_clk new_AGEMA_reg_buffer_2860 ( .C (CLK), .D (IN_plaintext_s2[54]), .Q (new_AGEMA_signal_5628) ) ;
    buf_clk new_AGEMA_reg_buffer_2864 ( .C (CLK), .D (IN_plaintext_s0[55]), .Q (new_AGEMA_signal_5632) ) ;
    buf_clk new_AGEMA_reg_buffer_2868 ( .C (CLK), .D (IN_plaintext_s1[55]), .Q (new_AGEMA_signal_5636) ) ;
    buf_clk new_AGEMA_reg_buffer_2872 ( .C (CLK), .D (IN_plaintext_s2[55]), .Q (new_AGEMA_signal_5640) ) ;
    buf_clk new_AGEMA_reg_buffer_2876 ( .C (CLK), .D (IN_plaintext_s0[56]), .Q (new_AGEMA_signal_5644) ) ;
    buf_clk new_AGEMA_reg_buffer_2880 ( .C (CLK), .D (IN_plaintext_s1[56]), .Q (new_AGEMA_signal_5648) ) ;
    buf_clk new_AGEMA_reg_buffer_2884 ( .C (CLK), .D (IN_plaintext_s2[56]), .Q (new_AGEMA_signal_5652) ) ;
    buf_clk new_AGEMA_reg_buffer_2888 ( .C (CLK), .D (IN_plaintext_s0[57]), .Q (new_AGEMA_signal_5656) ) ;
    buf_clk new_AGEMA_reg_buffer_2892 ( .C (CLK), .D (IN_plaintext_s1[57]), .Q (new_AGEMA_signal_5660) ) ;
    buf_clk new_AGEMA_reg_buffer_2896 ( .C (CLK), .D (IN_plaintext_s2[57]), .Q (new_AGEMA_signal_5664) ) ;
    buf_clk new_AGEMA_reg_buffer_2900 ( .C (CLK), .D (IN_plaintext_s0[58]), .Q (new_AGEMA_signal_5668) ) ;
    buf_clk new_AGEMA_reg_buffer_2904 ( .C (CLK), .D (IN_plaintext_s1[58]), .Q (new_AGEMA_signal_5672) ) ;
    buf_clk new_AGEMA_reg_buffer_2908 ( .C (CLK), .D (IN_plaintext_s2[58]), .Q (new_AGEMA_signal_5676) ) ;
    buf_clk new_AGEMA_reg_buffer_2912 ( .C (CLK), .D (IN_plaintext_s0[59]), .Q (new_AGEMA_signal_5680) ) ;
    buf_clk new_AGEMA_reg_buffer_2916 ( .C (CLK), .D (IN_plaintext_s1[59]), .Q (new_AGEMA_signal_5684) ) ;
    buf_clk new_AGEMA_reg_buffer_2920 ( .C (CLK), .D (IN_plaintext_s2[59]), .Q (new_AGEMA_signal_5688) ) ;
    buf_clk new_AGEMA_reg_buffer_2924 ( .C (CLK), .D (IN_plaintext_s0[60]), .Q (new_AGEMA_signal_5692) ) ;
    buf_clk new_AGEMA_reg_buffer_2928 ( .C (CLK), .D (IN_plaintext_s1[60]), .Q (new_AGEMA_signal_5696) ) ;
    buf_clk new_AGEMA_reg_buffer_2932 ( .C (CLK), .D (IN_plaintext_s2[60]), .Q (new_AGEMA_signal_5700) ) ;
    buf_clk new_AGEMA_reg_buffer_2936 ( .C (CLK), .D (IN_plaintext_s0[61]), .Q (new_AGEMA_signal_5704) ) ;
    buf_clk new_AGEMA_reg_buffer_2940 ( .C (CLK), .D (IN_plaintext_s1[61]), .Q (new_AGEMA_signal_5708) ) ;
    buf_clk new_AGEMA_reg_buffer_2944 ( .C (CLK), .D (IN_plaintext_s2[61]), .Q (new_AGEMA_signal_5712) ) ;
    buf_clk new_AGEMA_reg_buffer_2948 ( .C (CLK), .D (IN_plaintext_s0[62]), .Q (new_AGEMA_signal_5716) ) ;
    buf_clk new_AGEMA_reg_buffer_2952 ( .C (CLK), .D (IN_plaintext_s1[62]), .Q (new_AGEMA_signal_5720) ) ;
    buf_clk new_AGEMA_reg_buffer_2956 ( .C (CLK), .D (IN_plaintext_s2[62]), .Q (new_AGEMA_signal_5724) ) ;
    buf_clk new_AGEMA_reg_buffer_2960 ( .C (CLK), .D (IN_plaintext_s0[63]), .Q (new_AGEMA_signal_5728) ) ;
    buf_clk new_AGEMA_reg_buffer_2964 ( .C (CLK), .D (IN_plaintext_s1[63]), .Q (new_AGEMA_signal_5732) ) ;
    buf_clk new_AGEMA_reg_buffer_2968 ( .C (CLK), .D (IN_plaintext_s2[63]), .Q (new_AGEMA_signal_5736) ) ;
    buf_clk new_AGEMA_reg_buffer_2972 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_0_Q3), .Q (new_AGEMA_signal_5740) ) ;
    buf_clk new_AGEMA_reg_buffer_2974 ( .C (CLK), .D (new_AGEMA_signal_2428), .Q (new_AGEMA_signal_5742) ) ;
    buf_clk new_AGEMA_reg_buffer_2976 ( .C (CLK), .D (new_AGEMA_signal_2429), .Q (new_AGEMA_signal_5744) ) ;
    buf_clk new_AGEMA_reg_buffer_2978 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_0_Q7), .Q (new_AGEMA_signal_5746) ) ;
    buf_clk new_AGEMA_reg_buffer_2980 ( .C (CLK), .D (new_AGEMA_signal_2430), .Q (new_AGEMA_signal_5748) ) ;
    buf_clk new_AGEMA_reg_buffer_2982 ( .C (CLK), .D (new_AGEMA_signal_2431), .Q (new_AGEMA_signal_5750) ) ;
    buf_clk new_AGEMA_reg_buffer_2990 ( .C (CLK), .D (LED_128_Instance_addconst_out[0]), .Q (new_AGEMA_signal_5758) ) ;
    buf_clk new_AGEMA_reg_buffer_2994 ( .C (CLK), .D (new_AGEMA_signal_2002), .Q (new_AGEMA_signal_5762) ) ;
    buf_clk new_AGEMA_reg_buffer_2998 ( .C (CLK), .D (new_AGEMA_signal_2003), .Q (new_AGEMA_signal_5766) ) ;
    buf_clk new_AGEMA_reg_buffer_3002 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_0_L1), .Q (new_AGEMA_signal_5770) ) ;
    buf_clk new_AGEMA_reg_buffer_3006 ( .C (CLK), .D (new_AGEMA_signal_2274), .Q (new_AGEMA_signal_5774) ) ;
    buf_clk new_AGEMA_reg_buffer_3010 ( .C (CLK), .D (new_AGEMA_signal_2275), .Q (new_AGEMA_signal_5778) ) ;
    buf_clk new_AGEMA_reg_buffer_3020 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_1_Q3), .Q (new_AGEMA_signal_5788) ) ;
    buf_clk new_AGEMA_reg_buffer_3022 ( .C (CLK), .D (new_AGEMA_signal_2438), .Q (new_AGEMA_signal_5790) ) ;
    buf_clk new_AGEMA_reg_buffer_3024 ( .C (CLK), .D (new_AGEMA_signal_2439), .Q (new_AGEMA_signal_5792) ) ;
    buf_clk new_AGEMA_reg_buffer_3026 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_1_Q7), .Q (new_AGEMA_signal_5794) ) ;
    buf_clk new_AGEMA_reg_buffer_3028 ( .C (CLK), .D (new_AGEMA_signal_2440), .Q (new_AGEMA_signal_5796) ) ;
    buf_clk new_AGEMA_reg_buffer_3030 ( .C (CLK), .D (new_AGEMA_signal_2441), .Q (new_AGEMA_signal_5798) ) ;
    buf_clk new_AGEMA_reg_buffer_3038 ( .C (CLK), .D (LED_128_Instance_addconst_out[4]), .Q (new_AGEMA_signal_5806) ) ;
    buf_clk new_AGEMA_reg_buffer_3042 ( .C (CLK), .D (new_AGEMA_signal_2138), .Q (new_AGEMA_signal_5810) ) ;
    buf_clk new_AGEMA_reg_buffer_3046 ( .C (CLK), .D (new_AGEMA_signal_2139), .Q (new_AGEMA_signal_5814) ) ;
    buf_clk new_AGEMA_reg_buffer_3050 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_1_L1), .Q (new_AGEMA_signal_5818) ) ;
    buf_clk new_AGEMA_reg_buffer_3054 ( .C (CLK), .D (new_AGEMA_signal_2282), .Q (new_AGEMA_signal_5822) ) ;
    buf_clk new_AGEMA_reg_buffer_3058 ( .C (CLK), .D (new_AGEMA_signal_2283), .Q (new_AGEMA_signal_5826) ) ;
    buf_clk new_AGEMA_reg_buffer_3068 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_2_Q3), .Q (new_AGEMA_signal_5836) ) ;
    buf_clk new_AGEMA_reg_buffer_3070 ( .C (CLK), .D (new_AGEMA_signal_2292), .Q (new_AGEMA_signal_5838) ) ;
    buf_clk new_AGEMA_reg_buffer_3072 ( .C (CLK), .D (new_AGEMA_signal_2293), .Q (new_AGEMA_signal_5840) ) ;
    buf_clk new_AGEMA_reg_buffer_3074 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_2_Q7), .Q (new_AGEMA_signal_5842) ) ;
    buf_clk new_AGEMA_reg_buffer_3076 ( .C (CLK), .D (new_AGEMA_signal_2294), .Q (new_AGEMA_signal_5844) ) ;
    buf_clk new_AGEMA_reg_buffer_3078 ( .C (CLK), .D (new_AGEMA_signal_2295), .Q (new_AGEMA_signal_5846) ) ;
    buf_clk new_AGEMA_reg_buffer_3086 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_2_L1), .Q (new_AGEMA_signal_5854) ) ;
    buf_clk new_AGEMA_reg_buffer_3090 ( .C (CLK), .D (new_AGEMA_signal_2170), .Q (new_AGEMA_signal_5858) ) ;
    buf_clk new_AGEMA_reg_buffer_3094 ( .C (CLK), .D (new_AGEMA_signal_2171), .Q (new_AGEMA_signal_5862) ) ;
    buf_clk new_AGEMA_reg_buffer_3104 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_3_Q3), .Q (new_AGEMA_signal_5872) ) ;
    buf_clk new_AGEMA_reg_buffer_3106 ( .C (CLK), .D (new_AGEMA_signal_2302), .Q (new_AGEMA_signal_5874) ) ;
    buf_clk new_AGEMA_reg_buffer_3108 ( .C (CLK), .D (new_AGEMA_signal_2303), .Q (new_AGEMA_signal_5876) ) ;
    buf_clk new_AGEMA_reg_buffer_3110 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_3_Q7), .Q (new_AGEMA_signal_5878) ) ;
    buf_clk new_AGEMA_reg_buffer_3112 ( .C (CLK), .D (new_AGEMA_signal_2304), .Q (new_AGEMA_signal_5880) ) ;
    buf_clk new_AGEMA_reg_buffer_3114 ( .C (CLK), .D (new_AGEMA_signal_2305), .Q (new_AGEMA_signal_5882) ) ;
    buf_clk new_AGEMA_reg_buffer_3122 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_3_L1), .Q (new_AGEMA_signal_5890) ) ;
    buf_clk new_AGEMA_reg_buffer_3126 ( .C (CLK), .D (new_AGEMA_signal_2182), .Q (new_AGEMA_signal_5894) ) ;
    buf_clk new_AGEMA_reg_buffer_3130 ( .C (CLK), .D (new_AGEMA_signal_2183), .Q (new_AGEMA_signal_5898) ) ;
    buf_clk new_AGEMA_reg_buffer_3140 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_4_Q3), .Q (new_AGEMA_signal_5908) ) ;
    buf_clk new_AGEMA_reg_buffer_3142 ( .C (CLK), .D (new_AGEMA_signal_2456), .Q (new_AGEMA_signal_5910) ) ;
    buf_clk new_AGEMA_reg_buffer_3144 ( .C (CLK), .D (new_AGEMA_signal_2457), .Q (new_AGEMA_signal_5912) ) ;
    buf_clk new_AGEMA_reg_buffer_3146 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_4_Q7), .Q (new_AGEMA_signal_5914) ) ;
    buf_clk new_AGEMA_reg_buffer_3148 ( .C (CLK), .D (new_AGEMA_signal_2458), .Q (new_AGEMA_signal_5916) ) ;
    buf_clk new_AGEMA_reg_buffer_3150 ( .C (CLK), .D (new_AGEMA_signal_2459), .Q (new_AGEMA_signal_5918) ) ;
    buf_clk new_AGEMA_reg_buffer_3158 ( .C (CLK), .D (LED_128_Instance_addconst_out[16]), .Q (new_AGEMA_signal_5926) ) ;
    buf_clk new_AGEMA_reg_buffer_3162 ( .C (CLK), .D (new_AGEMA_signal_2000), .Q (new_AGEMA_signal_5930) ) ;
    buf_clk new_AGEMA_reg_buffer_3166 ( .C (CLK), .D (new_AGEMA_signal_2001), .Q (new_AGEMA_signal_5934) ) ;
    buf_clk new_AGEMA_reg_buffer_3170 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_4_L1), .Q (new_AGEMA_signal_5938) ) ;
    buf_clk new_AGEMA_reg_buffer_3174 ( .C (CLK), .D (new_AGEMA_signal_2312), .Q (new_AGEMA_signal_5942) ) ;
    buf_clk new_AGEMA_reg_buffer_3178 ( .C (CLK), .D (new_AGEMA_signal_2313), .Q (new_AGEMA_signal_5946) ) ;
    buf_clk new_AGEMA_reg_buffer_3188 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_5_Q3), .Q (new_AGEMA_signal_5956) ) ;
    buf_clk new_AGEMA_reg_buffer_3190 ( .C (CLK), .D (new_AGEMA_signal_2466), .Q (new_AGEMA_signal_5958) ) ;
    buf_clk new_AGEMA_reg_buffer_3192 ( .C (CLK), .D (new_AGEMA_signal_2467), .Q (new_AGEMA_signal_5960) ) ;
    buf_clk new_AGEMA_reg_buffer_3194 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_5_Q7), .Q (new_AGEMA_signal_5962) ) ;
    buf_clk new_AGEMA_reg_buffer_3196 ( .C (CLK), .D (new_AGEMA_signal_2468), .Q (new_AGEMA_signal_5964) ) ;
    buf_clk new_AGEMA_reg_buffer_3198 ( .C (CLK), .D (new_AGEMA_signal_2469), .Q (new_AGEMA_signal_5966) ) ;
    buf_clk new_AGEMA_reg_buffer_3206 ( .C (CLK), .D (LED_128_Instance_addconst_out[20]), .Q (new_AGEMA_signal_5974) ) ;
    buf_clk new_AGEMA_reg_buffer_3210 ( .C (CLK), .D (new_AGEMA_signal_2154), .Q (new_AGEMA_signal_5978) ) ;
    buf_clk new_AGEMA_reg_buffer_3214 ( .C (CLK), .D (new_AGEMA_signal_2155), .Q (new_AGEMA_signal_5982) ) ;
    buf_clk new_AGEMA_reg_buffer_3218 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_5_L1), .Q (new_AGEMA_signal_5986) ) ;
    buf_clk new_AGEMA_reg_buffer_3222 ( .C (CLK), .D (new_AGEMA_signal_2320), .Q (new_AGEMA_signal_5990) ) ;
    buf_clk new_AGEMA_reg_buffer_3226 ( .C (CLK), .D (new_AGEMA_signal_2321), .Q (new_AGEMA_signal_5994) ) ;
    buf_clk new_AGEMA_reg_buffer_3236 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_6_Q3), .Q (new_AGEMA_signal_6004) ) ;
    buf_clk new_AGEMA_reg_buffer_3238 ( .C (CLK), .D (new_AGEMA_signal_2330), .Q (new_AGEMA_signal_6006) ) ;
    buf_clk new_AGEMA_reg_buffer_3240 ( .C (CLK), .D (new_AGEMA_signal_2331), .Q (new_AGEMA_signal_6008) ) ;
    buf_clk new_AGEMA_reg_buffer_3242 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_6_Q7), .Q (new_AGEMA_signal_6010) ) ;
    buf_clk new_AGEMA_reg_buffer_3244 ( .C (CLK), .D (new_AGEMA_signal_2332), .Q (new_AGEMA_signal_6012) ) ;
    buf_clk new_AGEMA_reg_buffer_3246 ( .C (CLK), .D (new_AGEMA_signal_2333), .Q (new_AGEMA_signal_6014) ) ;
    buf_clk new_AGEMA_reg_buffer_3254 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_6_L1), .Q (new_AGEMA_signal_6022) ) ;
    buf_clk new_AGEMA_reg_buffer_3258 ( .C (CLK), .D (new_AGEMA_signal_2196), .Q (new_AGEMA_signal_6026) ) ;
    buf_clk new_AGEMA_reg_buffer_3262 ( .C (CLK), .D (new_AGEMA_signal_2197), .Q (new_AGEMA_signal_6030) ) ;
    buf_clk new_AGEMA_reg_buffer_3272 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_7_Q3), .Q (new_AGEMA_signal_6040) ) ;
    buf_clk new_AGEMA_reg_buffer_3274 ( .C (CLK), .D (new_AGEMA_signal_2340), .Q (new_AGEMA_signal_6042) ) ;
    buf_clk new_AGEMA_reg_buffer_3276 ( .C (CLK), .D (new_AGEMA_signal_2341), .Q (new_AGEMA_signal_6044) ) ;
    buf_clk new_AGEMA_reg_buffer_3278 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_7_Q7), .Q (new_AGEMA_signal_6046) ) ;
    buf_clk new_AGEMA_reg_buffer_3280 ( .C (CLK), .D (new_AGEMA_signal_2342), .Q (new_AGEMA_signal_6048) ) ;
    buf_clk new_AGEMA_reg_buffer_3282 ( .C (CLK), .D (new_AGEMA_signal_2343), .Q (new_AGEMA_signal_6050) ) ;
    buf_clk new_AGEMA_reg_buffer_3290 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_7_L1), .Q (new_AGEMA_signal_6058) ) ;
    buf_clk new_AGEMA_reg_buffer_3294 ( .C (CLK), .D (new_AGEMA_signal_2208), .Q (new_AGEMA_signal_6062) ) ;
    buf_clk new_AGEMA_reg_buffer_3298 ( .C (CLK), .D (new_AGEMA_signal_2209), .Q (new_AGEMA_signal_6066) ) ;
    buf_clk new_AGEMA_reg_buffer_3308 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_8_Q3), .Q (new_AGEMA_signal_6076) ) ;
    buf_clk new_AGEMA_reg_buffer_3310 ( .C (CLK), .D (new_AGEMA_signal_2484), .Q (new_AGEMA_signal_6078) ) ;
    buf_clk new_AGEMA_reg_buffer_3312 ( .C (CLK), .D (new_AGEMA_signal_2485), .Q (new_AGEMA_signal_6080) ) ;
    buf_clk new_AGEMA_reg_buffer_3314 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_8_Q7), .Q (new_AGEMA_signal_6082) ) ;
    buf_clk new_AGEMA_reg_buffer_3316 ( .C (CLK), .D (new_AGEMA_signal_2486), .Q (new_AGEMA_signal_6084) ) ;
    buf_clk new_AGEMA_reg_buffer_3318 ( .C (CLK), .D (new_AGEMA_signal_2487), .Q (new_AGEMA_signal_6086) ) ;
    buf_clk new_AGEMA_reg_buffer_3326 ( .C (CLK), .D (LED_128_Instance_addconst_out[32]), .Q (new_AGEMA_signal_6094) ) ;
    buf_clk new_AGEMA_reg_buffer_3330 ( .C (CLK), .D (new_AGEMA_signal_2112), .Q (new_AGEMA_signal_6098) ) ;
    buf_clk new_AGEMA_reg_buffer_3334 ( .C (CLK), .D (new_AGEMA_signal_2113), .Q (new_AGEMA_signal_6102) ) ;
    buf_clk new_AGEMA_reg_buffer_3338 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_8_L1), .Q (new_AGEMA_signal_6106) ) ;
    buf_clk new_AGEMA_reg_buffer_3342 ( .C (CLK), .D (new_AGEMA_signal_2350), .Q (new_AGEMA_signal_6110) ) ;
    buf_clk new_AGEMA_reg_buffer_3346 ( .C (CLK), .D (new_AGEMA_signal_2351), .Q (new_AGEMA_signal_6114) ) ;
    buf_clk new_AGEMA_reg_buffer_3356 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_9_Q3), .Q (new_AGEMA_signal_6124) ) ;
    buf_clk new_AGEMA_reg_buffer_3358 ( .C (CLK), .D (new_AGEMA_signal_2494), .Q (new_AGEMA_signal_6126) ) ;
    buf_clk new_AGEMA_reg_buffer_3360 ( .C (CLK), .D (new_AGEMA_signal_2495), .Q (new_AGEMA_signal_6128) ) ;
    buf_clk new_AGEMA_reg_buffer_3362 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_9_Q7), .Q (new_AGEMA_signal_6130) ) ;
    buf_clk new_AGEMA_reg_buffer_3364 ( .C (CLK), .D (new_AGEMA_signal_2496), .Q (new_AGEMA_signal_6132) ) ;
    buf_clk new_AGEMA_reg_buffer_3366 ( .C (CLK), .D (new_AGEMA_signal_2497), .Q (new_AGEMA_signal_6134) ) ;
    buf_clk new_AGEMA_reg_buffer_3374 ( .C (CLK), .D (LED_128_Instance_addconst_out[36]), .Q (new_AGEMA_signal_6142) ) ;
    buf_clk new_AGEMA_reg_buffer_3378 ( .C (CLK), .D (new_AGEMA_signal_2106), .Q (new_AGEMA_signal_6146) ) ;
    buf_clk new_AGEMA_reg_buffer_3382 ( .C (CLK), .D (new_AGEMA_signal_2107), .Q (new_AGEMA_signal_6150) ) ;
    buf_clk new_AGEMA_reg_buffer_3386 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_9_L1), .Q (new_AGEMA_signal_6154) ) ;
    buf_clk new_AGEMA_reg_buffer_3390 ( .C (CLK), .D (new_AGEMA_signal_2358), .Q (new_AGEMA_signal_6158) ) ;
    buf_clk new_AGEMA_reg_buffer_3394 ( .C (CLK), .D (new_AGEMA_signal_2359), .Q (new_AGEMA_signal_6162) ) ;
    buf_clk new_AGEMA_reg_buffer_3404 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_10_Q3), .Q (new_AGEMA_signal_6172) ) ;
    buf_clk new_AGEMA_reg_buffer_3406 ( .C (CLK), .D (new_AGEMA_signal_2366), .Q (new_AGEMA_signal_6174) ) ;
    buf_clk new_AGEMA_reg_buffer_3408 ( .C (CLK), .D (new_AGEMA_signal_2367), .Q (new_AGEMA_signal_6176) ) ;
    buf_clk new_AGEMA_reg_buffer_3410 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_10_Q7), .Q (new_AGEMA_signal_6178) ) ;
    buf_clk new_AGEMA_reg_buffer_3412 ( .C (CLK), .D (new_AGEMA_signal_2368), .Q (new_AGEMA_signal_6180) ) ;
    buf_clk new_AGEMA_reg_buffer_3414 ( .C (CLK), .D (new_AGEMA_signal_2369), .Q (new_AGEMA_signal_6182) ) ;
    buf_clk new_AGEMA_reg_buffer_3422 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_10_L1), .Q (new_AGEMA_signal_6190) ) ;
    buf_clk new_AGEMA_reg_buffer_3426 ( .C (CLK), .D (new_AGEMA_signal_2226), .Q (new_AGEMA_signal_6194) ) ;
    buf_clk new_AGEMA_reg_buffer_3430 ( .C (CLK), .D (new_AGEMA_signal_2227), .Q (new_AGEMA_signal_6198) ) ;
    buf_clk new_AGEMA_reg_buffer_3440 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_11_Q3), .Q (new_AGEMA_signal_6208) ) ;
    buf_clk new_AGEMA_reg_buffer_3442 ( .C (CLK), .D (new_AGEMA_signal_2376), .Q (new_AGEMA_signal_6210) ) ;
    buf_clk new_AGEMA_reg_buffer_3444 ( .C (CLK), .D (new_AGEMA_signal_2377), .Q (new_AGEMA_signal_6212) ) ;
    buf_clk new_AGEMA_reg_buffer_3446 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_11_Q7), .Q (new_AGEMA_signal_6214) ) ;
    buf_clk new_AGEMA_reg_buffer_3448 ( .C (CLK), .D (new_AGEMA_signal_2378), .Q (new_AGEMA_signal_6216) ) ;
    buf_clk new_AGEMA_reg_buffer_3450 ( .C (CLK), .D (new_AGEMA_signal_2379), .Q (new_AGEMA_signal_6218) ) ;
    buf_clk new_AGEMA_reg_buffer_3458 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_11_L1), .Q (new_AGEMA_signal_6226) ) ;
    buf_clk new_AGEMA_reg_buffer_3462 ( .C (CLK), .D (new_AGEMA_signal_2238), .Q (new_AGEMA_signal_6230) ) ;
    buf_clk new_AGEMA_reg_buffer_3466 ( .C (CLK), .D (new_AGEMA_signal_2239), .Q (new_AGEMA_signal_6234) ) ;
    buf_clk new_AGEMA_reg_buffer_3476 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_12_Q3), .Q (new_AGEMA_signal_6244) ) ;
    buf_clk new_AGEMA_reg_buffer_3478 ( .C (CLK), .D (new_AGEMA_signal_2512), .Q (new_AGEMA_signal_6246) ) ;
    buf_clk new_AGEMA_reg_buffer_3480 ( .C (CLK), .D (new_AGEMA_signal_2513), .Q (new_AGEMA_signal_6248) ) ;
    buf_clk new_AGEMA_reg_buffer_3482 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_12_Q7), .Q (new_AGEMA_signal_6250) ) ;
    buf_clk new_AGEMA_reg_buffer_3484 ( .C (CLK), .D (new_AGEMA_signal_2514), .Q (new_AGEMA_signal_6252) ) ;
    buf_clk new_AGEMA_reg_buffer_3486 ( .C (CLK), .D (new_AGEMA_signal_2515), .Q (new_AGEMA_signal_6254) ) ;
    buf_clk new_AGEMA_reg_buffer_3494 ( .C (CLK), .D (LED_128_Instance_addconst_out[48]), .Q (new_AGEMA_signal_6262) ) ;
    buf_clk new_AGEMA_reg_buffer_3498 ( .C (CLK), .D (new_AGEMA_signal_2142), .Q (new_AGEMA_signal_6266) ) ;
    buf_clk new_AGEMA_reg_buffer_3502 ( .C (CLK), .D (new_AGEMA_signal_2143), .Q (new_AGEMA_signal_6270) ) ;
    buf_clk new_AGEMA_reg_buffer_3506 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_12_L1), .Q (new_AGEMA_signal_6274) ) ;
    buf_clk new_AGEMA_reg_buffer_3510 ( .C (CLK), .D (new_AGEMA_signal_2388), .Q (new_AGEMA_signal_6278) ) ;
    buf_clk new_AGEMA_reg_buffer_3514 ( .C (CLK), .D (new_AGEMA_signal_2389), .Q (new_AGEMA_signal_6282) ) ;
    buf_clk new_AGEMA_reg_buffer_3524 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_13_Q3), .Q (new_AGEMA_signal_6292) ) ;
    buf_clk new_AGEMA_reg_buffer_3526 ( .C (CLK), .D (new_AGEMA_signal_2522), .Q (new_AGEMA_signal_6294) ) ;
    buf_clk new_AGEMA_reg_buffer_3528 ( .C (CLK), .D (new_AGEMA_signal_2523), .Q (new_AGEMA_signal_6296) ) ;
    buf_clk new_AGEMA_reg_buffer_3530 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_13_Q7), .Q (new_AGEMA_signal_6298) ) ;
    buf_clk new_AGEMA_reg_buffer_3532 ( .C (CLK), .D (new_AGEMA_signal_2524), .Q (new_AGEMA_signal_6300) ) ;
    buf_clk new_AGEMA_reg_buffer_3534 ( .C (CLK), .D (new_AGEMA_signal_2525), .Q (new_AGEMA_signal_6302) ) ;
    buf_clk new_AGEMA_reg_buffer_3542 ( .C (CLK), .D (LED_128_Instance_addconst_out[52]), .Q (new_AGEMA_signal_6310) ) ;
    buf_clk new_AGEMA_reg_buffer_3546 ( .C (CLK), .D (new_AGEMA_signal_2132), .Q (new_AGEMA_signal_6314) ) ;
    buf_clk new_AGEMA_reg_buffer_3550 ( .C (CLK), .D (new_AGEMA_signal_2133), .Q (new_AGEMA_signal_6318) ) ;
    buf_clk new_AGEMA_reg_buffer_3554 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_13_L1), .Q (new_AGEMA_signal_6322) ) ;
    buf_clk new_AGEMA_reg_buffer_3558 ( .C (CLK), .D (new_AGEMA_signal_2398), .Q (new_AGEMA_signal_6326) ) ;
    buf_clk new_AGEMA_reg_buffer_3562 ( .C (CLK), .D (new_AGEMA_signal_2399), .Q (new_AGEMA_signal_6330) ) ;
    buf_clk new_AGEMA_reg_buffer_3572 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_14_Q3), .Q (new_AGEMA_signal_6340) ) ;
    buf_clk new_AGEMA_reg_buffer_3574 ( .C (CLK), .D (new_AGEMA_signal_2408), .Q (new_AGEMA_signal_6342) ) ;
    buf_clk new_AGEMA_reg_buffer_3576 ( .C (CLK), .D (new_AGEMA_signal_2409), .Q (new_AGEMA_signal_6344) ) ;
    buf_clk new_AGEMA_reg_buffer_3578 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_14_Q7), .Q (new_AGEMA_signal_6346) ) ;
    buf_clk new_AGEMA_reg_buffer_3580 ( .C (CLK), .D (new_AGEMA_signal_2410), .Q (new_AGEMA_signal_6348) ) ;
    buf_clk new_AGEMA_reg_buffer_3582 ( .C (CLK), .D (new_AGEMA_signal_2411), .Q (new_AGEMA_signal_6350) ) ;
    buf_clk new_AGEMA_reg_buffer_3590 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_14_L1), .Q (new_AGEMA_signal_6358) ) ;
    buf_clk new_AGEMA_reg_buffer_3594 ( .C (CLK), .D (new_AGEMA_signal_2252), .Q (new_AGEMA_signal_6362) ) ;
    buf_clk new_AGEMA_reg_buffer_3598 ( .C (CLK), .D (new_AGEMA_signal_2253), .Q (new_AGEMA_signal_6366) ) ;
    buf_clk new_AGEMA_reg_buffer_3608 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_15_Q3), .Q (new_AGEMA_signal_6376) ) ;
    buf_clk new_AGEMA_reg_buffer_3610 ( .C (CLK), .D (new_AGEMA_signal_2418), .Q (new_AGEMA_signal_6378) ) ;
    buf_clk new_AGEMA_reg_buffer_3612 ( .C (CLK), .D (new_AGEMA_signal_2419), .Q (new_AGEMA_signal_6380) ) ;
    buf_clk new_AGEMA_reg_buffer_3614 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_15_Q7), .Q (new_AGEMA_signal_6382) ) ;
    buf_clk new_AGEMA_reg_buffer_3616 ( .C (CLK), .D (new_AGEMA_signal_2420), .Q (new_AGEMA_signal_6384) ) ;
    buf_clk new_AGEMA_reg_buffer_3618 ( .C (CLK), .D (new_AGEMA_signal_2421), .Q (new_AGEMA_signal_6386) ) ;
    buf_clk new_AGEMA_reg_buffer_3626 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_15_L1), .Q (new_AGEMA_signal_6394) ) ;
    buf_clk new_AGEMA_reg_buffer_3630 ( .C (CLK), .D (new_AGEMA_signal_2264), .Q (new_AGEMA_signal_6398) ) ;
    buf_clk new_AGEMA_reg_buffer_3634 ( .C (CLK), .D (new_AGEMA_signal_2265), .Q (new_AGEMA_signal_6402) ) ;
    buf_clk new_AGEMA_reg_buffer_3740 ( .C (CLK), .D (LED_128_Instance_N10), .Q (new_AGEMA_signal_6508) ) ;
    buf_clk new_AGEMA_reg_buffer_3744 ( .C (CLK), .D (LED_128_Instance_N11), .Q (new_AGEMA_signal_6512) ) ;
    buf_clk new_AGEMA_reg_buffer_3748 ( .C (CLK), .D (LED_128_Instance_N12), .Q (new_AGEMA_signal_6516) ) ;
    buf_clk new_AGEMA_reg_buffer_3752 ( .C (CLK), .D (LED_128_Instance_N13), .Q (new_AGEMA_signal_6520) ) ;
    buf_clk new_AGEMA_reg_buffer_3756 ( .C (CLK), .D (LED_128_Instance_N4), .Q (new_AGEMA_signal_6524) ) ;
    buf_clk new_AGEMA_reg_buffer_3760 ( .C (CLK), .D (LED_128_Instance_N5), .Q (new_AGEMA_signal_6528) ) ;
    buf_clk new_AGEMA_reg_buffer_3764 ( .C (CLK), .D (LED_128_Instance_N6), .Q (new_AGEMA_signal_6532) ) ;
    buf_clk new_AGEMA_reg_buffer_3768 ( .C (CLK), .D (LED_128_Instance_N7), .Q (new_AGEMA_signal_6536) ) ;
    buf_clk new_AGEMA_reg_buffer_3772 ( .C (CLK), .D (LED_128_Instance_N8), .Q (new_AGEMA_signal_6540) ) ;
    buf_clk new_AGEMA_reg_buffer_3776 ( .C (CLK), .D (LED_128_Instance_N9), .Q (new_AGEMA_signal_6544) ) ;
    buf_clk new_AGEMA_reg_buffer_3780 ( .C (CLK), .D (n15), .Q (new_AGEMA_signal_6548) ) ;

    /* cells in depth 2 */
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR16_U1 ( .a ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, LED_128_Instance_SBox_Instance_0_T0}), .b ({new_AGEMA_signal_3901, new_AGEMA_signal_3899, new_AGEMA_signal_3897}), .c ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, LED_128_Instance_SBox_Instance_0_Q2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR7_U1 ( .a ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, LED_128_Instance_SBox_Instance_0_T0}), .b ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, LED_128_Instance_SBox_Instance_0_T2}), .c ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, LED_128_Instance_SBox_Instance_0_L5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR8_U1 ( .a ({new_AGEMA_signal_3907, new_AGEMA_signal_3905, new_AGEMA_signal_3903}), .b ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, LED_128_Instance_SBox_Instance_0_L5}), .c ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, LED_128_Instance_SBox_Instance_0_Q6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_AND1_U1 ( .a ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, LED_128_Instance_SBox_Instance_0_n1}), .b ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, LED_128_Instance_SBox_Instance_0_n2}), .clk (CLK), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, LED_128_Instance_SBox_Instance_0_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_AND3_U1 ( .a ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, LED_128_Instance_SBox_Instance_0_n3}), .b ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, LED_128_Instance_addconst_out[2]}), .clk (CLK), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, LED_128_Instance_SBox_Instance_0_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR15_U1 ( .a ({new_AGEMA_signal_3913, new_AGEMA_signal_3911, new_AGEMA_signal_3909}), .b ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, LED_128_Instance_SBox_Instance_0_T2}), .c ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, LED_128_Instance_subcells_out[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR16_U1 ( .a ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, LED_128_Instance_SBox_Instance_1_T0}), .b ({new_AGEMA_signal_3919, new_AGEMA_signal_3917, new_AGEMA_signal_3915}), .c ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, LED_128_Instance_SBox_Instance_1_Q2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR7_U1 ( .a ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, LED_128_Instance_SBox_Instance_1_T0}), .b ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, LED_128_Instance_SBox_Instance_1_T2}), .c ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, LED_128_Instance_SBox_Instance_1_L5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR8_U1 ( .a ({new_AGEMA_signal_3925, new_AGEMA_signal_3923, new_AGEMA_signal_3921}), .b ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, LED_128_Instance_SBox_Instance_1_L5}), .c ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, LED_128_Instance_SBox_Instance_1_Q6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_AND1_U1 ( .a ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, LED_128_Instance_SBox_Instance_1_n1}), .b ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, LED_128_Instance_SBox_Instance_1_n2}), .clk (CLK), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, LED_128_Instance_SBox_Instance_1_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_AND3_U1 ( .a ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, LED_128_Instance_SBox_Instance_1_n3}), .b ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, LED_128_Instance_addconst_out[6]}), .clk (CLK), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, LED_128_Instance_SBox_Instance_1_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR15_U1 ( .a ({new_AGEMA_signal_3931, new_AGEMA_signal_3929, new_AGEMA_signal_3927}), .b ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, LED_128_Instance_SBox_Instance_1_T2}), .c ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, LED_128_Instance_subcells_out[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR16_U1 ( .a ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, LED_128_Instance_SBox_Instance_2_T0}), .b ({new_AGEMA_signal_3937, new_AGEMA_signal_3935, new_AGEMA_signal_3933}), .c ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, LED_128_Instance_SBox_Instance_2_Q2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR7_U1 ( .a ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, LED_128_Instance_SBox_Instance_2_T0}), .b ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, LED_128_Instance_SBox_Instance_2_T2}), .c ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, LED_128_Instance_SBox_Instance_2_L5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR8_U1 ( .a ({new_AGEMA_signal_3943, new_AGEMA_signal_3941, new_AGEMA_signal_3939}), .b ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, LED_128_Instance_SBox_Instance_2_L5}), .c ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, LED_128_Instance_SBox_Instance_2_Q6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_AND1_U1 ( .a ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, LED_128_Instance_SBox_Instance_2_n1}), .b ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, LED_128_Instance_SBox_Instance_2_n2}), .clk (CLK), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, LED_128_Instance_SBox_Instance_2_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_AND3_U1 ( .a ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, LED_128_Instance_SBox_Instance_2_n3}), .b ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, LED_128_Instance_addconst_out[10]}), .clk (CLK), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, LED_128_Instance_SBox_Instance_2_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR15_U1 ( .a ({new_AGEMA_signal_3949, new_AGEMA_signal_3947, new_AGEMA_signal_3945}), .b ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, LED_128_Instance_SBox_Instance_2_T2}), .c ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, LED_128_Instance_subcells_out[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR16_U1 ( .a ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, LED_128_Instance_SBox_Instance_3_T0}), .b ({new_AGEMA_signal_3955, new_AGEMA_signal_3953, new_AGEMA_signal_3951}), .c ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, LED_128_Instance_SBox_Instance_3_Q2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR7_U1 ( .a ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, LED_128_Instance_SBox_Instance_3_T0}), .b ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, LED_128_Instance_SBox_Instance_3_T2}), .c ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, LED_128_Instance_SBox_Instance_3_L5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR8_U1 ( .a ({new_AGEMA_signal_3961, new_AGEMA_signal_3959, new_AGEMA_signal_3957}), .b ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, LED_128_Instance_SBox_Instance_3_L5}), .c ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, LED_128_Instance_SBox_Instance_3_Q6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_AND1_U1 ( .a ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, LED_128_Instance_SBox_Instance_3_n1}), .b ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, LED_128_Instance_SBox_Instance_3_n2}), .clk (CLK), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, LED_128_Instance_SBox_Instance_3_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_AND3_U1 ( .a ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, LED_128_Instance_SBox_Instance_3_n3}), .b ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, LED_128_Instance_addconst_out[14]}), .clk (CLK), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, LED_128_Instance_SBox_Instance_3_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR15_U1 ( .a ({new_AGEMA_signal_3967, new_AGEMA_signal_3965, new_AGEMA_signal_3963}), .b ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, LED_128_Instance_SBox_Instance_3_T2}), .c ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, LED_128_Instance_subcells_out[12]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR16_U1 ( .a ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, LED_128_Instance_SBox_Instance_4_T0}), .b ({new_AGEMA_signal_3973, new_AGEMA_signal_3971, new_AGEMA_signal_3969}), .c ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, LED_128_Instance_SBox_Instance_4_Q2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR7_U1 ( .a ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, LED_128_Instance_SBox_Instance_4_T0}), .b ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, LED_128_Instance_SBox_Instance_4_T2}), .c ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, LED_128_Instance_SBox_Instance_4_L5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR8_U1 ( .a ({new_AGEMA_signal_3979, new_AGEMA_signal_3977, new_AGEMA_signal_3975}), .b ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, LED_128_Instance_SBox_Instance_4_L5}), .c ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, LED_128_Instance_SBox_Instance_4_Q6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_AND1_U1 ( .a ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, LED_128_Instance_SBox_Instance_4_n1}), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, LED_128_Instance_SBox_Instance_4_n2}), .clk (CLK), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, LED_128_Instance_SBox_Instance_4_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_AND3_U1 ( .a ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, LED_128_Instance_SBox_Instance_4_n3}), .b ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, LED_128_Instance_addconst_out[18]}), .clk (CLK), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, LED_128_Instance_SBox_Instance_4_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR15_U1 ( .a ({new_AGEMA_signal_3985, new_AGEMA_signal_3983, new_AGEMA_signal_3981}), .b ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, LED_128_Instance_SBox_Instance_4_T2}), .c ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, LED_128_Instance_subcells_out[16]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR16_U1 ( .a ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, LED_128_Instance_SBox_Instance_5_T0}), .b ({new_AGEMA_signal_3991, new_AGEMA_signal_3989, new_AGEMA_signal_3987}), .c ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, LED_128_Instance_SBox_Instance_5_Q2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR7_U1 ( .a ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, LED_128_Instance_SBox_Instance_5_T0}), .b ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, LED_128_Instance_SBox_Instance_5_T2}), .c ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, LED_128_Instance_SBox_Instance_5_L5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR8_U1 ( .a ({new_AGEMA_signal_3997, new_AGEMA_signal_3995, new_AGEMA_signal_3993}), .b ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, LED_128_Instance_SBox_Instance_5_L5}), .c ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, LED_128_Instance_SBox_Instance_5_Q6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_AND1_U1 ( .a ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, LED_128_Instance_SBox_Instance_5_n1}), .b ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, LED_128_Instance_SBox_Instance_5_n2}), .clk (CLK), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, LED_128_Instance_SBox_Instance_5_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_AND3_U1 ( .a ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, LED_128_Instance_SBox_Instance_5_n3}), .b ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_addconst_out[22]}), .clk (CLK), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, LED_128_Instance_SBox_Instance_5_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR15_U1 ( .a ({new_AGEMA_signal_4003, new_AGEMA_signal_4001, new_AGEMA_signal_3999}), .b ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, LED_128_Instance_SBox_Instance_5_T2}), .c ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, LED_128_Instance_subcells_out[20]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR16_U1 ( .a ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, LED_128_Instance_SBox_Instance_6_T0}), .b ({new_AGEMA_signal_4009, new_AGEMA_signal_4007, new_AGEMA_signal_4005}), .c ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, LED_128_Instance_SBox_Instance_6_Q2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR7_U1 ( .a ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, LED_128_Instance_SBox_Instance_6_T0}), .b ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, LED_128_Instance_SBox_Instance_6_T2}), .c ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, LED_128_Instance_SBox_Instance_6_L5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR8_U1 ( .a ({new_AGEMA_signal_4015, new_AGEMA_signal_4013, new_AGEMA_signal_4011}), .b ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, LED_128_Instance_SBox_Instance_6_L5}), .c ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, LED_128_Instance_SBox_Instance_6_Q6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_AND1_U1 ( .a ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, LED_128_Instance_SBox_Instance_6_n1}), .b ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, LED_128_Instance_SBox_Instance_6_n2}), .clk (CLK), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, LED_128_Instance_SBox_Instance_6_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_AND3_U1 ( .a ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, LED_128_Instance_SBox_Instance_6_n3}), .b ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_addconst_out[26]}), .clk (CLK), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, LED_128_Instance_SBox_Instance_6_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR15_U1 ( .a ({new_AGEMA_signal_4021, new_AGEMA_signal_4019, new_AGEMA_signal_4017}), .b ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, LED_128_Instance_SBox_Instance_6_T2}), .c ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, LED_128_Instance_subcells_out[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR16_U1 ( .a ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, LED_128_Instance_SBox_Instance_7_T0}), .b ({new_AGEMA_signal_4027, new_AGEMA_signal_4025, new_AGEMA_signal_4023}), .c ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, LED_128_Instance_SBox_Instance_7_Q2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR7_U1 ( .a ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, LED_128_Instance_SBox_Instance_7_T0}), .b ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, LED_128_Instance_SBox_Instance_7_T2}), .c ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, LED_128_Instance_SBox_Instance_7_L5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR8_U1 ( .a ({new_AGEMA_signal_4033, new_AGEMA_signal_4031, new_AGEMA_signal_4029}), .b ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, LED_128_Instance_SBox_Instance_7_L5}), .c ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, LED_128_Instance_SBox_Instance_7_Q6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_AND1_U1 ( .a ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, LED_128_Instance_SBox_Instance_7_n1}), .b ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, LED_128_Instance_SBox_Instance_7_n2}), .clk (CLK), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, LED_128_Instance_SBox_Instance_7_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_AND3_U1 ( .a ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, LED_128_Instance_SBox_Instance_7_n3}), .b ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, LED_128_Instance_addconst_out[30]}), .clk (CLK), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, LED_128_Instance_SBox_Instance_7_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR15_U1 ( .a ({new_AGEMA_signal_4039, new_AGEMA_signal_4037, new_AGEMA_signal_4035}), .b ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, LED_128_Instance_SBox_Instance_7_T2}), .c ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, LED_128_Instance_subcells_out[28]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR16_U1 ( .a ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, LED_128_Instance_SBox_Instance_8_T0}), .b ({new_AGEMA_signal_4045, new_AGEMA_signal_4043, new_AGEMA_signal_4041}), .c ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, LED_128_Instance_SBox_Instance_8_Q2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR7_U1 ( .a ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, LED_128_Instance_SBox_Instance_8_T0}), .b ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, LED_128_Instance_SBox_Instance_8_T2}), .c ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, LED_128_Instance_SBox_Instance_8_L5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR8_U1 ( .a ({new_AGEMA_signal_4051, new_AGEMA_signal_4049, new_AGEMA_signal_4047}), .b ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, LED_128_Instance_SBox_Instance_8_L5}), .c ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, LED_128_Instance_SBox_Instance_8_Q6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_AND1_U1 ( .a ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, LED_128_Instance_SBox_Instance_8_n1}), .b ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, LED_128_Instance_SBox_Instance_8_n2}), .clk (CLK), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, LED_128_Instance_SBox_Instance_8_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_AND3_U1 ( .a ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, LED_128_Instance_SBox_Instance_8_n3}), .b ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, LED_128_Instance_addconst_out[34]}), .clk (CLK), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, LED_128_Instance_SBox_Instance_8_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR15_U1 ( .a ({new_AGEMA_signal_4057, new_AGEMA_signal_4055, new_AGEMA_signal_4053}), .b ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, LED_128_Instance_SBox_Instance_8_T2}), .c ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, LED_128_Instance_subcells_out[32]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR16_U1 ( .a ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, LED_128_Instance_SBox_Instance_9_T0}), .b ({new_AGEMA_signal_4063, new_AGEMA_signal_4061, new_AGEMA_signal_4059}), .c ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, LED_128_Instance_SBox_Instance_9_Q2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR7_U1 ( .a ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, LED_128_Instance_SBox_Instance_9_T0}), .b ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, LED_128_Instance_SBox_Instance_9_T2}), .c ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, LED_128_Instance_SBox_Instance_9_L5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR8_U1 ( .a ({new_AGEMA_signal_4069, new_AGEMA_signal_4067, new_AGEMA_signal_4065}), .b ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, LED_128_Instance_SBox_Instance_9_L5}), .c ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, LED_128_Instance_SBox_Instance_9_Q6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_AND1_U1 ( .a ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, LED_128_Instance_SBox_Instance_9_n1}), .b ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, LED_128_Instance_SBox_Instance_9_n2}), .clk (CLK), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, LED_128_Instance_SBox_Instance_9_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_AND3_U1 ( .a ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, LED_128_Instance_SBox_Instance_9_n3}), .b ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, LED_128_Instance_addconst_out[38]}), .clk (CLK), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, LED_128_Instance_SBox_Instance_9_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR15_U1 ( .a ({new_AGEMA_signal_4075, new_AGEMA_signal_4073, new_AGEMA_signal_4071}), .b ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, LED_128_Instance_SBox_Instance_9_T2}), .c ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, LED_128_Instance_subcells_out[36]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR16_U1 ( .a ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, LED_128_Instance_SBox_Instance_10_T0}), .b ({new_AGEMA_signal_4081, new_AGEMA_signal_4079, new_AGEMA_signal_4077}), .c ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, LED_128_Instance_SBox_Instance_10_Q2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR7_U1 ( .a ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, LED_128_Instance_SBox_Instance_10_T0}), .b ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, LED_128_Instance_SBox_Instance_10_T2}), .c ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, LED_128_Instance_SBox_Instance_10_L5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR8_U1 ( .a ({new_AGEMA_signal_4087, new_AGEMA_signal_4085, new_AGEMA_signal_4083}), .b ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, LED_128_Instance_SBox_Instance_10_L5}), .c ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, LED_128_Instance_SBox_Instance_10_Q6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_AND1_U1 ( .a ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, LED_128_Instance_SBox_Instance_10_n1}), .b ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, LED_128_Instance_SBox_Instance_10_n2}), .clk (CLK), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, LED_128_Instance_SBox_Instance_10_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_AND3_U1 ( .a ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, LED_128_Instance_SBox_Instance_10_n3}), .b ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, LED_128_Instance_addconst_out[42]}), .clk (CLK), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, LED_128_Instance_SBox_Instance_10_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR15_U1 ( .a ({new_AGEMA_signal_4093, new_AGEMA_signal_4091, new_AGEMA_signal_4089}), .b ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, LED_128_Instance_SBox_Instance_10_T2}), .c ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, LED_128_Instance_subcells_out[40]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR16_U1 ( .a ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, LED_128_Instance_SBox_Instance_11_T0}), .b ({new_AGEMA_signal_4099, new_AGEMA_signal_4097, new_AGEMA_signal_4095}), .c ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, LED_128_Instance_SBox_Instance_11_Q2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR7_U1 ( .a ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, LED_128_Instance_SBox_Instance_11_T0}), .b ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, LED_128_Instance_SBox_Instance_11_T2}), .c ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, LED_128_Instance_SBox_Instance_11_L5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR8_U1 ( .a ({new_AGEMA_signal_4105, new_AGEMA_signal_4103, new_AGEMA_signal_4101}), .b ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, LED_128_Instance_SBox_Instance_11_L5}), .c ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, LED_128_Instance_SBox_Instance_11_Q6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_AND1_U1 ( .a ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, LED_128_Instance_SBox_Instance_11_n1}), .b ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, LED_128_Instance_SBox_Instance_11_n2}), .clk (CLK), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, LED_128_Instance_SBox_Instance_11_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_AND3_U1 ( .a ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, LED_128_Instance_SBox_Instance_11_n3}), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, LED_128_Instance_addconst_out[46]}), .clk (CLK), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, LED_128_Instance_SBox_Instance_11_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR15_U1 ( .a ({new_AGEMA_signal_4111, new_AGEMA_signal_4109, new_AGEMA_signal_4107}), .b ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, LED_128_Instance_SBox_Instance_11_T2}), .c ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, LED_128_Instance_subcells_out[44]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR16_U1 ( .a ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, LED_128_Instance_SBox_Instance_12_T0}), .b ({new_AGEMA_signal_4117, new_AGEMA_signal_4115, new_AGEMA_signal_4113}), .c ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, LED_128_Instance_SBox_Instance_12_Q2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR7_U1 ( .a ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, LED_128_Instance_SBox_Instance_12_T0}), .b ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, LED_128_Instance_SBox_Instance_12_T2}), .c ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, LED_128_Instance_SBox_Instance_12_L5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR8_U1 ( .a ({new_AGEMA_signal_4123, new_AGEMA_signal_4121, new_AGEMA_signal_4119}), .b ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, LED_128_Instance_SBox_Instance_12_L5}), .c ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, LED_128_Instance_SBox_Instance_12_Q6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_AND1_U1 ( .a ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, LED_128_Instance_SBox_Instance_12_n1}), .b ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, LED_128_Instance_SBox_Instance_12_n2}), .clk (CLK), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, LED_128_Instance_SBox_Instance_12_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_AND3_U1 ( .a ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, LED_128_Instance_SBox_Instance_12_n3}), .b ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, LED_128_Instance_addconst_out[50]}), .clk (CLK), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, LED_128_Instance_SBox_Instance_12_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR15_U1 ( .a ({new_AGEMA_signal_4129, new_AGEMA_signal_4127, new_AGEMA_signal_4125}), .b ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, LED_128_Instance_SBox_Instance_12_T2}), .c ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, LED_128_Instance_subcells_out[48]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR16_U1 ( .a ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, LED_128_Instance_SBox_Instance_13_T0}), .b ({new_AGEMA_signal_4135, new_AGEMA_signal_4133, new_AGEMA_signal_4131}), .c ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, LED_128_Instance_SBox_Instance_13_Q2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR7_U1 ( .a ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, LED_128_Instance_SBox_Instance_13_T0}), .b ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, LED_128_Instance_SBox_Instance_13_T2}), .c ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, LED_128_Instance_SBox_Instance_13_L5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR8_U1 ( .a ({new_AGEMA_signal_4141, new_AGEMA_signal_4139, new_AGEMA_signal_4137}), .b ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, LED_128_Instance_SBox_Instance_13_L5}), .c ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, LED_128_Instance_SBox_Instance_13_Q6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_AND1_U1 ( .a ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, LED_128_Instance_SBox_Instance_13_n1}), .b ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, LED_128_Instance_SBox_Instance_13_n2}), .clk (CLK), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, LED_128_Instance_SBox_Instance_13_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_AND3_U1 ( .a ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, LED_128_Instance_SBox_Instance_13_n3}), .b ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, LED_128_Instance_addconst_out[54]}), .clk (CLK), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, LED_128_Instance_SBox_Instance_13_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR15_U1 ( .a ({new_AGEMA_signal_4147, new_AGEMA_signal_4145, new_AGEMA_signal_4143}), .b ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, LED_128_Instance_SBox_Instance_13_T2}), .c ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, LED_128_Instance_subcells_out[52]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR16_U1 ( .a ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, LED_128_Instance_SBox_Instance_14_T0}), .b ({new_AGEMA_signal_4153, new_AGEMA_signal_4151, new_AGEMA_signal_4149}), .c ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, LED_128_Instance_SBox_Instance_14_Q2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR7_U1 ( .a ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, LED_128_Instance_SBox_Instance_14_T0}), .b ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, LED_128_Instance_SBox_Instance_14_T2}), .c ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, LED_128_Instance_SBox_Instance_14_L5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR8_U1 ( .a ({new_AGEMA_signal_4159, new_AGEMA_signal_4157, new_AGEMA_signal_4155}), .b ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, LED_128_Instance_SBox_Instance_14_L5}), .c ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, LED_128_Instance_SBox_Instance_14_Q6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_AND1_U1 ( .a ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, LED_128_Instance_SBox_Instance_14_n1}), .b ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, LED_128_Instance_SBox_Instance_14_n2}), .clk (CLK), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, LED_128_Instance_SBox_Instance_14_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_AND3_U1 ( .a ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, LED_128_Instance_SBox_Instance_14_n3}), .b ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, LED_128_Instance_addconst_out[58]}), .clk (CLK), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, LED_128_Instance_SBox_Instance_14_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR15_U1 ( .a ({new_AGEMA_signal_4165, new_AGEMA_signal_4163, new_AGEMA_signal_4161}), .b ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, LED_128_Instance_SBox_Instance_14_T2}), .c ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, LED_128_Instance_subcells_out[56]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR16_U1 ( .a ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, LED_128_Instance_SBox_Instance_15_T0}), .b ({new_AGEMA_signal_4171, new_AGEMA_signal_4169, new_AGEMA_signal_4167}), .c ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, LED_128_Instance_SBox_Instance_15_Q2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR7_U1 ( .a ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, LED_128_Instance_SBox_Instance_15_T0}), .b ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, LED_128_Instance_SBox_Instance_15_T2}), .c ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, LED_128_Instance_SBox_Instance_15_L5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR8_U1 ( .a ({new_AGEMA_signal_4177, new_AGEMA_signal_4175, new_AGEMA_signal_4173}), .b ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, LED_128_Instance_SBox_Instance_15_L5}), .c ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, LED_128_Instance_SBox_Instance_15_Q6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_AND1_U1 ( .a ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, LED_128_Instance_SBox_Instance_15_n1}), .b ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, LED_128_Instance_SBox_Instance_15_n2}), .clk (CLK), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, LED_128_Instance_SBox_Instance_15_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_AND3_U1 ( .a ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, LED_128_Instance_SBox_Instance_15_n3}), .b ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, LED_128_Instance_addconst_out[62]}), .clk (CLK), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, LED_128_Instance_SBox_Instance_15_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR15_U1 ( .a ({new_AGEMA_signal_4183, new_AGEMA_signal_4181, new_AGEMA_signal_4179}), .b ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, LED_128_Instance_SBox_Instance_15_T2}), .c ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, LED_128_Instance_subcells_out[60]}) ) ;
    buf_clk new_AGEMA_reg_buffer_1129 ( .C (CLK), .D (new_AGEMA_signal_3896), .Q (new_AGEMA_signal_3897) ) ;
    buf_clk new_AGEMA_reg_buffer_1131 ( .C (CLK), .D (new_AGEMA_signal_3898), .Q (new_AGEMA_signal_3899) ) ;
    buf_clk new_AGEMA_reg_buffer_1133 ( .C (CLK), .D (new_AGEMA_signal_3900), .Q (new_AGEMA_signal_3901) ) ;
    buf_clk new_AGEMA_reg_buffer_1135 ( .C (CLK), .D (new_AGEMA_signal_3902), .Q (new_AGEMA_signal_3903) ) ;
    buf_clk new_AGEMA_reg_buffer_1137 ( .C (CLK), .D (new_AGEMA_signal_3904), .Q (new_AGEMA_signal_3905) ) ;
    buf_clk new_AGEMA_reg_buffer_1139 ( .C (CLK), .D (new_AGEMA_signal_3906), .Q (new_AGEMA_signal_3907) ) ;
    buf_clk new_AGEMA_reg_buffer_1141 ( .C (CLK), .D (new_AGEMA_signal_3908), .Q (new_AGEMA_signal_3909) ) ;
    buf_clk new_AGEMA_reg_buffer_1143 ( .C (CLK), .D (new_AGEMA_signal_3910), .Q (new_AGEMA_signal_3911) ) ;
    buf_clk new_AGEMA_reg_buffer_1145 ( .C (CLK), .D (new_AGEMA_signal_3912), .Q (new_AGEMA_signal_3913) ) ;
    buf_clk new_AGEMA_reg_buffer_1147 ( .C (CLK), .D (new_AGEMA_signal_3914), .Q (new_AGEMA_signal_3915) ) ;
    buf_clk new_AGEMA_reg_buffer_1149 ( .C (CLK), .D (new_AGEMA_signal_3916), .Q (new_AGEMA_signal_3917) ) ;
    buf_clk new_AGEMA_reg_buffer_1151 ( .C (CLK), .D (new_AGEMA_signal_3918), .Q (new_AGEMA_signal_3919) ) ;
    buf_clk new_AGEMA_reg_buffer_1153 ( .C (CLK), .D (new_AGEMA_signal_3920), .Q (new_AGEMA_signal_3921) ) ;
    buf_clk new_AGEMA_reg_buffer_1155 ( .C (CLK), .D (new_AGEMA_signal_3922), .Q (new_AGEMA_signal_3923) ) ;
    buf_clk new_AGEMA_reg_buffer_1157 ( .C (CLK), .D (new_AGEMA_signal_3924), .Q (new_AGEMA_signal_3925) ) ;
    buf_clk new_AGEMA_reg_buffer_1159 ( .C (CLK), .D (new_AGEMA_signal_3926), .Q (new_AGEMA_signal_3927) ) ;
    buf_clk new_AGEMA_reg_buffer_1161 ( .C (CLK), .D (new_AGEMA_signal_3928), .Q (new_AGEMA_signal_3929) ) ;
    buf_clk new_AGEMA_reg_buffer_1163 ( .C (CLK), .D (new_AGEMA_signal_3930), .Q (new_AGEMA_signal_3931) ) ;
    buf_clk new_AGEMA_reg_buffer_1165 ( .C (CLK), .D (new_AGEMA_signal_3932), .Q (new_AGEMA_signal_3933) ) ;
    buf_clk new_AGEMA_reg_buffer_1167 ( .C (CLK), .D (new_AGEMA_signal_3934), .Q (new_AGEMA_signal_3935) ) ;
    buf_clk new_AGEMA_reg_buffer_1169 ( .C (CLK), .D (new_AGEMA_signal_3936), .Q (new_AGEMA_signal_3937) ) ;
    buf_clk new_AGEMA_reg_buffer_1171 ( .C (CLK), .D (new_AGEMA_signal_3938), .Q (new_AGEMA_signal_3939) ) ;
    buf_clk new_AGEMA_reg_buffer_1173 ( .C (CLK), .D (new_AGEMA_signal_3940), .Q (new_AGEMA_signal_3941) ) ;
    buf_clk new_AGEMA_reg_buffer_1175 ( .C (CLK), .D (new_AGEMA_signal_3942), .Q (new_AGEMA_signal_3943) ) ;
    buf_clk new_AGEMA_reg_buffer_1177 ( .C (CLK), .D (new_AGEMA_signal_3944), .Q (new_AGEMA_signal_3945) ) ;
    buf_clk new_AGEMA_reg_buffer_1179 ( .C (CLK), .D (new_AGEMA_signal_3946), .Q (new_AGEMA_signal_3947) ) ;
    buf_clk new_AGEMA_reg_buffer_1181 ( .C (CLK), .D (new_AGEMA_signal_3948), .Q (new_AGEMA_signal_3949) ) ;
    buf_clk new_AGEMA_reg_buffer_1183 ( .C (CLK), .D (new_AGEMA_signal_3950), .Q (new_AGEMA_signal_3951) ) ;
    buf_clk new_AGEMA_reg_buffer_1185 ( .C (CLK), .D (new_AGEMA_signal_3952), .Q (new_AGEMA_signal_3953) ) ;
    buf_clk new_AGEMA_reg_buffer_1187 ( .C (CLK), .D (new_AGEMA_signal_3954), .Q (new_AGEMA_signal_3955) ) ;
    buf_clk new_AGEMA_reg_buffer_1189 ( .C (CLK), .D (new_AGEMA_signal_3956), .Q (new_AGEMA_signal_3957) ) ;
    buf_clk new_AGEMA_reg_buffer_1191 ( .C (CLK), .D (new_AGEMA_signal_3958), .Q (new_AGEMA_signal_3959) ) ;
    buf_clk new_AGEMA_reg_buffer_1193 ( .C (CLK), .D (new_AGEMA_signal_3960), .Q (new_AGEMA_signal_3961) ) ;
    buf_clk new_AGEMA_reg_buffer_1195 ( .C (CLK), .D (new_AGEMA_signal_3962), .Q (new_AGEMA_signal_3963) ) ;
    buf_clk new_AGEMA_reg_buffer_1197 ( .C (CLK), .D (new_AGEMA_signal_3964), .Q (new_AGEMA_signal_3965) ) ;
    buf_clk new_AGEMA_reg_buffer_1199 ( .C (CLK), .D (new_AGEMA_signal_3966), .Q (new_AGEMA_signal_3967) ) ;
    buf_clk new_AGEMA_reg_buffer_1201 ( .C (CLK), .D (new_AGEMA_signal_3968), .Q (new_AGEMA_signal_3969) ) ;
    buf_clk new_AGEMA_reg_buffer_1203 ( .C (CLK), .D (new_AGEMA_signal_3970), .Q (new_AGEMA_signal_3971) ) ;
    buf_clk new_AGEMA_reg_buffer_1205 ( .C (CLK), .D (new_AGEMA_signal_3972), .Q (new_AGEMA_signal_3973) ) ;
    buf_clk new_AGEMA_reg_buffer_1207 ( .C (CLK), .D (new_AGEMA_signal_3974), .Q (new_AGEMA_signal_3975) ) ;
    buf_clk new_AGEMA_reg_buffer_1209 ( .C (CLK), .D (new_AGEMA_signal_3976), .Q (new_AGEMA_signal_3977) ) ;
    buf_clk new_AGEMA_reg_buffer_1211 ( .C (CLK), .D (new_AGEMA_signal_3978), .Q (new_AGEMA_signal_3979) ) ;
    buf_clk new_AGEMA_reg_buffer_1213 ( .C (CLK), .D (new_AGEMA_signal_3980), .Q (new_AGEMA_signal_3981) ) ;
    buf_clk new_AGEMA_reg_buffer_1215 ( .C (CLK), .D (new_AGEMA_signal_3982), .Q (new_AGEMA_signal_3983) ) ;
    buf_clk new_AGEMA_reg_buffer_1217 ( .C (CLK), .D (new_AGEMA_signal_3984), .Q (new_AGEMA_signal_3985) ) ;
    buf_clk new_AGEMA_reg_buffer_1219 ( .C (CLK), .D (new_AGEMA_signal_3986), .Q (new_AGEMA_signal_3987) ) ;
    buf_clk new_AGEMA_reg_buffer_1221 ( .C (CLK), .D (new_AGEMA_signal_3988), .Q (new_AGEMA_signal_3989) ) ;
    buf_clk new_AGEMA_reg_buffer_1223 ( .C (CLK), .D (new_AGEMA_signal_3990), .Q (new_AGEMA_signal_3991) ) ;
    buf_clk new_AGEMA_reg_buffer_1225 ( .C (CLK), .D (new_AGEMA_signal_3992), .Q (new_AGEMA_signal_3993) ) ;
    buf_clk new_AGEMA_reg_buffer_1227 ( .C (CLK), .D (new_AGEMA_signal_3994), .Q (new_AGEMA_signal_3995) ) ;
    buf_clk new_AGEMA_reg_buffer_1229 ( .C (CLK), .D (new_AGEMA_signal_3996), .Q (new_AGEMA_signal_3997) ) ;
    buf_clk new_AGEMA_reg_buffer_1231 ( .C (CLK), .D (new_AGEMA_signal_3998), .Q (new_AGEMA_signal_3999) ) ;
    buf_clk new_AGEMA_reg_buffer_1233 ( .C (CLK), .D (new_AGEMA_signal_4000), .Q (new_AGEMA_signal_4001) ) ;
    buf_clk new_AGEMA_reg_buffer_1235 ( .C (CLK), .D (new_AGEMA_signal_4002), .Q (new_AGEMA_signal_4003) ) ;
    buf_clk new_AGEMA_reg_buffer_1237 ( .C (CLK), .D (new_AGEMA_signal_4004), .Q (new_AGEMA_signal_4005) ) ;
    buf_clk new_AGEMA_reg_buffer_1239 ( .C (CLK), .D (new_AGEMA_signal_4006), .Q (new_AGEMA_signal_4007) ) ;
    buf_clk new_AGEMA_reg_buffer_1241 ( .C (CLK), .D (new_AGEMA_signal_4008), .Q (new_AGEMA_signal_4009) ) ;
    buf_clk new_AGEMA_reg_buffer_1243 ( .C (CLK), .D (new_AGEMA_signal_4010), .Q (new_AGEMA_signal_4011) ) ;
    buf_clk new_AGEMA_reg_buffer_1245 ( .C (CLK), .D (new_AGEMA_signal_4012), .Q (new_AGEMA_signal_4013) ) ;
    buf_clk new_AGEMA_reg_buffer_1247 ( .C (CLK), .D (new_AGEMA_signal_4014), .Q (new_AGEMA_signal_4015) ) ;
    buf_clk new_AGEMA_reg_buffer_1249 ( .C (CLK), .D (new_AGEMA_signal_4016), .Q (new_AGEMA_signal_4017) ) ;
    buf_clk new_AGEMA_reg_buffer_1251 ( .C (CLK), .D (new_AGEMA_signal_4018), .Q (new_AGEMA_signal_4019) ) ;
    buf_clk new_AGEMA_reg_buffer_1253 ( .C (CLK), .D (new_AGEMA_signal_4020), .Q (new_AGEMA_signal_4021) ) ;
    buf_clk new_AGEMA_reg_buffer_1255 ( .C (CLK), .D (new_AGEMA_signal_4022), .Q (new_AGEMA_signal_4023) ) ;
    buf_clk new_AGEMA_reg_buffer_1257 ( .C (CLK), .D (new_AGEMA_signal_4024), .Q (new_AGEMA_signal_4025) ) ;
    buf_clk new_AGEMA_reg_buffer_1259 ( .C (CLK), .D (new_AGEMA_signal_4026), .Q (new_AGEMA_signal_4027) ) ;
    buf_clk new_AGEMA_reg_buffer_1261 ( .C (CLK), .D (new_AGEMA_signal_4028), .Q (new_AGEMA_signal_4029) ) ;
    buf_clk new_AGEMA_reg_buffer_1263 ( .C (CLK), .D (new_AGEMA_signal_4030), .Q (new_AGEMA_signal_4031) ) ;
    buf_clk new_AGEMA_reg_buffer_1265 ( .C (CLK), .D (new_AGEMA_signal_4032), .Q (new_AGEMA_signal_4033) ) ;
    buf_clk new_AGEMA_reg_buffer_1267 ( .C (CLK), .D (new_AGEMA_signal_4034), .Q (new_AGEMA_signal_4035) ) ;
    buf_clk new_AGEMA_reg_buffer_1269 ( .C (CLK), .D (new_AGEMA_signal_4036), .Q (new_AGEMA_signal_4037) ) ;
    buf_clk new_AGEMA_reg_buffer_1271 ( .C (CLK), .D (new_AGEMA_signal_4038), .Q (new_AGEMA_signal_4039) ) ;
    buf_clk new_AGEMA_reg_buffer_1273 ( .C (CLK), .D (new_AGEMA_signal_4040), .Q (new_AGEMA_signal_4041) ) ;
    buf_clk new_AGEMA_reg_buffer_1275 ( .C (CLK), .D (new_AGEMA_signal_4042), .Q (new_AGEMA_signal_4043) ) ;
    buf_clk new_AGEMA_reg_buffer_1277 ( .C (CLK), .D (new_AGEMA_signal_4044), .Q (new_AGEMA_signal_4045) ) ;
    buf_clk new_AGEMA_reg_buffer_1279 ( .C (CLK), .D (new_AGEMA_signal_4046), .Q (new_AGEMA_signal_4047) ) ;
    buf_clk new_AGEMA_reg_buffer_1281 ( .C (CLK), .D (new_AGEMA_signal_4048), .Q (new_AGEMA_signal_4049) ) ;
    buf_clk new_AGEMA_reg_buffer_1283 ( .C (CLK), .D (new_AGEMA_signal_4050), .Q (new_AGEMA_signal_4051) ) ;
    buf_clk new_AGEMA_reg_buffer_1285 ( .C (CLK), .D (new_AGEMA_signal_4052), .Q (new_AGEMA_signal_4053) ) ;
    buf_clk new_AGEMA_reg_buffer_1287 ( .C (CLK), .D (new_AGEMA_signal_4054), .Q (new_AGEMA_signal_4055) ) ;
    buf_clk new_AGEMA_reg_buffer_1289 ( .C (CLK), .D (new_AGEMA_signal_4056), .Q (new_AGEMA_signal_4057) ) ;
    buf_clk new_AGEMA_reg_buffer_1291 ( .C (CLK), .D (new_AGEMA_signal_4058), .Q (new_AGEMA_signal_4059) ) ;
    buf_clk new_AGEMA_reg_buffer_1293 ( .C (CLK), .D (new_AGEMA_signal_4060), .Q (new_AGEMA_signal_4061) ) ;
    buf_clk new_AGEMA_reg_buffer_1295 ( .C (CLK), .D (new_AGEMA_signal_4062), .Q (new_AGEMA_signal_4063) ) ;
    buf_clk new_AGEMA_reg_buffer_1297 ( .C (CLK), .D (new_AGEMA_signal_4064), .Q (new_AGEMA_signal_4065) ) ;
    buf_clk new_AGEMA_reg_buffer_1299 ( .C (CLK), .D (new_AGEMA_signal_4066), .Q (new_AGEMA_signal_4067) ) ;
    buf_clk new_AGEMA_reg_buffer_1301 ( .C (CLK), .D (new_AGEMA_signal_4068), .Q (new_AGEMA_signal_4069) ) ;
    buf_clk new_AGEMA_reg_buffer_1303 ( .C (CLK), .D (new_AGEMA_signal_4070), .Q (new_AGEMA_signal_4071) ) ;
    buf_clk new_AGEMA_reg_buffer_1305 ( .C (CLK), .D (new_AGEMA_signal_4072), .Q (new_AGEMA_signal_4073) ) ;
    buf_clk new_AGEMA_reg_buffer_1307 ( .C (CLK), .D (new_AGEMA_signal_4074), .Q (new_AGEMA_signal_4075) ) ;
    buf_clk new_AGEMA_reg_buffer_1309 ( .C (CLK), .D (new_AGEMA_signal_4076), .Q (new_AGEMA_signal_4077) ) ;
    buf_clk new_AGEMA_reg_buffer_1311 ( .C (CLK), .D (new_AGEMA_signal_4078), .Q (new_AGEMA_signal_4079) ) ;
    buf_clk new_AGEMA_reg_buffer_1313 ( .C (CLK), .D (new_AGEMA_signal_4080), .Q (new_AGEMA_signal_4081) ) ;
    buf_clk new_AGEMA_reg_buffer_1315 ( .C (CLK), .D (new_AGEMA_signal_4082), .Q (new_AGEMA_signal_4083) ) ;
    buf_clk new_AGEMA_reg_buffer_1317 ( .C (CLK), .D (new_AGEMA_signal_4084), .Q (new_AGEMA_signal_4085) ) ;
    buf_clk new_AGEMA_reg_buffer_1319 ( .C (CLK), .D (new_AGEMA_signal_4086), .Q (new_AGEMA_signal_4087) ) ;
    buf_clk new_AGEMA_reg_buffer_1321 ( .C (CLK), .D (new_AGEMA_signal_4088), .Q (new_AGEMA_signal_4089) ) ;
    buf_clk new_AGEMA_reg_buffer_1323 ( .C (CLK), .D (new_AGEMA_signal_4090), .Q (new_AGEMA_signal_4091) ) ;
    buf_clk new_AGEMA_reg_buffer_1325 ( .C (CLK), .D (new_AGEMA_signal_4092), .Q (new_AGEMA_signal_4093) ) ;
    buf_clk new_AGEMA_reg_buffer_1327 ( .C (CLK), .D (new_AGEMA_signal_4094), .Q (new_AGEMA_signal_4095) ) ;
    buf_clk new_AGEMA_reg_buffer_1329 ( .C (CLK), .D (new_AGEMA_signal_4096), .Q (new_AGEMA_signal_4097) ) ;
    buf_clk new_AGEMA_reg_buffer_1331 ( .C (CLK), .D (new_AGEMA_signal_4098), .Q (new_AGEMA_signal_4099) ) ;
    buf_clk new_AGEMA_reg_buffer_1333 ( .C (CLK), .D (new_AGEMA_signal_4100), .Q (new_AGEMA_signal_4101) ) ;
    buf_clk new_AGEMA_reg_buffer_1335 ( .C (CLK), .D (new_AGEMA_signal_4102), .Q (new_AGEMA_signal_4103) ) ;
    buf_clk new_AGEMA_reg_buffer_1337 ( .C (CLK), .D (new_AGEMA_signal_4104), .Q (new_AGEMA_signal_4105) ) ;
    buf_clk new_AGEMA_reg_buffer_1339 ( .C (CLK), .D (new_AGEMA_signal_4106), .Q (new_AGEMA_signal_4107) ) ;
    buf_clk new_AGEMA_reg_buffer_1341 ( .C (CLK), .D (new_AGEMA_signal_4108), .Q (new_AGEMA_signal_4109) ) ;
    buf_clk new_AGEMA_reg_buffer_1343 ( .C (CLK), .D (new_AGEMA_signal_4110), .Q (new_AGEMA_signal_4111) ) ;
    buf_clk new_AGEMA_reg_buffer_1345 ( .C (CLK), .D (new_AGEMA_signal_4112), .Q (new_AGEMA_signal_4113) ) ;
    buf_clk new_AGEMA_reg_buffer_1347 ( .C (CLK), .D (new_AGEMA_signal_4114), .Q (new_AGEMA_signal_4115) ) ;
    buf_clk new_AGEMA_reg_buffer_1349 ( .C (CLK), .D (new_AGEMA_signal_4116), .Q (new_AGEMA_signal_4117) ) ;
    buf_clk new_AGEMA_reg_buffer_1351 ( .C (CLK), .D (new_AGEMA_signal_4118), .Q (new_AGEMA_signal_4119) ) ;
    buf_clk new_AGEMA_reg_buffer_1353 ( .C (CLK), .D (new_AGEMA_signal_4120), .Q (new_AGEMA_signal_4121) ) ;
    buf_clk new_AGEMA_reg_buffer_1355 ( .C (CLK), .D (new_AGEMA_signal_4122), .Q (new_AGEMA_signal_4123) ) ;
    buf_clk new_AGEMA_reg_buffer_1357 ( .C (CLK), .D (new_AGEMA_signal_4124), .Q (new_AGEMA_signal_4125) ) ;
    buf_clk new_AGEMA_reg_buffer_1359 ( .C (CLK), .D (new_AGEMA_signal_4126), .Q (new_AGEMA_signal_4127) ) ;
    buf_clk new_AGEMA_reg_buffer_1361 ( .C (CLK), .D (new_AGEMA_signal_4128), .Q (new_AGEMA_signal_4129) ) ;
    buf_clk new_AGEMA_reg_buffer_1363 ( .C (CLK), .D (new_AGEMA_signal_4130), .Q (new_AGEMA_signal_4131) ) ;
    buf_clk new_AGEMA_reg_buffer_1365 ( .C (CLK), .D (new_AGEMA_signal_4132), .Q (new_AGEMA_signal_4133) ) ;
    buf_clk new_AGEMA_reg_buffer_1367 ( .C (CLK), .D (new_AGEMA_signal_4134), .Q (new_AGEMA_signal_4135) ) ;
    buf_clk new_AGEMA_reg_buffer_1369 ( .C (CLK), .D (new_AGEMA_signal_4136), .Q (new_AGEMA_signal_4137) ) ;
    buf_clk new_AGEMA_reg_buffer_1371 ( .C (CLK), .D (new_AGEMA_signal_4138), .Q (new_AGEMA_signal_4139) ) ;
    buf_clk new_AGEMA_reg_buffer_1373 ( .C (CLK), .D (new_AGEMA_signal_4140), .Q (new_AGEMA_signal_4141) ) ;
    buf_clk new_AGEMA_reg_buffer_1375 ( .C (CLK), .D (new_AGEMA_signal_4142), .Q (new_AGEMA_signal_4143) ) ;
    buf_clk new_AGEMA_reg_buffer_1377 ( .C (CLK), .D (new_AGEMA_signal_4144), .Q (new_AGEMA_signal_4145) ) ;
    buf_clk new_AGEMA_reg_buffer_1379 ( .C (CLK), .D (new_AGEMA_signal_4146), .Q (new_AGEMA_signal_4147) ) ;
    buf_clk new_AGEMA_reg_buffer_1381 ( .C (CLK), .D (new_AGEMA_signal_4148), .Q (new_AGEMA_signal_4149) ) ;
    buf_clk new_AGEMA_reg_buffer_1383 ( .C (CLK), .D (new_AGEMA_signal_4150), .Q (new_AGEMA_signal_4151) ) ;
    buf_clk new_AGEMA_reg_buffer_1385 ( .C (CLK), .D (new_AGEMA_signal_4152), .Q (new_AGEMA_signal_4153) ) ;
    buf_clk new_AGEMA_reg_buffer_1387 ( .C (CLK), .D (new_AGEMA_signal_4154), .Q (new_AGEMA_signal_4155) ) ;
    buf_clk new_AGEMA_reg_buffer_1389 ( .C (CLK), .D (new_AGEMA_signal_4156), .Q (new_AGEMA_signal_4157) ) ;
    buf_clk new_AGEMA_reg_buffer_1391 ( .C (CLK), .D (new_AGEMA_signal_4158), .Q (new_AGEMA_signal_4159) ) ;
    buf_clk new_AGEMA_reg_buffer_1393 ( .C (CLK), .D (new_AGEMA_signal_4160), .Q (new_AGEMA_signal_4161) ) ;
    buf_clk new_AGEMA_reg_buffer_1395 ( .C (CLK), .D (new_AGEMA_signal_4162), .Q (new_AGEMA_signal_4163) ) ;
    buf_clk new_AGEMA_reg_buffer_1397 ( .C (CLK), .D (new_AGEMA_signal_4164), .Q (new_AGEMA_signal_4165) ) ;
    buf_clk new_AGEMA_reg_buffer_1399 ( .C (CLK), .D (new_AGEMA_signal_4166), .Q (new_AGEMA_signal_4167) ) ;
    buf_clk new_AGEMA_reg_buffer_1401 ( .C (CLK), .D (new_AGEMA_signal_4168), .Q (new_AGEMA_signal_4169) ) ;
    buf_clk new_AGEMA_reg_buffer_1403 ( .C (CLK), .D (new_AGEMA_signal_4170), .Q (new_AGEMA_signal_4171) ) ;
    buf_clk new_AGEMA_reg_buffer_1405 ( .C (CLK), .D (new_AGEMA_signal_4172), .Q (new_AGEMA_signal_4173) ) ;
    buf_clk new_AGEMA_reg_buffer_1407 ( .C (CLK), .D (new_AGEMA_signal_4174), .Q (new_AGEMA_signal_4175) ) ;
    buf_clk new_AGEMA_reg_buffer_1409 ( .C (CLK), .D (new_AGEMA_signal_4176), .Q (new_AGEMA_signal_4177) ) ;
    buf_clk new_AGEMA_reg_buffer_1411 ( .C (CLK), .D (new_AGEMA_signal_4178), .Q (new_AGEMA_signal_4179) ) ;
    buf_clk new_AGEMA_reg_buffer_1413 ( .C (CLK), .D (new_AGEMA_signal_4180), .Q (new_AGEMA_signal_4181) ) ;
    buf_clk new_AGEMA_reg_buffer_1415 ( .C (CLK), .D (new_AGEMA_signal_4182), .Q (new_AGEMA_signal_4183) ) ;
    buf_clk new_AGEMA_reg_buffer_1417 ( .C (CLK), .D (new_AGEMA_signal_4184), .Q (new_AGEMA_signal_4185) ) ;
    buf_clk new_AGEMA_reg_buffer_1421 ( .C (CLK), .D (new_AGEMA_signal_4188), .Q (new_AGEMA_signal_4189) ) ;
    buf_clk new_AGEMA_reg_buffer_1425 ( .C (CLK), .D (new_AGEMA_signal_4192), .Q (new_AGEMA_signal_4193) ) ;
    buf_clk new_AGEMA_reg_buffer_1429 ( .C (CLK), .D (new_AGEMA_signal_4196), .Q (new_AGEMA_signal_4197) ) ;
    buf_clk new_AGEMA_reg_buffer_1433 ( .C (CLK), .D (new_AGEMA_signal_4200), .Q (new_AGEMA_signal_4201) ) ;
    buf_clk new_AGEMA_reg_buffer_1437 ( .C (CLK), .D (new_AGEMA_signal_4204), .Q (new_AGEMA_signal_4205) ) ;
    buf_clk new_AGEMA_reg_buffer_1441 ( .C (CLK), .D (new_AGEMA_signal_4208), .Q (new_AGEMA_signal_4209) ) ;
    buf_clk new_AGEMA_reg_buffer_1445 ( .C (CLK), .D (new_AGEMA_signal_4212), .Q (new_AGEMA_signal_4213) ) ;
    buf_clk new_AGEMA_reg_buffer_1449 ( .C (CLK), .D (new_AGEMA_signal_4216), .Q (new_AGEMA_signal_4217) ) ;
    buf_clk new_AGEMA_reg_buffer_1453 ( .C (CLK), .D (new_AGEMA_signal_4220), .Q (new_AGEMA_signal_4221) ) ;
    buf_clk new_AGEMA_reg_buffer_1457 ( .C (CLK), .D (new_AGEMA_signal_4224), .Q (new_AGEMA_signal_4225) ) ;
    buf_clk new_AGEMA_reg_buffer_1461 ( .C (CLK), .D (new_AGEMA_signal_4228), .Q (new_AGEMA_signal_4229) ) ;
    buf_clk new_AGEMA_reg_buffer_1465 ( .C (CLK), .D (new_AGEMA_signal_4232), .Q (new_AGEMA_signal_4233) ) ;
    buf_clk new_AGEMA_reg_buffer_1469 ( .C (CLK), .D (new_AGEMA_signal_4236), .Q (new_AGEMA_signal_4237) ) ;
    buf_clk new_AGEMA_reg_buffer_1473 ( .C (CLK), .D (new_AGEMA_signal_4240), .Q (new_AGEMA_signal_4241) ) ;
    buf_clk new_AGEMA_reg_buffer_1477 ( .C (CLK), .D (new_AGEMA_signal_4244), .Q (new_AGEMA_signal_4245) ) ;
    buf_clk new_AGEMA_reg_buffer_1481 ( .C (CLK), .D (new_AGEMA_signal_4248), .Q (new_AGEMA_signal_4249) ) ;
    buf_clk new_AGEMA_reg_buffer_1485 ( .C (CLK), .D (new_AGEMA_signal_4252), .Q (new_AGEMA_signal_4253) ) ;
    buf_clk new_AGEMA_reg_buffer_1489 ( .C (CLK), .D (new_AGEMA_signal_4256), .Q (new_AGEMA_signal_4257) ) ;
    buf_clk new_AGEMA_reg_buffer_1493 ( .C (CLK), .D (new_AGEMA_signal_4260), .Q (new_AGEMA_signal_4261) ) ;
    buf_clk new_AGEMA_reg_buffer_1497 ( .C (CLK), .D (new_AGEMA_signal_4264), .Q (new_AGEMA_signal_4265) ) ;
    buf_clk new_AGEMA_reg_buffer_1501 ( .C (CLK), .D (new_AGEMA_signal_4268), .Q (new_AGEMA_signal_4269) ) ;
    buf_clk new_AGEMA_reg_buffer_1505 ( .C (CLK), .D (new_AGEMA_signal_4272), .Q (new_AGEMA_signal_4273) ) ;
    buf_clk new_AGEMA_reg_buffer_1509 ( .C (CLK), .D (new_AGEMA_signal_4276), .Q (new_AGEMA_signal_4277) ) ;
    buf_clk new_AGEMA_reg_buffer_1513 ( .C (CLK), .D (new_AGEMA_signal_4280), .Q (new_AGEMA_signal_4281) ) ;
    buf_clk new_AGEMA_reg_buffer_1517 ( .C (CLK), .D (new_AGEMA_signal_4284), .Q (new_AGEMA_signal_4285) ) ;
    buf_clk new_AGEMA_reg_buffer_1521 ( .C (CLK), .D (new_AGEMA_signal_4288), .Q (new_AGEMA_signal_4289) ) ;
    buf_clk new_AGEMA_reg_buffer_1525 ( .C (CLK), .D (new_AGEMA_signal_4292), .Q (new_AGEMA_signal_4293) ) ;
    buf_clk new_AGEMA_reg_buffer_1529 ( .C (CLK), .D (new_AGEMA_signal_4296), .Q (new_AGEMA_signal_4297) ) ;
    buf_clk new_AGEMA_reg_buffer_1533 ( .C (CLK), .D (new_AGEMA_signal_4300), .Q (new_AGEMA_signal_4301) ) ;
    buf_clk new_AGEMA_reg_buffer_1537 ( .C (CLK), .D (new_AGEMA_signal_4304), .Q (new_AGEMA_signal_4305) ) ;
    buf_clk new_AGEMA_reg_buffer_1541 ( .C (CLK), .D (new_AGEMA_signal_4308), .Q (new_AGEMA_signal_4309) ) ;
    buf_clk new_AGEMA_reg_buffer_1545 ( .C (CLK), .D (new_AGEMA_signal_4312), .Q (new_AGEMA_signal_4313) ) ;
    buf_clk new_AGEMA_reg_buffer_1549 ( .C (CLK), .D (new_AGEMA_signal_4316), .Q (new_AGEMA_signal_4317) ) ;
    buf_clk new_AGEMA_reg_buffer_1553 ( .C (CLK), .D (new_AGEMA_signal_4320), .Q (new_AGEMA_signal_4321) ) ;
    buf_clk new_AGEMA_reg_buffer_1557 ( .C (CLK), .D (new_AGEMA_signal_4324), .Q (new_AGEMA_signal_4325) ) ;
    buf_clk new_AGEMA_reg_buffer_1561 ( .C (CLK), .D (new_AGEMA_signal_4328), .Q (new_AGEMA_signal_4329) ) ;
    buf_clk new_AGEMA_reg_buffer_1565 ( .C (CLK), .D (new_AGEMA_signal_4332), .Q (new_AGEMA_signal_4333) ) ;
    buf_clk new_AGEMA_reg_buffer_1569 ( .C (CLK), .D (new_AGEMA_signal_4336), .Q (new_AGEMA_signal_4337) ) ;
    buf_clk new_AGEMA_reg_buffer_1573 ( .C (CLK), .D (new_AGEMA_signal_4340), .Q (new_AGEMA_signal_4341) ) ;
    buf_clk new_AGEMA_reg_buffer_1577 ( .C (CLK), .D (new_AGEMA_signal_4344), .Q (new_AGEMA_signal_4345) ) ;
    buf_clk new_AGEMA_reg_buffer_1581 ( .C (CLK), .D (new_AGEMA_signal_4348), .Q (new_AGEMA_signal_4349) ) ;
    buf_clk new_AGEMA_reg_buffer_1585 ( .C (CLK), .D (new_AGEMA_signal_4352), .Q (new_AGEMA_signal_4353) ) ;
    buf_clk new_AGEMA_reg_buffer_1589 ( .C (CLK), .D (new_AGEMA_signal_4356), .Q (new_AGEMA_signal_4357) ) ;
    buf_clk new_AGEMA_reg_buffer_1593 ( .C (CLK), .D (new_AGEMA_signal_4360), .Q (new_AGEMA_signal_4361) ) ;
    buf_clk new_AGEMA_reg_buffer_1597 ( .C (CLK), .D (new_AGEMA_signal_4364), .Q (new_AGEMA_signal_4365) ) ;
    buf_clk new_AGEMA_reg_buffer_1601 ( .C (CLK), .D (new_AGEMA_signal_4368), .Q (new_AGEMA_signal_4369) ) ;
    buf_clk new_AGEMA_reg_buffer_1605 ( .C (CLK), .D (new_AGEMA_signal_4372), .Q (new_AGEMA_signal_4373) ) ;
    buf_clk new_AGEMA_reg_buffer_1609 ( .C (CLK), .D (new_AGEMA_signal_4376), .Q (new_AGEMA_signal_4377) ) ;
    buf_clk new_AGEMA_reg_buffer_1613 ( .C (CLK), .D (new_AGEMA_signal_4380), .Q (new_AGEMA_signal_4381) ) ;
    buf_clk new_AGEMA_reg_buffer_1617 ( .C (CLK), .D (new_AGEMA_signal_4384), .Q (new_AGEMA_signal_4385) ) ;
    buf_clk new_AGEMA_reg_buffer_1621 ( .C (CLK), .D (new_AGEMA_signal_4388), .Q (new_AGEMA_signal_4389) ) ;
    buf_clk new_AGEMA_reg_buffer_1625 ( .C (CLK), .D (new_AGEMA_signal_4392), .Q (new_AGEMA_signal_4393) ) ;
    buf_clk new_AGEMA_reg_buffer_1629 ( .C (CLK), .D (new_AGEMA_signal_4396), .Q (new_AGEMA_signal_4397) ) ;
    buf_clk new_AGEMA_reg_buffer_1633 ( .C (CLK), .D (new_AGEMA_signal_4400), .Q (new_AGEMA_signal_4401) ) ;
    buf_clk new_AGEMA_reg_buffer_1637 ( .C (CLK), .D (new_AGEMA_signal_4404), .Q (new_AGEMA_signal_4405) ) ;
    buf_clk new_AGEMA_reg_buffer_1641 ( .C (CLK), .D (new_AGEMA_signal_4408), .Q (new_AGEMA_signal_4409) ) ;
    buf_clk new_AGEMA_reg_buffer_1645 ( .C (CLK), .D (new_AGEMA_signal_4412), .Q (new_AGEMA_signal_4413) ) ;
    buf_clk new_AGEMA_reg_buffer_1649 ( .C (CLK), .D (new_AGEMA_signal_4416), .Q (new_AGEMA_signal_4417) ) ;
    buf_clk new_AGEMA_reg_buffer_1653 ( .C (CLK), .D (new_AGEMA_signal_4420), .Q (new_AGEMA_signal_4421) ) ;
    buf_clk new_AGEMA_reg_buffer_1657 ( .C (CLK), .D (new_AGEMA_signal_4424), .Q (new_AGEMA_signal_4425) ) ;
    buf_clk new_AGEMA_reg_buffer_1661 ( .C (CLK), .D (new_AGEMA_signal_4428), .Q (new_AGEMA_signal_4429) ) ;
    buf_clk new_AGEMA_reg_buffer_1665 ( .C (CLK), .D (new_AGEMA_signal_4432), .Q (new_AGEMA_signal_4433) ) ;
    buf_clk new_AGEMA_reg_buffer_1669 ( .C (CLK), .D (new_AGEMA_signal_4436), .Q (new_AGEMA_signal_4437) ) ;
    buf_clk new_AGEMA_reg_buffer_1673 ( .C (CLK), .D (new_AGEMA_signal_4440), .Q (new_AGEMA_signal_4441) ) ;
    buf_clk new_AGEMA_reg_buffer_1677 ( .C (CLK), .D (new_AGEMA_signal_4444), .Q (new_AGEMA_signal_4445) ) ;
    buf_clk new_AGEMA_reg_buffer_1681 ( .C (CLK), .D (new_AGEMA_signal_4448), .Q (new_AGEMA_signal_4449) ) ;
    buf_clk new_AGEMA_reg_buffer_1685 ( .C (CLK), .D (new_AGEMA_signal_4452), .Q (new_AGEMA_signal_4453) ) ;
    buf_clk new_AGEMA_reg_buffer_1689 ( .C (CLK), .D (new_AGEMA_signal_4456), .Q (new_AGEMA_signal_4457) ) ;
    buf_clk new_AGEMA_reg_buffer_1693 ( .C (CLK), .D (new_AGEMA_signal_4460), .Q (new_AGEMA_signal_4461) ) ;
    buf_clk new_AGEMA_reg_buffer_1697 ( .C (CLK), .D (new_AGEMA_signal_4464), .Q (new_AGEMA_signal_4465) ) ;
    buf_clk new_AGEMA_reg_buffer_1701 ( .C (CLK), .D (new_AGEMA_signal_4468), .Q (new_AGEMA_signal_4469) ) ;
    buf_clk new_AGEMA_reg_buffer_1705 ( .C (CLK), .D (new_AGEMA_signal_4472), .Q (new_AGEMA_signal_4473) ) ;
    buf_clk new_AGEMA_reg_buffer_1709 ( .C (CLK), .D (new_AGEMA_signal_4476), .Q (new_AGEMA_signal_4477) ) ;
    buf_clk new_AGEMA_reg_buffer_1713 ( .C (CLK), .D (new_AGEMA_signal_4480), .Q (new_AGEMA_signal_4481) ) ;
    buf_clk new_AGEMA_reg_buffer_1717 ( .C (CLK), .D (new_AGEMA_signal_4484), .Q (new_AGEMA_signal_4485) ) ;
    buf_clk new_AGEMA_reg_buffer_1721 ( .C (CLK), .D (new_AGEMA_signal_4488), .Q (new_AGEMA_signal_4489) ) ;
    buf_clk new_AGEMA_reg_buffer_1725 ( .C (CLK), .D (new_AGEMA_signal_4492), .Q (new_AGEMA_signal_4493) ) ;
    buf_clk new_AGEMA_reg_buffer_1729 ( .C (CLK), .D (new_AGEMA_signal_4496), .Q (new_AGEMA_signal_4497) ) ;
    buf_clk new_AGEMA_reg_buffer_1733 ( .C (CLK), .D (new_AGEMA_signal_4500), .Q (new_AGEMA_signal_4501) ) ;
    buf_clk new_AGEMA_reg_buffer_1737 ( .C (CLK), .D (new_AGEMA_signal_4504), .Q (new_AGEMA_signal_4505) ) ;
    buf_clk new_AGEMA_reg_buffer_1741 ( .C (CLK), .D (new_AGEMA_signal_4508), .Q (new_AGEMA_signal_4509) ) ;
    buf_clk new_AGEMA_reg_buffer_1745 ( .C (CLK), .D (new_AGEMA_signal_4512), .Q (new_AGEMA_signal_4513) ) ;
    buf_clk new_AGEMA_reg_buffer_1749 ( .C (CLK), .D (new_AGEMA_signal_4516), .Q (new_AGEMA_signal_4517) ) ;
    buf_clk new_AGEMA_reg_buffer_1753 ( .C (CLK), .D (new_AGEMA_signal_4520), .Q (new_AGEMA_signal_4521) ) ;
    buf_clk new_AGEMA_reg_buffer_1757 ( .C (CLK), .D (new_AGEMA_signal_4524), .Q (new_AGEMA_signal_4525) ) ;
    buf_clk new_AGEMA_reg_buffer_1761 ( .C (CLK), .D (new_AGEMA_signal_4528), .Q (new_AGEMA_signal_4529) ) ;
    buf_clk new_AGEMA_reg_buffer_1765 ( .C (CLK), .D (new_AGEMA_signal_4532), .Q (new_AGEMA_signal_4533) ) ;
    buf_clk new_AGEMA_reg_buffer_1769 ( .C (CLK), .D (new_AGEMA_signal_4536), .Q (new_AGEMA_signal_4537) ) ;
    buf_clk new_AGEMA_reg_buffer_1773 ( .C (CLK), .D (new_AGEMA_signal_4540), .Q (new_AGEMA_signal_4541) ) ;
    buf_clk new_AGEMA_reg_buffer_1777 ( .C (CLK), .D (new_AGEMA_signal_4544), .Q (new_AGEMA_signal_4545) ) ;
    buf_clk new_AGEMA_reg_buffer_1781 ( .C (CLK), .D (new_AGEMA_signal_4548), .Q (new_AGEMA_signal_4549) ) ;
    buf_clk new_AGEMA_reg_buffer_1785 ( .C (CLK), .D (new_AGEMA_signal_4552), .Q (new_AGEMA_signal_4553) ) ;
    buf_clk new_AGEMA_reg_buffer_1789 ( .C (CLK), .D (new_AGEMA_signal_4556), .Q (new_AGEMA_signal_4557) ) ;
    buf_clk new_AGEMA_reg_buffer_1793 ( .C (CLK), .D (new_AGEMA_signal_4560), .Q (new_AGEMA_signal_4561) ) ;
    buf_clk new_AGEMA_reg_buffer_1797 ( .C (CLK), .D (new_AGEMA_signal_4564), .Q (new_AGEMA_signal_4565) ) ;
    buf_clk new_AGEMA_reg_buffer_1801 ( .C (CLK), .D (new_AGEMA_signal_4568), .Q (new_AGEMA_signal_4569) ) ;
    buf_clk new_AGEMA_reg_buffer_1805 ( .C (CLK), .D (new_AGEMA_signal_4572), .Q (new_AGEMA_signal_4573) ) ;
    buf_clk new_AGEMA_reg_buffer_1809 ( .C (CLK), .D (new_AGEMA_signal_4576), .Q (new_AGEMA_signal_4577) ) ;
    buf_clk new_AGEMA_reg_buffer_1813 ( .C (CLK), .D (new_AGEMA_signal_4580), .Q (new_AGEMA_signal_4581) ) ;
    buf_clk new_AGEMA_reg_buffer_1817 ( .C (CLK), .D (new_AGEMA_signal_4584), .Q (new_AGEMA_signal_4585) ) ;
    buf_clk new_AGEMA_reg_buffer_1821 ( .C (CLK), .D (new_AGEMA_signal_4588), .Q (new_AGEMA_signal_4589) ) ;
    buf_clk new_AGEMA_reg_buffer_1825 ( .C (CLK), .D (new_AGEMA_signal_4592), .Q (new_AGEMA_signal_4593) ) ;
    buf_clk new_AGEMA_reg_buffer_1829 ( .C (CLK), .D (new_AGEMA_signal_4596), .Q (new_AGEMA_signal_4597) ) ;
    buf_clk new_AGEMA_reg_buffer_1833 ( .C (CLK), .D (new_AGEMA_signal_4600), .Q (new_AGEMA_signal_4601) ) ;
    buf_clk new_AGEMA_reg_buffer_1837 ( .C (CLK), .D (new_AGEMA_signal_4604), .Q (new_AGEMA_signal_4605) ) ;
    buf_clk new_AGEMA_reg_buffer_1841 ( .C (CLK), .D (new_AGEMA_signal_4608), .Q (new_AGEMA_signal_4609) ) ;
    buf_clk new_AGEMA_reg_buffer_1845 ( .C (CLK), .D (new_AGEMA_signal_4612), .Q (new_AGEMA_signal_4613) ) ;
    buf_clk new_AGEMA_reg_buffer_1849 ( .C (CLK), .D (new_AGEMA_signal_4616), .Q (new_AGEMA_signal_4617) ) ;
    buf_clk new_AGEMA_reg_buffer_1853 ( .C (CLK), .D (new_AGEMA_signal_4620), .Q (new_AGEMA_signal_4621) ) ;
    buf_clk new_AGEMA_reg_buffer_1857 ( .C (CLK), .D (new_AGEMA_signal_4624), .Q (new_AGEMA_signal_4625) ) ;
    buf_clk new_AGEMA_reg_buffer_1861 ( .C (CLK), .D (new_AGEMA_signal_4628), .Q (new_AGEMA_signal_4629) ) ;
    buf_clk new_AGEMA_reg_buffer_1865 ( .C (CLK), .D (new_AGEMA_signal_4632), .Q (new_AGEMA_signal_4633) ) ;
    buf_clk new_AGEMA_reg_buffer_1869 ( .C (CLK), .D (new_AGEMA_signal_4636), .Q (new_AGEMA_signal_4637) ) ;
    buf_clk new_AGEMA_reg_buffer_1873 ( .C (CLK), .D (new_AGEMA_signal_4640), .Q (new_AGEMA_signal_4641) ) ;
    buf_clk new_AGEMA_reg_buffer_1877 ( .C (CLK), .D (new_AGEMA_signal_4644), .Q (new_AGEMA_signal_4645) ) ;
    buf_clk new_AGEMA_reg_buffer_1881 ( .C (CLK), .D (new_AGEMA_signal_4648), .Q (new_AGEMA_signal_4649) ) ;
    buf_clk new_AGEMA_reg_buffer_1885 ( .C (CLK), .D (new_AGEMA_signal_4652), .Q (new_AGEMA_signal_4653) ) ;
    buf_clk new_AGEMA_reg_buffer_1889 ( .C (CLK), .D (new_AGEMA_signal_4656), .Q (new_AGEMA_signal_4657) ) ;
    buf_clk new_AGEMA_reg_buffer_1893 ( .C (CLK), .D (new_AGEMA_signal_4660), .Q (new_AGEMA_signal_4661) ) ;
    buf_clk new_AGEMA_reg_buffer_1897 ( .C (CLK), .D (new_AGEMA_signal_4664), .Q (new_AGEMA_signal_4665) ) ;
    buf_clk new_AGEMA_reg_buffer_1901 ( .C (CLK), .D (new_AGEMA_signal_4668), .Q (new_AGEMA_signal_4669) ) ;
    buf_clk new_AGEMA_reg_buffer_1905 ( .C (CLK), .D (new_AGEMA_signal_4672), .Q (new_AGEMA_signal_4673) ) ;
    buf_clk new_AGEMA_reg_buffer_1909 ( .C (CLK), .D (new_AGEMA_signal_4676), .Q (new_AGEMA_signal_4677) ) ;
    buf_clk new_AGEMA_reg_buffer_1913 ( .C (CLK), .D (new_AGEMA_signal_4680), .Q (new_AGEMA_signal_4681) ) ;
    buf_clk new_AGEMA_reg_buffer_1917 ( .C (CLK), .D (new_AGEMA_signal_4684), .Q (new_AGEMA_signal_4685) ) ;
    buf_clk new_AGEMA_reg_buffer_1921 ( .C (CLK), .D (new_AGEMA_signal_4688), .Q (new_AGEMA_signal_4689) ) ;
    buf_clk new_AGEMA_reg_buffer_1925 ( .C (CLK), .D (new_AGEMA_signal_4692), .Q (new_AGEMA_signal_4693) ) ;
    buf_clk new_AGEMA_reg_buffer_1929 ( .C (CLK), .D (new_AGEMA_signal_4696), .Q (new_AGEMA_signal_4697) ) ;
    buf_clk new_AGEMA_reg_buffer_1933 ( .C (CLK), .D (new_AGEMA_signal_4700), .Q (new_AGEMA_signal_4701) ) ;
    buf_clk new_AGEMA_reg_buffer_1937 ( .C (CLK), .D (new_AGEMA_signal_4704), .Q (new_AGEMA_signal_4705) ) ;
    buf_clk new_AGEMA_reg_buffer_1941 ( .C (CLK), .D (new_AGEMA_signal_4708), .Q (new_AGEMA_signal_4709) ) ;
    buf_clk new_AGEMA_reg_buffer_1945 ( .C (CLK), .D (new_AGEMA_signal_4712), .Q (new_AGEMA_signal_4713) ) ;
    buf_clk new_AGEMA_reg_buffer_1949 ( .C (CLK), .D (new_AGEMA_signal_4716), .Q (new_AGEMA_signal_4717) ) ;
    buf_clk new_AGEMA_reg_buffer_1953 ( .C (CLK), .D (new_AGEMA_signal_4720), .Q (new_AGEMA_signal_4721) ) ;
    buf_clk new_AGEMA_reg_buffer_1957 ( .C (CLK), .D (new_AGEMA_signal_4724), .Q (new_AGEMA_signal_4725) ) ;
    buf_clk new_AGEMA_reg_buffer_1961 ( .C (CLK), .D (new_AGEMA_signal_4728), .Q (new_AGEMA_signal_4729) ) ;
    buf_clk new_AGEMA_reg_buffer_1965 ( .C (CLK), .D (new_AGEMA_signal_4732), .Q (new_AGEMA_signal_4733) ) ;
    buf_clk new_AGEMA_reg_buffer_1969 ( .C (CLK), .D (new_AGEMA_signal_4736), .Q (new_AGEMA_signal_4737) ) ;
    buf_clk new_AGEMA_reg_buffer_1973 ( .C (CLK), .D (new_AGEMA_signal_4740), .Q (new_AGEMA_signal_4741) ) ;
    buf_clk new_AGEMA_reg_buffer_1977 ( .C (CLK), .D (new_AGEMA_signal_4744), .Q (new_AGEMA_signal_4745) ) ;
    buf_clk new_AGEMA_reg_buffer_1981 ( .C (CLK), .D (new_AGEMA_signal_4748), .Q (new_AGEMA_signal_4749) ) ;
    buf_clk new_AGEMA_reg_buffer_1985 ( .C (CLK), .D (new_AGEMA_signal_4752), .Q (new_AGEMA_signal_4753) ) ;
    buf_clk new_AGEMA_reg_buffer_1989 ( .C (CLK), .D (new_AGEMA_signal_4756), .Q (new_AGEMA_signal_4757) ) ;
    buf_clk new_AGEMA_reg_buffer_1993 ( .C (CLK), .D (new_AGEMA_signal_4760), .Q (new_AGEMA_signal_4761) ) ;
    buf_clk new_AGEMA_reg_buffer_1997 ( .C (CLK), .D (new_AGEMA_signal_4764), .Q (new_AGEMA_signal_4765) ) ;
    buf_clk new_AGEMA_reg_buffer_2001 ( .C (CLK), .D (new_AGEMA_signal_4768), .Q (new_AGEMA_signal_4769) ) ;
    buf_clk new_AGEMA_reg_buffer_2005 ( .C (CLK), .D (new_AGEMA_signal_4772), .Q (new_AGEMA_signal_4773) ) ;
    buf_clk new_AGEMA_reg_buffer_2009 ( .C (CLK), .D (new_AGEMA_signal_4776), .Q (new_AGEMA_signal_4777) ) ;
    buf_clk new_AGEMA_reg_buffer_2013 ( .C (CLK), .D (new_AGEMA_signal_4780), .Q (new_AGEMA_signal_4781) ) ;
    buf_clk new_AGEMA_reg_buffer_2017 ( .C (CLK), .D (new_AGEMA_signal_4784), .Q (new_AGEMA_signal_4785) ) ;
    buf_clk new_AGEMA_reg_buffer_2021 ( .C (CLK), .D (new_AGEMA_signal_4788), .Q (new_AGEMA_signal_4789) ) ;
    buf_clk new_AGEMA_reg_buffer_2025 ( .C (CLK), .D (new_AGEMA_signal_4792), .Q (new_AGEMA_signal_4793) ) ;
    buf_clk new_AGEMA_reg_buffer_2029 ( .C (CLK), .D (new_AGEMA_signal_4796), .Q (new_AGEMA_signal_4797) ) ;
    buf_clk new_AGEMA_reg_buffer_2033 ( .C (CLK), .D (new_AGEMA_signal_4800), .Q (new_AGEMA_signal_4801) ) ;
    buf_clk new_AGEMA_reg_buffer_2037 ( .C (CLK), .D (new_AGEMA_signal_4804), .Q (new_AGEMA_signal_4805) ) ;
    buf_clk new_AGEMA_reg_buffer_2041 ( .C (CLK), .D (new_AGEMA_signal_4808), .Q (new_AGEMA_signal_4809) ) ;
    buf_clk new_AGEMA_reg_buffer_2045 ( .C (CLK), .D (new_AGEMA_signal_4812), .Q (new_AGEMA_signal_4813) ) ;
    buf_clk new_AGEMA_reg_buffer_2049 ( .C (CLK), .D (new_AGEMA_signal_4816), .Q (new_AGEMA_signal_4817) ) ;
    buf_clk new_AGEMA_reg_buffer_2053 ( .C (CLK), .D (new_AGEMA_signal_4820), .Q (new_AGEMA_signal_4821) ) ;
    buf_clk new_AGEMA_reg_buffer_2057 ( .C (CLK), .D (new_AGEMA_signal_4824), .Q (new_AGEMA_signal_4825) ) ;
    buf_clk new_AGEMA_reg_buffer_2061 ( .C (CLK), .D (new_AGEMA_signal_4828), .Q (new_AGEMA_signal_4829) ) ;
    buf_clk new_AGEMA_reg_buffer_2065 ( .C (CLK), .D (new_AGEMA_signal_4832), .Q (new_AGEMA_signal_4833) ) ;
    buf_clk new_AGEMA_reg_buffer_2069 ( .C (CLK), .D (new_AGEMA_signal_4836), .Q (new_AGEMA_signal_4837) ) ;
    buf_clk new_AGEMA_reg_buffer_2073 ( .C (CLK), .D (new_AGEMA_signal_4840), .Q (new_AGEMA_signal_4841) ) ;
    buf_clk new_AGEMA_reg_buffer_2077 ( .C (CLK), .D (new_AGEMA_signal_4844), .Q (new_AGEMA_signal_4845) ) ;
    buf_clk new_AGEMA_reg_buffer_2081 ( .C (CLK), .D (new_AGEMA_signal_4848), .Q (new_AGEMA_signal_4849) ) ;
    buf_clk new_AGEMA_reg_buffer_2085 ( .C (CLK), .D (new_AGEMA_signal_4852), .Q (new_AGEMA_signal_4853) ) ;
    buf_clk new_AGEMA_reg_buffer_2089 ( .C (CLK), .D (new_AGEMA_signal_4856), .Q (new_AGEMA_signal_4857) ) ;
    buf_clk new_AGEMA_reg_buffer_2093 ( .C (CLK), .D (new_AGEMA_signal_4860), .Q (new_AGEMA_signal_4861) ) ;
    buf_clk new_AGEMA_reg_buffer_2097 ( .C (CLK), .D (new_AGEMA_signal_4864), .Q (new_AGEMA_signal_4865) ) ;
    buf_clk new_AGEMA_reg_buffer_2101 ( .C (CLK), .D (new_AGEMA_signal_4868), .Q (new_AGEMA_signal_4869) ) ;
    buf_clk new_AGEMA_reg_buffer_2105 ( .C (CLK), .D (new_AGEMA_signal_4872), .Q (new_AGEMA_signal_4873) ) ;
    buf_clk new_AGEMA_reg_buffer_2109 ( .C (CLK), .D (new_AGEMA_signal_4876), .Q (new_AGEMA_signal_4877) ) ;
    buf_clk new_AGEMA_reg_buffer_2113 ( .C (CLK), .D (new_AGEMA_signal_4880), .Q (new_AGEMA_signal_4881) ) ;
    buf_clk new_AGEMA_reg_buffer_2117 ( .C (CLK), .D (new_AGEMA_signal_4884), .Q (new_AGEMA_signal_4885) ) ;
    buf_clk new_AGEMA_reg_buffer_2121 ( .C (CLK), .D (new_AGEMA_signal_4888), .Q (new_AGEMA_signal_4889) ) ;
    buf_clk new_AGEMA_reg_buffer_2125 ( .C (CLK), .D (new_AGEMA_signal_4892), .Q (new_AGEMA_signal_4893) ) ;
    buf_clk new_AGEMA_reg_buffer_2129 ( .C (CLK), .D (new_AGEMA_signal_4896), .Q (new_AGEMA_signal_4897) ) ;
    buf_clk new_AGEMA_reg_buffer_2133 ( .C (CLK), .D (new_AGEMA_signal_4900), .Q (new_AGEMA_signal_4901) ) ;
    buf_clk new_AGEMA_reg_buffer_2137 ( .C (CLK), .D (new_AGEMA_signal_4904), .Q (new_AGEMA_signal_4905) ) ;
    buf_clk new_AGEMA_reg_buffer_2141 ( .C (CLK), .D (new_AGEMA_signal_4908), .Q (new_AGEMA_signal_4909) ) ;
    buf_clk new_AGEMA_reg_buffer_2145 ( .C (CLK), .D (new_AGEMA_signal_4912), .Q (new_AGEMA_signal_4913) ) ;
    buf_clk new_AGEMA_reg_buffer_2149 ( .C (CLK), .D (new_AGEMA_signal_4916), .Q (new_AGEMA_signal_4917) ) ;
    buf_clk new_AGEMA_reg_buffer_2153 ( .C (CLK), .D (new_AGEMA_signal_4920), .Q (new_AGEMA_signal_4921) ) ;
    buf_clk new_AGEMA_reg_buffer_2157 ( .C (CLK), .D (new_AGEMA_signal_4924), .Q (new_AGEMA_signal_4925) ) ;
    buf_clk new_AGEMA_reg_buffer_2161 ( .C (CLK), .D (new_AGEMA_signal_4928), .Q (new_AGEMA_signal_4929) ) ;
    buf_clk new_AGEMA_reg_buffer_2165 ( .C (CLK), .D (new_AGEMA_signal_4932), .Q (new_AGEMA_signal_4933) ) ;
    buf_clk new_AGEMA_reg_buffer_2169 ( .C (CLK), .D (new_AGEMA_signal_4936), .Q (new_AGEMA_signal_4937) ) ;
    buf_clk new_AGEMA_reg_buffer_2173 ( .C (CLK), .D (new_AGEMA_signal_4940), .Q (new_AGEMA_signal_4941) ) ;
    buf_clk new_AGEMA_reg_buffer_2177 ( .C (CLK), .D (new_AGEMA_signal_4944), .Q (new_AGEMA_signal_4945) ) ;
    buf_clk new_AGEMA_reg_buffer_2181 ( .C (CLK), .D (new_AGEMA_signal_4948), .Q (new_AGEMA_signal_4949) ) ;
    buf_clk new_AGEMA_reg_buffer_2185 ( .C (CLK), .D (new_AGEMA_signal_4952), .Q (new_AGEMA_signal_4953) ) ;
    buf_clk new_AGEMA_reg_buffer_2189 ( .C (CLK), .D (new_AGEMA_signal_4956), .Q (new_AGEMA_signal_4957) ) ;
    buf_clk new_AGEMA_reg_buffer_2193 ( .C (CLK), .D (new_AGEMA_signal_4960), .Q (new_AGEMA_signal_4961) ) ;
    buf_clk new_AGEMA_reg_buffer_2197 ( .C (CLK), .D (new_AGEMA_signal_4964), .Q (new_AGEMA_signal_4965) ) ;
    buf_clk new_AGEMA_reg_buffer_2201 ( .C (CLK), .D (new_AGEMA_signal_4968), .Q (new_AGEMA_signal_4969) ) ;
    buf_clk new_AGEMA_reg_buffer_2205 ( .C (CLK), .D (new_AGEMA_signal_4972), .Q (new_AGEMA_signal_4973) ) ;
    buf_clk new_AGEMA_reg_buffer_2209 ( .C (CLK), .D (new_AGEMA_signal_4976), .Q (new_AGEMA_signal_4977) ) ;
    buf_clk new_AGEMA_reg_buffer_2213 ( .C (CLK), .D (new_AGEMA_signal_4980), .Q (new_AGEMA_signal_4981) ) ;
    buf_clk new_AGEMA_reg_buffer_2217 ( .C (CLK), .D (new_AGEMA_signal_4984), .Q (new_AGEMA_signal_4985) ) ;
    buf_clk new_AGEMA_reg_buffer_2221 ( .C (CLK), .D (new_AGEMA_signal_4988), .Q (new_AGEMA_signal_4989) ) ;
    buf_clk new_AGEMA_reg_buffer_2225 ( .C (CLK), .D (new_AGEMA_signal_4992), .Q (new_AGEMA_signal_4993) ) ;
    buf_clk new_AGEMA_reg_buffer_2229 ( .C (CLK), .D (new_AGEMA_signal_4996), .Q (new_AGEMA_signal_4997) ) ;
    buf_clk new_AGEMA_reg_buffer_2233 ( .C (CLK), .D (new_AGEMA_signal_5000), .Q (new_AGEMA_signal_5001) ) ;
    buf_clk new_AGEMA_reg_buffer_2237 ( .C (CLK), .D (new_AGEMA_signal_5004), .Q (new_AGEMA_signal_5005) ) ;
    buf_clk new_AGEMA_reg_buffer_2241 ( .C (CLK), .D (new_AGEMA_signal_5008), .Q (new_AGEMA_signal_5009) ) ;
    buf_clk new_AGEMA_reg_buffer_2245 ( .C (CLK), .D (new_AGEMA_signal_5012), .Q (new_AGEMA_signal_5013) ) ;
    buf_clk new_AGEMA_reg_buffer_2249 ( .C (CLK), .D (new_AGEMA_signal_5016), .Q (new_AGEMA_signal_5017) ) ;
    buf_clk new_AGEMA_reg_buffer_2253 ( .C (CLK), .D (new_AGEMA_signal_5020), .Q (new_AGEMA_signal_5021) ) ;
    buf_clk new_AGEMA_reg_buffer_2257 ( .C (CLK), .D (new_AGEMA_signal_5024), .Q (new_AGEMA_signal_5025) ) ;
    buf_clk new_AGEMA_reg_buffer_2261 ( .C (CLK), .D (new_AGEMA_signal_5028), .Q (new_AGEMA_signal_5029) ) ;
    buf_clk new_AGEMA_reg_buffer_2265 ( .C (CLK), .D (new_AGEMA_signal_5032), .Q (new_AGEMA_signal_5033) ) ;
    buf_clk new_AGEMA_reg_buffer_2269 ( .C (CLK), .D (new_AGEMA_signal_5036), .Q (new_AGEMA_signal_5037) ) ;
    buf_clk new_AGEMA_reg_buffer_2273 ( .C (CLK), .D (new_AGEMA_signal_5040), .Q (new_AGEMA_signal_5041) ) ;
    buf_clk new_AGEMA_reg_buffer_2277 ( .C (CLK), .D (new_AGEMA_signal_5044), .Q (new_AGEMA_signal_5045) ) ;
    buf_clk new_AGEMA_reg_buffer_2281 ( .C (CLK), .D (new_AGEMA_signal_5048), .Q (new_AGEMA_signal_5049) ) ;
    buf_clk new_AGEMA_reg_buffer_2285 ( .C (CLK), .D (new_AGEMA_signal_5052), .Q (new_AGEMA_signal_5053) ) ;
    buf_clk new_AGEMA_reg_buffer_2289 ( .C (CLK), .D (new_AGEMA_signal_5056), .Q (new_AGEMA_signal_5057) ) ;
    buf_clk new_AGEMA_reg_buffer_2293 ( .C (CLK), .D (new_AGEMA_signal_5060), .Q (new_AGEMA_signal_5061) ) ;
    buf_clk new_AGEMA_reg_buffer_2297 ( .C (CLK), .D (new_AGEMA_signal_5064), .Q (new_AGEMA_signal_5065) ) ;
    buf_clk new_AGEMA_reg_buffer_2301 ( .C (CLK), .D (new_AGEMA_signal_5068), .Q (new_AGEMA_signal_5069) ) ;
    buf_clk new_AGEMA_reg_buffer_2305 ( .C (CLK), .D (new_AGEMA_signal_5072), .Q (new_AGEMA_signal_5073) ) ;
    buf_clk new_AGEMA_reg_buffer_2309 ( .C (CLK), .D (new_AGEMA_signal_5076), .Q (new_AGEMA_signal_5077) ) ;
    buf_clk new_AGEMA_reg_buffer_2313 ( .C (CLK), .D (new_AGEMA_signal_5080), .Q (new_AGEMA_signal_5081) ) ;
    buf_clk new_AGEMA_reg_buffer_2317 ( .C (CLK), .D (new_AGEMA_signal_5084), .Q (new_AGEMA_signal_5085) ) ;
    buf_clk new_AGEMA_reg_buffer_2321 ( .C (CLK), .D (new_AGEMA_signal_5088), .Q (new_AGEMA_signal_5089) ) ;
    buf_clk new_AGEMA_reg_buffer_2325 ( .C (CLK), .D (new_AGEMA_signal_5092), .Q (new_AGEMA_signal_5093) ) ;
    buf_clk new_AGEMA_reg_buffer_2329 ( .C (CLK), .D (new_AGEMA_signal_5096), .Q (new_AGEMA_signal_5097) ) ;
    buf_clk new_AGEMA_reg_buffer_2333 ( .C (CLK), .D (new_AGEMA_signal_5100), .Q (new_AGEMA_signal_5101) ) ;
    buf_clk new_AGEMA_reg_buffer_2337 ( .C (CLK), .D (new_AGEMA_signal_5104), .Q (new_AGEMA_signal_5105) ) ;
    buf_clk new_AGEMA_reg_buffer_2341 ( .C (CLK), .D (new_AGEMA_signal_5108), .Q (new_AGEMA_signal_5109) ) ;
    buf_clk new_AGEMA_reg_buffer_2345 ( .C (CLK), .D (new_AGEMA_signal_5112), .Q (new_AGEMA_signal_5113) ) ;
    buf_clk new_AGEMA_reg_buffer_2349 ( .C (CLK), .D (new_AGEMA_signal_5116), .Q (new_AGEMA_signal_5117) ) ;
    buf_clk new_AGEMA_reg_buffer_2353 ( .C (CLK), .D (new_AGEMA_signal_5120), .Q (new_AGEMA_signal_5121) ) ;
    buf_clk new_AGEMA_reg_buffer_2357 ( .C (CLK), .D (new_AGEMA_signal_5124), .Q (new_AGEMA_signal_5125) ) ;
    buf_clk new_AGEMA_reg_buffer_2361 ( .C (CLK), .D (new_AGEMA_signal_5128), .Q (new_AGEMA_signal_5129) ) ;
    buf_clk new_AGEMA_reg_buffer_2365 ( .C (CLK), .D (new_AGEMA_signal_5132), .Q (new_AGEMA_signal_5133) ) ;
    buf_clk new_AGEMA_reg_buffer_2369 ( .C (CLK), .D (new_AGEMA_signal_5136), .Q (new_AGEMA_signal_5137) ) ;
    buf_clk new_AGEMA_reg_buffer_2373 ( .C (CLK), .D (new_AGEMA_signal_5140), .Q (new_AGEMA_signal_5141) ) ;
    buf_clk new_AGEMA_reg_buffer_2377 ( .C (CLK), .D (new_AGEMA_signal_5144), .Q (new_AGEMA_signal_5145) ) ;
    buf_clk new_AGEMA_reg_buffer_2381 ( .C (CLK), .D (new_AGEMA_signal_5148), .Q (new_AGEMA_signal_5149) ) ;
    buf_clk new_AGEMA_reg_buffer_2385 ( .C (CLK), .D (new_AGEMA_signal_5152), .Q (new_AGEMA_signal_5153) ) ;
    buf_clk new_AGEMA_reg_buffer_2389 ( .C (CLK), .D (new_AGEMA_signal_5156), .Q (new_AGEMA_signal_5157) ) ;
    buf_clk new_AGEMA_reg_buffer_2393 ( .C (CLK), .D (new_AGEMA_signal_5160), .Q (new_AGEMA_signal_5161) ) ;
    buf_clk new_AGEMA_reg_buffer_2397 ( .C (CLK), .D (new_AGEMA_signal_5164), .Q (new_AGEMA_signal_5165) ) ;
    buf_clk new_AGEMA_reg_buffer_2401 ( .C (CLK), .D (new_AGEMA_signal_5168), .Q (new_AGEMA_signal_5169) ) ;
    buf_clk new_AGEMA_reg_buffer_2405 ( .C (CLK), .D (new_AGEMA_signal_5172), .Q (new_AGEMA_signal_5173) ) ;
    buf_clk new_AGEMA_reg_buffer_2409 ( .C (CLK), .D (new_AGEMA_signal_5176), .Q (new_AGEMA_signal_5177) ) ;
    buf_clk new_AGEMA_reg_buffer_2413 ( .C (CLK), .D (new_AGEMA_signal_5180), .Q (new_AGEMA_signal_5181) ) ;
    buf_clk new_AGEMA_reg_buffer_2417 ( .C (CLK), .D (new_AGEMA_signal_5184), .Q (new_AGEMA_signal_5185) ) ;
    buf_clk new_AGEMA_reg_buffer_2421 ( .C (CLK), .D (new_AGEMA_signal_5188), .Q (new_AGEMA_signal_5189) ) ;
    buf_clk new_AGEMA_reg_buffer_2425 ( .C (CLK), .D (new_AGEMA_signal_5192), .Q (new_AGEMA_signal_5193) ) ;
    buf_clk new_AGEMA_reg_buffer_2429 ( .C (CLK), .D (new_AGEMA_signal_5196), .Q (new_AGEMA_signal_5197) ) ;
    buf_clk new_AGEMA_reg_buffer_2433 ( .C (CLK), .D (new_AGEMA_signal_5200), .Q (new_AGEMA_signal_5201) ) ;
    buf_clk new_AGEMA_reg_buffer_2437 ( .C (CLK), .D (new_AGEMA_signal_5204), .Q (new_AGEMA_signal_5205) ) ;
    buf_clk new_AGEMA_reg_buffer_2441 ( .C (CLK), .D (new_AGEMA_signal_5208), .Q (new_AGEMA_signal_5209) ) ;
    buf_clk new_AGEMA_reg_buffer_2445 ( .C (CLK), .D (new_AGEMA_signal_5212), .Q (new_AGEMA_signal_5213) ) ;
    buf_clk new_AGEMA_reg_buffer_2449 ( .C (CLK), .D (new_AGEMA_signal_5216), .Q (new_AGEMA_signal_5217) ) ;
    buf_clk new_AGEMA_reg_buffer_2453 ( .C (CLK), .D (new_AGEMA_signal_5220), .Q (new_AGEMA_signal_5221) ) ;
    buf_clk new_AGEMA_reg_buffer_2457 ( .C (CLK), .D (new_AGEMA_signal_5224), .Q (new_AGEMA_signal_5225) ) ;
    buf_clk new_AGEMA_reg_buffer_2461 ( .C (CLK), .D (new_AGEMA_signal_5228), .Q (new_AGEMA_signal_5229) ) ;
    buf_clk new_AGEMA_reg_buffer_2465 ( .C (CLK), .D (new_AGEMA_signal_5232), .Q (new_AGEMA_signal_5233) ) ;
    buf_clk new_AGEMA_reg_buffer_2469 ( .C (CLK), .D (new_AGEMA_signal_5236), .Q (new_AGEMA_signal_5237) ) ;
    buf_clk new_AGEMA_reg_buffer_2473 ( .C (CLK), .D (new_AGEMA_signal_5240), .Q (new_AGEMA_signal_5241) ) ;
    buf_clk new_AGEMA_reg_buffer_2477 ( .C (CLK), .D (new_AGEMA_signal_5244), .Q (new_AGEMA_signal_5245) ) ;
    buf_clk new_AGEMA_reg_buffer_2481 ( .C (CLK), .D (new_AGEMA_signal_5248), .Q (new_AGEMA_signal_5249) ) ;
    buf_clk new_AGEMA_reg_buffer_2485 ( .C (CLK), .D (new_AGEMA_signal_5252), .Q (new_AGEMA_signal_5253) ) ;
    buf_clk new_AGEMA_reg_buffer_2489 ( .C (CLK), .D (new_AGEMA_signal_5256), .Q (new_AGEMA_signal_5257) ) ;
    buf_clk new_AGEMA_reg_buffer_2493 ( .C (CLK), .D (new_AGEMA_signal_5260), .Q (new_AGEMA_signal_5261) ) ;
    buf_clk new_AGEMA_reg_buffer_2497 ( .C (CLK), .D (new_AGEMA_signal_5264), .Q (new_AGEMA_signal_5265) ) ;
    buf_clk new_AGEMA_reg_buffer_2501 ( .C (CLK), .D (new_AGEMA_signal_5268), .Q (new_AGEMA_signal_5269) ) ;
    buf_clk new_AGEMA_reg_buffer_2505 ( .C (CLK), .D (new_AGEMA_signal_5272), .Q (new_AGEMA_signal_5273) ) ;
    buf_clk new_AGEMA_reg_buffer_2509 ( .C (CLK), .D (new_AGEMA_signal_5276), .Q (new_AGEMA_signal_5277) ) ;
    buf_clk new_AGEMA_reg_buffer_2513 ( .C (CLK), .D (new_AGEMA_signal_5280), .Q (new_AGEMA_signal_5281) ) ;
    buf_clk new_AGEMA_reg_buffer_2517 ( .C (CLK), .D (new_AGEMA_signal_5284), .Q (new_AGEMA_signal_5285) ) ;
    buf_clk new_AGEMA_reg_buffer_2521 ( .C (CLK), .D (new_AGEMA_signal_5288), .Q (new_AGEMA_signal_5289) ) ;
    buf_clk new_AGEMA_reg_buffer_2525 ( .C (CLK), .D (new_AGEMA_signal_5292), .Q (new_AGEMA_signal_5293) ) ;
    buf_clk new_AGEMA_reg_buffer_2529 ( .C (CLK), .D (new_AGEMA_signal_5296), .Q (new_AGEMA_signal_5297) ) ;
    buf_clk new_AGEMA_reg_buffer_2533 ( .C (CLK), .D (new_AGEMA_signal_5300), .Q (new_AGEMA_signal_5301) ) ;
    buf_clk new_AGEMA_reg_buffer_2537 ( .C (CLK), .D (new_AGEMA_signal_5304), .Q (new_AGEMA_signal_5305) ) ;
    buf_clk new_AGEMA_reg_buffer_2541 ( .C (CLK), .D (new_AGEMA_signal_5308), .Q (new_AGEMA_signal_5309) ) ;
    buf_clk new_AGEMA_reg_buffer_2545 ( .C (CLK), .D (new_AGEMA_signal_5312), .Q (new_AGEMA_signal_5313) ) ;
    buf_clk new_AGEMA_reg_buffer_2549 ( .C (CLK), .D (new_AGEMA_signal_5316), .Q (new_AGEMA_signal_5317) ) ;
    buf_clk new_AGEMA_reg_buffer_2553 ( .C (CLK), .D (new_AGEMA_signal_5320), .Q (new_AGEMA_signal_5321) ) ;
    buf_clk new_AGEMA_reg_buffer_2557 ( .C (CLK), .D (new_AGEMA_signal_5324), .Q (new_AGEMA_signal_5325) ) ;
    buf_clk new_AGEMA_reg_buffer_2561 ( .C (CLK), .D (new_AGEMA_signal_5328), .Q (new_AGEMA_signal_5329) ) ;
    buf_clk new_AGEMA_reg_buffer_2565 ( .C (CLK), .D (new_AGEMA_signal_5332), .Q (new_AGEMA_signal_5333) ) ;
    buf_clk new_AGEMA_reg_buffer_2569 ( .C (CLK), .D (new_AGEMA_signal_5336), .Q (new_AGEMA_signal_5337) ) ;
    buf_clk new_AGEMA_reg_buffer_2573 ( .C (CLK), .D (new_AGEMA_signal_5340), .Q (new_AGEMA_signal_5341) ) ;
    buf_clk new_AGEMA_reg_buffer_2577 ( .C (CLK), .D (new_AGEMA_signal_5344), .Q (new_AGEMA_signal_5345) ) ;
    buf_clk new_AGEMA_reg_buffer_2581 ( .C (CLK), .D (new_AGEMA_signal_5348), .Q (new_AGEMA_signal_5349) ) ;
    buf_clk new_AGEMA_reg_buffer_2585 ( .C (CLK), .D (new_AGEMA_signal_5352), .Q (new_AGEMA_signal_5353) ) ;
    buf_clk new_AGEMA_reg_buffer_2589 ( .C (CLK), .D (new_AGEMA_signal_5356), .Q (new_AGEMA_signal_5357) ) ;
    buf_clk new_AGEMA_reg_buffer_2593 ( .C (CLK), .D (new_AGEMA_signal_5360), .Q (new_AGEMA_signal_5361) ) ;
    buf_clk new_AGEMA_reg_buffer_2597 ( .C (CLK), .D (new_AGEMA_signal_5364), .Q (new_AGEMA_signal_5365) ) ;
    buf_clk new_AGEMA_reg_buffer_2601 ( .C (CLK), .D (new_AGEMA_signal_5368), .Q (new_AGEMA_signal_5369) ) ;
    buf_clk new_AGEMA_reg_buffer_2605 ( .C (CLK), .D (new_AGEMA_signal_5372), .Q (new_AGEMA_signal_5373) ) ;
    buf_clk new_AGEMA_reg_buffer_2609 ( .C (CLK), .D (new_AGEMA_signal_5376), .Q (new_AGEMA_signal_5377) ) ;
    buf_clk new_AGEMA_reg_buffer_2613 ( .C (CLK), .D (new_AGEMA_signal_5380), .Q (new_AGEMA_signal_5381) ) ;
    buf_clk new_AGEMA_reg_buffer_2617 ( .C (CLK), .D (new_AGEMA_signal_5384), .Q (new_AGEMA_signal_5385) ) ;
    buf_clk new_AGEMA_reg_buffer_2621 ( .C (CLK), .D (new_AGEMA_signal_5388), .Q (new_AGEMA_signal_5389) ) ;
    buf_clk new_AGEMA_reg_buffer_2625 ( .C (CLK), .D (new_AGEMA_signal_5392), .Q (new_AGEMA_signal_5393) ) ;
    buf_clk new_AGEMA_reg_buffer_2629 ( .C (CLK), .D (new_AGEMA_signal_5396), .Q (new_AGEMA_signal_5397) ) ;
    buf_clk new_AGEMA_reg_buffer_2633 ( .C (CLK), .D (new_AGEMA_signal_5400), .Q (new_AGEMA_signal_5401) ) ;
    buf_clk new_AGEMA_reg_buffer_2637 ( .C (CLK), .D (new_AGEMA_signal_5404), .Q (new_AGEMA_signal_5405) ) ;
    buf_clk new_AGEMA_reg_buffer_2641 ( .C (CLK), .D (new_AGEMA_signal_5408), .Q (new_AGEMA_signal_5409) ) ;
    buf_clk new_AGEMA_reg_buffer_2645 ( .C (CLK), .D (new_AGEMA_signal_5412), .Q (new_AGEMA_signal_5413) ) ;
    buf_clk new_AGEMA_reg_buffer_2649 ( .C (CLK), .D (new_AGEMA_signal_5416), .Q (new_AGEMA_signal_5417) ) ;
    buf_clk new_AGEMA_reg_buffer_2653 ( .C (CLK), .D (new_AGEMA_signal_5420), .Q (new_AGEMA_signal_5421) ) ;
    buf_clk new_AGEMA_reg_buffer_2657 ( .C (CLK), .D (new_AGEMA_signal_5424), .Q (new_AGEMA_signal_5425) ) ;
    buf_clk new_AGEMA_reg_buffer_2661 ( .C (CLK), .D (new_AGEMA_signal_5428), .Q (new_AGEMA_signal_5429) ) ;
    buf_clk new_AGEMA_reg_buffer_2665 ( .C (CLK), .D (new_AGEMA_signal_5432), .Q (new_AGEMA_signal_5433) ) ;
    buf_clk new_AGEMA_reg_buffer_2669 ( .C (CLK), .D (new_AGEMA_signal_5436), .Q (new_AGEMA_signal_5437) ) ;
    buf_clk new_AGEMA_reg_buffer_2673 ( .C (CLK), .D (new_AGEMA_signal_5440), .Q (new_AGEMA_signal_5441) ) ;
    buf_clk new_AGEMA_reg_buffer_2677 ( .C (CLK), .D (new_AGEMA_signal_5444), .Q (new_AGEMA_signal_5445) ) ;
    buf_clk new_AGEMA_reg_buffer_2681 ( .C (CLK), .D (new_AGEMA_signal_5448), .Q (new_AGEMA_signal_5449) ) ;
    buf_clk new_AGEMA_reg_buffer_2685 ( .C (CLK), .D (new_AGEMA_signal_5452), .Q (new_AGEMA_signal_5453) ) ;
    buf_clk new_AGEMA_reg_buffer_2689 ( .C (CLK), .D (new_AGEMA_signal_5456), .Q (new_AGEMA_signal_5457) ) ;
    buf_clk new_AGEMA_reg_buffer_2693 ( .C (CLK), .D (new_AGEMA_signal_5460), .Q (new_AGEMA_signal_5461) ) ;
    buf_clk new_AGEMA_reg_buffer_2697 ( .C (CLK), .D (new_AGEMA_signal_5464), .Q (new_AGEMA_signal_5465) ) ;
    buf_clk new_AGEMA_reg_buffer_2701 ( .C (CLK), .D (new_AGEMA_signal_5468), .Q (new_AGEMA_signal_5469) ) ;
    buf_clk new_AGEMA_reg_buffer_2705 ( .C (CLK), .D (new_AGEMA_signal_5472), .Q (new_AGEMA_signal_5473) ) ;
    buf_clk new_AGEMA_reg_buffer_2709 ( .C (CLK), .D (new_AGEMA_signal_5476), .Q (new_AGEMA_signal_5477) ) ;
    buf_clk new_AGEMA_reg_buffer_2713 ( .C (CLK), .D (new_AGEMA_signal_5480), .Q (new_AGEMA_signal_5481) ) ;
    buf_clk new_AGEMA_reg_buffer_2717 ( .C (CLK), .D (new_AGEMA_signal_5484), .Q (new_AGEMA_signal_5485) ) ;
    buf_clk new_AGEMA_reg_buffer_2721 ( .C (CLK), .D (new_AGEMA_signal_5488), .Q (new_AGEMA_signal_5489) ) ;
    buf_clk new_AGEMA_reg_buffer_2725 ( .C (CLK), .D (new_AGEMA_signal_5492), .Q (new_AGEMA_signal_5493) ) ;
    buf_clk new_AGEMA_reg_buffer_2729 ( .C (CLK), .D (new_AGEMA_signal_5496), .Q (new_AGEMA_signal_5497) ) ;
    buf_clk new_AGEMA_reg_buffer_2733 ( .C (CLK), .D (new_AGEMA_signal_5500), .Q (new_AGEMA_signal_5501) ) ;
    buf_clk new_AGEMA_reg_buffer_2737 ( .C (CLK), .D (new_AGEMA_signal_5504), .Q (new_AGEMA_signal_5505) ) ;
    buf_clk new_AGEMA_reg_buffer_2741 ( .C (CLK), .D (new_AGEMA_signal_5508), .Q (new_AGEMA_signal_5509) ) ;
    buf_clk new_AGEMA_reg_buffer_2745 ( .C (CLK), .D (new_AGEMA_signal_5512), .Q (new_AGEMA_signal_5513) ) ;
    buf_clk new_AGEMA_reg_buffer_2749 ( .C (CLK), .D (new_AGEMA_signal_5516), .Q (new_AGEMA_signal_5517) ) ;
    buf_clk new_AGEMA_reg_buffer_2753 ( .C (CLK), .D (new_AGEMA_signal_5520), .Q (new_AGEMA_signal_5521) ) ;
    buf_clk new_AGEMA_reg_buffer_2757 ( .C (CLK), .D (new_AGEMA_signal_5524), .Q (new_AGEMA_signal_5525) ) ;
    buf_clk new_AGEMA_reg_buffer_2761 ( .C (CLK), .D (new_AGEMA_signal_5528), .Q (new_AGEMA_signal_5529) ) ;
    buf_clk new_AGEMA_reg_buffer_2765 ( .C (CLK), .D (new_AGEMA_signal_5532), .Q (new_AGEMA_signal_5533) ) ;
    buf_clk new_AGEMA_reg_buffer_2769 ( .C (CLK), .D (new_AGEMA_signal_5536), .Q (new_AGEMA_signal_5537) ) ;
    buf_clk new_AGEMA_reg_buffer_2773 ( .C (CLK), .D (new_AGEMA_signal_5540), .Q (new_AGEMA_signal_5541) ) ;
    buf_clk new_AGEMA_reg_buffer_2777 ( .C (CLK), .D (new_AGEMA_signal_5544), .Q (new_AGEMA_signal_5545) ) ;
    buf_clk new_AGEMA_reg_buffer_2781 ( .C (CLK), .D (new_AGEMA_signal_5548), .Q (new_AGEMA_signal_5549) ) ;
    buf_clk new_AGEMA_reg_buffer_2785 ( .C (CLK), .D (new_AGEMA_signal_5552), .Q (new_AGEMA_signal_5553) ) ;
    buf_clk new_AGEMA_reg_buffer_2789 ( .C (CLK), .D (new_AGEMA_signal_5556), .Q (new_AGEMA_signal_5557) ) ;
    buf_clk new_AGEMA_reg_buffer_2793 ( .C (CLK), .D (new_AGEMA_signal_5560), .Q (new_AGEMA_signal_5561) ) ;
    buf_clk new_AGEMA_reg_buffer_2797 ( .C (CLK), .D (new_AGEMA_signal_5564), .Q (new_AGEMA_signal_5565) ) ;
    buf_clk new_AGEMA_reg_buffer_2801 ( .C (CLK), .D (new_AGEMA_signal_5568), .Q (new_AGEMA_signal_5569) ) ;
    buf_clk new_AGEMA_reg_buffer_2805 ( .C (CLK), .D (new_AGEMA_signal_5572), .Q (new_AGEMA_signal_5573) ) ;
    buf_clk new_AGEMA_reg_buffer_2809 ( .C (CLK), .D (new_AGEMA_signal_5576), .Q (new_AGEMA_signal_5577) ) ;
    buf_clk new_AGEMA_reg_buffer_2813 ( .C (CLK), .D (new_AGEMA_signal_5580), .Q (new_AGEMA_signal_5581) ) ;
    buf_clk new_AGEMA_reg_buffer_2817 ( .C (CLK), .D (new_AGEMA_signal_5584), .Q (new_AGEMA_signal_5585) ) ;
    buf_clk new_AGEMA_reg_buffer_2821 ( .C (CLK), .D (new_AGEMA_signal_5588), .Q (new_AGEMA_signal_5589) ) ;
    buf_clk new_AGEMA_reg_buffer_2825 ( .C (CLK), .D (new_AGEMA_signal_5592), .Q (new_AGEMA_signal_5593) ) ;
    buf_clk new_AGEMA_reg_buffer_2829 ( .C (CLK), .D (new_AGEMA_signal_5596), .Q (new_AGEMA_signal_5597) ) ;
    buf_clk new_AGEMA_reg_buffer_2833 ( .C (CLK), .D (new_AGEMA_signal_5600), .Q (new_AGEMA_signal_5601) ) ;
    buf_clk new_AGEMA_reg_buffer_2837 ( .C (CLK), .D (new_AGEMA_signal_5604), .Q (new_AGEMA_signal_5605) ) ;
    buf_clk new_AGEMA_reg_buffer_2841 ( .C (CLK), .D (new_AGEMA_signal_5608), .Q (new_AGEMA_signal_5609) ) ;
    buf_clk new_AGEMA_reg_buffer_2845 ( .C (CLK), .D (new_AGEMA_signal_5612), .Q (new_AGEMA_signal_5613) ) ;
    buf_clk new_AGEMA_reg_buffer_2849 ( .C (CLK), .D (new_AGEMA_signal_5616), .Q (new_AGEMA_signal_5617) ) ;
    buf_clk new_AGEMA_reg_buffer_2853 ( .C (CLK), .D (new_AGEMA_signal_5620), .Q (new_AGEMA_signal_5621) ) ;
    buf_clk new_AGEMA_reg_buffer_2857 ( .C (CLK), .D (new_AGEMA_signal_5624), .Q (new_AGEMA_signal_5625) ) ;
    buf_clk new_AGEMA_reg_buffer_2861 ( .C (CLK), .D (new_AGEMA_signal_5628), .Q (new_AGEMA_signal_5629) ) ;
    buf_clk new_AGEMA_reg_buffer_2865 ( .C (CLK), .D (new_AGEMA_signal_5632), .Q (new_AGEMA_signal_5633) ) ;
    buf_clk new_AGEMA_reg_buffer_2869 ( .C (CLK), .D (new_AGEMA_signal_5636), .Q (new_AGEMA_signal_5637) ) ;
    buf_clk new_AGEMA_reg_buffer_2873 ( .C (CLK), .D (new_AGEMA_signal_5640), .Q (new_AGEMA_signal_5641) ) ;
    buf_clk new_AGEMA_reg_buffer_2877 ( .C (CLK), .D (new_AGEMA_signal_5644), .Q (new_AGEMA_signal_5645) ) ;
    buf_clk new_AGEMA_reg_buffer_2881 ( .C (CLK), .D (new_AGEMA_signal_5648), .Q (new_AGEMA_signal_5649) ) ;
    buf_clk new_AGEMA_reg_buffer_2885 ( .C (CLK), .D (new_AGEMA_signal_5652), .Q (new_AGEMA_signal_5653) ) ;
    buf_clk new_AGEMA_reg_buffer_2889 ( .C (CLK), .D (new_AGEMA_signal_5656), .Q (new_AGEMA_signal_5657) ) ;
    buf_clk new_AGEMA_reg_buffer_2893 ( .C (CLK), .D (new_AGEMA_signal_5660), .Q (new_AGEMA_signal_5661) ) ;
    buf_clk new_AGEMA_reg_buffer_2897 ( .C (CLK), .D (new_AGEMA_signal_5664), .Q (new_AGEMA_signal_5665) ) ;
    buf_clk new_AGEMA_reg_buffer_2901 ( .C (CLK), .D (new_AGEMA_signal_5668), .Q (new_AGEMA_signal_5669) ) ;
    buf_clk new_AGEMA_reg_buffer_2905 ( .C (CLK), .D (new_AGEMA_signal_5672), .Q (new_AGEMA_signal_5673) ) ;
    buf_clk new_AGEMA_reg_buffer_2909 ( .C (CLK), .D (new_AGEMA_signal_5676), .Q (new_AGEMA_signal_5677) ) ;
    buf_clk new_AGEMA_reg_buffer_2913 ( .C (CLK), .D (new_AGEMA_signal_5680), .Q (new_AGEMA_signal_5681) ) ;
    buf_clk new_AGEMA_reg_buffer_2917 ( .C (CLK), .D (new_AGEMA_signal_5684), .Q (new_AGEMA_signal_5685) ) ;
    buf_clk new_AGEMA_reg_buffer_2921 ( .C (CLK), .D (new_AGEMA_signal_5688), .Q (new_AGEMA_signal_5689) ) ;
    buf_clk new_AGEMA_reg_buffer_2925 ( .C (CLK), .D (new_AGEMA_signal_5692), .Q (new_AGEMA_signal_5693) ) ;
    buf_clk new_AGEMA_reg_buffer_2929 ( .C (CLK), .D (new_AGEMA_signal_5696), .Q (new_AGEMA_signal_5697) ) ;
    buf_clk new_AGEMA_reg_buffer_2933 ( .C (CLK), .D (new_AGEMA_signal_5700), .Q (new_AGEMA_signal_5701) ) ;
    buf_clk new_AGEMA_reg_buffer_2937 ( .C (CLK), .D (new_AGEMA_signal_5704), .Q (new_AGEMA_signal_5705) ) ;
    buf_clk new_AGEMA_reg_buffer_2941 ( .C (CLK), .D (new_AGEMA_signal_5708), .Q (new_AGEMA_signal_5709) ) ;
    buf_clk new_AGEMA_reg_buffer_2945 ( .C (CLK), .D (new_AGEMA_signal_5712), .Q (new_AGEMA_signal_5713) ) ;
    buf_clk new_AGEMA_reg_buffer_2949 ( .C (CLK), .D (new_AGEMA_signal_5716), .Q (new_AGEMA_signal_5717) ) ;
    buf_clk new_AGEMA_reg_buffer_2953 ( .C (CLK), .D (new_AGEMA_signal_5720), .Q (new_AGEMA_signal_5721) ) ;
    buf_clk new_AGEMA_reg_buffer_2957 ( .C (CLK), .D (new_AGEMA_signal_5724), .Q (new_AGEMA_signal_5725) ) ;
    buf_clk new_AGEMA_reg_buffer_2961 ( .C (CLK), .D (new_AGEMA_signal_5728), .Q (new_AGEMA_signal_5729) ) ;
    buf_clk new_AGEMA_reg_buffer_2965 ( .C (CLK), .D (new_AGEMA_signal_5732), .Q (new_AGEMA_signal_5733) ) ;
    buf_clk new_AGEMA_reg_buffer_2969 ( .C (CLK), .D (new_AGEMA_signal_5736), .Q (new_AGEMA_signal_5737) ) ;
    buf_clk new_AGEMA_reg_buffer_2973 ( .C (CLK), .D (new_AGEMA_signal_5740), .Q (new_AGEMA_signal_5741) ) ;
    buf_clk new_AGEMA_reg_buffer_2975 ( .C (CLK), .D (new_AGEMA_signal_5742), .Q (new_AGEMA_signal_5743) ) ;
    buf_clk new_AGEMA_reg_buffer_2977 ( .C (CLK), .D (new_AGEMA_signal_5744), .Q (new_AGEMA_signal_5745) ) ;
    buf_clk new_AGEMA_reg_buffer_2979 ( .C (CLK), .D (new_AGEMA_signal_5746), .Q (new_AGEMA_signal_5747) ) ;
    buf_clk new_AGEMA_reg_buffer_2981 ( .C (CLK), .D (new_AGEMA_signal_5748), .Q (new_AGEMA_signal_5749) ) ;
    buf_clk new_AGEMA_reg_buffer_2983 ( .C (CLK), .D (new_AGEMA_signal_5750), .Q (new_AGEMA_signal_5751) ) ;
    buf_clk new_AGEMA_reg_buffer_2991 ( .C (CLK), .D (new_AGEMA_signal_5758), .Q (new_AGEMA_signal_5759) ) ;
    buf_clk new_AGEMA_reg_buffer_2995 ( .C (CLK), .D (new_AGEMA_signal_5762), .Q (new_AGEMA_signal_5763) ) ;
    buf_clk new_AGEMA_reg_buffer_2999 ( .C (CLK), .D (new_AGEMA_signal_5766), .Q (new_AGEMA_signal_5767) ) ;
    buf_clk new_AGEMA_reg_buffer_3003 ( .C (CLK), .D (new_AGEMA_signal_5770), .Q (new_AGEMA_signal_5771) ) ;
    buf_clk new_AGEMA_reg_buffer_3007 ( .C (CLK), .D (new_AGEMA_signal_5774), .Q (new_AGEMA_signal_5775) ) ;
    buf_clk new_AGEMA_reg_buffer_3011 ( .C (CLK), .D (new_AGEMA_signal_5778), .Q (new_AGEMA_signal_5779) ) ;
    buf_clk new_AGEMA_reg_buffer_3021 ( .C (CLK), .D (new_AGEMA_signal_5788), .Q (new_AGEMA_signal_5789) ) ;
    buf_clk new_AGEMA_reg_buffer_3023 ( .C (CLK), .D (new_AGEMA_signal_5790), .Q (new_AGEMA_signal_5791) ) ;
    buf_clk new_AGEMA_reg_buffer_3025 ( .C (CLK), .D (new_AGEMA_signal_5792), .Q (new_AGEMA_signal_5793) ) ;
    buf_clk new_AGEMA_reg_buffer_3027 ( .C (CLK), .D (new_AGEMA_signal_5794), .Q (new_AGEMA_signal_5795) ) ;
    buf_clk new_AGEMA_reg_buffer_3029 ( .C (CLK), .D (new_AGEMA_signal_5796), .Q (new_AGEMA_signal_5797) ) ;
    buf_clk new_AGEMA_reg_buffer_3031 ( .C (CLK), .D (new_AGEMA_signal_5798), .Q (new_AGEMA_signal_5799) ) ;
    buf_clk new_AGEMA_reg_buffer_3039 ( .C (CLK), .D (new_AGEMA_signal_5806), .Q (new_AGEMA_signal_5807) ) ;
    buf_clk new_AGEMA_reg_buffer_3043 ( .C (CLK), .D (new_AGEMA_signal_5810), .Q (new_AGEMA_signal_5811) ) ;
    buf_clk new_AGEMA_reg_buffer_3047 ( .C (CLK), .D (new_AGEMA_signal_5814), .Q (new_AGEMA_signal_5815) ) ;
    buf_clk new_AGEMA_reg_buffer_3051 ( .C (CLK), .D (new_AGEMA_signal_5818), .Q (new_AGEMA_signal_5819) ) ;
    buf_clk new_AGEMA_reg_buffer_3055 ( .C (CLK), .D (new_AGEMA_signal_5822), .Q (new_AGEMA_signal_5823) ) ;
    buf_clk new_AGEMA_reg_buffer_3059 ( .C (CLK), .D (new_AGEMA_signal_5826), .Q (new_AGEMA_signal_5827) ) ;
    buf_clk new_AGEMA_reg_buffer_3069 ( .C (CLK), .D (new_AGEMA_signal_5836), .Q (new_AGEMA_signal_5837) ) ;
    buf_clk new_AGEMA_reg_buffer_3071 ( .C (CLK), .D (new_AGEMA_signal_5838), .Q (new_AGEMA_signal_5839) ) ;
    buf_clk new_AGEMA_reg_buffer_3073 ( .C (CLK), .D (new_AGEMA_signal_5840), .Q (new_AGEMA_signal_5841) ) ;
    buf_clk new_AGEMA_reg_buffer_3075 ( .C (CLK), .D (new_AGEMA_signal_5842), .Q (new_AGEMA_signal_5843) ) ;
    buf_clk new_AGEMA_reg_buffer_3077 ( .C (CLK), .D (new_AGEMA_signal_5844), .Q (new_AGEMA_signal_5845) ) ;
    buf_clk new_AGEMA_reg_buffer_3079 ( .C (CLK), .D (new_AGEMA_signal_5846), .Q (new_AGEMA_signal_5847) ) ;
    buf_clk new_AGEMA_reg_buffer_3087 ( .C (CLK), .D (new_AGEMA_signal_5854), .Q (new_AGEMA_signal_5855) ) ;
    buf_clk new_AGEMA_reg_buffer_3091 ( .C (CLK), .D (new_AGEMA_signal_5858), .Q (new_AGEMA_signal_5859) ) ;
    buf_clk new_AGEMA_reg_buffer_3095 ( .C (CLK), .D (new_AGEMA_signal_5862), .Q (new_AGEMA_signal_5863) ) ;
    buf_clk new_AGEMA_reg_buffer_3105 ( .C (CLK), .D (new_AGEMA_signal_5872), .Q (new_AGEMA_signal_5873) ) ;
    buf_clk new_AGEMA_reg_buffer_3107 ( .C (CLK), .D (new_AGEMA_signal_5874), .Q (new_AGEMA_signal_5875) ) ;
    buf_clk new_AGEMA_reg_buffer_3109 ( .C (CLK), .D (new_AGEMA_signal_5876), .Q (new_AGEMA_signal_5877) ) ;
    buf_clk new_AGEMA_reg_buffer_3111 ( .C (CLK), .D (new_AGEMA_signal_5878), .Q (new_AGEMA_signal_5879) ) ;
    buf_clk new_AGEMA_reg_buffer_3113 ( .C (CLK), .D (new_AGEMA_signal_5880), .Q (new_AGEMA_signal_5881) ) ;
    buf_clk new_AGEMA_reg_buffer_3115 ( .C (CLK), .D (new_AGEMA_signal_5882), .Q (new_AGEMA_signal_5883) ) ;
    buf_clk new_AGEMA_reg_buffer_3123 ( .C (CLK), .D (new_AGEMA_signal_5890), .Q (new_AGEMA_signal_5891) ) ;
    buf_clk new_AGEMA_reg_buffer_3127 ( .C (CLK), .D (new_AGEMA_signal_5894), .Q (new_AGEMA_signal_5895) ) ;
    buf_clk new_AGEMA_reg_buffer_3131 ( .C (CLK), .D (new_AGEMA_signal_5898), .Q (new_AGEMA_signal_5899) ) ;
    buf_clk new_AGEMA_reg_buffer_3141 ( .C (CLK), .D (new_AGEMA_signal_5908), .Q (new_AGEMA_signal_5909) ) ;
    buf_clk new_AGEMA_reg_buffer_3143 ( .C (CLK), .D (new_AGEMA_signal_5910), .Q (new_AGEMA_signal_5911) ) ;
    buf_clk new_AGEMA_reg_buffer_3145 ( .C (CLK), .D (new_AGEMA_signal_5912), .Q (new_AGEMA_signal_5913) ) ;
    buf_clk new_AGEMA_reg_buffer_3147 ( .C (CLK), .D (new_AGEMA_signal_5914), .Q (new_AGEMA_signal_5915) ) ;
    buf_clk new_AGEMA_reg_buffer_3149 ( .C (CLK), .D (new_AGEMA_signal_5916), .Q (new_AGEMA_signal_5917) ) ;
    buf_clk new_AGEMA_reg_buffer_3151 ( .C (CLK), .D (new_AGEMA_signal_5918), .Q (new_AGEMA_signal_5919) ) ;
    buf_clk new_AGEMA_reg_buffer_3159 ( .C (CLK), .D (new_AGEMA_signal_5926), .Q (new_AGEMA_signal_5927) ) ;
    buf_clk new_AGEMA_reg_buffer_3163 ( .C (CLK), .D (new_AGEMA_signal_5930), .Q (new_AGEMA_signal_5931) ) ;
    buf_clk new_AGEMA_reg_buffer_3167 ( .C (CLK), .D (new_AGEMA_signal_5934), .Q (new_AGEMA_signal_5935) ) ;
    buf_clk new_AGEMA_reg_buffer_3171 ( .C (CLK), .D (new_AGEMA_signal_5938), .Q (new_AGEMA_signal_5939) ) ;
    buf_clk new_AGEMA_reg_buffer_3175 ( .C (CLK), .D (new_AGEMA_signal_5942), .Q (new_AGEMA_signal_5943) ) ;
    buf_clk new_AGEMA_reg_buffer_3179 ( .C (CLK), .D (new_AGEMA_signal_5946), .Q (new_AGEMA_signal_5947) ) ;
    buf_clk new_AGEMA_reg_buffer_3189 ( .C (CLK), .D (new_AGEMA_signal_5956), .Q (new_AGEMA_signal_5957) ) ;
    buf_clk new_AGEMA_reg_buffer_3191 ( .C (CLK), .D (new_AGEMA_signal_5958), .Q (new_AGEMA_signal_5959) ) ;
    buf_clk new_AGEMA_reg_buffer_3193 ( .C (CLK), .D (new_AGEMA_signal_5960), .Q (new_AGEMA_signal_5961) ) ;
    buf_clk new_AGEMA_reg_buffer_3195 ( .C (CLK), .D (new_AGEMA_signal_5962), .Q (new_AGEMA_signal_5963) ) ;
    buf_clk new_AGEMA_reg_buffer_3197 ( .C (CLK), .D (new_AGEMA_signal_5964), .Q (new_AGEMA_signal_5965) ) ;
    buf_clk new_AGEMA_reg_buffer_3199 ( .C (CLK), .D (new_AGEMA_signal_5966), .Q (new_AGEMA_signal_5967) ) ;
    buf_clk new_AGEMA_reg_buffer_3207 ( .C (CLK), .D (new_AGEMA_signal_5974), .Q (new_AGEMA_signal_5975) ) ;
    buf_clk new_AGEMA_reg_buffer_3211 ( .C (CLK), .D (new_AGEMA_signal_5978), .Q (new_AGEMA_signal_5979) ) ;
    buf_clk new_AGEMA_reg_buffer_3215 ( .C (CLK), .D (new_AGEMA_signal_5982), .Q (new_AGEMA_signal_5983) ) ;
    buf_clk new_AGEMA_reg_buffer_3219 ( .C (CLK), .D (new_AGEMA_signal_5986), .Q (new_AGEMA_signal_5987) ) ;
    buf_clk new_AGEMA_reg_buffer_3223 ( .C (CLK), .D (new_AGEMA_signal_5990), .Q (new_AGEMA_signal_5991) ) ;
    buf_clk new_AGEMA_reg_buffer_3227 ( .C (CLK), .D (new_AGEMA_signal_5994), .Q (new_AGEMA_signal_5995) ) ;
    buf_clk new_AGEMA_reg_buffer_3237 ( .C (CLK), .D (new_AGEMA_signal_6004), .Q (new_AGEMA_signal_6005) ) ;
    buf_clk new_AGEMA_reg_buffer_3239 ( .C (CLK), .D (new_AGEMA_signal_6006), .Q (new_AGEMA_signal_6007) ) ;
    buf_clk new_AGEMA_reg_buffer_3241 ( .C (CLK), .D (new_AGEMA_signal_6008), .Q (new_AGEMA_signal_6009) ) ;
    buf_clk new_AGEMA_reg_buffer_3243 ( .C (CLK), .D (new_AGEMA_signal_6010), .Q (new_AGEMA_signal_6011) ) ;
    buf_clk new_AGEMA_reg_buffer_3245 ( .C (CLK), .D (new_AGEMA_signal_6012), .Q (new_AGEMA_signal_6013) ) ;
    buf_clk new_AGEMA_reg_buffer_3247 ( .C (CLK), .D (new_AGEMA_signal_6014), .Q (new_AGEMA_signal_6015) ) ;
    buf_clk new_AGEMA_reg_buffer_3255 ( .C (CLK), .D (new_AGEMA_signal_6022), .Q (new_AGEMA_signal_6023) ) ;
    buf_clk new_AGEMA_reg_buffer_3259 ( .C (CLK), .D (new_AGEMA_signal_6026), .Q (new_AGEMA_signal_6027) ) ;
    buf_clk new_AGEMA_reg_buffer_3263 ( .C (CLK), .D (new_AGEMA_signal_6030), .Q (new_AGEMA_signal_6031) ) ;
    buf_clk new_AGEMA_reg_buffer_3273 ( .C (CLK), .D (new_AGEMA_signal_6040), .Q (new_AGEMA_signal_6041) ) ;
    buf_clk new_AGEMA_reg_buffer_3275 ( .C (CLK), .D (new_AGEMA_signal_6042), .Q (new_AGEMA_signal_6043) ) ;
    buf_clk new_AGEMA_reg_buffer_3277 ( .C (CLK), .D (new_AGEMA_signal_6044), .Q (new_AGEMA_signal_6045) ) ;
    buf_clk new_AGEMA_reg_buffer_3279 ( .C (CLK), .D (new_AGEMA_signal_6046), .Q (new_AGEMA_signal_6047) ) ;
    buf_clk new_AGEMA_reg_buffer_3281 ( .C (CLK), .D (new_AGEMA_signal_6048), .Q (new_AGEMA_signal_6049) ) ;
    buf_clk new_AGEMA_reg_buffer_3283 ( .C (CLK), .D (new_AGEMA_signal_6050), .Q (new_AGEMA_signal_6051) ) ;
    buf_clk new_AGEMA_reg_buffer_3291 ( .C (CLK), .D (new_AGEMA_signal_6058), .Q (new_AGEMA_signal_6059) ) ;
    buf_clk new_AGEMA_reg_buffer_3295 ( .C (CLK), .D (new_AGEMA_signal_6062), .Q (new_AGEMA_signal_6063) ) ;
    buf_clk new_AGEMA_reg_buffer_3299 ( .C (CLK), .D (new_AGEMA_signal_6066), .Q (new_AGEMA_signal_6067) ) ;
    buf_clk new_AGEMA_reg_buffer_3309 ( .C (CLK), .D (new_AGEMA_signal_6076), .Q (new_AGEMA_signal_6077) ) ;
    buf_clk new_AGEMA_reg_buffer_3311 ( .C (CLK), .D (new_AGEMA_signal_6078), .Q (new_AGEMA_signal_6079) ) ;
    buf_clk new_AGEMA_reg_buffer_3313 ( .C (CLK), .D (new_AGEMA_signal_6080), .Q (new_AGEMA_signal_6081) ) ;
    buf_clk new_AGEMA_reg_buffer_3315 ( .C (CLK), .D (new_AGEMA_signal_6082), .Q (new_AGEMA_signal_6083) ) ;
    buf_clk new_AGEMA_reg_buffer_3317 ( .C (CLK), .D (new_AGEMA_signal_6084), .Q (new_AGEMA_signal_6085) ) ;
    buf_clk new_AGEMA_reg_buffer_3319 ( .C (CLK), .D (new_AGEMA_signal_6086), .Q (new_AGEMA_signal_6087) ) ;
    buf_clk new_AGEMA_reg_buffer_3327 ( .C (CLK), .D (new_AGEMA_signal_6094), .Q (new_AGEMA_signal_6095) ) ;
    buf_clk new_AGEMA_reg_buffer_3331 ( .C (CLK), .D (new_AGEMA_signal_6098), .Q (new_AGEMA_signal_6099) ) ;
    buf_clk new_AGEMA_reg_buffer_3335 ( .C (CLK), .D (new_AGEMA_signal_6102), .Q (new_AGEMA_signal_6103) ) ;
    buf_clk new_AGEMA_reg_buffer_3339 ( .C (CLK), .D (new_AGEMA_signal_6106), .Q (new_AGEMA_signal_6107) ) ;
    buf_clk new_AGEMA_reg_buffer_3343 ( .C (CLK), .D (new_AGEMA_signal_6110), .Q (new_AGEMA_signal_6111) ) ;
    buf_clk new_AGEMA_reg_buffer_3347 ( .C (CLK), .D (new_AGEMA_signal_6114), .Q (new_AGEMA_signal_6115) ) ;
    buf_clk new_AGEMA_reg_buffer_3357 ( .C (CLK), .D (new_AGEMA_signal_6124), .Q (new_AGEMA_signal_6125) ) ;
    buf_clk new_AGEMA_reg_buffer_3359 ( .C (CLK), .D (new_AGEMA_signal_6126), .Q (new_AGEMA_signal_6127) ) ;
    buf_clk new_AGEMA_reg_buffer_3361 ( .C (CLK), .D (new_AGEMA_signal_6128), .Q (new_AGEMA_signal_6129) ) ;
    buf_clk new_AGEMA_reg_buffer_3363 ( .C (CLK), .D (new_AGEMA_signal_6130), .Q (new_AGEMA_signal_6131) ) ;
    buf_clk new_AGEMA_reg_buffer_3365 ( .C (CLK), .D (new_AGEMA_signal_6132), .Q (new_AGEMA_signal_6133) ) ;
    buf_clk new_AGEMA_reg_buffer_3367 ( .C (CLK), .D (new_AGEMA_signal_6134), .Q (new_AGEMA_signal_6135) ) ;
    buf_clk new_AGEMA_reg_buffer_3375 ( .C (CLK), .D (new_AGEMA_signal_6142), .Q (new_AGEMA_signal_6143) ) ;
    buf_clk new_AGEMA_reg_buffer_3379 ( .C (CLK), .D (new_AGEMA_signal_6146), .Q (new_AGEMA_signal_6147) ) ;
    buf_clk new_AGEMA_reg_buffer_3383 ( .C (CLK), .D (new_AGEMA_signal_6150), .Q (new_AGEMA_signal_6151) ) ;
    buf_clk new_AGEMA_reg_buffer_3387 ( .C (CLK), .D (new_AGEMA_signal_6154), .Q (new_AGEMA_signal_6155) ) ;
    buf_clk new_AGEMA_reg_buffer_3391 ( .C (CLK), .D (new_AGEMA_signal_6158), .Q (new_AGEMA_signal_6159) ) ;
    buf_clk new_AGEMA_reg_buffer_3395 ( .C (CLK), .D (new_AGEMA_signal_6162), .Q (new_AGEMA_signal_6163) ) ;
    buf_clk new_AGEMA_reg_buffer_3405 ( .C (CLK), .D (new_AGEMA_signal_6172), .Q (new_AGEMA_signal_6173) ) ;
    buf_clk new_AGEMA_reg_buffer_3407 ( .C (CLK), .D (new_AGEMA_signal_6174), .Q (new_AGEMA_signal_6175) ) ;
    buf_clk new_AGEMA_reg_buffer_3409 ( .C (CLK), .D (new_AGEMA_signal_6176), .Q (new_AGEMA_signal_6177) ) ;
    buf_clk new_AGEMA_reg_buffer_3411 ( .C (CLK), .D (new_AGEMA_signal_6178), .Q (new_AGEMA_signal_6179) ) ;
    buf_clk new_AGEMA_reg_buffer_3413 ( .C (CLK), .D (new_AGEMA_signal_6180), .Q (new_AGEMA_signal_6181) ) ;
    buf_clk new_AGEMA_reg_buffer_3415 ( .C (CLK), .D (new_AGEMA_signal_6182), .Q (new_AGEMA_signal_6183) ) ;
    buf_clk new_AGEMA_reg_buffer_3423 ( .C (CLK), .D (new_AGEMA_signal_6190), .Q (new_AGEMA_signal_6191) ) ;
    buf_clk new_AGEMA_reg_buffer_3427 ( .C (CLK), .D (new_AGEMA_signal_6194), .Q (new_AGEMA_signal_6195) ) ;
    buf_clk new_AGEMA_reg_buffer_3431 ( .C (CLK), .D (new_AGEMA_signal_6198), .Q (new_AGEMA_signal_6199) ) ;
    buf_clk new_AGEMA_reg_buffer_3441 ( .C (CLK), .D (new_AGEMA_signal_6208), .Q (new_AGEMA_signal_6209) ) ;
    buf_clk new_AGEMA_reg_buffer_3443 ( .C (CLK), .D (new_AGEMA_signal_6210), .Q (new_AGEMA_signal_6211) ) ;
    buf_clk new_AGEMA_reg_buffer_3445 ( .C (CLK), .D (new_AGEMA_signal_6212), .Q (new_AGEMA_signal_6213) ) ;
    buf_clk new_AGEMA_reg_buffer_3447 ( .C (CLK), .D (new_AGEMA_signal_6214), .Q (new_AGEMA_signal_6215) ) ;
    buf_clk new_AGEMA_reg_buffer_3449 ( .C (CLK), .D (new_AGEMA_signal_6216), .Q (new_AGEMA_signal_6217) ) ;
    buf_clk new_AGEMA_reg_buffer_3451 ( .C (CLK), .D (new_AGEMA_signal_6218), .Q (new_AGEMA_signal_6219) ) ;
    buf_clk new_AGEMA_reg_buffer_3459 ( .C (CLK), .D (new_AGEMA_signal_6226), .Q (new_AGEMA_signal_6227) ) ;
    buf_clk new_AGEMA_reg_buffer_3463 ( .C (CLK), .D (new_AGEMA_signal_6230), .Q (new_AGEMA_signal_6231) ) ;
    buf_clk new_AGEMA_reg_buffer_3467 ( .C (CLK), .D (new_AGEMA_signal_6234), .Q (new_AGEMA_signal_6235) ) ;
    buf_clk new_AGEMA_reg_buffer_3477 ( .C (CLK), .D (new_AGEMA_signal_6244), .Q (new_AGEMA_signal_6245) ) ;
    buf_clk new_AGEMA_reg_buffer_3479 ( .C (CLK), .D (new_AGEMA_signal_6246), .Q (new_AGEMA_signal_6247) ) ;
    buf_clk new_AGEMA_reg_buffer_3481 ( .C (CLK), .D (new_AGEMA_signal_6248), .Q (new_AGEMA_signal_6249) ) ;
    buf_clk new_AGEMA_reg_buffer_3483 ( .C (CLK), .D (new_AGEMA_signal_6250), .Q (new_AGEMA_signal_6251) ) ;
    buf_clk new_AGEMA_reg_buffer_3485 ( .C (CLK), .D (new_AGEMA_signal_6252), .Q (new_AGEMA_signal_6253) ) ;
    buf_clk new_AGEMA_reg_buffer_3487 ( .C (CLK), .D (new_AGEMA_signal_6254), .Q (new_AGEMA_signal_6255) ) ;
    buf_clk new_AGEMA_reg_buffer_3495 ( .C (CLK), .D (new_AGEMA_signal_6262), .Q (new_AGEMA_signal_6263) ) ;
    buf_clk new_AGEMA_reg_buffer_3499 ( .C (CLK), .D (new_AGEMA_signal_6266), .Q (new_AGEMA_signal_6267) ) ;
    buf_clk new_AGEMA_reg_buffer_3503 ( .C (CLK), .D (new_AGEMA_signal_6270), .Q (new_AGEMA_signal_6271) ) ;
    buf_clk new_AGEMA_reg_buffer_3507 ( .C (CLK), .D (new_AGEMA_signal_6274), .Q (new_AGEMA_signal_6275) ) ;
    buf_clk new_AGEMA_reg_buffer_3511 ( .C (CLK), .D (new_AGEMA_signal_6278), .Q (new_AGEMA_signal_6279) ) ;
    buf_clk new_AGEMA_reg_buffer_3515 ( .C (CLK), .D (new_AGEMA_signal_6282), .Q (new_AGEMA_signal_6283) ) ;
    buf_clk new_AGEMA_reg_buffer_3525 ( .C (CLK), .D (new_AGEMA_signal_6292), .Q (new_AGEMA_signal_6293) ) ;
    buf_clk new_AGEMA_reg_buffer_3527 ( .C (CLK), .D (new_AGEMA_signal_6294), .Q (new_AGEMA_signal_6295) ) ;
    buf_clk new_AGEMA_reg_buffer_3529 ( .C (CLK), .D (new_AGEMA_signal_6296), .Q (new_AGEMA_signal_6297) ) ;
    buf_clk new_AGEMA_reg_buffer_3531 ( .C (CLK), .D (new_AGEMA_signal_6298), .Q (new_AGEMA_signal_6299) ) ;
    buf_clk new_AGEMA_reg_buffer_3533 ( .C (CLK), .D (new_AGEMA_signal_6300), .Q (new_AGEMA_signal_6301) ) ;
    buf_clk new_AGEMA_reg_buffer_3535 ( .C (CLK), .D (new_AGEMA_signal_6302), .Q (new_AGEMA_signal_6303) ) ;
    buf_clk new_AGEMA_reg_buffer_3543 ( .C (CLK), .D (new_AGEMA_signal_6310), .Q (new_AGEMA_signal_6311) ) ;
    buf_clk new_AGEMA_reg_buffer_3547 ( .C (CLK), .D (new_AGEMA_signal_6314), .Q (new_AGEMA_signal_6315) ) ;
    buf_clk new_AGEMA_reg_buffer_3551 ( .C (CLK), .D (new_AGEMA_signal_6318), .Q (new_AGEMA_signal_6319) ) ;
    buf_clk new_AGEMA_reg_buffer_3555 ( .C (CLK), .D (new_AGEMA_signal_6322), .Q (new_AGEMA_signal_6323) ) ;
    buf_clk new_AGEMA_reg_buffer_3559 ( .C (CLK), .D (new_AGEMA_signal_6326), .Q (new_AGEMA_signal_6327) ) ;
    buf_clk new_AGEMA_reg_buffer_3563 ( .C (CLK), .D (new_AGEMA_signal_6330), .Q (new_AGEMA_signal_6331) ) ;
    buf_clk new_AGEMA_reg_buffer_3573 ( .C (CLK), .D (new_AGEMA_signal_6340), .Q (new_AGEMA_signal_6341) ) ;
    buf_clk new_AGEMA_reg_buffer_3575 ( .C (CLK), .D (new_AGEMA_signal_6342), .Q (new_AGEMA_signal_6343) ) ;
    buf_clk new_AGEMA_reg_buffer_3577 ( .C (CLK), .D (new_AGEMA_signal_6344), .Q (new_AGEMA_signal_6345) ) ;
    buf_clk new_AGEMA_reg_buffer_3579 ( .C (CLK), .D (new_AGEMA_signal_6346), .Q (new_AGEMA_signal_6347) ) ;
    buf_clk new_AGEMA_reg_buffer_3581 ( .C (CLK), .D (new_AGEMA_signal_6348), .Q (new_AGEMA_signal_6349) ) ;
    buf_clk new_AGEMA_reg_buffer_3583 ( .C (CLK), .D (new_AGEMA_signal_6350), .Q (new_AGEMA_signal_6351) ) ;
    buf_clk new_AGEMA_reg_buffer_3591 ( .C (CLK), .D (new_AGEMA_signal_6358), .Q (new_AGEMA_signal_6359) ) ;
    buf_clk new_AGEMA_reg_buffer_3595 ( .C (CLK), .D (new_AGEMA_signal_6362), .Q (new_AGEMA_signal_6363) ) ;
    buf_clk new_AGEMA_reg_buffer_3599 ( .C (CLK), .D (new_AGEMA_signal_6366), .Q (new_AGEMA_signal_6367) ) ;
    buf_clk new_AGEMA_reg_buffer_3609 ( .C (CLK), .D (new_AGEMA_signal_6376), .Q (new_AGEMA_signal_6377) ) ;
    buf_clk new_AGEMA_reg_buffer_3611 ( .C (CLK), .D (new_AGEMA_signal_6378), .Q (new_AGEMA_signal_6379) ) ;
    buf_clk new_AGEMA_reg_buffer_3613 ( .C (CLK), .D (new_AGEMA_signal_6380), .Q (new_AGEMA_signal_6381) ) ;
    buf_clk new_AGEMA_reg_buffer_3615 ( .C (CLK), .D (new_AGEMA_signal_6382), .Q (new_AGEMA_signal_6383) ) ;
    buf_clk new_AGEMA_reg_buffer_3617 ( .C (CLK), .D (new_AGEMA_signal_6384), .Q (new_AGEMA_signal_6385) ) ;
    buf_clk new_AGEMA_reg_buffer_3619 ( .C (CLK), .D (new_AGEMA_signal_6386), .Q (new_AGEMA_signal_6387) ) ;
    buf_clk new_AGEMA_reg_buffer_3627 ( .C (CLK), .D (new_AGEMA_signal_6394), .Q (new_AGEMA_signal_6395) ) ;
    buf_clk new_AGEMA_reg_buffer_3631 ( .C (CLK), .D (new_AGEMA_signal_6398), .Q (new_AGEMA_signal_6399) ) ;
    buf_clk new_AGEMA_reg_buffer_3635 ( .C (CLK), .D (new_AGEMA_signal_6402), .Q (new_AGEMA_signal_6403) ) ;
    buf_clk new_AGEMA_reg_buffer_3741 ( .C (CLK), .D (new_AGEMA_signal_6508), .Q (new_AGEMA_signal_6509) ) ;
    buf_clk new_AGEMA_reg_buffer_3745 ( .C (CLK), .D (new_AGEMA_signal_6512), .Q (new_AGEMA_signal_6513) ) ;
    buf_clk new_AGEMA_reg_buffer_3749 ( .C (CLK), .D (new_AGEMA_signal_6516), .Q (new_AGEMA_signal_6517) ) ;
    buf_clk new_AGEMA_reg_buffer_3753 ( .C (CLK), .D (new_AGEMA_signal_6520), .Q (new_AGEMA_signal_6521) ) ;
    buf_clk new_AGEMA_reg_buffer_3757 ( .C (CLK), .D (new_AGEMA_signal_6524), .Q (new_AGEMA_signal_6525) ) ;
    buf_clk new_AGEMA_reg_buffer_3761 ( .C (CLK), .D (new_AGEMA_signal_6528), .Q (new_AGEMA_signal_6529) ) ;
    buf_clk new_AGEMA_reg_buffer_3765 ( .C (CLK), .D (new_AGEMA_signal_6532), .Q (new_AGEMA_signal_6533) ) ;
    buf_clk new_AGEMA_reg_buffer_3769 ( .C (CLK), .D (new_AGEMA_signal_6536), .Q (new_AGEMA_signal_6537) ) ;
    buf_clk new_AGEMA_reg_buffer_3773 ( .C (CLK), .D (new_AGEMA_signal_6540), .Q (new_AGEMA_signal_6541) ) ;
    buf_clk new_AGEMA_reg_buffer_3777 ( .C (CLK), .D (new_AGEMA_signal_6544), .Q (new_AGEMA_signal_6545) ) ;
    buf_clk new_AGEMA_reg_buffer_3781 ( .C (CLK), .D (new_AGEMA_signal_6548), .Q (new_AGEMA_signal_6549) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_1418 ( .C (CLK), .D (new_AGEMA_signal_4185), .Q (new_AGEMA_signal_4186) ) ;
    buf_clk new_AGEMA_reg_buffer_1422 ( .C (CLK), .D (new_AGEMA_signal_4189), .Q (new_AGEMA_signal_4190) ) ;
    buf_clk new_AGEMA_reg_buffer_1426 ( .C (CLK), .D (new_AGEMA_signal_4193), .Q (new_AGEMA_signal_4194) ) ;
    buf_clk new_AGEMA_reg_buffer_1430 ( .C (CLK), .D (new_AGEMA_signal_4197), .Q (new_AGEMA_signal_4198) ) ;
    buf_clk new_AGEMA_reg_buffer_1434 ( .C (CLK), .D (new_AGEMA_signal_4201), .Q (new_AGEMA_signal_4202) ) ;
    buf_clk new_AGEMA_reg_buffer_1438 ( .C (CLK), .D (new_AGEMA_signal_4205), .Q (new_AGEMA_signal_4206) ) ;
    buf_clk new_AGEMA_reg_buffer_1442 ( .C (CLK), .D (new_AGEMA_signal_4209), .Q (new_AGEMA_signal_4210) ) ;
    buf_clk new_AGEMA_reg_buffer_1446 ( .C (CLK), .D (new_AGEMA_signal_4213), .Q (new_AGEMA_signal_4214) ) ;
    buf_clk new_AGEMA_reg_buffer_1450 ( .C (CLK), .D (new_AGEMA_signal_4217), .Q (new_AGEMA_signal_4218) ) ;
    buf_clk new_AGEMA_reg_buffer_1454 ( .C (CLK), .D (new_AGEMA_signal_4221), .Q (new_AGEMA_signal_4222) ) ;
    buf_clk new_AGEMA_reg_buffer_1458 ( .C (CLK), .D (new_AGEMA_signal_4225), .Q (new_AGEMA_signal_4226) ) ;
    buf_clk new_AGEMA_reg_buffer_1462 ( .C (CLK), .D (new_AGEMA_signal_4229), .Q (new_AGEMA_signal_4230) ) ;
    buf_clk new_AGEMA_reg_buffer_1466 ( .C (CLK), .D (new_AGEMA_signal_4233), .Q (new_AGEMA_signal_4234) ) ;
    buf_clk new_AGEMA_reg_buffer_1470 ( .C (CLK), .D (new_AGEMA_signal_4237), .Q (new_AGEMA_signal_4238) ) ;
    buf_clk new_AGEMA_reg_buffer_1474 ( .C (CLK), .D (new_AGEMA_signal_4241), .Q (new_AGEMA_signal_4242) ) ;
    buf_clk new_AGEMA_reg_buffer_1478 ( .C (CLK), .D (new_AGEMA_signal_4245), .Q (new_AGEMA_signal_4246) ) ;
    buf_clk new_AGEMA_reg_buffer_1482 ( .C (CLK), .D (new_AGEMA_signal_4249), .Q (new_AGEMA_signal_4250) ) ;
    buf_clk new_AGEMA_reg_buffer_1486 ( .C (CLK), .D (new_AGEMA_signal_4253), .Q (new_AGEMA_signal_4254) ) ;
    buf_clk new_AGEMA_reg_buffer_1490 ( .C (CLK), .D (new_AGEMA_signal_4257), .Q (new_AGEMA_signal_4258) ) ;
    buf_clk new_AGEMA_reg_buffer_1494 ( .C (CLK), .D (new_AGEMA_signal_4261), .Q (new_AGEMA_signal_4262) ) ;
    buf_clk new_AGEMA_reg_buffer_1498 ( .C (CLK), .D (new_AGEMA_signal_4265), .Q (new_AGEMA_signal_4266) ) ;
    buf_clk new_AGEMA_reg_buffer_1502 ( .C (CLK), .D (new_AGEMA_signal_4269), .Q (new_AGEMA_signal_4270) ) ;
    buf_clk new_AGEMA_reg_buffer_1506 ( .C (CLK), .D (new_AGEMA_signal_4273), .Q (new_AGEMA_signal_4274) ) ;
    buf_clk new_AGEMA_reg_buffer_1510 ( .C (CLK), .D (new_AGEMA_signal_4277), .Q (new_AGEMA_signal_4278) ) ;
    buf_clk new_AGEMA_reg_buffer_1514 ( .C (CLK), .D (new_AGEMA_signal_4281), .Q (new_AGEMA_signal_4282) ) ;
    buf_clk new_AGEMA_reg_buffer_1518 ( .C (CLK), .D (new_AGEMA_signal_4285), .Q (new_AGEMA_signal_4286) ) ;
    buf_clk new_AGEMA_reg_buffer_1522 ( .C (CLK), .D (new_AGEMA_signal_4289), .Q (new_AGEMA_signal_4290) ) ;
    buf_clk new_AGEMA_reg_buffer_1526 ( .C (CLK), .D (new_AGEMA_signal_4293), .Q (new_AGEMA_signal_4294) ) ;
    buf_clk new_AGEMA_reg_buffer_1530 ( .C (CLK), .D (new_AGEMA_signal_4297), .Q (new_AGEMA_signal_4298) ) ;
    buf_clk new_AGEMA_reg_buffer_1534 ( .C (CLK), .D (new_AGEMA_signal_4301), .Q (new_AGEMA_signal_4302) ) ;
    buf_clk new_AGEMA_reg_buffer_1538 ( .C (CLK), .D (new_AGEMA_signal_4305), .Q (new_AGEMA_signal_4306) ) ;
    buf_clk new_AGEMA_reg_buffer_1542 ( .C (CLK), .D (new_AGEMA_signal_4309), .Q (new_AGEMA_signal_4310) ) ;
    buf_clk new_AGEMA_reg_buffer_1546 ( .C (CLK), .D (new_AGEMA_signal_4313), .Q (new_AGEMA_signal_4314) ) ;
    buf_clk new_AGEMA_reg_buffer_1550 ( .C (CLK), .D (new_AGEMA_signal_4317), .Q (new_AGEMA_signal_4318) ) ;
    buf_clk new_AGEMA_reg_buffer_1554 ( .C (CLK), .D (new_AGEMA_signal_4321), .Q (new_AGEMA_signal_4322) ) ;
    buf_clk new_AGEMA_reg_buffer_1558 ( .C (CLK), .D (new_AGEMA_signal_4325), .Q (new_AGEMA_signal_4326) ) ;
    buf_clk new_AGEMA_reg_buffer_1562 ( .C (CLK), .D (new_AGEMA_signal_4329), .Q (new_AGEMA_signal_4330) ) ;
    buf_clk new_AGEMA_reg_buffer_1566 ( .C (CLK), .D (new_AGEMA_signal_4333), .Q (new_AGEMA_signal_4334) ) ;
    buf_clk new_AGEMA_reg_buffer_1570 ( .C (CLK), .D (new_AGEMA_signal_4337), .Q (new_AGEMA_signal_4338) ) ;
    buf_clk new_AGEMA_reg_buffer_1574 ( .C (CLK), .D (new_AGEMA_signal_4341), .Q (new_AGEMA_signal_4342) ) ;
    buf_clk new_AGEMA_reg_buffer_1578 ( .C (CLK), .D (new_AGEMA_signal_4345), .Q (new_AGEMA_signal_4346) ) ;
    buf_clk new_AGEMA_reg_buffer_1582 ( .C (CLK), .D (new_AGEMA_signal_4349), .Q (new_AGEMA_signal_4350) ) ;
    buf_clk new_AGEMA_reg_buffer_1586 ( .C (CLK), .D (new_AGEMA_signal_4353), .Q (new_AGEMA_signal_4354) ) ;
    buf_clk new_AGEMA_reg_buffer_1590 ( .C (CLK), .D (new_AGEMA_signal_4357), .Q (new_AGEMA_signal_4358) ) ;
    buf_clk new_AGEMA_reg_buffer_1594 ( .C (CLK), .D (new_AGEMA_signal_4361), .Q (new_AGEMA_signal_4362) ) ;
    buf_clk new_AGEMA_reg_buffer_1598 ( .C (CLK), .D (new_AGEMA_signal_4365), .Q (new_AGEMA_signal_4366) ) ;
    buf_clk new_AGEMA_reg_buffer_1602 ( .C (CLK), .D (new_AGEMA_signal_4369), .Q (new_AGEMA_signal_4370) ) ;
    buf_clk new_AGEMA_reg_buffer_1606 ( .C (CLK), .D (new_AGEMA_signal_4373), .Q (new_AGEMA_signal_4374) ) ;
    buf_clk new_AGEMA_reg_buffer_1610 ( .C (CLK), .D (new_AGEMA_signal_4377), .Q (new_AGEMA_signal_4378) ) ;
    buf_clk new_AGEMA_reg_buffer_1614 ( .C (CLK), .D (new_AGEMA_signal_4381), .Q (new_AGEMA_signal_4382) ) ;
    buf_clk new_AGEMA_reg_buffer_1618 ( .C (CLK), .D (new_AGEMA_signal_4385), .Q (new_AGEMA_signal_4386) ) ;
    buf_clk new_AGEMA_reg_buffer_1622 ( .C (CLK), .D (new_AGEMA_signal_4389), .Q (new_AGEMA_signal_4390) ) ;
    buf_clk new_AGEMA_reg_buffer_1626 ( .C (CLK), .D (new_AGEMA_signal_4393), .Q (new_AGEMA_signal_4394) ) ;
    buf_clk new_AGEMA_reg_buffer_1630 ( .C (CLK), .D (new_AGEMA_signal_4397), .Q (new_AGEMA_signal_4398) ) ;
    buf_clk new_AGEMA_reg_buffer_1634 ( .C (CLK), .D (new_AGEMA_signal_4401), .Q (new_AGEMA_signal_4402) ) ;
    buf_clk new_AGEMA_reg_buffer_1638 ( .C (CLK), .D (new_AGEMA_signal_4405), .Q (new_AGEMA_signal_4406) ) ;
    buf_clk new_AGEMA_reg_buffer_1642 ( .C (CLK), .D (new_AGEMA_signal_4409), .Q (new_AGEMA_signal_4410) ) ;
    buf_clk new_AGEMA_reg_buffer_1646 ( .C (CLK), .D (new_AGEMA_signal_4413), .Q (new_AGEMA_signal_4414) ) ;
    buf_clk new_AGEMA_reg_buffer_1650 ( .C (CLK), .D (new_AGEMA_signal_4417), .Q (new_AGEMA_signal_4418) ) ;
    buf_clk new_AGEMA_reg_buffer_1654 ( .C (CLK), .D (new_AGEMA_signal_4421), .Q (new_AGEMA_signal_4422) ) ;
    buf_clk new_AGEMA_reg_buffer_1658 ( .C (CLK), .D (new_AGEMA_signal_4425), .Q (new_AGEMA_signal_4426) ) ;
    buf_clk new_AGEMA_reg_buffer_1662 ( .C (CLK), .D (new_AGEMA_signal_4429), .Q (new_AGEMA_signal_4430) ) ;
    buf_clk new_AGEMA_reg_buffer_1666 ( .C (CLK), .D (new_AGEMA_signal_4433), .Q (new_AGEMA_signal_4434) ) ;
    buf_clk new_AGEMA_reg_buffer_1670 ( .C (CLK), .D (new_AGEMA_signal_4437), .Q (new_AGEMA_signal_4438) ) ;
    buf_clk new_AGEMA_reg_buffer_1674 ( .C (CLK), .D (new_AGEMA_signal_4441), .Q (new_AGEMA_signal_4442) ) ;
    buf_clk new_AGEMA_reg_buffer_1678 ( .C (CLK), .D (new_AGEMA_signal_4445), .Q (new_AGEMA_signal_4446) ) ;
    buf_clk new_AGEMA_reg_buffer_1682 ( .C (CLK), .D (new_AGEMA_signal_4449), .Q (new_AGEMA_signal_4450) ) ;
    buf_clk new_AGEMA_reg_buffer_1686 ( .C (CLK), .D (new_AGEMA_signal_4453), .Q (new_AGEMA_signal_4454) ) ;
    buf_clk new_AGEMA_reg_buffer_1690 ( .C (CLK), .D (new_AGEMA_signal_4457), .Q (new_AGEMA_signal_4458) ) ;
    buf_clk new_AGEMA_reg_buffer_1694 ( .C (CLK), .D (new_AGEMA_signal_4461), .Q (new_AGEMA_signal_4462) ) ;
    buf_clk new_AGEMA_reg_buffer_1698 ( .C (CLK), .D (new_AGEMA_signal_4465), .Q (new_AGEMA_signal_4466) ) ;
    buf_clk new_AGEMA_reg_buffer_1702 ( .C (CLK), .D (new_AGEMA_signal_4469), .Q (new_AGEMA_signal_4470) ) ;
    buf_clk new_AGEMA_reg_buffer_1706 ( .C (CLK), .D (new_AGEMA_signal_4473), .Q (new_AGEMA_signal_4474) ) ;
    buf_clk new_AGEMA_reg_buffer_1710 ( .C (CLK), .D (new_AGEMA_signal_4477), .Q (new_AGEMA_signal_4478) ) ;
    buf_clk new_AGEMA_reg_buffer_1714 ( .C (CLK), .D (new_AGEMA_signal_4481), .Q (new_AGEMA_signal_4482) ) ;
    buf_clk new_AGEMA_reg_buffer_1718 ( .C (CLK), .D (new_AGEMA_signal_4485), .Q (new_AGEMA_signal_4486) ) ;
    buf_clk new_AGEMA_reg_buffer_1722 ( .C (CLK), .D (new_AGEMA_signal_4489), .Q (new_AGEMA_signal_4490) ) ;
    buf_clk new_AGEMA_reg_buffer_1726 ( .C (CLK), .D (new_AGEMA_signal_4493), .Q (new_AGEMA_signal_4494) ) ;
    buf_clk new_AGEMA_reg_buffer_1730 ( .C (CLK), .D (new_AGEMA_signal_4497), .Q (new_AGEMA_signal_4498) ) ;
    buf_clk new_AGEMA_reg_buffer_1734 ( .C (CLK), .D (new_AGEMA_signal_4501), .Q (new_AGEMA_signal_4502) ) ;
    buf_clk new_AGEMA_reg_buffer_1738 ( .C (CLK), .D (new_AGEMA_signal_4505), .Q (new_AGEMA_signal_4506) ) ;
    buf_clk new_AGEMA_reg_buffer_1742 ( .C (CLK), .D (new_AGEMA_signal_4509), .Q (new_AGEMA_signal_4510) ) ;
    buf_clk new_AGEMA_reg_buffer_1746 ( .C (CLK), .D (new_AGEMA_signal_4513), .Q (new_AGEMA_signal_4514) ) ;
    buf_clk new_AGEMA_reg_buffer_1750 ( .C (CLK), .D (new_AGEMA_signal_4517), .Q (new_AGEMA_signal_4518) ) ;
    buf_clk new_AGEMA_reg_buffer_1754 ( .C (CLK), .D (new_AGEMA_signal_4521), .Q (new_AGEMA_signal_4522) ) ;
    buf_clk new_AGEMA_reg_buffer_1758 ( .C (CLK), .D (new_AGEMA_signal_4525), .Q (new_AGEMA_signal_4526) ) ;
    buf_clk new_AGEMA_reg_buffer_1762 ( .C (CLK), .D (new_AGEMA_signal_4529), .Q (new_AGEMA_signal_4530) ) ;
    buf_clk new_AGEMA_reg_buffer_1766 ( .C (CLK), .D (new_AGEMA_signal_4533), .Q (new_AGEMA_signal_4534) ) ;
    buf_clk new_AGEMA_reg_buffer_1770 ( .C (CLK), .D (new_AGEMA_signal_4537), .Q (new_AGEMA_signal_4538) ) ;
    buf_clk new_AGEMA_reg_buffer_1774 ( .C (CLK), .D (new_AGEMA_signal_4541), .Q (new_AGEMA_signal_4542) ) ;
    buf_clk new_AGEMA_reg_buffer_1778 ( .C (CLK), .D (new_AGEMA_signal_4545), .Q (new_AGEMA_signal_4546) ) ;
    buf_clk new_AGEMA_reg_buffer_1782 ( .C (CLK), .D (new_AGEMA_signal_4549), .Q (new_AGEMA_signal_4550) ) ;
    buf_clk new_AGEMA_reg_buffer_1786 ( .C (CLK), .D (new_AGEMA_signal_4553), .Q (new_AGEMA_signal_4554) ) ;
    buf_clk new_AGEMA_reg_buffer_1790 ( .C (CLK), .D (new_AGEMA_signal_4557), .Q (new_AGEMA_signal_4558) ) ;
    buf_clk new_AGEMA_reg_buffer_1794 ( .C (CLK), .D (new_AGEMA_signal_4561), .Q (new_AGEMA_signal_4562) ) ;
    buf_clk new_AGEMA_reg_buffer_1798 ( .C (CLK), .D (new_AGEMA_signal_4565), .Q (new_AGEMA_signal_4566) ) ;
    buf_clk new_AGEMA_reg_buffer_1802 ( .C (CLK), .D (new_AGEMA_signal_4569), .Q (new_AGEMA_signal_4570) ) ;
    buf_clk new_AGEMA_reg_buffer_1806 ( .C (CLK), .D (new_AGEMA_signal_4573), .Q (new_AGEMA_signal_4574) ) ;
    buf_clk new_AGEMA_reg_buffer_1810 ( .C (CLK), .D (new_AGEMA_signal_4577), .Q (new_AGEMA_signal_4578) ) ;
    buf_clk new_AGEMA_reg_buffer_1814 ( .C (CLK), .D (new_AGEMA_signal_4581), .Q (new_AGEMA_signal_4582) ) ;
    buf_clk new_AGEMA_reg_buffer_1818 ( .C (CLK), .D (new_AGEMA_signal_4585), .Q (new_AGEMA_signal_4586) ) ;
    buf_clk new_AGEMA_reg_buffer_1822 ( .C (CLK), .D (new_AGEMA_signal_4589), .Q (new_AGEMA_signal_4590) ) ;
    buf_clk new_AGEMA_reg_buffer_1826 ( .C (CLK), .D (new_AGEMA_signal_4593), .Q (new_AGEMA_signal_4594) ) ;
    buf_clk new_AGEMA_reg_buffer_1830 ( .C (CLK), .D (new_AGEMA_signal_4597), .Q (new_AGEMA_signal_4598) ) ;
    buf_clk new_AGEMA_reg_buffer_1834 ( .C (CLK), .D (new_AGEMA_signal_4601), .Q (new_AGEMA_signal_4602) ) ;
    buf_clk new_AGEMA_reg_buffer_1838 ( .C (CLK), .D (new_AGEMA_signal_4605), .Q (new_AGEMA_signal_4606) ) ;
    buf_clk new_AGEMA_reg_buffer_1842 ( .C (CLK), .D (new_AGEMA_signal_4609), .Q (new_AGEMA_signal_4610) ) ;
    buf_clk new_AGEMA_reg_buffer_1846 ( .C (CLK), .D (new_AGEMA_signal_4613), .Q (new_AGEMA_signal_4614) ) ;
    buf_clk new_AGEMA_reg_buffer_1850 ( .C (CLK), .D (new_AGEMA_signal_4617), .Q (new_AGEMA_signal_4618) ) ;
    buf_clk new_AGEMA_reg_buffer_1854 ( .C (CLK), .D (new_AGEMA_signal_4621), .Q (new_AGEMA_signal_4622) ) ;
    buf_clk new_AGEMA_reg_buffer_1858 ( .C (CLK), .D (new_AGEMA_signal_4625), .Q (new_AGEMA_signal_4626) ) ;
    buf_clk new_AGEMA_reg_buffer_1862 ( .C (CLK), .D (new_AGEMA_signal_4629), .Q (new_AGEMA_signal_4630) ) ;
    buf_clk new_AGEMA_reg_buffer_1866 ( .C (CLK), .D (new_AGEMA_signal_4633), .Q (new_AGEMA_signal_4634) ) ;
    buf_clk new_AGEMA_reg_buffer_1870 ( .C (CLK), .D (new_AGEMA_signal_4637), .Q (new_AGEMA_signal_4638) ) ;
    buf_clk new_AGEMA_reg_buffer_1874 ( .C (CLK), .D (new_AGEMA_signal_4641), .Q (new_AGEMA_signal_4642) ) ;
    buf_clk new_AGEMA_reg_buffer_1878 ( .C (CLK), .D (new_AGEMA_signal_4645), .Q (new_AGEMA_signal_4646) ) ;
    buf_clk new_AGEMA_reg_buffer_1882 ( .C (CLK), .D (new_AGEMA_signal_4649), .Q (new_AGEMA_signal_4650) ) ;
    buf_clk new_AGEMA_reg_buffer_1886 ( .C (CLK), .D (new_AGEMA_signal_4653), .Q (new_AGEMA_signal_4654) ) ;
    buf_clk new_AGEMA_reg_buffer_1890 ( .C (CLK), .D (new_AGEMA_signal_4657), .Q (new_AGEMA_signal_4658) ) ;
    buf_clk new_AGEMA_reg_buffer_1894 ( .C (CLK), .D (new_AGEMA_signal_4661), .Q (new_AGEMA_signal_4662) ) ;
    buf_clk new_AGEMA_reg_buffer_1898 ( .C (CLK), .D (new_AGEMA_signal_4665), .Q (new_AGEMA_signal_4666) ) ;
    buf_clk new_AGEMA_reg_buffer_1902 ( .C (CLK), .D (new_AGEMA_signal_4669), .Q (new_AGEMA_signal_4670) ) ;
    buf_clk new_AGEMA_reg_buffer_1906 ( .C (CLK), .D (new_AGEMA_signal_4673), .Q (new_AGEMA_signal_4674) ) ;
    buf_clk new_AGEMA_reg_buffer_1910 ( .C (CLK), .D (new_AGEMA_signal_4677), .Q (new_AGEMA_signal_4678) ) ;
    buf_clk new_AGEMA_reg_buffer_1914 ( .C (CLK), .D (new_AGEMA_signal_4681), .Q (new_AGEMA_signal_4682) ) ;
    buf_clk new_AGEMA_reg_buffer_1918 ( .C (CLK), .D (new_AGEMA_signal_4685), .Q (new_AGEMA_signal_4686) ) ;
    buf_clk new_AGEMA_reg_buffer_1922 ( .C (CLK), .D (new_AGEMA_signal_4689), .Q (new_AGEMA_signal_4690) ) ;
    buf_clk new_AGEMA_reg_buffer_1926 ( .C (CLK), .D (new_AGEMA_signal_4693), .Q (new_AGEMA_signal_4694) ) ;
    buf_clk new_AGEMA_reg_buffer_1930 ( .C (CLK), .D (new_AGEMA_signal_4697), .Q (new_AGEMA_signal_4698) ) ;
    buf_clk new_AGEMA_reg_buffer_1934 ( .C (CLK), .D (new_AGEMA_signal_4701), .Q (new_AGEMA_signal_4702) ) ;
    buf_clk new_AGEMA_reg_buffer_1938 ( .C (CLK), .D (new_AGEMA_signal_4705), .Q (new_AGEMA_signal_4706) ) ;
    buf_clk new_AGEMA_reg_buffer_1942 ( .C (CLK), .D (new_AGEMA_signal_4709), .Q (new_AGEMA_signal_4710) ) ;
    buf_clk new_AGEMA_reg_buffer_1946 ( .C (CLK), .D (new_AGEMA_signal_4713), .Q (new_AGEMA_signal_4714) ) ;
    buf_clk new_AGEMA_reg_buffer_1950 ( .C (CLK), .D (new_AGEMA_signal_4717), .Q (new_AGEMA_signal_4718) ) ;
    buf_clk new_AGEMA_reg_buffer_1954 ( .C (CLK), .D (new_AGEMA_signal_4721), .Q (new_AGEMA_signal_4722) ) ;
    buf_clk new_AGEMA_reg_buffer_1958 ( .C (CLK), .D (new_AGEMA_signal_4725), .Q (new_AGEMA_signal_4726) ) ;
    buf_clk new_AGEMA_reg_buffer_1962 ( .C (CLK), .D (new_AGEMA_signal_4729), .Q (new_AGEMA_signal_4730) ) ;
    buf_clk new_AGEMA_reg_buffer_1966 ( .C (CLK), .D (new_AGEMA_signal_4733), .Q (new_AGEMA_signal_4734) ) ;
    buf_clk new_AGEMA_reg_buffer_1970 ( .C (CLK), .D (new_AGEMA_signal_4737), .Q (new_AGEMA_signal_4738) ) ;
    buf_clk new_AGEMA_reg_buffer_1974 ( .C (CLK), .D (new_AGEMA_signal_4741), .Q (new_AGEMA_signal_4742) ) ;
    buf_clk new_AGEMA_reg_buffer_1978 ( .C (CLK), .D (new_AGEMA_signal_4745), .Q (new_AGEMA_signal_4746) ) ;
    buf_clk new_AGEMA_reg_buffer_1982 ( .C (CLK), .D (new_AGEMA_signal_4749), .Q (new_AGEMA_signal_4750) ) ;
    buf_clk new_AGEMA_reg_buffer_1986 ( .C (CLK), .D (new_AGEMA_signal_4753), .Q (new_AGEMA_signal_4754) ) ;
    buf_clk new_AGEMA_reg_buffer_1990 ( .C (CLK), .D (new_AGEMA_signal_4757), .Q (new_AGEMA_signal_4758) ) ;
    buf_clk new_AGEMA_reg_buffer_1994 ( .C (CLK), .D (new_AGEMA_signal_4761), .Q (new_AGEMA_signal_4762) ) ;
    buf_clk new_AGEMA_reg_buffer_1998 ( .C (CLK), .D (new_AGEMA_signal_4765), .Q (new_AGEMA_signal_4766) ) ;
    buf_clk new_AGEMA_reg_buffer_2002 ( .C (CLK), .D (new_AGEMA_signal_4769), .Q (new_AGEMA_signal_4770) ) ;
    buf_clk new_AGEMA_reg_buffer_2006 ( .C (CLK), .D (new_AGEMA_signal_4773), .Q (new_AGEMA_signal_4774) ) ;
    buf_clk new_AGEMA_reg_buffer_2010 ( .C (CLK), .D (new_AGEMA_signal_4777), .Q (new_AGEMA_signal_4778) ) ;
    buf_clk new_AGEMA_reg_buffer_2014 ( .C (CLK), .D (new_AGEMA_signal_4781), .Q (new_AGEMA_signal_4782) ) ;
    buf_clk new_AGEMA_reg_buffer_2018 ( .C (CLK), .D (new_AGEMA_signal_4785), .Q (new_AGEMA_signal_4786) ) ;
    buf_clk new_AGEMA_reg_buffer_2022 ( .C (CLK), .D (new_AGEMA_signal_4789), .Q (new_AGEMA_signal_4790) ) ;
    buf_clk new_AGEMA_reg_buffer_2026 ( .C (CLK), .D (new_AGEMA_signal_4793), .Q (new_AGEMA_signal_4794) ) ;
    buf_clk new_AGEMA_reg_buffer_2030 ( .C (CLK), .D (new_AGEMA_signal_4797), .Q (new_AGEMA_signal_4798) ) ;
    buf_clk new_AGEMA_reg_buffer_2034 ( .C (CLK), .D (new_AGEMA_signal_4801), .Q (new_AGEMA_signal_4802) ) ;
    buf_clk new_AGEMA_reg_buffer_2038 ( .C (CLK), .D (new_AGEMA_signal_4805), .Q (new_AGEMA_signal_4806) ) ;
    buf_clk new_AGEMA_reg_buffer_2042 ( .C (CLK), .D (new_AGEMA_signal_4809), .Q (new_AGEMA_signal_4810) ) ;
    buf_clk new_AGEMA_reg_buffer_2046 ( .C (CLK), .D (new_AGEMA_signal_4813), .Q (new_AGEMA_signal_4814) ) ;
    buf_clk new_AGEMA_reg_buffer_2050 ( .C (CLK), .D (new_AGEMA_signal_4817), .Q (new_AGEMA_signal_4818) ) ;
    buf_clk new_AGEMA_reg_buffer_2054 ( .C (CLK), .D (new_AGEMA_signal_4821), .Q (new_AGEMA_signal_4822) ) ;
    buf_clk new_AGEMA_reg_buffer_2058 ( .C (CLK), .D (new_AGEMA_signal_4825), .Q (new_AGEMA_signal_4826) ) ;
    buf_clk new_AGEMA_reg_buffer_2062 ( .C (CLK), .D (new_AGEMA_signal_4829), .Q (new_AGEMA_signal_4830) ) ;
    buf_clk new_AGEMA_reg_buffer_2066 ( .C (CLK), .D (new_AGEMA_signal_4833), .Q (new_AGEMA_signal_4834) ) ;
    buf_clk new_AGEMA_reg_buffer_2070 ( .C (CLK), .D (new_AGEMA_signal_4837), .Q (new_AGEMA_signal_4838) ) ;
    buf_clk new_AGEMA_reg_buffer_2074 ( .C (CLK), .D (new_AGEMA_signal_4841), .Q (new_AGEMA_signal_4842) ) ;
    buf_clk new_AGEMA_reg_buffer_2078 ( .C (CLK), .D (new_AGEMA_signal_4845), .Q (new_AGEMA_signal_4846) ) ;
    buf_clk new_AGEMA_reg_buffer_2082 ( .C (CLK), .D (new_AGEMA_signal_4849), .Q (new_AGEMA_signal_4850) ) ;
    buf_clk new_AGEMA_reg_buffer_2086 ( .C (CLK), .D (new_AGEMA_signal_4853), .Q (new_AGEMA_signal_4854) ) ;
    buf_clk new_AGEMA_reg_buffer_2090 ( .C (CLK), .D (new_AGEMA_signal_4857), .Q (new_AGEMA_signal_4858) ) ;
    buf_clk new_AGEMA_reg_buffer_2094 ( .C (CLK), .D (new_AGEMA_signal_4861), .Q (new_AGEMA_signal_4862) ) ;
    buf_clk new_AGEMA_reg_buffer_2098 ( .C (CLK), .D (new_AGEMA_signal_4865), .Q (new_AGEMA_signal_4866) ) ;
    buf_clk new_AGEMA_reg_buffer_2102 ( .C (CLK), .D (new_AGEMA_signal_4869), .Q (new_AGEMA_signal_4870) ) ;
    buf_clk new_AGEMA_reg_buffer_2106 ( .C (CLK), .D (new_AGEMA_signal_4873), .Q (new_AGEMA_signal_4874) ) ;
    buf_clk new_AGEMA_reg_buffer_2110 ( .C (CLK), .D (new_AGEMA_signal_4877), .Q (new_AGEMA_signal_4878) ) ;
    buf_clk new_AGEMA_reg_buffer_2114 ( .C (CLK), .D (new_AGEMA_signal_4881), .Q (new_AGEMA_signal_4882) ) ;
    buf_clk new_AGEMA_reg_buffer_2118 ( .C (CLK), .D (new_AGEMA_signal_4885), .Q (new_AGEMA_signal_4886) ) ;
    buf_clk new_AGEMA_reg_buffer_2122 ( .C (CLK), .D (new_AGEMA_signal_4889), .Q (new_AGEMA_signal_4890) ) ;
    buf_clk new_AGEMA_reg_buffer_2126 ( .C (CLK), .D (new_AGEMA_signal_4893), .Q (new_AGEMA_signal_4894) ) ;
    buf_clk new_AGEMA_reg_buffer_2130 ( .C (CLK), .D (new_AGEMA_signal_4897), .Q (new_AGEMA_signal_4898) ) ;
    buf_clk new_AGEMA_reg_buffer_2134 ( .C (CLK), .D (new_AGEMA_signal_4901), .Q (new_AGEMA_signal_4902) ) ;
    buf_clk new_AGEMA_reg_buffer_2138 ( .C (CLK), .D (new_AGEMA_signal_4905), .Q (new_AGEMA_signal_4906) ) ;
    buf_clk new_AGEMA_reg_buffer_2142 ( .C (CLK), .D (new_AGEMA_signal_4909), .Q (new_AGEMA_signal_4910) ) ;
    buf_clk new_AGEMA_reg_buffer_2146 ( .C (CLK), .D (new_AGEMA_signal_4913), .Q (new_AGEMA_signal_4914) ) ;
    buf_clk new_AGEMA_reg_buffer_2150 ( .C (CLK), .D (new_AGEMA_signal_4917), .Q (new_AGEMA_signal_4918) ) ;
    buf_clk new_AGEMA_reg_buffer_2154 ( .C (CLK), .D (new_AGEMA_signal_4921), .Q (new_AGEMA_signal_4922) ) ;
    buf_clk new_AGEMA_reg_buffer_2158 ( .C (CLK), .D (new_AGEMA_signal_4925), .Q (new_AGEMA_signal_4926) ) ;
    buf_clk new_AGEMA_reg_buffer_2162 ( .C (CLK), .D (new_AGEMA_signal_4929), .Q (new_AGEMA_signal_4930) ) ;
    buf_clk new_AGEMA_reg_buffer_2166 ( .C (CLK), .D (new_AGEMA_signal_4933), .Q (new_AGEMA_signal_4934) ) ;
    buf_clk new_AGEMA_reg_buffer_2170 ( .C (CLK), .D (new_AGEMA_signal_4937), .Q (new_AGEMA_signal_4938) ) ;
    buf_clk new_AGEMA_reg_buffer_2174 ( .C (CLK), .D (new_AGEMA_signal_4941), .Q (new_AGEMA_signal_4942) ) ;
    buf_clk new_AGEMA_reg_buffer_2178 ( .C (CLK), .D (new_AGEMA_signal_4945), .Q (new_AGEMA_signal_4946) ) ;
    buf_clk new_AGEMA_reg_buffer_2182 ( .C (CLK), .D (new_AGEMA_signal_4949), .Q (new_AGEMA_signal_4950) ) ;
    buf_clk new_AGEMA_reg_buffer_2186 ( .C (CLK), .D (new_AGEMA_signal_4953), .Q (new_AGEMA_signal_4954) ) ;
    buf_clk new_AGEMA_reg_buffer_2190 ( .C (CLK), .D (new_AGEMA_signal_4957), .Q (new_AGEMA_signal_4958) ) ;
    buf_clk new_AGEMA_reg_buffer_2194 ( .C (CLK), .D (new_AGEMA_signal_4961), .Q (new_AGEMA_signal_4962) ) ;
    buf_clk new_AGEMA_reg_buffer_2198 ( .C (CLK), .D (new_AGEMA_signal_4965), .Q (new_AGEMA_signal_4966) ) ;
    buf_clk new_AGEMA_reg_buffer_2202 ( .C (CLK), .D (new_AGEMA_signal_4969), .Q (new_AGEMA_signal_4970) ) ;
    buf_clk new_AGEMA_reg_buffer_2206 ( .C (CLK), .D (new_AGEMA_signal_4973), .Q (new_AGEMA_signal_4974) ) ;
    buf_clk new_AGEMA_reg_buffer_2210 ( .C (CLK), .D (new_AGEMA_signal_4977), .Q (new_AGEMA_signal_4978) ) ;
    buf_clk new_AGEMA_reg_buffer_2214 ( .C (CLK), .D (new_AGEMA_signal_4981), .Q (new_AGEMA_signal_4982) ) ;
    buf_clk new_AGEMA_reg_buffer_2218 ( .C (CLK), .D (new_AGEMA_signal_4985), .Q (new_AGEMA_signal_4986) ) ;
    buf_clk new_AGEMA_reg_buffer_2222 ( .C (CLK), .D (new_AGEMA_signal_4989), .Q (new_AGEMA_signal_4990) ) ;
    buf_clk new_AGEMA_reg_buffer_2226 ( .C (CLK), .D (new_AGEMA_signal_4993), .Q (new_AGEMA_signal_4994) ) ;
    buf_clk new_AGEMA_reg_buffer_2230 ( .C (CLK), .D (new_AGEMA_signal_4997), .Q (new_AGEMA_signal_4998) ) ;
    buf_clk new_AGEMA_reg_buffer_2234 ( .C (CLK), .D (new_AGEMA_signal_5001), .Q (new_AGEMA_signal_5002) ) ;
    buf_clk new_AGEMA_reg_buffer_2238 ( .C (CLK), .D (new_AGEMA_signal_5005), .Q (new_AGEMA_signal_5006) ) ;
    buf_clk new_AGEMA_reg_buffer_2242 ( .C (CLK), .D (new_AGEMA_signal_5009), .Q (new_AGEMA_signal_5010) ) ;
    buf_clk new_AGEMA_reg_buffer_2246 ( .C (CLK), .D (new_AGEMA_signal_5013), .Q (new_AGEMA_signal_5014) ) ;
    buf_clk new_AGEMA_reg_buffer_2250 ( .C (CLK), .D (new_AGEMA_signal_5017), .Q (new_AGEMA_signal_5018) ) ;
    buf_clk new_AGEMA_reg_buffer_2254 ( .C (CLK), .D (new_AGEMA_signal_5021), .Q (new_AGEMA_signal_5022) ) ;
    buf_clk new_AGEMA_reg_buffer_2258 ( .C (CLK), .D (new_AGEMA_signal_5025), .Q (new_AGEMA_signal_5026) ) ;
    buf_clk new_AGEMA_reg_buffer_2262 ( .C (CLK), .D (new_AGEMA_signal_5029), .Q (new_AGEMA_signal_5030) ) ;
    buf_clk new_AGEMA_reg_buffer_2266 ( .C (CLK), .D (new_AGEMA_signal_5033), .Q (new_AGEMA_signal_5034) ) ;
    buf_clk new_AGEMA_reg_buffer_2270 ( .C (CLK), .D (new_AGEMA_signal_5037), .Q (new_AGEMA_signal_5038) ) ;
    buf_clk new_AGEMA_reg_buffer_2274 ( .C (CLK), .D (new_AGEMA_signal_5041), .Q (new_AGEMA_signal_5042) ) ;
    buf_clk new_AGEMA_reg_buffer_2278 ( .C (CLK), .D (new_AGEMA_signal_5045), .Q (new_AGEMA_signal_5046) ) ;
    buf_clk new_AGEMA_reg_buffer_2282 ( .C (CLK), .D (new_AGEMA_signal_5049), .Q (new_AGEMA_signal_5050) ) ;
    buf_clk new_AGEMA_reg_buffer_2286 ( .C (CLK), .D (new_AGEMA_signal_5053), .Q (new_AGEMA_signal_5054) ) ;
    buf_clk new_AGEMA_reg_buffer_2290 ( .C (CLK), .D (new_AGEMA_signal_5057), .Q (new_AGEMA_signal_5058) ) ;
    buf_clk new_AGEMA_reg_buffer_2294 ( .C (CLK), .D (new_AGEMA_signal_5061), .Q (new_AGEMA_signal_5062) ) ;
    buf_clk new_AGEMA_reg_buffer_2298 ( .C (CLK), .D (new_AGEMA_signal_5065), .Q (new_AGEMA_signal_5066) ) ;
    buf_clk new_AGEMA_reg_buffer_2302 ( .C (CLK), .D (new_AGEMA_signal_5069), .Q (new_AGEMA_signal_5070) ) ;
    buf_clk new_AGEMA_reg_buffer_2306 ( .C (CLK), .D (new_AGEMA_signal_5073), .Q (new_AGEMA_signal_5074) ) ;
    buf_clk new_AGEMA_reg_buffer_2310 ( .C (CLK), .D (new_AGEMA_signal_5077), .Q (new_AGEMA_signal_5078) ) ;
    buf_clk new_AGEMA_reg_buffer_2314 ( .C (CLK), .D (new_AGEMA_signal_5081), .Q (new_AGEMA_signal_5082) ) ;
    buf_clk new_AGEMA_reg_buffer_2318 ( .C (CLK), .D (new_AGEMA_signal_5085), .Q (new_AGEMA_signal_5086) ) ;
    buf_clk new_AGEMA_reg_buffer_2322 ( .C (CLK), .D (new_AGEMA_signal_5089), .Q (new_AGEMA_signal_5090) ) ;
    buf_clk new_AGEMA_reg_buffer_2326 ( .C (CLK), .D (new_AGEMA_signal_5093), .Q (new_AGEMA_signal_5094) ) ;
    buf_clk new_AGEMA_reg_buffer_2330 ( .C (CLK), .D (new_AGEMA_signal_5097), .Q (new_AGEMA_signal_5098) ) ;
    buf_clk new_AGEMA_reg_buffer_2334 ( .C (CLK), .D (new_AGEMA_signal_5101), .Q (new_AGEMA_signal_5102) ) ;
    buf_clk new_AGEMA_reg_buffer_2338 ( .C (CLK), .D (new_AGEMA_signal_5105), .Q (new_AGEMA_signal_5106) ) ;
    buf_clk new_AGEMA_reg_buffer_2342 ( .C (CLK), .D (new_AGEMA_signal_5109), .Q (new_AGEMA_signal_5110) ) ;
    buf_clk new_AGEMA_reg_buffer_2346 ( .C (CLK), .D (new_AGEMA_signal_5113), .Q (new_AGEMA_signal_5114) ) ;
    buf_clk new_AGEMA_reg_buffer_2350 ( .C (CLK), .D (new_AGEMA_signal_5117), .Q (new_AGEMA_signal_5118) ) ;
    buf_clk new_AGEMA_reg_buffer_2354 ( .C (CLK), .D (new_AGEMA_signal_5121), .Q (new_AGEMA_signal_5122) ) ;
    buf_clk new_AGEMA_reg_buffer_2358 ( .C (CLK), .D (new_AGEMA_signal_5125), .Q (new_AGEMA_signal_5126) ) ;
    buf_clk new_AGEMA_reg_buffer_2362 ( .C (CLK), .D (new_AGEMA_signal_5129), .Q (new_AGEMA_signal_5130) ) ;
    buf_clk new_AGEMA_reg_buffer_2366 ( .C (CLK), .D (new_AGEMA_signal_5133), .Q (new_AGEMA_signal_5134) ) ;
    buf_clk new_AGEMA_reg_buffer_2370 ( .C (CLK), .D (new_AGEMA_signal_5137), .Q (new_AGEMA_signal_5138) ) ;
    buf_clk new_AGEMA_reg_buffer_2374 ( .C (CLK), .D (new_AGEMA_signal_5141), .Q (new_AGEMA_signal_5142) ) ;
    buf_clk new_AGEMA_reg_buffer_2378 ( .C (CLK), .D (new_AGEMA_signal_5145), .Q (new_AGEMA_signal_5146) ) ;
    buf_clk new_AGEMA_reg_buffer_2382 ( .C (CLK), .D (new_AGEMA_signal_5149), .Q (new_AGEMA_signal_5150) ) ;
    buf_clk new_AGEMA_reg_buffer_2386 ( .C (CLK), .D (new_AGEMA_signal_5153), .Q (new_AGEMA_signal_5154) ) ;
    buf_clk new_AGEMA_reg_buffer_2390 ( .C (CLK), .D (new_AGEMA_signal_5157), .Q (new_AGEMA_signal_5158) ) ;
    buf_clk new_AGEMA_reg_buffer_2394 ( .C (CLK), .D (new_AGEMA_signal_5161), .Q (new_AGEMA_signal_5162) ) ;
    buf_clk new_AGEMA_reg_buffer_2398 ( .C (CLK), .D (new_AGEMA_signal_5165), .Q (new_AGEMA_signal_5166) ) ;
    buf_clk new_AGEMA_reg_buffer_2402 ( .C (CLK), .D (new_AGEMA_signal_5169), .Q (new_AGEMA_signal_5170) ) ;
    buf_clk new_AGEMA_reg_buffer_2406 ( .C (CLK), .D (new_AGEMA_signal_5173), .Q (new_AGEMA_signal_5174) ) ;
    buf_clk new_AGEMA_reg_buffer_2410 ( .C (CLK), .D (new_AGEMA_signal_5177), .Q (new_AGEMA_signal_5178) ) ;
    buf_clk new_AGEMA_reg_buffer_2414 ( .C (CLK), .D (new_AGEMA_signal_5181), .Q (new_AGEMA_signal_5182) ) ;
    buf_clk new_AGEMA_reg_buffer_2418 ( .C (CLK), .D (new_AGEMA_signal_5185), .Q (new_AGEMA_signal_5186) ) ;
    buf_clk new_AGEMA_reg_buffer_2422 ( .C (CLK), .D (new_AGEMA_signal_5189), .Q (new_AGEMA_signal_5190) ) ;
    buf_clk new_AGEMA_reg_buffer_2426 ( .C (CLK), .D (new_AGEMA_signal_5193), .Q (new_AGEMA_signal_5194) ) ;
    buf_clk new_AGEMA_reg_buffer_2430 ( .C (CLK), .D (new_AGEMA_signal_5197), .Q (new_AGEMA_signal_5198) ) ;
    buf_clk new_AGEMA_reg_buffer_2434 ( .C (CLK), .D (new_AGEMA_signal_5201), .Q (new_AGEMA_signal_5202) ) ;
    buf_clk new_AGEMA_reg_buffer_2438 ( .C (CLK), .D (new_AGEMA_signal_5205), .Q (new_AGEMA_signal_5206) ) ;
    buf_clk new_AGEMA_reg_buffer_2442 ( .C (CLK), .D (new_AGEMA_signal_5209), .Q (new_AGEMA_signal_5210) ) ;
    buf_clk new_AGEMA_reg_buffer_2446 ( .C (CLK), .D (new_AGEMA_signal_5213), .Q (new_AGEMA_signal_5214) ) ;
    buf_clk new_AGEMA_reg_buffer_2450 ( .C (CLK), .D (new_AGEMA_signal_5217), .Q (new_AGEMA_signal_5218) ) ;
    buf_clk new_AGEMA_reg_buffer_2454 ( .C (CLK), .D (new_AGEMA_signal_5221), .Q (new_AGEMA_signal_5222) ) ;
    buf_clk new_AGEMA_reg_buffer_2458 ( .C (CLK), .D (new_AGEMA_signal_5225), .Q (new_AGEMA_signal_5226) ) ;
    buf_clk new_AGEMA_reg_buffer_2462 ( .C (CLK), .D (new_AGEMA_signal_5229), .Q (new_AGEMA_signal_5230) ) ;
    buf_clk new_AGEMA_reg_buffer_2466 ( .C (CLK), .D (new_AGEMA_signal_5233), .Q (new_AGEMA_signal_5234) ) ;
    buf_clk new_AGEMA_reg_buffer_2470 ( .C (CLK), .D (new_AGEMA_signal_5237), .Q (new_AGEMA_signal_5238) ) ;
    buf_clk new_AGEMA_reg_buffer_2474 ( .C (CLK), .D (new_AGEMA_signal_5241), .Q (new_AGEMA_signal_5242) ) ;
    buf_clk new_AGEMA_reg_buffer_2478 ( .C (CLK), .D (new_AGEMA_signal_5245), .Q (new_AGEMA_signal_5246) ) ;
    buf_clk new_AGEMA_reg_buffer_2482 ( .C (CLK), .D (new_AGEMA_signal_5249), .Q (new_AGEMA_signal_5250) ) ;
    buf_clk new_AGEMA_reg_buffer_2486 ( .C (CLK), .D (new_AGEMA_signal_5253), .Q (new_AGEMA_signal_5254) ) ;
    buf_clk new_AGEMA_reg_buffer_2490 ( .C (CLK), .D (new_AGEMA_signal_5257), .Q (new_AGEMA_signal_5258) ) ;
    buf_clk new_AGEMA_reg_buffer_2494 ( .C (CLK), .D (new_AGEMA_signal_5261), .Q (new_AGEMA_signal_5262) ) ;
    buf_clk new_AGEMA_reg_buffer_2498 ( .C (CLK), .D (new_AGEMA_signal_5265), .Q (new_AGEMA_signal_5266) ) ;
    buf_clk new_AGEMA_reg_buffer_2502 ( .C (CLK), .D (new_AGEMA_signal_5269), .Q (new_AGEMA_signal_5270) ) ;
    buf_clk new_AGEMA_reg_buffer_2506 ( .C (CLK), .D (new_AGEMA_signal_5273), .Q (new_AGEMA_signal_5274) ) ;
    buf_clk new_AGEMA_reg_buffer_2510 ( .C (CLK), .D (new_AGEMA_signal_5277), .Q (new_AGEMA_signal_5278) ) ;
    buf_clk new_AGEMA_reg_buffer_2514 ( .C (CLK), .D (new_AGEMA_signal_5281), .Q (new_AGEMA_signal_5282) ) ;
    buf_clk new_AGEMA_reg_buffer_2518 ( .C (CLK), .D (new_AGEMA_signal_5285), .Q (new_AGEMA_signal_5286) ) ;
    buf_clk new_AGEMA_reg_buffer_2522 ( .C (CLK), .D (new_AGEMA_signal_5289), .Q (new_AGEMA_signal_5290) ) ;
    buf_clk new_AGEMA_reg_buffer_2526 ( .C (CLK), .D (new_AGEMA_signal_5293), .Q (new_AGEMA_signal_5294) ) ;
    buf_clk new_AGEMA_reg_buffer_2530 ( .C (CLK), .D (new_AGEMA_signal_5297), .Q (new_AGEMA_signal_5298) ) ;
    buf_clk new_AGEMA_reg_buffer_2534 ( .C (CLK), .D (new_AGEMA_signal_5301), .Q (new_AGEMA_signal_5302) ) ;
    buf_clk new_AGEMA_reg_buffer_2538 ( .C (CLK), .D (new_AGEMA_signal_5305), .Q (new_AGEMA_signal_5306) ) ;
    buf_clk new_AGEMA_reg_buffer_2542 ( .C (CLK), .D (new_AGEMA_signal_5309), .Q (new_AGEMA_signal_5310) ) ;
    buf_clk new_AGEMA_reg_buffer_2546 ( .C (CLK), .D (new_AGEMA_signal_5313), .Q (new_AGEMA_signal_5314) ) ;
    buf_clk new_AGEMA_reg_buffer_2550 ( .C (CLK), .D (new_AGEMA_signal_5317), .Q (new_AGEMA_signal_5318) ) ;
    buf_clk new_AGEMA_reg_buffer_2554 ( .C (CLK), .D (new_AGEMA_signal_5321), .Q (new_AGEMA_signal_5322) ) ;
    buf_clk new_AGEMA_reg_buffer_2558 ( .C (CLK), .D (new_AGEMA_signal_5325), .Q (new_AGEMA_signal_5326) ) ;
    buf_clk new_AGEMA_reg_buffer_2562 ( .C (CLK), .D (new_AGEMA_signal_5329), .Q (new_AGEMA_signal_5330) ) ;
    buf_clk new_AGEMA_reg_buffer_2566 ( .C (CLK), .D (new_AGEMA_signal_5333), .Q (new_AGEMA_signal_5334) ) ;
    buf_clk new_AGEMA_reg_buffer_2570 ( .C (CLK), .D (new_AGEMA_signal_5337), .Q (new_AGEMA_signal_5338) ) ;
    buf_clk new_AGEMA_reg_buffer_2574 ( .C (CLK), .D (new_AGEMA_signal_5341), .Q (new_AGEMA_signal_5342) ) ;
    buf_clk new_AGEMA_reg_buffer_2578 ( .C (CLK), .D (new_AGEMA_signal_5345), .Q (new_AGEMA_signal_5346) ) ;
    buf_clk new_AGEMA_reg_buffer_2582 ( .C (CLK), .D (new_AGEMA_signal_5349), .Q (new_AGEMA_signal_5350) ) ;
    buf_clk new_AGEMA_reg_buffer_2586 ( .C (CLK), .D (new_AGEMA_signal_5353), .Q (new_AGEMA_signal_5354) ) ;
    buf_clk new_AGEMA_reg_buffer_2590 ( .C (CLK), .D (new_AGEMA_signal_5357), .Q (new_AGEMA_signal_5358) ) ;
    buf_clk new_AGEMA_reg_buffer_2594 ( .C (CLK), .D (new_AGEMA_signal_5361), .Q (new_AGEMA_signal_5362) ) ;
    buf_clk new_AGEMA_reg_buffer_2598 ( .C (CLK), .D (new_AGEMA_signal_5365), .Q (new_AGEMA_signal_5366) ) ;
    buf_clk new_AGEMA_reg_buffer_2602 ( .C (CLK), .D (new_AGEMA_signal_5369), .Q (new_AGEMA_signal_5370) ) ;
    buf_clk new_AGEMA_reg_buffer_2606 ( .C (CLK), .D (new_AGEMA_signal_5373), .Q (new_AGEMA_signal_5374) ) ;
    buf_clk new_AGEMA_reg_buffer_2610 ( .C (CLK), .D (new_AGEMA_signal_5377), .Q (new_AGEMA_signal_5378) ) ;
    buf_clk new_AGEMA_reg_buffer_2614 ( .C (CLK), .D (new_AGEMA_signal_5381), .Q (new_AGEMA_signal_5382) ) ;
    buf_clk new_AGEMA_reg_buffer_2618 ( .C (CLK), .D (new_AGEMA_signal_5385), .Q (new_AGEMA_signal_5386) ) ;
    buf_clk new_AGEMA_reg_buffer_2622 ( .C (CLK), .D (new_AGEMA_signal_5389), .Q (new_AGEMA_signal_5390) ) ;
    buf_clk new_AGEMA_reg_buffer_2626 ( .C (CLK), .D (new_AGEMA_signal_5393), .Q (new_AGEMA_signal_5394) ) ;
    buf_clk new_AGEMA_reg_buffer_2630 ( .C (CLK), .D (new_AGEMA_signal_5397), .Q (new_AGEMA_signal_5398) ) ;
    buf_clk new_AGEMA_reg_buffer_2634 ( .C (CLK), .D (new_AGEMA_signal_5401), .Q (new_AGEMA_signal_5402) ) ;
    buf_clk new_AGEMA_reg_buffer_2638 ( .C (CLK), .D (new_AGEMA_signal_5405), .Q (new_AGEMA_signal_5406) ) ;
    buf_clk new_AGEMA_reg_buffer_2642 ( .C (CLK), .D (new_AGEMA_signal_5409), .Q (new_AGEMA_signal_5410) ) ;
    buf_clk new_AGEMA_reg_buffer_2646 ( .C (CLK), .D (new_AGEMA_signal_5413), .Q (new_AGEMA_signal_5414) ) ;
    buf_clk new_AGEMA_reg_buffer_2650 ( .C (CLK), .D (new_AGEMA_signal_5417), .Q (new_AGEMA_signal_5418) ) ;
    buf_clk new_AGEMA_reg_buffer_2654 ( .C (CLK), .D (new_AGEMA_signal_5421), .Q (new_AGEMA_signal_5422) ) ;
    buf_clk new_AGEMA_reg_buffer_2658 ( .C (CLK), .D (new_AGEMA_signal_5425), .Q (new_AGEMA_signal_5426) ) ;
    buf_clk new_AGEMA_reg_buffer_2662 ( .C (CLK), .D (new_AGEMA_signal_5429), .Q (new_AGEMA_signal_5430) ) ;
    buf_clk new_AGEMA_reg_buffer_2666 ( .C (CLK), .D (new_AGEMA_signal_5433), .Q (new_AGEMA_signal_5434) ) ;
    buf_clk new_AGEMA_reg_buffer_2670 ( .C (CLK), .D (new_AGEMA_signal_5437), .Q (new_AGEMA_signal_5438) ) ;
    buf_clk new_AGEMA_reg_buffer_2674 ( .C (CLK), .D (new_AGEMA_signal_5441), .Q (new_AGEMA_signal_5442) ) ;
    buf_clk new_AGEMA_reg_buffer_2678 ( .C (CLK), .D (new_AGEMA_signal_5445), .Q (new_AGEMA_signal_5446) ) ;
    buf_clk new_AGEMA_reg_buffer_2682 ( .C (CLK), .D (new_AGEMA_signal_5449), .Q (new_AGEMA_signal_5450) ) ;
    buf_clk new_AGEMA_reg_buffer_2686 ( .C (CLK), .D (new_AGEMA_signal_5453), .Q (new_AGEMA_signal_5454) ) ;
    buf_clk new_AGEMA_reg_buffer_2690 ( .C (CLK), .D (new_AGEMA_signal_5457), .Q (new_AGEMA_signal_5458) ) ;
    buf_clk new_AGEMA_reg_buffer_2694 ( .C (CLK), .D (new_AGEMA_signal_5461), .Q (new_AGEMA_signal_5462) ) ;
    buf_clk new_AGEMA_reg_buffer_2698 ( .C (CLK), .D (new_AGEMA_signal_5465), .Q (new_AGEMA_signal_5466) ) ;
    buf_clk new_AGEMA_reg_buffer_2702 ( .C (CLK), .D (new_AGEMA_signal_5469), .Q (new_AGEMA_signal_5470) ) ;
    buf_clk new_AGEMA_reg_buffer_2706 ( .C (CLK), .D (new_AGEMA_signal_5473), .Q (new_AGEMA_signal_5474) ) ;
    buf_clk new_AGEMA_reg_buffer_2710 ( .C (CLK), .D (new_AGEMA_signal_5477), .Q (new_AGEMA_signal_5478) ) ;
    buf_clk new_AGEMA_reg_buffer_2714 ( .C (CLK), .D (new_AGEMA_signal_5481), .Q (new_AGEMA_signal_5482) ) ;
    buf_clk new_AGEMA_reg_buffer_2718 ( .C (CLK), .D (new_AGEMA_signal_5485), .Q (new_AGEMA_signal_5486) ) ;
    buf_clk new_AGEMA_reg_buffer_2722 ( .C (CLK), .D (new_AGEMA_signal_5489), .Q (new_AGEMA_signal_5490) ) ;
    buf_clk new_AGEMA_reg_buffer_2726 ( .C (CLK), .D (new_AGEMA_signal_5493), .Q (new_AGEMA_signal_5494) ) ;
    buf_clk new_AGEMA_reg_buffer_2730 ( .C (CLK), .D (new_AGEMA_signal_5497), .Q (new_AGEMA_signal_5498) ) ;
    buf_clk new_AGEMA_reg_buffer_2734 ( .C (CLK), .D (new_AGEMA_signal_5501), .Q (new_AGEMA_signal_5502) ) ;
    buf_clk new_AGEMA_reg_buffer_2738 ( .C (CLK), .D (new_AGEMA_signal_5505), .Q (new_AGEMA_signal_5506) ) ;
    buf_clk new_AGEMA_reg_buffer_2742 ( .C (CLK), .D (new_AGEMA_signal_5509), .Q (new_AGEMA_signal_5510) ) ;
    buf_clk new_AGEMA_reg_buffer_2746 ( .C (CLK), .D (new_AGEMA_signal_5513), .Q (new_AGEMA_signal_5514) ) ;
    buf_clk new_AGEMA_reg_buffer_2750 ( .C (CLK), .D (new_AGEMA_signal_5517), .Q (new_AGEMA_signal_5518) ) ;
    buf_clk new_AGEMA_reg_buffer_2754 ( .C (CLK), .D (new_AGEMA_signal_5521), .Q (new_AGEMA_signal_5522) ) ;
    buf_clk new_AGEMA_reg_buffer_2758 ( .C (CLK), .D (new_AGEMA_signal_5525), .Q (new_AGEMA_signal_5526) ) ;
    buf_clk new_AGEMA_reg_buffer_2762 ( .C (CLK), .D (new_AGEMA_signal_5529), .Q (new_AGEMA_signal_5530) ) ;
    buf_clk new_AGEMA_reg_buffer_2766 ( .C (CLK), .D (new_AGEMA_signal_5533), .Q (new_AGEMA_signal_5534) ) ;
    buf_clk new_AGEMA_reg_buffer_2770 ( .C (CLK), .D (new_AGEMA_signal_5537), .Q (new_AGEMA_signal_5538) ) ;
    buf_clk new_AGEMA_reg_buffer_2774 ( .C (CLK), .D (new_AGEMA_signal_5541), .Q (new_AGEMA_signal_5542) ) ;
    buf_clk new_AGEMA_reg_buffer_2778 ( .C (CLK), .D (new_AGEMA_signal_5545), .Q (new_AGEMA_signal_5546) ) ;
    buf_clk new_AGEMA_reg_buffer_2782 ( .C (CLK), .D (new_AGEMA_signal_5549), .Q (new_AGEMA_signal_5550) ) ;
    buf_clk new_AGEMA_reg_buffer_2786 ( .C (CLK), .D (new_AGEMA_signal_5553), .Q (new_AGEMA_signal_5554) ) ;
    buf_clk new_AGEMA_reg_buffer_2790 ( .C (CLK), .D (new_AGEMA_signal_5557), .Q (new_AGEMA_signal_5558) ) ;
    buf_clk new_AGEMA_reg_buffer_2794 ( .C (CLK), .D (new_AGEMA_signal_5561), .Q (new_AGEMA_signal_5562) ) ;
    buf_clk new_AGEMA_reg_buffer_2798 ( .C (CLK), .D (new_AGEMA_signal_5565), .Q (new_AGEMA_signal_5566) ) ;
    buf_clk new_AGEMA_reg_buffer_2802 ( .C (CLK), .D (new_AGEMA_signal_5569), .Q (new_AGEMA_signal_5570) ) ;
    buf_clk new_AGEMA_reg_buffer_2806 ( .C (CLK), .D (new_AGEMA_signal_5573), .Q (new_AGEMA_signal_5574) ) ;
    buf_clk new_AGEMA_reg_buffer_2810 ( .C (CLK), .D (new_AGEMA_signal_5577), .Q (new_AGEMA_signal_5578) ) ;
    buf_clk new_AGEMA_reg_buffer_2814 ( .C (CLK), .D (new_AGEMA_signal_5581), .Q (new_AGEMA_signal_5582) ) ;
    buf_clk new_AGEMA_reg_buffer_2818 ( .C (CLK), .D (new_AGEMA_signal_5585), .Q (new_AGEMA_signal_5586) ) ;
    buf_clk new_AGEMA_reg_buffer_2822 ( .C (CLK), .D (new_AGEMA_signal_5589), .Q (new_AGEMA_signal_5590) ) ;
    buf_clk new_AGEMA_reg_buffer_2826 ( .C (CLK), .D (new_AGEMA_signal_5593), .Q (new_AGEMA_signal_5594) ) ;
    buf_clk new_AGEMA_reg_buffer_2830 ( .C (CLK), .D (new_AGEMA_signal_5597), .Q (new_AGEMA_signal_5598) ) ;
    buf_clk new_AGEMA_reg_buffer_2834 ( .C (CLK), .D (new_AGEMA_signal_5601), .Q (new_AGEMA_signal_5602) ) ;
    buf_clk new_AGEMA_reg_buffer_2838 ( .C (CLK), .D (new_AGEMA_signal_5605), .Q (new_AGEMA_signal_5606) ) ;
    buf_clk new_AGEMA_reg_buffer_2842 ( .C (CLK), .D (new_AGEMA_signal_5609), .Q (new_AGEMA_signal_5610) ) ;
    buf_clk new_AGEMA_reg_buffer_2846 ( .C (CLK), .D (new_AGEMA_signal_5613), .Q (new_AGEMA_signal_5614) ) ;
    buf_clk new_AGEMA_reg_buffer_2850 ( .C (CLK), .D (new_AGEMA_signal_5617), .Q (new_AGEMA_signal_5618) ) ;
    buf_clk new_AGEMA_reg_buffer_2854 ( .C (CLK), .D (new_AGEMA_signal_5621), .Q (new_AGEMA_signal_5622) ) ;
    buf_clk new_AGEMA_reg_buffer_2858 ( .C (CLK), .D (new_AGEMA_signal_5625), .Q (new_AGEMA_signal_5626) ) ;
    buf_clk new_AGEMA_reg_buffer_2862 ( .C (CLK), .D (new_AGEMA_signal_5629), .Q (new_AGEMA_signal_5630) ) ;
    buf_clk new_AGEMA_reg_buffer_2866 ( .C (CLK), .D (new_AGEMA_signal_5633), .Q (new_AGEMA_signal_5634) ) ;
    buf_clk new_AGEMA_reg_buffer_2870 ( .C (CLK), .D (new_AGEMA_signal_5637), .Q (new_AGEMA_signal_5638) ) ;
    buf_clk new_AGEMA_reg_buffer_2874 ( .C (CLK), .D (new_AGEMA_signal_5641), .Q (new_AGEMA_signal_5642) ) ;
    buf_clk new_AGEMA_reg_buffer_2878 ( .C (CLK), .D (new_AGEMA_signal_5645), .Q (new_AGEMA_signal_5646) ) ;
    buf_clk new_AGEMA_reg_buffer_2882 ( .C (CLK), .D (new_AGEMA_signal_5649), .Q (new_AGEMA_signal_5650) ) ;
    buf_clk new_AGEMA_reg_buffer_2886 ( .C (CLK), .D (new_AGEMA_signal_5653), .Q (new_AGEMA_signal_5654) ) ;
    buf_clk new_AGEMA_reg_buffer_2890 ( .C (CLK), .D (new_AGEMA_signal_5657), .Q (new_AGEMA_signal_5658) ) ;
    buf_clk new_AGEMA_reg_buffer_2894 ( .C (CLK), .D (new_AGEMA_signal_5661), .Q (new_AGEMA_signal_5662) ) ;
    buf_clk new_AGEMA_reg_buffer_2898 ( .C (CLK), .D (new_AGEMA_signal_5665), .Q (new_AGEMA_signal_5666) ) ;
    buf_clk new_AGEMA_reg_buffer_2902 ( .C (CLK), .D (new_AGEMA_signal_5669), .Q (new_AGEMA_signal_5670) ) ;
    buf_clk new_AGEMA_reg_buffer_2906 ( .C (CLK), .D (new_AGEMA_signal_5673), .Q (new_AGEMA_signal_5674) ) ;
    buf_clk new_AGEMA_reg_buffer_2910 ( .C (CLK), .D (new_AGEMA_signal_5677), .Q (new_AGEMA_signal_5678) ) ;
    buf_clk new_AGEMA_reg_buffer_2914 ( .C (CLK), .D (new_AGEMA_signal_5681), .Q (new_AGEMA_signal_5682) ) ;
    buf_clk new_AGEMA_reg_buffer_2918 ( .C (CLK), .D (new_AGEMA_signal_5685), .Q (new_AGEMA_signal_5686) ) ;
    buf_clk new_AGEMA_reg_buffer_2922 ( .C (CLK), .D (new_AGEMA_signal_5689), .Q (new_AGEMA_signal_5690) ) ;
    buf_clk new_AGEMA_reg_buffer_2926 ( .C (CLK), .D (new_AGEMA_signal_5693), .Q (new_AGEMA_signal_5694) ) ;
    buf_clk new_AGEMA_reg_buffer_2930 ( .C (CLK), .D (new_AGEMA_signal_5697), .Q (new_AGEMA_signal_5698) ) ;
    buf_clk new_AGEMA_reg_buffer_2934 ( .C (CLK), .D (new_AGEMA_signal_5701), .Q (new_AGEMA_signal_5702) ) ;
    buf_clk new_AGEMA_reg_buffer_2938 ( .C (CLK), .D (new_AGEMA_signal_5705), .Q (new_AGEMA_signal_5706) ) ;
    buf_clk new_AGEMA_reg_buffer_2942 ( .C (CLK), .D (new_AGEMA_signal_5709), .Q (new_AGEMA_signal_5710) ) ;
    buf_clk new_AGEMA_reg_buffer_2946 ( .C (CLK), .D (new_AGEMA_signal_5713), .Q (new_AGEMA_signal_5714) ) ;
    buf_clk new_AGEMA_reg_buffer_2950 ( .C (CLK), .D (new_AGEMA_signal_5717), .Q (new_AGEMA_signal_5718) ) ;
    buf_clk new_AGEMA_reg_buffer_2954 ( .C (CLK), .D (new_AGEMA_signal_5721), .Q (new_AGEMA_signal_5722) ) ;
    buf_clk new_AGEMA_reg_buffer_2958 ( .C (CLK), .D (new_AGEMA_signal_5725), .Q (new_AGEMA_signal_5726) ) ;
    buf_clk new_AGEMA_reg_buffer_2962 ( .C (CLK), .D (new_AGEMA_signal_5729), .Q (new_AGEMA_signal_5730) ) ;
    buf_clk new_AGEMA_reg_buffer_2966 ( .C (CLK), .D (new_AGEMA_signal_5733), .Q (new_AGEMA_signal_5734) ) ;
    buf_clk new_AGEMA_reg_buffer_2970 ( .C (CLK), .D (new_AGEMA_signal_5737), .Q (new_AGEMA_signal_5738) ) ;
    buf_clk new_AGEMA_reg_buffer_2984 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_0_L5), .Q (new_AGEMA_signal_5752) ) ;
    buf_clk new_AGEMA_reg_buffer_2986 ( .C (CLK), .D (new_AGEMA_signal_2602), .Q (new_AGEMA_signal_5754) ) ;
    buf_clk new_AGEMA_reg_buffer_2988 ( .C (CLK), .D (new_AGEMA_signal_2603), .Q (new_AGEMA_signal_5756) ) ;
    buf_clk new_AGEMA_reg_buffer_2992 ( .C (CLK), .D (new_AGEMA_signal_5759), .Q (new_AGEMA_signal_5760) ) ;
    buf_clk new_AGEMA_reg_buffer_2996 ( .C (CLK), .D (new_AGEMA_signal_5763), .Q (new_AGEMA_signal_5764) ) ;
    buf_clk new_AGEMA_reg_buffer_3000 ( .C (CLK), .D (new_AGEMA_signal_5767), .Q (new_AGEMA_signal_5768) ) ;
    buf_clk new_AGEMA_reg_buffer_3004 ( .C (CLK), .D (new_AGEMA_signal_5771), .Q (new_AGEMA_signal_5772) ) ;
    buf_clk new_AGEMA_reg_buffer_3008 ( .C (CLK), .D (new_AGEMA_signal_5775), .Q (new_AGEMA_signal_5776) ) ;
    buf_clk new_AGEMA_reg_buffer_3012 ( .C (CLK), .D (new_AGEMA_signal_5779), .Q (new_AGEMA_signal_5780) ) ;
    buf_clk new_AGEMA_reg_buffer_3014 ( .C (CLK), .D (new_AGEMA_signal_3903), .Q (new_AGEMA_signal_5782) ) ;
    buf_clk new_AGEMA_reg_buffer_3016 ( .C (CLK), .D (new_AGEMA_signal_3905), .Q (new_AGEMA_signal_5784) ) ;
    buf_clk new_AGEMA_reg_buffer_3018 ( .C (CLK), .D (new_AGEMA_signal_3907), .Q (new_AGEMA_signal_5786) ) ;
    buf_clk new_AGEMA_reg_buffer_3032 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_1_L5), .Q (new_AGEMA_signal_5800) ) ;
    buf_clk new_AGEMA_reg_buffer_3034 ( .C (CLK), .D (new_AGEMA_signal_2606), .Q (new_AGEMA_signal_5802) ) ;
    buf_clk new_AGEMA_reg_buffer_3036 ( .C (CLK), .D (new_AGEMA_signal_2607), .Q (new_AGEMA_signal_5804) ) ;
    buf_clk new_AGEMA_reg_buffer_3040 ( .C (CLK), .D (new_AGEMA_signal_5807), .Q (new_AGEMA_signal_5808) ) ;
    buf_clk new_AGEMA_reg_buffer_3044 ( .C (CLK), .D (new_AGEMA_signal_5811), .Q (new_AGEMA_signal_5812) ) ;
    buf_clk new_AGEMA_reg_buffer_3048 ( .C (CLK), .D (new_AGEMA_signal_5815), .Q (new_AGEMA_signal_5816) ) ;
    buf_clk new_AGEMA_reg_buffer_3052 ( .C (CLK), .D (new_AGEMA_signal_5819), .Q (new_AGEMA_signal_5820) ) ;
    buf_clk new_AGEMA_reg_buffer_3056 ( .C (CLK), .D (new_AGEMA_signal_5823), .Q (new_AGEMA_signal_5824) ) ;
    buf_clk new_AGEMA_reg_buffer_3060 ( .C (CLK), .D (new_AGEMA_signal_5827), .Q (new_AGEMA_signal_5828) ) ;
    buf_clk new_AGEMA_reg_buffer_3062 ( .C (CLK), .D (new_AGEMA_signal_3921), .Q (new_AGEMA_signal_5830) ) ;
    buf_clk new_AGEMA_reg_buffer_3064 ( .C (CLK), .D (new_AGEMA_signal_3923), .Q (new_AGEMA_signal_5832) ) ;
    buf_clk new_AGEMA_reg_buffer_3066 ( .C (CLK), .D (new_AGEMA_signal_3925), .Q (new_AGEMA_signal_5834) ) ;
    buf_clk new_AGEMA_reg_buffer_3080 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_2_L5), .Q (new_AGEMA_signal_5848) ) ;
    buf_clk new_AGEMA_reg_buffer_3082 ( .C (CLK), .D (new_AGEMA_signal_2546), .Q (new_AGEMA_signal_5850) ) ;
    buf_clk new_AGEMA_reg_buffer_3084 ( .C (CLK), .D (new_AGEMA_signal_2547), .Q (new_AGEMA_signal_5852) ) ;
    buf_clk new_AGEMA_reg_buffer_3088 ( .C (CLK), .D (new_AGEMA_signal_5855), .Q (new_AGEMA_signal_5856) ) ;
    buf_clk new_AGEMA_reg_buffer_3092 ( .C (CLK), .D (new_AGEMA_signal_5859), .Q (new_AGEMA_signal_5860) ) ;
    buf_clk new_AGEMA_reg_buffer_3096 ( .C (CLK), .D (new_AGEMA_signal_5863), .Q (new_AGEMA_signal_5864) ) ;
    buf_clk new_AGEMA_reg_buffer_3098 ( .C (CLK), .D (new_AGEMA_signal_3939), .Q (new_AGEMA_signal_5866) ) ;
    buf_clk new_AGEMA_reg_buffer_3100 ( .C (CLK), .D (new_AGEMA_signal_3941), .Q (new_AGEMA_signal_5868) ) ;
    buf_clk new_AGEMA_reg_buffer_3102 ( .C (CLK), .D (new_AGEMA_signal_3943), .Q (new_AGEMA_signal_5870) ) ;
    buf_clk new_AGEMA_reg_buffer_3116 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_3_L5), .Q (new_AGEMA_signal_5884) ) ;
    buf_clk new_AGEMA_reg_buffer_3118 ( .C (CLK), .D (new_AGEMA_signal_2550), .Q (new_AGEMA_signal_5886) ) ;
    buf_clk new_AGEMA_reg_buffer_3120 ( .C (CLK), .D (new_AGEMA_signal_2551), .Q (new_AGEMA_signal_5888) ) ;
    buf_clk new_AGEMA_reg_buffer_3124 ( .C (CLK), .D (new_AGEMA_signal_5891), .Q (new_AGEMA_signal_5892) ) ;
    buf_clk new_AGEMA_reg_buffer_3128 ( .C (CLK), .D (new_AGEMA_signal_5895), .Q (new_AGEMA_signal_5896) ) ;
    buf_clk new_AGEMA_reg_buffer_3132 ( .C (CLK), .D (new_AGEMA_signal_5899), .Q (new_AGEMA_signal_5900) ) ;
    buf_clk new_AGEMA_reg_buffer_3134 ( .C (CLK), .D (new_AGEMA_signal_3957), .Q (new_AGEMA_signal_5902) ) ;
    buf_clk new_AGEMA_reg_buffer_3136 ( .C (CLK), .D (new_AGEMA_signal_3959), .Q (new_AGEMA_signal_5904) ) ;
    buf_clk new_AGEMA_reg_buffer_3138 ( .C (CLK), .D (new_AGEMA_signal_3961), .Q (new_AGEMA_signal_5906) ) ;
    buf_clk new_AGEMA_reg_buffer_3152 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_4_L5), .Q (new_AGEMA_signal_5920) ) ;
    buf_clk new_AGEMA_reg_buffer_3154 ( .C (CLK), .D (new_AGEMA_signal_2618), .Q (new_AGEMA_signal_5922) ) ;
    buf_clk new_AGEMA_reg_buffer_3156 ( .C (CLK), .D (new_AGEMA_signal_2619), .Q (new_AGEMA_signal_5924) ) ;
    buf_clk new_AGEMA_reg_buffer_3160 ( .C (CLK), .D (new_AGEMA_signal_5927), .Q (new_AGEMA_signal_5928) ) ;
    buf_clk new_AGEMA_reg_buffer_3164 ( .C (CLK), .D (new_AGEMA_signal_5931), .Q (new_AGEMA_signal_5932) ) ;
    buf_clk new_AGEMA_reg_buffer_3168 ( .C (CLK), .D (new_AGEMA_signal_5935), .Q (new_AGEMA_signal_5936) ) ;
    buf_clk new_AGEMA_reg_buffer_3172 ( .C (CLK), .D (new_AGEMA_signal_5939), .Q (new_AGEMA_signal_5940) ) ;
    buf_clk new_AGEMA_reg_buffer_3176 ( .C (CLK), .D (new_AGEMA_signal_5943), .Q (new_AGEMA_signal_5944) ) ;
    buf_clk new_AGEMA_reg_buffer_3180 ( .C (CLK), .D (new_AGEMA_signal_5947), .Q (new_AGEMA_signal_5948) ) ;
    buf_clk new_AGEMA_reg_buffer_3182 ( .C (CLK), .D (new_AGEMA_signal_3975), .Q (new_AGEMA_signal_5950) ) ;
    buf_clk new_AGEMA_reg_buffer_3184 ( .C (CLK), .D (new_AGEMA_signal_3977), .Q (new_AGEMA_signal_5952) ) ;
    buf_clk new_AGEMA_reg_buffer_3186 ( .C (CLK), .D (new_AGEMA_signal_3979), .Q (new_AGEMA_signal_5954) ) ;
    buf_clk new_AGEMA_reg_buffer_3200 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_5_L5), .Q (new_AGEMA_signal_5968) ) ;
    buf_clk new_AGEMA_reg_buffer_3202 ( .C (CLK), .D (new_AGEMA_signal_2622), .Q (new_AGEMA_signal_5970) ) ;
    buf_clk new_AGEMA_reg_buffer_3204 ( .C (CLK), .D (new_AGEMA_signal_2623), .Q (new_AGEMA_signal_5972) ) ;
    buf_clk new_AGEMA_reg_buffer_3208 ( .C (CLK), .D (new_AGEMA_signal_5975), .Q (new_AGEMA_signal_5976) ) ;
    buf_clk new_AGEMA_reg_buffer_3212 ( .C (CLK), .D (new_AGEMA_signal_5979), .Q (new_AGEMA_signal_5980) ) ;
    buf_clk new_AGEMA_reg_buffer_3216 ( .C (CLK), .D (new_AGEMA_signal_5983), .Q (new_AGEMA_signal_5984) ) ;
    buf_clk new_AGEMA_reg_buffer_3220 ( .C (CLK), .D (new_AGEMA_signal_5987), .Q (new_AGEMA_signal_5988) ) ;
    buf_clk new_AGEMA_reg_buffer_3224 ( .C (CLK), .D (new_AGEMA_signal_5991), .Q (new_AGEMA_signal_5992) ) ;
    buf_clk new_AGEMA_reg_buffer_3228 ( .C (CLK), .D (new_AGEMA_signal_5995), .Q (new_AGEMA_signal_5996) ) ;
    buf_clk new_AGEMA_reg_buffer_3230 ( .C (CLK), .D (new_AGEMA_signal_3993), .Q (new_AGEMA_signal_5998) ) ;
    buf_clk new_AGEMA_reg_buffer_3232 ( .C (CLK), .D (new_AGEMA_signal_3995), .Q (new_AGEMA_signal_6000) ) ;
    buf_clk new_AGEMA_reg_buffer_3234 ( .C (CLK), .D (new_AGEMA_signal_3997), .Q (new_AGEMA_signal_6002) ) ;
    buf_clk new_AGEMA_reg_buffer_3248 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_6_L5), .Q (new_AGEMA_signal_6016) ) ;
    buf_clk new_AGEMA_reg_buffer_3250 ( .C (CLK), .D (new_AGEMA_signal_2562), .Q (new_AGEMA_signal_6018) ) ;
    buf_clk new_AGEMA_reg_buffer_3252 ( .C (CLK), .D (new_AGEMA_signal_2563), .Q (new_AGEMA_signal_6020) ) ;
    buf_clk new_AGEMA_reg_buffer_3256 ( .C (CLK), .D (new_AGEMA_signal_6023), .Q (new_AGEMA_signal_6024) ) ;
    buf_clk new_AGEMA_reg_buffer_3260 ( .C (CLK), .D (new_AGEMA_signal_6027), .Q (new_AGEMA_signal_6028) ) ;
    buf_clk new_AGEMA_reg_buffer_3264 ( .C (CLK), .D (new_AGEMA_signal_6031), .Q (new_AGEMA_signal_6032) ) ;
    buf_clk new_AGEMA_reg_buffer_3266 ( .C (CLK), .D (new_AGEMA_signal_4011), .Q (new_AGEMA_signal_6034) ) ;
    buf_clk new_AGEMA_reg_buffer_3268 ( .C (CLK), .D (new_AGEMA_signal_4013), .Q (new_AGEMA_signal_6036) ) ;
    buf_clk new_AGEMA_reg_buffer_3270 ( .C (CLK), .D (new_AGEMA_signal_4015), .Q (new_AGEMA_signal_6038) ) ;
    buf_clk new_AGEMA_reg_buffer_3284 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_7_L5), .Q (new_AGEMA_signal_6052) ) ;
    buf_clk new_AGEMA_reg_buffer_3286 ( .C (CLK), .D (new_AGEMA_signal_2566), .Q (new_AGEMA_signal_6054) ) ;
    buf_clk new_AGEMA_reg_buffer_3288 ( .C (CLK), .D (new_AGEMA_signal_2567), .Q (new_AGEMA_signal_6056) ) ;
    buf_clk new_AGEMA_reg_buffer_3292 ( .C (CLK), .D (new_AGEMA_signal_6059), .Q (new_AGEMA_signal_6060) ) ;
    buf_clk new_AGEMA_reg_buffer_3296 ( .C (CLK), .D (new_AGEMA_signal_6063), .Q (new_AGEMA_signal_6064) ) ;
    buf_clk new_AGEMA_reg_buffer_3300 ( .C (CLK), .D (new_AGEMA_signal_6067), .Q (new_AGEMA_signal_6068) ) ;
    buf_clk new_AGEMA_reg_buffer_3302 ( .C (CLK), .D (new_AGEMA_signal_4029), .Q (new_AGEMA_signal_6070) ) ;
    buf_clk new_AGEMA_reg_buffer_3304 ( .C (CLK), .D (new_AGEMA_signal_4031), .Q (new_AGEMA_signal_6072) ) ;
    buf_clk new_AGEMA_reg_buffer_3306 ( .C (CLK), .D (new_AGEMA_signal_4033), .Q (new_AGEMA_signal_6074) ) ;
    buf_clk new_AGEMA_reg_buffer_3320 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_8_L5), .Q (new_AGEMA_signal_6088) ) ;
    buf_clk new_AGEMA_reg_buffer_3322 ( .C (CLK), .D (new_AGEMA_signal_2634), .Q (new_AGEMA_signal_6090) ) ;
    buf_clk new_AGEMA_reg_buffer_3324 ( .C (CLK), .D (new_AGEMA_signal_2635), .Q (new_AGEMA_signal_6092) ) ;
    buf_clk new_AGEMA_reg_buffer_3328 ( .C (CLK), .D (new_AGEMA_signal_6095), .Q (new_AGEMA_signal_6096) ) ;
    buf_clk new_AGEMA_reg_buffer_3332 ( .C (CLK), .D (new_AGEMA_signal_6099), .Q (new_AGEMA_signal_6100) ) ;
    buf_clk new_AGEMA_reg_buffer_3336 ( .C (CLK), .D (new_AGEMA_signal_6103), .Q (new_AGEMA_signal_6104) ) ;
    buf_clk new_AGEMA_reg_buffer_3340 ( .C (CLK), .D (new_AGEMA_signal_6107), .Q (new_AGEMA_signal_6108) ) ;
    buf_clk new_AGEMA_reg_buffer_3344 ( .C (CLK), .D (new_AGEMA_signal_6111), .Q (new_AGEMA_signal_6112) ) ;
    buf_clk new_AGEMA_reg_buffer_3348 ( .C (CLK), .D (new_AGEMA_signal_6115), .Q (new_AGEMA_signal_6116) ) ;
    buf_clk new_AGEMA_reg_buffer_3350 ( .C (CLK), .D (new_AGEMA_signal_4047), .Q (new_AGEMA_signal_6118) ) ;
    buf_clk new_AGEMA_reg_buffer_3352 ( .C (CLK), .D (new_AGEMA_signal_4049), .Q (new_AGEMA_signal_6120) ) ;
    buf_clk new_AGEMA_reg_buffer_3354 ( .C (CLK), .D (new_AGEMA_signal_4051), .Q (new_AGEMA_signal_6122) ) ;
    buf_clk new_AGEMA_reg_buffer_3368 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_9_L5), .Q (new_AGEMA_signal_6136) ) ;
    buf_clk new_AGEMA_reg_buffer_3370 ( .C (CLK), .D (new_AGEMA_signal_2638), .Q (new_AGEMA_signal_6138) ) ;
    buf_clk new_AGEMA_reg_buffer_3372 ( .C (CLK), .D (new_AGEMA_signal_2639), .Q (new_AGEMA_signal_6140) ) ;
    buf_clk new_AGEMA_reg_buffer_3376 ( .C (CLK), .D (new_AGEMA_signal_6143), .Q (new_AGEMA_signal_6144) ) ;
    buf_clk new_AGEMA_reg_buffer_3380 ( .C (CLK), .D (new_AGEMA_signal_6147), .Q (new_AGEMA_signal_6148) ) ;
    buf_clk new_AGEMA_reg_buffer_3384 ( .C (CLK), .D (new_AGEMA_signal_6151), .Q (new_AGEMA_signal_6152) ) ;
    buf_clk new_AGEMA_reg_buffer_3388 ( .C (CLK), .D (new_AGEMA_signal_6155), .Q (new_AGEMA_signal_6156) ) ;
    buf_clk new_AGEMA_reg_buffer_3392 ( .C (CLK), .D (new_AGEMA_signal_6159), .Q (new_AGEMA_signal_6160) ) ;
    buf_clk new_AGEMA_reg_buffer_3396 ( .C (CLK), .D (new_AGEMA_signal_6163), .Q (new_AGEMA_signal_6164) ) ;
    buf_clk new_AGEMA_reg_buffer_3398 ( .C (CLK), .D (new_AGEMA_signal_4065), .Q (new_AGEMA_signal_6166) ) ;
    buf_clk new_AGEMA_reg_buffer_3400 ( .C (CLK), .D (new_AGEMA_signal_4067), .Q (new_AGEMA_signal_6168) ) ;
    buf_clk new_AGEMA_reg_buffer_3402 ( .C (CLK), .D (new_AGEMA_signal_4069), .Q (new_AGEMA_signal_6170) ) ;
    buf_clk new_AGEMA_reg_buffer_3416 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_10_L5), .Q (new_AGEMA_signal_6184) ) ;
    buf_clk new_AGEMA_reg_buffer_3418 ( .C (CLK), .D (new_AGEMA_signal_2578), .Q (new_AGEMA_signal_6186) ) ;
    buf_clk new_AGEMA_reg_buffer_3420 ( .C (CLK), .D (new_AGEMA_signal_2579), .Q (new_AGEMA_signal_6188) ) ;
    buf_clk new_AGEMA_reg_buffer_3424 ( .C (CLK), .D (new_AGEMA_signal_6191), .Q (new_AGEMA_signal_6192) ) ;
    buf_clk new_AGEMA_reg_buffer_3428 ( .C (CLK), .D (new_AGEMA_signal_6195), .Q (new_AGEMA_signal_6196) ) ;
    buf_clk new_AGEMA_reg_buffer_3432 ( .C (CLK), .D (new_AGEMA_signal_6199), .Q (new_AGEMA_signal_6200) ) ;
    buf_clk new_AGEMA_reg_buffer_3434 ( .C (CLK), .D (new_AGEMA_signal_4083), .Q (new_AGEMA_signal_6202) ) ;
    buf_clk new_AGEMA_reg_buffer_3436 ( .C (CLK), .D (new_AGEMA_signal_4085), .Q (new_AGEMA_signal_6204) ) ;
    buf_clk new_AGEMA_reg_buffer_3438 ( .C (CLK), .D (new_AGEMA_signal_4087), .Q (new_AGEMA_signal_6206) ) ;
    buf_clk new_AGEMA_reg_buffer_3452 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_11_L5), .Q (new_AGEMA_signal_6220) ) ;
    buf_clk new_AGEMA_reg_buffer_3454 ( .C (CLK), .D (new_AGEMA_signal_2582), .Q (new_AGEMA_signal_6222) ) ;
    buf_clk new_AGEMA_reg_buffer_3456 ( .C (CLK), .D (new_AGEMA_signal_2583), .Q (new_AGEMA_signal_6224) ) ;
    buf_clk new_AGEMA_reg_buffer_3460 ( .C (CLK), .D (new_AGEMA_signal_6227), .Q (new_AGEMA_signal_6228) ) ;
    buf_clk new_AGEMA_reg_buffer_3464 ( .C (CLK), .D (new_AGEMA_signal_6231), .Q (new_AGEMA_signal_6232) ) ;
    buf_clk new_AGEMA_reg_buffer_3468 ( .C (CLK), .D (new_AGEMA_signal_6235), .Q (new_AGEMA_signal_6236) ) ;
    buf_clk new_AGEMA_reg_buffer_3470 ( .C (CLK), .D (new_AGEMA_signal_4101), .Q (new_AGEMA_signal_6238) ) ;
    buf_clk new_AGEMA_reg_buffer_3472 ( .C (CLK), .D (new_AGEMA_signal_4103), .Q (new_AGEMA_signal_6240) ) ;
    buf_clk new_AGEMA_reg_buffer_3474 ( .C (CLK), .D (new_AGEMA_signal_4105), .Q (new_AGEMA_signal_6242) ) ;
    buf_clk new_AGEMA_reg_buffer_3488 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_12_L5), .Q (new_AGEMA_signal_6256) ) ;
    buf_clk new_AGEMA_reg_buffer_3490 ( .C (CLK), .D (new_AGEMA_signal_2650), .Q (new_AGEMA_signal_6258) ) ;
    buf_clk new_AGEMA_reg_buffer_3492 ( .C (CLK), .D (new_AGEMA_signal_2651), .Q (new_AGEMA_signal_6260) ) ;
    buf_clk new_AGEMA_reg_buffer_3496 ( .C (CLK), .D (new_AGEMA_signal_6263), .Q (new_AGEMA_signal_6264) ) ;
    buf_clk new_AGEMA_reg_buffer_3500 ( .C (CLK), .D (new_AGEMA_signal_6267), .Q (new_AGEMA_signal_6268) ) ;
    buf_clk new_AGEMA_reg_buffer_3504 ( .C (CLK), .D (new_AGEMA_signal_6271), .Q (new_AGEMA_signal_6272) ) ;
    buf_clk new_AGEMA_reg_buffer_3508 ( .C (CLK), .D (new_AGEMA_signal_6275), .Q (new_AGEMA_signal_6276) ) ;
    buf_clk new_AGEMA_reg_buffer_3512 ( .C (CLK), .D (new_AGEMA_signal_6279), .Q (new_AGEMA_signal_6280) ) ;
    buf_clk new_AGEMA_reg_buffer_3516 ( .C (CLK), .D (new_AGEMA_signal_6283), .Q (new_AGEMA_signal_6284) ) ;
    buf_clk new_AGEMA_reg_buffer_3518 ( .C (CLK), .D (new_AGEMA_signal_4119), .Q (new_AGEMA_signal_6286) ) ;
    buf_clk new_AGEMA_reg_buffer_3520 ( .C (CLK), .D (new_AGEMA_signal_4121), .Q (new_AGEMA_signal_6288) ) ;
    buf_clk new_AGEMA_reg_buffer_3522 ( .C (CLK), .D (new_AGEMA_signal_4123), .Q (new_AGEMA_signal_6290) ) ;
    buf_clk new_AGEMA_reg_buffer_3536 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_13_L5), .Q (new_AGEMA_signal_6304) ) ;
    buf_clk new_AGEMA_reg_buffer_3538 ( .C (CLK), .D (new_AGEMA_signal_2654), .Q (new_AGEMA_signal_6306) ) ;
    buf_clk new_AGEMA_reg_buffer_3540 ( .C (CLK), .D (new_AGEMA_signal_2655), .Q (new_AGEMA_signal_6308) ) ;
    buf_clk new_AGEMA_reg_buffer_3544 ( .C (CLK), .D (new_AGEMA_signal_6311), .Q (new_AGEMA_signal_6312) ) ;
    buf_clk new_AGEMA_reg_buffer_3548 ( .C (CLK), .D (new_AGEMA_signal_6315), .Q (new_AGEMA_signal_6316) ) ;
    buf_clk new_AGEMA_reg_buffer_3552 ( .C (CLK), .D (new_AGEMA_signal_6319), .Q (new_AGEMA_signal_6320) ) ;
    buf_clk new_AGEMA_reg_buffer_3556 ( .C (CLK), .D (new_AGEMA_signal_6323), .Q (new_AGEMA_signal_6324) ) ;
    buf_clk new_AGEMA_reg_buffer_3560 ( .C (CLK), .D (new_AGEMA_signal_6327), .Q (new_AGEMA_signal_6328) ) ;
    buf_clk new_AGEMA_reg_buffer_3564 ( .C (CLK), .D (new_AGEMA_signal_6331), .Q (new_AGEMA_signal_6332) ) ;
    buf_clk new_AGEMA_reg_buffer_3566 ( .C (CLK), .D (new_AGEMA_signal_4137), .Q (new_AGEMA_signal_6334) ) ;
    buf_clk new_AGEMA_reg_buffer_3568 ( .C (CLK), .D (new_AGEMA_signal_4139), .Q (new_AGEMA_signal_6336) ) ;
    buf_clk new_AGEMA_reg_buffer_3570 ( .C (CLK), .D (new_AGEMA_signal_4141), .Q (new_AGEMA_signal_6338) ) ;
    buf_clk new_AGEMA_reg_buffer_3584 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_14_L5), .Q (new_AGEMA_signal_6352) ) ;
    buf_clk new_AGEMA_reg_buffer_3586 ( .C (CLK), .D (new_AGEMA_signal_2594), .Q (new_AGEMA_signal_6354) ) ;
    buf_clk new_AGEMA_reg_buffer_3588 ( .C (CLK), .D (new_AGEMA_signal_2595), .Q (new_AGEMA_signal_6356) ) ;
    buf_clk new_AGEMA_reg_buffer_3592 ( .C (CLK), .D (new_AGEMA_signal_6359), .Q (new_AGEMA_signal_6360) ) ;
    buf_clk new_AGEMA_reg_buffer_3596 ( .C (CLK), .D (new_AGEMA_signal_6363), .Q (new_AGEMA_signal_6364) ) ;
    buf_clk new_AGEMA_reg_buffer_3600 ( .C (CLK), .D (new_AGEMA_signal_6367), .Q (new_AGEMA_signal_6368) ) ;
    buf_clk new_AGEMA_reg_buffer_3602 ( .C (CLK), .D (new_AGEMA_signal_4155), .Q (new_AGEMA_signal_6370) ) ;
    buf_clk new_AGEMA_reg_buffer_3604 ( .C (CLK), .D (new_AGEMA_signal_4157), .Q (new_AGEMA_signal_6372) ) ;
    buf_clk new_AGEMA_reg_buffer_3606 ( .C (CLK), .D (new_AGEMA_signal_4159), .Q (new_AGEMA_signal_6374) ) ;
    buf_clk new_AGEMA_reg_buffer_3620 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_15_L5), .Q (new_AGEMA_signal_6388) ) ;
    buf_clk new_AGEMA_reg_buffer_3622 ( .C (CLK), .D (new_AGEMA_signal_2598), .Q (new_AGEMA_signal_6390) ) ;
    buf_clk new_AGEMA_reg_buffer_3624 ( .C (CLK), .D (new_AGEMA_signal_2599), .Q (new_AGEMA_signal_6392) ) ;
    buf_clk new_AGEMA_reg_buffer_3628 ( .C (CLK), .D (new_AGEMA_signal_6395), .Q (new_AGEMA_signal_6396) ) ;
    buf_clk new_AGEMA_reg_buffer_3632 ( .C (CLK), .D (new_AGEMA_signal_6399), .Q (new_AGEMA_signal_6400) ) ;
    buf_clk new_AGEMA_reg_buffer_3636 ( .C (CLK), .D (new_AGEMA_signal_6403), .Q (new_AGEMA_signal_6404) ) ;
    buf_clk new_AGEMA_reg_buffer_3638 ( .C (CLK), .D (new_AGEMA_signal_4173), .Q (new_AGEMA_signal_6406) ) ;
    buf_clk new_AGEMA_reg_buffer_3640 ( .C (CLK), .D (new_AGEMA_signal_4175), .Q (new_AGEMA_signal_6408) ) ;
    buf_clk new_AGEMA_reg_buffer_3642 ( .C (CLK), .D (new_AGEMA_signal_4177), .Q (new_AGEMA_signal_6410) ) ;
    buf_clk new_AGEMA_reg_buffer_3644 ( .C (CLK), .D (LED_128_Instance_subcells_out[60]), .Q (new_AGEMA_signal_6412) ) ;
    buf_clk new_AGEMA_reg_buffer_3646 ( .C (CLK), .D (new_AGEMA_signal_2534), .Q (new_AGEMA_signal_6414) ) ;
    buf_clk new_AGEMA_reg_buffer_3648 ( .C (CLK), .D (new_AGEMA_signal_2535), .Q (new_AGEMA_signal_6416) ) ;
    buf_clk new_AGEMA_reg_buffer_3650 ( .C (CLK), .D (LED_128_Instance_subcells_out[20]), .Q (new_AGEMA_signal_6418) ) ;
    buf_clk new_AGEMA_reg_buffer_3652 ( .C (CLK), .D (new_AGEMA_signal_2558), .Q (new_AGEMA_signal_6420) ) ;
    buf_clk new_AGEMA_reg_buffer_3654 ( .C (CLK), .D (new_AGEMA_signal_2559), .Q (new_AGEMA_signal_6422) ) ;
    buf_clk new_AGEMA_reg_buffer_3656 ( .C (CLK), .D (LED_128_Instance_subcells_out[40]), .Q (new_AGEMA_signal_6424) ) ;
    buf_clk new_AGEMA_reg_buffer_3658 ( .C (CLK), .D (new_AGEMA_signal_2502), .Q (new_AGEMA_signal_6426) ) ;
    buf_clk new_AGEMA_reg_buffer_3660 ( .C (CLK), .D (new_AGEMA_signal_2503), .Q (new_AGEMA_signal_6428) ) ;
    buf_clk new_AGEMA_reg_buffer_3662 ( .C (CLK), .D (LED_128_Instance_subcells_out[0]), .Q (new_AGEMA_signal_6430) ) ;
    buf_clk new_AGEMA_reg_buffer_3664 ( .C (CLK), .D (new_AGEMA_signal_2538), .Q (new_AGEMA_signal_6432) ) ;
    buf_clk new_AGEMA_reg_buffer_3666 ( .C (CLK), .D (new_AGEMA_signal_2539), .Q (new_AGEMA_signal_6434) ) ;
    buf_clk new_AGEMA_reg_buffer_3668 ( .C (CLK), .D (LED_128_Instance_subcells_out[48]), .Q (new_AGEMA_signal_6436) ) ;
    buf_clk new_AGEMA_reg_buffer_3670 ( .C (CLK), .D (new_AGEMA_signal_2586), .Q (new_AGEMA_signal_6438) ) ;
    buf_clk new_AGEMA_reg_buffer_3672 ( .C (CLK), .D (new_AGEMA_signal_2587), .Q (new_AGEMA_signal_6440) ) ;
    buf_clk new_AGEMA_reg_buffer_3674 ( .C (CLK), .D (LED_128_Instance_subcells_out[24]), .Q (new_AGEMA_signal_6442) ) ;
    buf_clk new_AGEMA_reg_buffer_3676 ( .C (CLK), .D (new_AGEMA_signal_2474), .Q (new_AGEMA_signal_6444) ) ;
    buf_clk new_AGEMA_reg_buffer_3678 ( .C (CLK), .D (new_AGEMA_signal_2475), .Q (new_AGEMA_signal_6446) ) ;
    buf_clk new_AGEMA_reg_buffer_3680 ( .C (CLK), .D (LED_128_Instance_subcells_out[44]), .Q (new_AGEMA_signal_6448) ) ;
    buf_clk new_AGEMA_reg_buffer_3682 ( .C (CLK), .D (new_AGEMA_signal_2506), .Q (new_AGEMA_signal_6450) ) ;
    buf_clk new_AGEMA_reg_buffer_3684 ( .C (CLK), .D (new_AGEMA_signal_2507), .Q (new_AGEMA_signal_6452) ) ;
    buf_clk new_AGEMA_reg_buffer_3686 ( .C (CLK), .D (LED_128_Instance_subcells_out[4]), .Q (new_AGEMA_signal_6454) ) ;
    buf_clk new_AGEMA_reg_buffer_3688 ( .C (CLK), .D (new_AGEMA_signal_2542), .Q (new_AGEMA_signal_6456) ) ;
    buf_clk new_AGEMA_reg_buffer_3690 ( .C (CLK), .D (new_AGEMA_signal_2543), .Q (new_AGEMA_signal_6458) ) ;
    buf_clk new_AGEMA_reg_buffer_3692 ( .C (CLK), .D (LED_128_Instance_subcells_out[52]), .Q (new_AGEMA_signal_6460) ) ;
    buf_clk new_AGEMA_reg_buffer_3694 ( .C (CLK), .D (new_AGEMA_signal_2590), .Q (new_AGEMA_signal_6462) ) ;
    buf_clk new_AGEMA_reg_buffer_3696 ( .C (CLK), .D (new_AGEMA_signal_2591), .Q (new_AGEMA_signal_6464) ) ;
    buf_clk new_AGEMA_reg_buffer_3698 ( .C (CLK), .D (LED_128_Instance_subcells_out[28]), .Q (new_AGEMA_signal_6466) ) ;
    buf_clk new_AGEMA_reg_buffer_3700 ( .C (CLK), .D (new_AGEMA_signal_2478), .Q (new_AGEMA_signal_6468) ) ;
    buf_clk new_AGEMA_reg_buffer_3702 ( .C (CLK), .D (new_AGEMA_signal_2479), .Q (new_AGEMA_signal_6470) ) ;
    buf_clk new_AGEMA_reg_buffer_3704 ( .C (CLK), .D (LED_128_Instance_subcells_out[32]), .Q (new_AGEMA_signal_6472) ) ;
    buf_clk new_AGEMA_reg_buffer_3706 ( .C (CLK), .D (new_AGEMA_signal_2570), .Q (new_AGEMA_signal_6474) ) ;
    buf_clk new_AGEMA_reg_buffer_3708 ( .C (CLK), .D (new_AGEMA_signal_2571), .Q (new_AGEMA_signal_6476) ) ;
    buf_clk new_AGEMA_reg_buffer_3710 ( .C (CLK), .D (LED_128_Instance_subcells_out[8]), .Q (new_AGEMA_signal_6478) ) ;
    buf_clk new_AGEMA_reg_buffer_3712 ( .C (CLK), .D (new_AGEMA_signal_2446), .Q (new_AGEMA_signal_6480) ) ;
    buf_clk new_AGEMA_reg_buffer_3714 ( .C (CLK), .D (new_AGEMA_signal_2447), .Q (new_AGEMA_signal_6482) ) ;
    buf_clk new_AGEMA_reg_buffer_3716 ( .C (CLK), .D (LED_128_Instance_subcells_out[56]), .Q (new_AGEMA_signal_6484) ) ;
    buf_clk new_AGEMA_reg_buffer_3718 ( .C (CLK), .D (new_AGEMA_signal_2530), .Q (new_AGEMA_signal_6486) ) ;
    buf_clk new_AGEMA_reg_buffer_3720 ( .C (CLK), .D (new_AGEMA_signal_2531), .Q (new_AGEMA_signal_6488) ) ;
    buf_clk new_AGEMA_reg_buffer_3722 ( .C (CLK), .D (LED_128_Instance_subcells_out[16]), .Q (new_AGEMA_signal_6490) ) ;
    buf_clk new_AGEMA_reg_buffer_3724 ( .C (CLK), .D (new_AGEMA_signal_2554), .Q (new_AGEMA_signal_6492) ) ;
    buf_clk new_AGEMA_reg_buffer_3726 ( .C (CLK), .D (new_AGEMA_signal_2555), .Q (new_AGEMA_signal_6494) ) ;
    buf_clk new_AGEMA_reg_buffer_3728 ( .C (CLK), .D (LED_128_Instance_subcells_out[36]), .Q (new_AGEMA_signal_6496) ) ;
    buf_clk new_AGEMA_reg_buffer_3730 ( .C (CLK), .D (new_AGEMA_signal_2574), .Q (new_AGEMA_signal_6498) ) ;
    buf_clk new_AGEMA_reg_buffer_3732 ( .C (CLK), .D (new_AGEMA_signal_2575), .Q (new_AGEMA_signal_6500) ) ;
    buf_clk new_AGEMA_reg_buffer_3734 ( .C (CLK), .D (LED_128_Instance_subcells_out[12]), .Q (new_AGEMA_signal_6502) ) ;
    buf_clk new_AGEMA_reg_buffer_3736 ( .C (CLK), .D (new_AGEMA_signal_2450), .Q (new_AGEMA_signal_6504) ) ;
    buf_clk new_AGEMA_reg_buffer_3738 ( .C (CLK), .D (new_AGEMA_signal_2451), .Q (new_AGEMA_signal_6506) ) ;
    buf_clk new_AGEMA_reg_buffer_3742 ( .C (CLK), .D (new_AGEMA_signal_6509), .Q (new_AGEMA_signal_6510) ) ;
    buf_clk new_AGEMA_reg_buffer_3746 ( .C (CLK), .D (new_AGEMA_signal_6513), .Q (new_AGEMA_signal_6514) ) ;
    buf_clk new_AGEMA_reg_buffer_3750 ( .C (CLK), .D (new_AGEMA_signal_6517), .Q (new_AGEMA_signal_6518) ) ;
    buf_clk new_AGEMA_reg_buffer_3754 ( .C (CLK), .D (new_AGEMA_signal_6521), .Q (new_AGEMA_signal_6522) ) ;
    buf_clk new_AGEMA_reg_buffer_3758 ( .C (CLK), .D (new_AGEMA_signal_6525), .Q (new_AGEMA_signal_6526) ) ;
    buf_clk new_AGEMA_reg_buffer_3762 ( .C (CLK), .D (new_AGEMA_signal_6529), .Q (new_AGEMA_signal_6530) ) ;
    buf_clk new_AGEMA_reg_buffer_3766 ( .C (CLK), .D (new_AGEMA_signal_6533), .Q (new_AGEMA_signal_6534) ) ;
    buf_clk new_AGEMA_reg_buffer_3770 ( .C (CLK), .D (new_AGEMA_signal_6537), .Q (new_AGEMA_signal_6538) ) ;
    buf_clk new_AGEMA_reg_buffer_3774 ( .C (CLK), .D (new_AGEMA_signal_6541), .Q (new_AGEMA_signal_6542) ) ;
    buf_clk new_AGEMA_reg_buffer_3778 ( .C (CLK), .D (new_AGEMA_signal_6545), .Q (new_AGEMA_signal_6546) ) ;
    buf_clk new_AGEMA_reg_buffer_3782 ( .C (CLK), .D (new_AGEMA_signal_6549), .Q (new_AGEMA_signal_6550) ) ;

    /* cells in depth 4 */
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_0_U1 ( .s (new_AGEMA_signal_4187), .b ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, LED_128_Instance_mixcolumns_out[0]}), .a ({new_AGEMA_signal_4199, new_AGEMA_signal_4195, new_AGEMA_signal_4191}), .c ({new_AGEMA_signal_3015, new_AGEMA_signal_3014, LED_128_Instance_state0[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_1_U1 ( .s (new_AGEMA_signal_4187), .b ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, LED_128_Instance_mixcolumns_out[1]}), .a ({new_AGEMA_signal_4211, new_AGEMA_signal_4207, new_AGEMA_signal_4203}), .c ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, LED_128_Instance_state0[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_2_U1 ( .s (new_AGEMA_signal_4215), .b ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, LED_128_Instance_mixcolumns_out[2]}), .a ({new_AGEMA_signal_4227, new_AGEMA_signal_4223, new_AGEMA_signal_4219}), .c ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, LED_128_Instance_state0[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_3_U1 ( .s (new_AGEMA_signal_4231), .b ({new_AGEMA_signal_3083, new_AGEMA_signal_3082, LED_128_Instance_mixcolumns_out[3]}), .a ({new_AGEMA_signal_4243, new_AGEMA_signal_4239, new_AGEMA_signal_4235}), .c ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, LED_128_Instance_state0[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_4_U1 ( .s (new_AGEMA_signal_4231), .b ({new_AGEMA_signal_3029, new_AGEMA_signal_3028, LED_128_Instance_mixcolumns_out[4]}), .a ({new_AGEMA_signal_4255, new_AGEMA_signal_4251, new_AGEMA_signal_4247}), .c ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, LED_128_Instance_state0[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_5_U1 ( .s (new_AGEMA_signal_4231), .b ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, LED_128_Instance_mixcolumns_out[5]}), .a ({new_AGEMA_signal_4267, new_AGEMA_signal_4263, new_AGEMA_signal_4259}), .c ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, LED_128_Instance_state0[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_6_U1 ( .s (new_AGEMA_signal_4231), .b ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, LED_128_Instance_mixcolumns_out[6]}), .a ({new_AGEMA_signal_4279, new_AGEMA_signal_4275, new_AGEMA_signal_4271}), .c ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, LED_128_Instance_state0[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_7_U1 ( .s (new_AGEMA_signal_4231), .b ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, LED_128_Instance_mixcolumns_out[7]}), .a ({new_AGEMA_signal_4291, new_AGEMA_signal_4287, new_AGEMA_signal_4283}), .c ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, LED_128_Instance_state0[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_8_U1 ( .s (new_AGEMA_signal_4231), .b ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, LED_128_Instance_mixcolumns_out[8]}), .a ({new_AGEMA_signal_4303, new_AGEMA_signal_4299, new_AGEMA_signal_4295}), .c ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, LED_128_Instance_state0[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_9_U1 ( .s (new_AGEMA_signal_4231), .b ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, LED_128_Instance_mixcolumns_out[9]}), .a ({new_AGEMA_signal_4315, new_AGEMA_signal_4311, new_AGEMA_signal_4307}), .c ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, LED_128_Instance_state0[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_10_U1 ( .s (new_AGEMA_signal_4231), .b ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, LED_128_Instance_mixcolumns_out[10]}), .a ({new_AGEMA_signal_4327, new_AGEMA_signal_4323, new_AGEMA_signal_4319}), .c ({new_AGEMA_signal_3065, new_AGEMA_signal_3064, LED_128_Instance_state0[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_11_U1 ( .s (new_AGEMA_signal_4231), .b ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, LED_128_Instance_mixcolumns_out[11]}), .a ({new_AGEMA_signal_4339, new_AGEMA_signal_4335, new_AGEMA_signal_4331}), .c ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, LED_128_Instance_state0[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_12_U1 ( .s (new_AGEMA_signal_4231), .b ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, LED_128_Instance_mixcolumns_out[12]}), .a ({new_AGEMA_signal_4351, new_AGEMA_signal_4347, new_AGEMA_signal_4343}), .c ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, LED_128_Instance_state0[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_13_U1 ( .s (new_AGEMA_signal_4231), .b ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, LED_128_Instance_mixcolumns_out[13]}), .a ({new_AGEMA_signal_4363, new_AGEMA_signal_4359, new_AGEMA_signal_4355}), .c ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, LED_128_Instance_state0[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_14_U1 ( .s (new_AGEMA_signal_4231), .b ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, LED_128_Instance_mixcolumns_out[14]}), .a ({new_AGEMA_signal_4375, new_AGEMA_signal_4371, new_AGEMA_signal_4367}), .c ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, LED_128_Instance_state0[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_15_U1 ( .s (new_AGEMA_signal_4231), .b ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, LED_128_Instance_mixcolumns_out[15]}), .a ({new_AGEMA_signal_4387, new_AGEMA_signal_4383, new_AGEMA_signal_4379}), .c ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, LED_128_Instance_state0[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_16_U1 ( .s (new_AGEMA_signal_4187), .b ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, LED_128_Instance_mixcolumns_out[16]}), .a ({new_AGEMA_signal_4399, new_AGEMA_signal_4395, new_AGEMA_signal_4391}), .c ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, LED_128_Instance_state0[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_17_U1 ( .s (new_AGEMA_signal_4187), .b ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, LED_128_Instance_mixcolumns_out[17]}), .a ({new_AGEMA_signal_4411, new_AGEMA_signal_4407, new_AGEMA_signal_4403}), .c ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, LED_128_Instance_state0[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_18_U1 ( .s (new_AGEMA_signal_4187), .b ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, LED_128_Instance_mixcolumns_out[18]}), .a ({new_AGEMA_signal_4423, new_AGEMA_signal_4419, new_AGEMA_signal_4415}), .c ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, LED_128_Instance_state0[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_19_U1 ( .s (new_AGEMA_signal_4187), .b ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, LED_128_Instance_mixcolumns_out[19]}), .a ({new_AGEMA_signal_4435, new_AGEMA_signal_4431, new_AGEMA_signal_4427}), .c ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, LED_128_Instance_state0[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_20_U1 ( .s (new_AGEMA_signal_4187), .b ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, LED_128_Instance_mixcolumns_out[20]}), .a ({new_AGEMA_signal_4447, new_AGEMA_signal_4443, new_AGEMA_signal_4439}), .c ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, LED_128_Instance_state0[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_21_U1 ( .s (new_AGEMA_signal_4187), .b ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, LED_128_Instance_mixcolumns_out[21]}), .a ({new_AGEMA_signal_4459, new_AGEMA_signal_4455, new_AGEMA_signal_4451}), .c ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, LED_128_Instance_state0[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_22_U1 ( .s (new_AGEMA_signal_4187), .b ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, LED_128_Instance_mixcolumns_out[22]}), .a ({new_AGEMA_signal_4471, new_AGEMA_signal_4467, new_AGEMA_signal_4463}), .c ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, LED_128_Instance_state0[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_23_U1 ( .s (new_AGEMA_signal_4187), .b ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, LED_128_Instance_mixcolumns_out[23]}), .a ({new_AGEMA_signal_4483, new_AGEMA_signal_4479, new_AGEMA_signal_4475}), .c ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, LED_128_Instance_state0[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_24_U1 ( .s (new_AGEMA_signal_4187), .b ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, LED_128_Instance_mixcolumns_out[24]}), .a ({new_AGEMA_signal_4495, new_AGEMA_signal_4491, new_AGEMA_signal_4487}), .c ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, LED_128_Instance_state0[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_25_U1 ( .s (new_AGEMA_signal_4187), .b ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, LED_128_Instance_mixcolumns_out[25]}), .a ({new_AGEMA_signal_4507, new_AGEMA_signal_4503, new_AGEMA_signal_4499}), .c ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, LED_128_Instance_state0[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_26_U1 ( .s (new_AGEMA_signal_4187), .b ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, LED_128_Instance_mixcolumns_out[26]}), .a ({new_AGEMA_signal_4519, new_AGEMA_signal_4515, new_AGEMA_signal_4511}), .c ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, LED_128_Instance_state0[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_27_U1 ( .s (new_AGEMA_signal_4187), .b ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, LED_128_Instance_mixcolumns_out[27]}), .a ({new_AGEMA_signal_4531, new_AGEMA_signal_4527, new_AGEMA_signal_4523}), .c ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, LED_128_Instance_state0[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_28_U1 ( .s (new_AGEMA_signal_4215), .b ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, LED_128_Instance_mixcolumns_out[28]}), .a ({new_AGEMA_signal_4543, new_AGEMA_signal_4539, new_AGEMA_signal_4535}), .c ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, LED_128_Instance_state0[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_29_U1 ( .s (new_AGEMA_signal_4215), .b ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, LED_128_Instance_mixcolumns_out[29]}), .a ({new_AGEMA_signal_4555, new_AGEMA_signal_4551, new_AGEMA_signal_4547}), .c ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, LED_128_Instance_state0[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_30_U1 ( .s (new_AGEMA_signal_4215), .b ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, LED_128_Instance_mixcolumns_out[30]}), .a ({new_AGEMA_signal_4567, new_AGEMA_signal_4563, new_AGEMA_signal_4559}), .c ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, LED_128_Instance_state0[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_31_U1 ( .s (new_AGEMA_signal_4215), .b ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, LED_128_Instance_mixcolumns_out[31]}), .a ({new_AGEMA_signal_4579, new_AGEMA_signal_4575, new_AGEMA_signal_4571}), .c ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, LED_128_Instance_state0[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_32_U1 ( .s (new_AGEMA_signal_4215), .b ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, LED_128_Instance_mixcolumns_out[32]}), .a ({new_AGEMA_signal_4591, new_AGEMA_signal_4587, new_AGEMA_signal_4583}), .c ({new_AGEMA_signal_3391, new_AGEMA_signal_3390, LED_128_Instance_state0[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_33_U1 ( .s (new_AGEMA_signal_4215), .b ({new_AGEMA_signal_3443, new_AGEMA_signal_3442, LED_128_Instance_mixcolumns_out[33]}), .a ({new_AGEMA_signal_4603, new_AGEMA_signal_4599, new_AGEMA_signal_4595}), .c ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, LED_128_Instance_state0[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_34_U1 ( .s (new_AGEMA_signal_4215), .b ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, LED_128_Instance_mixcolumns_out[34]}), .a ({new_AGEMA_signal_4615, new_AGEMA_signal_4611, new_AGEMA_signal_4607}), .c ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, LED_128_Instance_state0[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_35_U1 ( .s (new_AGEMA_signal_4215), .b ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, LED_128_Instance_mixcolumns_out[35]}), .a ({new_AGEMA_signal_4627, new_AGEMA_signal_4623, new_AGEMA_signal_4619}), .c ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, LED_128_Instance_state0[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_36_U1 ( .s (new_AGEMA_signal_4215), .b ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, LED_128_Instance_mixcolumns_out[36]}), .a ({new_AGEMA_signal_4639, new_AGEMA_signal_4635, new_AGEMA_signal_4631}), .c ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, LED_128_Instance_state0[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_37_U1 ( .s (new_AGEMA_signal_4215), .b ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, LED_128_Instance_mixcolumns_out[37]}), .a ({new_AGEMA_signal_4651, new_AGEMA_signal_4647, new_AGEMA_signal_4643}), .c ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, LED_128_Instance_state0[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_38_U1 ( .s (new_AGEMA_signal_4215), .b ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, LED_128_Instance_mixcolumns_out[38]}), .a ({new_AGEMA_signal_4663, new_AGEMA_signal_4659, new_AGEMA_signal_4655}), .c ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, LED_128_Instance_state0[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_39_U1 ( .s (new_AGEMA_signal_4215), .b ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, LED_128_Instance_mixcolumns_out[39]}), .a ({new_AGEMA_signal_4675, new_AGEMA_signal_4671, new_AGEMA_signal_4667}), .c ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, LED_128_Instance_state0[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_40_U1 ( .s (new_AGEMA_signal_4215), .b ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, LED_128_Instance_mixcolumns_out[40]}), .a ({new_AGEMA_signal_4687, new_AGEMA_signal_4683, new_AGEMA_signal_4679}), .c ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, LED_128_Instance_state0[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_41_U1 ( .s (new_AGEMA_signal_4187), .b ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, LED_128_Instance_mixcolumns_out[41]}), .a ({new_AGEMA_signal_4699, new_AGEMA_signal_4695, new_AGEMA_signal_4691}), .c ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, LED_128_Instance_state0[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_42_U1 ( .s (new_AGEMA_signal_4231), .b ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, LED_128_Instance_mixcolumns_out[42]}), .a ({new_AGEMA_signal_4711, new_AGEMA_signal_4707, new_AGEMA_signal_4703}), .c ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, LED_128_Instance_state0[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_43_U1 ( .s (new_AGEMA_signal_4715), .b ({new_AGEMA_signal_3455, new_AGEMA_signal_3454, LED_128_Instance_mixcolumns_out[43]}), .a ({new_AGEMA_signal_4727, new_AGEMA_signal_4723, new_AGEMA_signal_4719}), .c ({new_AGEMA_signal_3465, new_AGEMA_signal_3464, LED_128_Instance_state0[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_44_U1 ( .s (new_AGEMA_signal_4187), .b ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, LED_128_Instance_mixcolumns_out[44]}), .a ({new_AGEMA_signal_4739, new_AGEMA_signal_4735, new_AGEMA_signal_4731}), .c ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, LED_128_Instance_state0[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_45_U1 ( .s (new_AGEMA_signal_4231), .b ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, LED_128_Instance_mixcolumns_out[45]}), .a ({new_AGEMA_signal_4751, new_AGEMA_signal_4747, new_AGEMA_signal_4743}), .c ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, LED_128_Instance_state0[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_46_U1 ( .s (new_AGEMA_signal_4215), .b ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, LED_128_Instance_mixcolumns_out[46]}), .a ({new_AGEMA_signal_4763, new_AGEMA_signal_4759, new_AGEMA_signal_4755}), .c ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, LED_128_Instance_state0[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_47_U1 ( .s (new_AGEMA_signal_4715), .b ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, LED_128_Instance_mixcolumns_out[47]}), .a ({new_AGEMA_signal_4775, new_AGEMA_signal_4771, new_AGEMA_signal_4767}), .c ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, LED_128_Instance_state0[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_48_U1 ( .s (new_AGEMA_signal_4715), .b ({new_AGEMA_signal_3647, new_AGEMA_signal_3646, LED_128_Instance_mixcolumns_out[48]}), .a ({new_AGEMA_signal_4787, new_AGEMA_signal_4783, new_AGEMA_signal_4779}), .c ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, LED_128_Instance_state0[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_49_U1 ( .s (new_AGEMA_signal_4715), .b ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, LED_128_Instance_mixcolumns_out[49]}), .a ({new_AGEMA_signal_4799, new_AGEMA_signal_4795, new_AGEMA_signal_4791}), .c ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, LED_128_Instance_state0[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_50_U1 ( .s (new_AGEMA_signal_4715), .b ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, LED_128_Instance_mixcolumns_out[50]}), .a ({new_AGEMA_signal_4811, new_AGEMA_signal_4807, new_AGEMA_signal_4803}), .c ({new_AGEMA_signal_3547, new_AGEMA_signal_3546, LED_128_Instance_state0[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_51_U1 ( .s (new_AGEMA_signal_4715), .b ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, LED_128_Instance_mixcolumns_out[51]}), .a ({new_AGEMA_signal_4823, new_AGEMA_signal_4819, new_AGEMA_signal_4815}), .c ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, LED_128_Instance_state0[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_52_U1 ( .s (new_AGEMA_signal_4715), .b ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, LED_128_Instance_mixcolumns_out[52]}), .a ({new_AGEMA_signal_4835, new_AGEMA_signal_4831, new_AGEMA_signal_4827}), .c ({new_AGEMA_signal_3659, new_AGEMA_signal_3658, LED_128_Instance_state0[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_53_U1 ( .s (new_AGEMA_signal_4715), .b ({new_AGEMA_signal_3675, new_AGEMA_signal_3674, LED_128_Instance_mixcolumns_out[53]}), .a ({new_AGEMA_signal_4847, new_AGEMA_signal_4843, new_AGEMA_signal_4839}), .c ({new_AGEMA_signal_3679, new_AGEMA_signal_3678, LED_128_Instance_state0[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_54_U1 ( .s (new_AGEMA_signal_4215), .b ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, LED_128_Instance_mixcolumns_out[54]}), .a ({new_AGEMA_signal_4859, new_AGEMA_signal_4855, new_AGEMA_signal_4851}), .c ({new_AGEMA_signal_3471, new_AGEMA_signal_3470, LED_128_Instance_state0[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_55_U1 ( .s (new_AGEMA_signal_4187), .b ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, LED_128_Instance_mixcolumns_out[55]}), .a ({new_AGEMA_signal_4871, new_AGEMA_signal_4867, new_AGEMA_signal_4863}), .c ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, LED_128_Instance_state0[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_56_U1 ( .s (new_AGEMA_signal_4231), .b ({new_AGEMA_signal_3635, new_AGEMA_signal_3634, LED_128_Instance_mixcolumns_out[56]}), .a ({new_AGEMA_signal_4883, new_AGEMA_signal_4879, new_AGEMA_signal_4875}), .c ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, LED_128_Instance_state0[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_57_U1 ( .s (new_AGEMA_signal_4215), .b ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, LED_128_Instance_mixcolumns_out[57]}), .a ({new_AGEMA_signal_4895, new_AGEMA_signal_4891, new_AGEMA_signal_4887}), .c ({new_AGEMA_signal_3661, new_AGEMA_signal_3660, LED_128_Instance_state0[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_58_U1 ( .s (new_AGEMA_signal_4187), .b ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, LED_128_Instance_mixcolumns_out[58]}), .a ({new_AGEMA_signal_4907, new_AGEMA_signal_4903, new_AGEMA_signal_4899}), .c ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, LED_128_Instance_state0[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_59_U1 ( .s (new_AGEMA_signal_4231), .b ({new_AGEMA_signal_3451, new_AGEMA_signal_3450, LED_128_Instance_mixcolumns_out[59]}), .a ({new_AGEMA_signal_4919, new_AGEMA_signal_4915, new_AGEMA_signal_4911}), .c ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, LED_128_Instance_state0[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_60_U1 ( .s (new_AGEMA_signal_4187), .b ({new_AGEMA_signal_3639, new_AGEMA_signal_3638, LED_128_Instance_mixcolumns_out[60]}), .a ({new_AGEMA_signal_4931, new_AGEMA_signal_4927, new_AGEMA_signal_4923}), .c ({new_AGEMA_signal_3643, new_AGEMA_signal_3642, LED_128_Instance_state0[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_61_U1 ( .s (new_AGEMA_signal_4231), .b ({new_AGEMA_signal_3655, new_AGEMA_signal_3654, LED_128_Instance_mixcolumns_out[61]}), .a ({new_AGEMA_signal_4943, new_AGEMA_signal_4939, new_AGEMA_signal_4935}), .c ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, LED_128_Instance_state0[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_62_U1 ( .s (new_AGEMA_signal_4215), .b ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, LED_128_Instance_mixcolumns_out[62]}), .a ({new_AGEMA_signal_4955, new_AGEMA_signal_4951, new_AGEMA_signal_4947}), .c ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, LED_128_Instance_state0[62]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_63_U1 ( .s (new_AGEMA_signal_4215), .b ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, LED_128_Instance_mixcolumns_out[63]}), .a ({new_AGEMA_signal_4967, new_AGEMA_signal_4963, new_AGEMA_signal_4959}), .c ({new_AGEMA_signal_3555, new_AGEMA_signal_3554, LED_128_Instance_state0[63]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_0_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3015, new_AGEMA_signal_3014, LED_128_Instance_state0[0]}), .a ({new_AGEMA_signal_4983, new_AGEMA_signal_4979, new_AGEMA_signal_4975}), .c ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_state1[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_1_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, LED_128_Instance_state0[1]}), .a ({new_AGEMA_signal_4995, new_AGEMA_signal_4991, new_AGEMA_signal_4987}), .c ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, LED_128_Instance_state1[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_2_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, LED_128_Instance_state0[2]}), .a ({new_AGEMA_signal_5007, new_AGEMA_signal_5003, new_AGEMA_signal_4999}), .c ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, LED_128_Instance_state1[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_3_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, LED_128_Instance_state0[3]}), .a ({new_AGEMA_signal_5019, new_AGEMA_signal_5015, new_AGEMA_signal_5011}), .c ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, LED_128_Instance_state1[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_4_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, LED_128_Instance_state0[4]}), .a ({new_AGEMA_signal_5031, new_AGEMA_signal_5027, new_AGEMA_signal_5023}), .c ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, LED_128_Instance_state1[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_5_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, LED_128_Instance_state0[5]}), .a ({new_AGEMA_signal_5043, new_AGEMA_signal_5039, new_AGEMA_signal_5035}), .c ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, LED_128_Instance_state1[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_6_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, LED_128_Instance_state0[6]}), .a ({new_AGEMA_signal_5055, new_AGEMA_signal_5051, new_AGEMA_signal_5047}), .c ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, LED_128_Instance_state1[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_7_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, LED_128_Instance_state0[7]}), .a ({new_AGEMA_signal_5067, new_AGEMA_signal_5063, new_AGEMA_signal_5059}), .c ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, LED_128_Instance_state1[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_8_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, LED_128_Instance_state0[8]}), .a ({new_AGEMA_signal_5079, new_AGEMA_signal_5075, new_AGEMA_signal_5071}), .c ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, LED_128_Instance_state1[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_9_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, LED_128_Instance_state0[9]}), .a ({new_AGEMA_signal_5091, new_AGEMA_signal_5087, new_AGEMA_signal_5083}), .c ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, LED_128_Instance_state1[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_10_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3065, new_AGEMA_signal_3064, LED_128_Instance_state0[10]}), .a ({new_AGEMA_signal_5103, new_AGEMA_signal_5099, new_AGEMA_signal_5095}), .c ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, LED_128_Instance_state1[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_11_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, LED_128_Instance_state0[11]}), .a ({new_AGEMA_signal_5115, new_AGEMA_signal_5111, new_AGEMA_signal_5107}), .c ({new_AGEMA_signal_3151, new_AGEMA_signal_3150, LED_128_Instance_state1[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_12_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, LED_128_Instance_state0[12]}), .a ({new_AGEMA_signal_5127, new_AGEMA_signal_5123, new_AGEMA_signal_5119}), .c ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, LED_128_Instance_state1[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_13_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, LED_128_Instance_state0[13]}), .a ({new_AGEMA_signal_5139, new_AGEMA_signal_5135, new_AGEMA_signal_5131}), .c ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, LED_128_Instance_state1[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_14_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, LED_128_Instance_state0[14]}), .a ({new_AGEMA_signal_5151, new_AGEMA_signal_5147, new_AGEMA_signal_5143}), .c ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, LED_128_Instance_state1[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_15_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, LED_128_Instance_state0[15]}), .a ({new_AGEMA_signal_5163, new_AGEMA_signal_5159, new_AGEMA_signal_5155}), .c ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, LED_128_Instance_state1[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_16_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, LED_128_Instance_state0[16]}), .a ({new_AGEMA_signal_5175, new_AGEMA_signal_5171, new_AGEMA_signal_5167}), .c ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, LED_128_Instance_state1[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_17_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, LED_128_Instance_state0[17]}), .a ({new_AGEMA_signal_5187, new_AGEMA_signal_5183, new_AGEMA_signal_5179}), .c ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, LED_128_Instance_state1[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_18_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, LED_128_Instance_state0[18]}), .a ({new_AGEMA_signal_5199, new_AGEMA_signal_5195, new_AGEMA_signal_5191}), .c ({new_AGEMA_signal_3483, new_AGEMA_signal_3482, LED_128_Instance_state1[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_19_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, LED_128_Instance_state0[19]}), .a ({new_AGEMA_signal_5211, new_AGEMA_signal_5207, new_AGEMA_signal_5203}), .c ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, LED_128_Instance_state1[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_20_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, LED_128_Instance_state0[20]}), .a ({new_AGEMA_signal_5223, new_AGEMA_signal_5219, new_AGEMA_signal_5215}), .c ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, LED_128_Instance_state1[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_21_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, LED_128_Instance_state0[21]}), .a ({new_AGEMA_signal_5235, new_AGEMA_signal_5231, new_AGEMA_signal_5227}), .c ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, LED_128_Instance_state1[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_22_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, LED_128_Instance_state0[22]}), .a ({new_AGEMA_signal_5247, new_AGEMA_signal_5243, new_AGEMA_signal_5239}), .c ({new_AGEMA_signal_3487, new_AGEMA_signal_3486, LED_128_Instance_state1[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_23_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, LED_128_Instance_state0[23]}), .a ({new_AGEMA_signal_5259, new_AGEMA_signal_5255, new_AGEMA_signal_5251}), .c ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, LED_128_Instance_state1[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_24_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, LED_128_Instance_state0[24]}), .a ({new_AGEMA_signal_5271, new_AGEMA_signal_5267, new_AGEMA_signal_5263}), .c ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, LED_128_Instance_state1[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_25_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, LED_128_Instance_state0[25]}), .a ({new_AGEMA_signal_5283, new_AGEMA_signal_5279, new_AGEMA_signal_5275}), .c ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, LED_128_Instance_state1[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_26_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, LED_128_Instance_state0[26]}), .a ({new_AGEMA_signal_5295, new_AGEMA_signal_5291, new_AGEMA_signal_5287}), .c ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, LED_128_Instance_state1[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_27_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, LED_128_Instance_state0[27]}), .a ({new_AGEMA_signal_5307, new_AGEMA_signal_5303, new_AGEMA_signal_5299}), .c ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, LED_128_Instance_state1[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_28_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, LED_128_Instance_state0[28]}), .a ({new_AGEMA_signal_5319, new_AGEMA_signal_5315, new_AGEMA_signal_5311}), .c ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, LED_128_Instance_state1[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_29_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, LED_128_Instance_state0[29]}), .a ({new_AGEMA_signal_5331, new_AGEMA_signal_5327, new_AGEMA_signal_5323}), .c ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, LED_128_Instance_state1[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_30_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, LED_128_Instance_state0[30]}), .a ({new_AGEMA_signal_5343, new_AGEMA_signal_5339, new_AGEMA_signal_5335}), .c ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, LED_128_Instance_state1[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_31_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, LED_128_Instance_state0[31]}), .a ({new_AGEMA_signal_5355, new_AGEMA_signal_5351, new_AGEMA_signal_5347}), .c ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, LED_128_Instance_state1[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_32_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3391, new_AGEMA_signal_3390, LED_128_Instance_state0[32]}), .a ({new_AGEMA_signal_5367, new_AGEMA_signal_5363, new_AGEMA_signal_5359}), .c ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, LED_128_Instance_state1[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_33_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, LED_128_Instance_state0[33]}), .a ({new_AGEMA_signal_5379, new_AGEMA_signal_5375, new_AGEMA_signal_5371}), .c ({new_AGEMA_signal_3559, new_AGEMA_signal_3558, LED_128_Instance_state1[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_34_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, LED_128_Instance_state0[34]}), .a ({new_AGEMA_signal_5391, new_AGEMA_signal_5387, new_AGEMA_signal_5383}), .c ({new_AGEMA_signal_3499, new_AGEMA_signal_3498, LED_128_Instance_state1[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_35_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, LED_128_Instance_state0[35]}), .a ({new_AGEMA_signal_5403, new_AGEMA_signal_5399, new_AGEMA_signal_5395}), .c ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, LED_128_Instance_state1[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_36_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, LED_128_Instance_state0[36]}), .a ({new_AGEMA_signal_5415, new_AGEMA_signal_5411, new_AGEMA_signal_5407}), .c ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, LED_128_Instance_state1[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_37_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, LED_128_Instance_state0[37]}), .a ({new_AGEMA_signal_5427, new_AGEMA_signal_5423, new_AGEMA_signal_5419}), .c ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, LED_128_Instance_state1[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_38_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, LED_128_Instance_state0[38]}), .a ({new_AGEMA_signal_5439, new_AGEMA_signal_5435, new_AGEMA_signal_5431}), .c ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, LED_128_Instance_state1[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_39_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, LED_128_Instance_state0[39]}), .a ({new_AGEMA_signal_5451, new_AGEMA_signal_5447, new_AGEMA_signal_5443}), .c ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, LED_128_Instance_state1[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_40_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, LED_128_Instance_state0[40]}), .a ({new_AGEMA_signal_5463, new_AGEMA_signal_5459, new_AGEMA_signal_5455}), .c ({new_AGEMA_signal_3511, new_AGEMA_signal_3510, LED_128_Instance_state1[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_41_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, LED_128_Instance_state0[41]}), .a ({new_AGEMA_signal_5475, new_AGEMA_signal_5471, new_AGEMA_signal_5467}), .c ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, LED_128_Instance_state1[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_42_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, LED_128_Instance_state0[42]}), .a ({new_AGEMA_signal_5487, new_AGEMA_signal_5483, new_AGEMA_signal_5479}), .c ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, LED_128_Instance_state1[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_43_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3465, new_AGEMA_signal_3464, LED_128_Instance_state0[43]}), .a ({new_AGEMA_signal_5499, new_AGEMA_signal_5495, new_AGEMA_signal_5491}), .c ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, LED_128_Instance_state1[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_44_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, LED_128_Instance_state0[44]}), .a ({new_AGEMA_signal_5511, new_AGEMA_signal_5507, new_AGEMA_signal_5503}), .c ({new_AGEMA_signal_3519, new_AGEMA_signal_3518, LED_128_Instance_state1[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_45_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, LED_128_Instance_state0[45]}), .a ({new_AGEMA_signal_5523, new_AGEMA_signal_5519, new_AGEMA_signal_5515}), .c ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, LED_128_Instance_state1[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_46_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, LED_128_Instance_state0[46]}), .a ({new_AGEMA_signal_5535, new_AGEMA_signal_5531, new_AGEMA_signal_5527}), .c ({new_AGEMA_signal_3523, new_AGEMA_signal_3522, LED_128_Instance_state1[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_47_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, LED_128_Instance_state0[47]}), .a ({new_AGEMA_signal_5547, new_AGEMA_signal_5543, new_AGEMA_signal_5539}), .c ({new_AGEMA_signal_3571, new_AGEMA_signal_3570, LED_128_Instance_state1[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_48_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, LED_128_Instance_state0[48]}), .a ({new_AGEMA_signal_5559, new_AGEMA_signal_5555, new_AGEMA_signal_5551}), .c ({new_AGEMA_signal_3683, new_AGEMA_signal_3682, LED_128_Instance_state1[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_49_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, LED_128_Instance_state0[49]}), .a ({new_AGEMA_signal_5571, new_AGEMA_signal_5567, new_AGEMA_signal_5563}), .c ({new_AGEMA_signal_3699, new_AGEMA_signal_3698, LED_128_Instance_state1[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_50_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3547, new_AGEMA_signal_3546, LED_128_Instance_state0[50]}), .a ({new_AGEMA_signal_5583, new_AGEMA_signal_5579, new_AGEMA_signal_5575}), .c ({new_AGEMA_signal_3607, new_AGEMA_signal_3606, LED_128_Instance_state1[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_51_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, LED_128_Instance_state0[51]}), .a ({new_AGEMA_signal_5595, new_AGEMA_signal_5591, new_AGEMA_signal_5587}), .c ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, LED_128_Instance_state1[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_52_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3659, new_AGEMA_signal_3658, LED_128_Instance_state0[52]}), .a ({new_AGEMA_signal_5607, new_AGEMA_signal_5603, new_AGEMA_signal_5599}), .c ({new_AGEMA_signal_3687, new_AGEMA_signal_3686, LED_128_Instance_state1[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_53_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3679, new_AGEMA_signal_3678, LED_128_Instance_state0[53]}), .a ({new_AGEMA_signal_5619, new_AGEMA_signal_5615, new_AGEMA_signal_5611}), .c ({new_AGEMA_signal_3703, new_AGEMA_signal_3702, LED_128_Instance_state1[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_54_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3471, new_AGEMA_signal_3470, LED_128_Instance_state0[54]}), .a ({new_AGEMA_signal_5631, new_AGEMA_signal_5627, new_AGEMA_signal_5623}), .c ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, LED_128_Instance_state1[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_55_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, LED_128_Instance_state0[55]}), .a ({new_AGEMA_signal_5643, new_AGEMA_signal_5639, new_AGEMA_signal_5635}), .c ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, LED_128_Instance_state1[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_56_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, LED_128_Instance_state0[56]}), .a ({new_AGEMA_signal_5655, new_AGEMA_signal_5651, new_AGEMA_signal_5647}), .c ({new_AGEMA_signal_3667, new_AGEMA_signal_3666, LED_128_Instance_state1[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_57_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3661, new_AGEMA_signal_3660, LED_128_Instance_state0[57]}), .a ({new_AGEMA_signal_5667, new_AGEMA_signal_5663, new_AGEMA_signal_5659}), .c ({new_AGEMA_signal_3691, new_AGEMA_signal_3690, LED_128_Instance_state1[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_58_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, LED_128_Instance_state0[58]}), .a ({new_AGEMA_signal_5679, new_AGEMA_signal_5675, new_AGEMA_signal_5671}), .c ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, LED_128_Instance_state1[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_59_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, LED_128_Instance_state0[59]}), .a ({new_AGEMA_signal_5691, new_AGEMA_signal_5687, new_AGEMA_signal_5683}), .c ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, LED_128_Instance_state1[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_60_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3643, new_AGEMA_signal_3642, LED_128_Instance_state0[60]}), .a ({new_AGEMA_signal_5703, new_AGEMA_signal_5699, new_AGEMA_signal_5695}), .c ({new_AGEMA_signal_3671, new_AGEMA_signal_3670, LED_128_Instance_state1[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_61_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, LED_128_Instance_state0[61]}), .a ({new_AGEMA_signal_5715, new_AGEMA_signal_5711, new_AGEMA_signal_5707}), .c ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, LED_128_Instance_state1[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_62_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, LED_128_Instance_state0[62]}), .a ({new_AGEMA_signal_5727, new_AGEMA_signal_5723, new_AGEMA_signal_5719}), .c ({new_AGEMA_signal_3619, new_AGEMA_signal_3618, LED_128_Instance_state1[62]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_63_U1 ( .s (new_AGEMA_signal_4971), .b ({new_AGEMA_signal_3555, new_AGEMA_signal_3554, LED_128_Instance_state0[63]}), .a ({new_AGEMA_signal_5739, new_AGEMA_signal_5735, new_AGEMA_signal_5731}), .c ({new_AGEMA_signal_3623, new_AGEMA_signal_3622, LED_128_Instance_state1[63]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_AND2_U1 ( .a ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, LED_128_Instance_SBox_Instance_0_Q2}), .b ({new_AGEMA_signal_5745, new_AGEMA_signal_5743, new_AGEMA_signal_5741}), .clk (CLK), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, LED_128_Instance_SBox_Instance_0_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_AND4_U1 ( .a ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, LED_128_Instance_SBox_Instance_0_Q6}), .b ({new_AGEMA_signal_5751, new_AGEMA_signal_5749, new_AGEMA_signal_5747}), .clk (CLK), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, LED_128_Instance_SBox_Instance_0_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR10_U1 ( .a ({new_AGEMA_signal_5757, new_AGEMA_signal_5755, new_AGEMA_signal_5753}), .b ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, LED_128_Instance_SBox_Instance_0_T3}), .c ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, LED_128_Instance_SBox_Instance_0_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR11_U1 ( .a ({new_AGEMA_signal_5769, new_AGEMA_signal_5765, new_AGEMA_signal_5761}), .b ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, LED_128_Instance_SBox_Instance_0_L7}), .c ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, LED_128_Instance_subcells_out[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR12_U1 ( .a ({new_AGEMA_signal_5757, new_AGEMA_signal_5755, new_AGEMA_signal_5753}), .b ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, LED_128_Instance_SBox_Instance_0_T1}), .c ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, LED_128_Instance_SBox_Instance_0_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR13_U1 ( .a ({new_AGEMA_signal_5781, new_AGEMA_signal_5777, new_AGEMA_signal_5773}), .b ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, LED_128_Instance_SBox_Instance_0_L8}), .c ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, LED_128_Instance_subcells_out[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR14_U1 ( .a ({new_AGEMA_signal_5787, new_AGEMA_signal_5785, new_AGEMA_signal_5783}), .b ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, LED_128_Instance_SBox_Instance_0_T3}), .c ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, LED_128_Instance_subcells_out[1]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_AND2_U1 ( .a ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, LED_128_Instance_SBox_Instance_1_Q2}), .b ({new_AGEMA_signal_5793, new_AGEMA_signal_5791, new_AGEMA_signal_5789}), .clk (CLK), .r ({Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, LED_128_Instance_SBox_Instance_1_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_AND4_U1 ( .a ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, LED_128_Instance_SBox_Instance_1_Q6}), .b ({new_AGEMA_signal_5799, new_AGEMA_signal_5797, new_AGEMA_signal_5795}), .clk (CLK), .r ({Fresh[107], Fresh[106], Fresh[105]}), .c ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, LED_128_Instance_SBox_Instance_1_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR10_U1 ( .a ({new_AGEMA_signal_5805, new_AGEMA_signal_5803, new_AGEMA_signal_5801}), .b ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, LED_128_Instance_SBox_Instance_1_T3}), .c ({new_AGEMA_signal_2815, new_AGEMA_signal_2814, LED_128_Instance_SBox_Instance_1_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR11_U1 ( .a ({new_AGEMA_signal_5817, new_AGEMA_signal_5813, new_AGEMA_signal_5809}), .b ({new_AGEMA_signal_2815, new_AGEMA_signal_2814, LED_128_Instance_SBox_Instance_1_L7}), .c ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, LED_128_Instance_subcells_out[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR12_U1 ( .a ({new_AGEMA_signal_5805, new_AGEMA_signal_5803, new_AGEMA_signal_5801}), .b ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, LED_128_Instance_SBox_Instance_1_T1}), .c ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, LED_128_Instance_SBox_Instance_1_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR13_U1 ( .a ({new_AGEMA_signal_5829, new_AGEMA_signal_5825, new_AGEMA_signal_5821}), .b ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, LED_128_Instance_SBox_Instance_1_L8}), .c ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, LED_128_Instance_subcells_out[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR14_U1 ( .a ({new_AGEMA_signal_5835, new_AGEMA_signal_5833, new_AGEMA_signal_5831}), .b ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, LED_128_Instance_SBox_Instance_1_T3}), .c ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, LED_128_Instance_subcells_out[5]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_AND2_U1 ( .a ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, LED_128_Instance_SBox_Instance_2_Q2}), .b ({new_AGEMA_signal_5841, new_AGEMA_signal_5839, new_AGEMA_signal_5837}), .clk (CLK), .r ({Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, LED_128_Instance_SBox_Instance_2_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_AND4_U1 ( .a ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, LED_128_Instance_SBox_Instance_2_Q6}), .b ({new_AGEMA_signal_5847, new_AGEMA_signal_5845, new_AGEMA_signal_5843}), .clk (CLK), .r ({Fresh[113], Fresh[112], Fresh[111]}), .c ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, LED_128_Instance_SBox_Instance_2_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR10_U1 ( .a ({new_AGEMA_signal_5853, new_AGEMA_signal_5851, new_AGEMA_signal_5849}), .b ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, LED_128_Instance_SBox_Instance_2_T3}), .c ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, LED_128_Instance_SBox_Instance_2_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR11_U1 ( .a ({new_AGEMA_signal_4303, new_AGEMA_signal_4299, new_AGEMA_signal_4295}), .b ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, LED_128_Instance_SBox_Instance_2_L7}), .c ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, LED_128_Instance_subcells_out[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR12_U1 ( .a ({new_AGEMA_signal_5853, new_AGEMA_signal_5851, new_AGEMA_signal_5849}), .b ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, LED_128_Instance_SBox_Instance_2_T1}), .c ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, LED_128_Instance_SBox_Instance_2_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR13_U1 ( .a ({new_AGEMA_signal_5865, new_AGEMA_signal_5861, new_AGEMA_signal_5857}), .b ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, LED_128_Instance_SBox_Instance_2_L8}), .c ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, LED_128_Instance_subcells_out[10]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR14_U1 ( .a ({new_AGEMA_signal_5871, new_AGEMA_signal_5869, new_AGEMA_signal_5867}), .b ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, LED_128_Instance_SBox_Instance_2_T3}), .c ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, LED_128_Instance_subcells_out[9]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_AND2_U1 ( .a ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, LED_128_Instance_SBox_Instance_3_Q2}), .b ({new_AGEMA_signal_5877, new_AGEMA_signal_5875, new_AGEMA_signal_5873}), .clk (CLK), .r ({Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, LED_128_Instance_SBox_Instance_3_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_AND4_U1 ( .a ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, LED_128_Instance_SBox_Instance_3_Q6}), .b ({new_AGEMA_signal_5883, new_AGEMA_signal_5881, new_AGEMA_signal_5879}), .clk (CLK), .r ({Fresh[119], Fresh[118], Fresh[117]}), .c ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, LED_128_Instance_SBox_Instance_3_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR10_U1 ( .a ({new_AGEMA_signal_5889, new_AGEMA_signal_5887, new_AGEMA_signal_5885}), .b ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, LED_128_Instance_SBox_Instance_3_T3}), .c ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, LED_128_Instance_SBox_Instance_3_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR11_U1 ( .a ({new_AGEMA_signal_4351, new_AGEMA_signal_4347, new_AGEMA_signal_4343}), .b ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, LED_128_Instance_SBox_Instance_3_L7}), .c ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, LED_128_Instance_subcells_out[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR12_U1 ( .a ({new_AGEMA_signal_5889, new_AGEMA_signal_5887, new_AGEMA_signal_5885}), .b ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, LED_128_Instance_SBox_Instance_3_T1}), .c ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, LED_128_Instance_SBox_Instance_3_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR13_U1 ( .a ({new_AGEMA_signal_5901, new_AGEMA_signal_5897, new_AGEMA_signal_5893}), .b ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, LED_128_Instance_SBox_Instance_3_L8}), .c ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, LED_128_Instance_subcells_out[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR14_U1 ( .a ({new_AGEMA_signal_5907, new_AGEMA_signal_5905, new_AGEMA_signal_5903}), .b ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, LED_128_Instance_SBox_Instance_3_T3}), .c ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, LED_128_Instance_subcells_out[13]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_AND2_U1 ( .a ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, LED_128_Instance_SBox_Instance_4_Q2}), .b ({new_AGEMA_signal_5913, new_AGEMA_signal_5911, new_AGEMA_signal_5909}), .clk (CLK), .r ({Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, LED_128_Instance_SBox_Instance_4_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_AND4_U1 ( .a ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, LED_128_Instance_SBox_Instance_4_Q6}), .b ({new_AGEMA_signal_5919, new_AGEMA_signal_5917, new_AGEMA_signal_5915}), .clk (CLK), .r ({Fresh[125], Fresh[124], Fresh[123]}), .c ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, LED_128_Instance_SBox_Instance_4_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR10_U1 ( .a ({new_AGEMA_signal_5925, new_AGEMA_signal_5923, new_AGEMA_signal_5921}), .b ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, LED_128_Instance_SBox_Instance_4_T3}), .c ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, LED_128_Instance_SBox_Instance_4_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR11_U1 ( .a ({new_AGEMA_signal_5937, new_AGEMA_signal_5933, new_AGEMA_signal_5929}), .b ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, LED_128_Instance_SBox_Instance_4_L7}), .c ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, LED_128_Instance_subcells_out[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR12_U1 ( .a ({new_AGEMA_signal_5925, new_AGEMA_signal_5923, new_AGEMA_signal_5921}), .b ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, LED_128_Instance_SBox_Instance_4_T1}), .c ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, LED_128_Instance_SBox_Instance_4_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR13_U1 ( .a ({new_AGEMA_signal_5949, new_AGEMA_signal_5945, new_AGEMA_signal_5941}), .b ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, LED_128_Instance_SBox_Instance_4_L8}), .c ({new_AGEMA_signal_2827, new_AGEMA_signal_2826, LED_128_Instance_subcells_out[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR14_U1 ( .a ({new_AGEMA_signal_5955, new_AGEMA_signal_5953, new_AGEMA_signal_5951}), .b ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, LED_128_Instance_SBox_Instance_4_T3}), .c ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, LED_128_Instance_subcells_out[17]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_AND2_U1 ( .a ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, LED_128_Instance_SBox_Instance_5_Q2}), .b ({new_AGEMA_signal_5961, new_AGEMA_signal_5959, new_AGEMA_signal_5957}), .clk (CLK), .r ({Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, LED_128_Instance_SBox_Instance_5_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_AND4_U1 ( .a ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, LED_128_Instance_SBox_Instance_5_Q6}), .b ({new_AGEMA_signal_5967, new_AGEMA_signal_5965, new_AGEMA_signal_5963}), .clk (CLK), .r ({Fresh[131], Fresh[130], Fresh[129]}), .c ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, LED_128_Instance_SBox_Instance_5_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR10_U1 ( .a ({new_AGEMA_signal_5973, new_AGEMA_signal_5971, new_AGEMA_signal_5969}), .b ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, LED_128_Instance_SBox_Instance_5_T3}), .c ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, LED_128_Instance_SBox_Instance_5_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR11_U1 ( .a ({new_AGEMA_signal_5985, new_AGEMA_signal_5981, new_AGEMA_signal_5977}), .b ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, LED_128_Instance_SBox_Instance_5_L7}), .c ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, LED_128_Instance_subcells_out[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR12_U1 ( .a ({new_AGEMA_signal_5973, new_AGEMA_signal_5971, new_AGEMA_signal_5969}), .b ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, LED_128_Instance_SBox_Instance_5_T1}), .c ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, LED_128_Instance_SBox_Instance_5_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR13_U1 ( .a ({new_AGEMA_signal_5997, new_AGEMA_signal_5993, new_AGEMA_signal_5989}), .b ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, LED_128_Instance_SBox_Instance_5_L8}), .c ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, LED_128_Instance_subcells_out[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR14_U1 ( .a ({new_AGEMA_signal_6003, new_AGEMA_signal_6001, new_AGEMA_signal_5999}), .b ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, LED_128_Instance_SBox_Instance_5_T3}), .c ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, LED_128_Instance_subcells_out[21]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_AND2_U1 ( .a ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, LED_128_Instance_SBox_Instance_6_Q2}), .b ({new_AGEMA_signal_6009, new_AGEMA_signal_6007, new_AGEMA_signal_6005}), .clk (CLK), .r ({Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, LED_128_Instance_SBox_Instance_6_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_AND4_U1 ( .a ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, LED_128_Instance_SBox_Instance_6_Q6}), .b ({new_AGEMA_signal_6015, new_AGEMA_signal_6013, new_AGEMA_signal_6011}), .clk (CLK), .r ({Fresh[137], Fresh[136], Fresh[135]}), .c ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, LED_128_Instance_SBox_Instance_6_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR10_U1 ( .a ({new_AGEMA_signal_6021, new_AGEMA_signal_6019, new_AGEMA_signal_6017}), .b ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, LED_128_Instance_SBox_Instance_6_T3}), .c ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, LED_128_Instance_SBox_Instance_6_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR11_U1 ( .a ({new_AGEMA_signal_4495, new_AGEMA_signal_4491, new_AGEMA_signal_4487}), .b ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, LED_128_Instance_SBox_Instance_6_L7}), .c ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, LED_128_Instance_subcells_out[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR12_U1 ( .a ({new_AGEMA_signal_6021, new_AGEMA_signal_6019, new_AGEMA_signal_6017}), .b ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, LED_128_Instance_SBox_Instance_6_T1}), .c ({new_AGEMA_signal_2691, new_AGEMA_signal_2690, LED_128_Instance_SBox_Instance_6_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR13_U1 ( .a ({new_AGEMA_signal_6033, new_AGEMA_signal_6029, new_AGEMA_signal_6025}), .b ({new_AGEMA_signal_2691, new_AGEMA_signal_2690, LED_128_Instance_SBox_Instance_6_L8}), .c ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, LED_128_Instance_subcells_out[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR14_U1 ( .a ({new_AGEMA_signal_6039, new_AGEMA_signal_6037, new_AGEMA_signal_6035}), .b ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, LED_128_Instance_SBox_Instance_6_T3}), .c ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, LED_128_Instance_subcells_out[25]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_AND2_U1 ( .a ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, LED_128_Instance_SBox_Instance_7_Q2}), .b ({new_AGEMA_signal_6045, new_AGEMA_signal_6043, new_AGEMA_signal_6041}), .clk (CLK), .r ({Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, LED_128_Instance_SBox_Instance_7_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_AND4_U1 ( .a ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, LED_128_Instance_SBox_Instance_7_Q6}), .b ({new_AGEMA_signal_6051, new_AGEMA_signal_6049, new_AGEMA_signal_6047}), .clk (CLK), .r ({Fresh[143], Fresh[142], Fresh[141]}), .c ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, LED_128_Instance_SBox_Instance_7_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR10_U1 ( .a ({new_AGEMA_signal_6057, new_AGEMA_signal_6055, new_AGEMA_signal_6053}), .b ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, LED_128_Instance_SBox_Instance_7_T3}), .c ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, LED_128_Instance_SBox_Instance_7_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR11_U1 ( .a ({new_AGEMA_signal_4543, new_AGEMA_signal_4539, new_AGEMA_signal_4535}), .b ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, LED_128_Instance_SBox_Instance_7_L7}), .c ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, LED_128_Instance_subcells_out[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR12_U1 ( .a ({new_AGEMA_signal_6057, new_AGEMA_signal_6055, new_AGEMA_signal_6053}), .b ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, LED_128_Instance_SBox_Instance_7_T1}), .c ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, LED_128_Instance_SBox_Instance_7_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR13_U1 ( .a ({new_AGEMA_signal_6069, new_AGEMA_signal_6065, new_AGEMA_signal_6061}), .b ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, LED_128_Instance_SBox_Instance_7_L8}), .c ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, LED_128_Instance_subcells_out[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR14_U1 ( .a ({new_AGEMA_signal_6075, new_AGEMA_signal_6073, new_AGEMA_signal_6071}), .b ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, LED_128_Instance_SBox_Instance_7_T3}), .c ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, LED_128_Instance_subcells_out[29]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_AND2_U1 ( .a ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, LED_128_Instance_SBox_Instance_8_Q2}), .b ({new_AGEMA_signal_6081, new_AGEMA_signal_6079, new_AGEMA_signal_6077}), .clk (CLK), .r ({Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, LED_128_Instance_SBox_Instance_8_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_AND4_U1 ( .a ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, LED_128_Instance_SBox_Instance_8_Q6}), .b ({new_AGEMA_signal_6087, new_AGEMA_signal_6085, new_AGEMA_signal_6083}), .clk (CLK), .r ({Fresh[149], Fresh[148], Fresh[147]}), .c ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, LED_128_Instance_SBox_Instance_8_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR10_U1 ( .a ({new_AGEMA_signal_6093, new_AGEMA_signal_6091, new_AGEMA_signal_6089}), .b ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, LED_128_Instance_SBox_Instance_8_T3}), .c ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, LED_128_Instance_SBox_Instance_8_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR11_U1 ( .a ({new_AGEMA_signal_6105, new_AGEMA_signal_6101, new_AGEMA_signal_6097}), .b ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, LED_128_Instance_SBox_Instance_8_L7}), .c ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, LED_128_Instance_subcells_out[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR12_U1 ( .a ({new_AGEMA_signal_6093, new_AGEMA_signal_6091, new_AGEMA_signal_6089}), .b ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, LED_128_Instance_SBox_Instance_8_T1}), .c ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, LED_128_Instance_SBox_Instance_8_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR13_U1 ( .a ({new_AGEMA_signal_6117, new_AGEMA_signal_6113, new_AGEMA_signal_6109}), .b ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, LED_128_Instance_SBox_Instance_8_L8}), .c ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, LED_128_Instance_subcells_out[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR14_U1 ( .a ({new_AGEMA_signal_6123, new_AGEMA_signal_6121, new_AGEMA_signal_6119}), .b ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, LED_128_Instance_SBox_Instance_8_T3}), .c ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, LED_128_Instance_subcells_out[33]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_AND2_U1 ( .a ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, LED_128_Instance_SBox_Instance_9_Q2}), .b ({new_AGEMA_signal_6129, new_AGEMA_signal_6127, new_AGEMA_signal_6125}), .clk (CLK), .r ({Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, LED_128_Instance_SBox_Instance_9_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_AND4_U1 ( .a ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, LED_128_Instance_SBox_Instance_9_Q6}), .b ({new_AGEMA_signal_6135, new_AGEMA_signal_6133, new_AGEMA_signal_6131}), .clk (CLK), .r ({Fresh[155], Fresh[154], Fresh[153]}), .c ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, LED_128_Instance_SBox_Instance_9_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR10_U1 ( .a ({new_AGEMA_signal_6141, new_AGEMA_signal_6139, new_AGEMA_signal_6137}), .b ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, LED_128_Instance_SBox_Instance_9_T3}), .c ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, LED_128_Instance_SBox_Instance_9_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR11_U1 ( .a ({new_AGEMA_signal_6153, new_AGEMA_signal_6149, new_AGEMA_signal_6145}), .b ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, LED_128_Instance_SBox_Instance_9_L7}), .c ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, LED_128_Instance_subcells_out[39]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR12_U1 ( .a ({new_AGEMA_signal_6141, new_AGEMA_signal_6139, new_AGEMA_signal_6137}), .b ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, LED_128_Instance_SBox_Instance_9_T1}), .c ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, LED_128_Instance_SBox_Instance_9_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR13_U1 ( .a ({new_AGEMA_signal_6165, new_AGEMA_signal_6161, new_AGEMA_signal_6157}), .b ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, LED_128_Instance_SBox_Instance_9_L8}), .c ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, LED_128_Instance_subcells_out[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR14_U1 ( .a ({new_AGEMA_signal_6171, new_AGEMA_signal_6169, new_AGEMA_signal_6167}), .b ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, LED_128_Instance_SBox_Instance_9_T3}), .c ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, LED_128_Instance_subcells_out[37]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_AND2_U1 ( .a ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, LED_128_Instance_SBox_Instance_10_Q2}), .b ({new_AGEMA_signal_6177, new_AGEMA_signal_6175, new_AGEMA_signal_6173}), .clk (CLK), .r ({Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, LED_128_Instance_SBox_Instance_10_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_AND4_U1 ( .a ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, LED_128_Instance_SBox_Instance_10_Q6}), .b ({new_AGEMA_signal_6183, new_AGEMA_signal_6181, new_AGEMA_signal_6179}), .clk (CLK), .r ({Fresh[161], Fresh[160], Fresh[159]}), .c ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, LED_128_Instance_SBox_Instance_10_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR10_U1 ( .a ({new_AGEMA_signal_6189, new_AGEMA_signal_6187, new_AGEMA_signal_6185}), .b ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, LED_128_Instance_SBox_Instance_10_T3}), .c ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, LED_128_Instance_SBox_Instance_10_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR11_U1 ( .a ({new_AGEMA_signal_4687, new_AGEMA_signal_4683, new_AGEMA_signal_4679}), .b ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, LED_128_Instance_SBox_Instance_10_L7}), .c ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, LED_128_Instance_subcells_out[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR12_U1 ( .a ({new_AGEMA_signal_6189, new_AGEMA_signal_6187, new_AGEMA_signal_6185}), .b ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, LED_128_Instance_SBox_Instance_10_T1}), .c ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, LED_128_Instance_SBox_Instance_10_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR13_U1 ( .a ({new_AGEMA_signal_6201, new_AGEMA_signal_6197, new_AGEMA_signal_6193}), .b ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, LED_128_Instance_SBox_Instance_10_L8}), .c ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, LED_128_Instance_subcells_out[42]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR14_U1 ( .a ({new_AGEMA_signal_6207, new_AGEMA_signal_6205, new_AGEMA_signal_6203}), .b ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, LED_128_Instance_SBox_Instance_10_T3}), .c ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, LED_128_Instance_subcells_out[41]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_AND2_U1 ( .a ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, LED_128_Instance_SBox_Instance_11_Q2}), .b ({new_AGEMA_signal_6213, new_AGEMA_signal_6211, new_AGEMA_signal_6209}), .clk (CLK), .r ({Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, LED_128_Instance_SBox_Instance_11_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_AND4_U1 ( .a ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, LED_128_Instance_SBox_Instance_11_Q6}), .b ({new_AGEMA_signal_6219, new_AGEMA_signal_6217, new_AGEMA_signal_6215}), .clk (CLK), .r ({Fresh[167], Fresh[166], Fresh[165]}), .c ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, LED_128_Instance_SBox_Instance_11_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR10_U1 ( .a ({new_AGEMA_signal_6225, new_AGEMA_signal_6223, new_AGEMA_signal_6221}), .b ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, LED_128_Instance_SBox_Instance_11_T3}), .c ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, LED_128_Instance_SBox_Instance_11_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR11_U1 ( .a ({new_AGEMA_signal_4739, new_AGEMA_signal_4735, new_AGEMA_signal_4731}), .b ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, LED_128_Instance_SBox_Instance_11_L7}), .c ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, LED_128_Instance_subcells_out[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR12_U1 ( .a ({new_AGEMA_signal_6225, new_AGEMA_signal_6223, new_AGEMA_signal_6221}), .b ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, LED_128_Instance_SBox_Instance_11_T1}), .c ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, LED_128_Instance_SBox_Instance_11_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR13_U1 ( .a ({new_AGEMA_signal_6237, new_AGEMA_signal_6233, new_AGEMA_signal_6229}), .b ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, LED_128_Instance_SBox_Instance_11_L8}), .c ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, LED_128_Instance_subcells_out[46]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR14_U1 ( .a ({new_AGEMA_signal_6243, new_AGEMA_signal_6241, new_AGEMA_signal_6239}), .b ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, LED_128_Instance_SBox_Instance_11_T3}), .c ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, LED_128_Instance_subcells_out[45]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_AND2_U1 ( .a ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, LED_128_Instance_SBox_Instance_12_Q2}), .b ({new_AGEMA_signal_6249, new_AGEMA_signal_6247, new_AGEMA_signal_6245}), .clk (CLK), .r ({Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, LED_128_Instance_SBox_Instance_12_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_AND4_U1 ( .a ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, LED_128_Instance_SBox_Instance_12_Q6}), .b ({new_AGEMA_signal_6255, new_AGEMA_signal_6253, new_AGEMA_signal_6251}), .clk (CLK), .r ({Fresh[173], Fresh[172], Fresh[171]}), .c ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, LED_128_Instance_SBox_Instance_12_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR10_U1 ( .a ({new_AGEMA_signal_6261, new_AGEMA_signal_6259, new_AGEMA_signal_6257}), .b ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, LED_128_Instance_SBox_Instance_12_T3}), .c ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, LED_128_Instance_SBox_Instance_12_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR11_U1 ( .a ({new_AGEMA_signal_6273, new_AGEMA_signal_6269, new_AGEMA_signal_6265}), .b ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, LED_128_Instance_SBox_Instance_12_L7}), .c ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, LED_128_Instance_subcells_out[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR12_U1 ( .a ({new_AGEMA_signal_6261, new_AGEMA_signal_6259, new_AGEMA_signal_6257}), .b ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, LED_128_Instance_SBox_Instance_12_T1}), .c ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, LED_128_Instance_SBox_Instance_12_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR13_U1 ( .a ({new_AGEMA_signal_6285, new_AGEMA_signal_6281, new_AGEMA_signal_6277}), .b ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, LED_128_Instance_SBox_Instance_12_L8}), .c ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, LED_128_Instance_subcells_out[50]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR14_U1 ( .a ({new_AGEMA_signal_6291, new_AGEMA_signal_6289, new_AGEMA_signal_6287}), .b ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, LED_128_Instance_SBox_Instance_12_T3}), .c ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, LED_128_Instance_subcells_out[49]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_AND2_U1 ( .a ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, LED_128_Instance_SBox_Instance_13_Q2}), .b ({new_AGEMA_signal_6297, new_AGEMA_signal_6295, new_AGEMA_signal_6293}), .clk (CLK), .r ({Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, LED_128_Instance_SBox_Instance_13_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_AND4_U1 ( .a ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, LED_128_Instance_SBox_Instance_13_Q6}), .b ({new_AGEMA_signal_6303, new_AGEMA_signal_6301, new_AGEMA_signal_6299}), .clk (CLK), .r ({Fresh[179], Fresh[178], Fresh[177]}), .c ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, LED_128_Instance_SBox_Instance_13_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR10_U1 ( .a ({new_AGEMA_signal_6309, new_AGEMA_signal_6307, new_AGEMA_signal_6305}), .b ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, LED_128_Instance_SBox_Instance_13_T3}), .c ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, LED_128_Instance_SBox_Instance_13_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR11_U1 ( .a ({new_AGEMA_signal_6321, new_AGEMA_signal_6317, new_AGEMA_signal_6313}), .b ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, LED_128_Instance_SBox_Instance_13_L7}), .c ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, LED_128_Instance_subcells_out[55]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR12_U1 ( .a ({new_AGEMA_signal_6309, new_AGEMA_signal_6307, new_AGEMA_signal_6305}), .b ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, LED_128_Instance_SBox_Instance_13_T1}), .c ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, LED_128_Instance_SBox_Instance_13_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR13_U1 ( .a ({new_AGEMA_signal_6333, new_AGEMA_signal_6329, new_AGEMA_signal_6325}), .b ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, LED_128_Instance_SBox_Instance_13_L8}), .c ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, LED_128_Instance_subcells_out[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR14_U1 ( .a ({new_AGEMA_signal_6339, new_AGEMA_signal_6337, new_AGEMA_signal_6335}), .b ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, LED_128_Instance_SBox_Instance_13_T3}), .c ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, LED_128_Instance_subcells_out[53]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_AND2_U1 ( .a ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, LED_128_Instance_SBox_Instance_14_Q2}), .b ({new_AGEMA_signal_6345, new_AGEMA_signal_6343, new_AGEMA_signal_6341}), .clk (CLK), .r ({Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, LED_128_Instance_SBox_Instance_14_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_AND4_U1 ( .a ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, LED_128_Instance_SBox_Instance_14_Q6}), .b ({new_AGEMA_signal_6351, new_AGEMA_signal_6349, new_AGEMA_signal_6347}), .clk (CLK), .r ({Fresh[185], Fresh[184], Fresh[183]}), .c ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, LED_128_Instance_SBox_Instance_14_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR10_U1 ( .a ({new_AGEMA_signal_6357, new_AGEMA_signal_6355, new_AGEMA_signal_6353}), .b ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, LED_128_Instance_SBox_Instance_14_T3}), .c ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, LED_128_Instance_SBox_Instance_14_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR11_U1 ( .a ({new_AGEMA_signal_4883, new_AGEMA_signal_4879, new_AGEMA_signal_4875}), .b ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, LED_128_Instance_SBox_Instance_14_L7}), .c ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, LED_128_Instance_subcells_out[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR12_U1 ( .a ({new_AGEMA_signal_6357, new_AGEMA_signal_6355, new_AGEMA_signal_6353}), .b ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, LED_128_Instance_SBox_Instance_14_T1}), .c ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, LED_128_Instance_SBox_Instance_14_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR13_U1 ( .a ({new_AGEMA_signal_6369, new_AGEMA_signal_6365, new_AGEMA_signal_6361}), .b ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, LED_128_Instance_SBox_Instance_14_L8}), .c ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, LED_128_Instance_subcells_out[58]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR14_U1 ( .a ({new_AGEMA_signal_6375, new_AGEMA_signal_6373, new_AGEMA_signal_6371}), .b ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, LED_128_Instance_SBox_Instance_14_T3}), .c ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, LED_128_Instance_subcells_out[57]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_AND2_U1 ( .a ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, LED_128_Instance_SBox_Instance_15_Q2}), .b ({new_AGEMA_signal_6381, new_AGEMA_signal_6379, new_AGEMA_signal_6377}), .clk (CLK), .r ({Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, LED_128_Instance_SBox_Instance_15_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_AND4_U1 ( .a ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, LED_128_Instance_SBox_Instance_15_Q6}), .b ({new_AGEMA_signal_6387, new_AGEMA_signal_6385, new_AGEMA_signal_6383}), .clk (CLK), .r ({Fresh[191], Fresh[190], Fresh[189]}), .c ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, LED_128_Instance_SBox_Instance_15_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR10_U1 ( .a ({new_AGEMA_signal_6393, new_AGEMA_signal_6391, new_AGEMA_signal_6389}), .b ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, LED_128_Instance_SBox_Instance_15_T3}), .c ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, LED_128_Instance_SBox_Instance_15_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR11_U1 ( .a ({new_AGEMA_signal_4931, new_AGEMA_signal_4927, new_AGEMA_signal_4923}), .b ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, LED_128_Instance_SBox_Instance_15_L7}), .c ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, LED_128_Instance_subcells_out[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR12_U1 ( .a ({new_AGEMA_signal_6393, new_AGEMA_signal_6391, new_AGEMA_signal_6389}), .b ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, LED_128_Instance_SBox_Instance_15_T1}), .c ({new_AGEMA_signal_2727, new_AGEMA_signal_2726, LED_128_Instance_SBox_Instance_15_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR13_U1 ( .a ({new_AGEMA_signal_6405, new_AGEMA_signal_6401, new_AGEMA_signal_6397}), .b ({new_AGEMA_signal_2727, new_AGEMA_signal_2726, LED_128_Instance_SBox_Instance_15_L8}), .c ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, LED_128_Instance_subcells_out[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR14_U1 ( .a ({new_AGEMA_signal_6411, new_AGEMA_signal_6409, new_AGEMA_signal_6407}), .b ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, LED_128_Instance_SBox_Instance_15_T3}), .c ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, LED_128_Instance_subcells_out[61]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U54 ( .a ({new_AGEMA_signal_3439, new_AGEMA_signal_3438, LED_128_Instance_MCS_Instance_0_n38}), .b ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, LED_128_Instance_MCS_Instance_0_n37}), .c ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, LED_128_Instance_mixcolumns_out[51]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U53 ( .a ({new_AGEMA_signal_3083, new_AGEMA_signal_3082, LED_128_Instance_mixcolumns_out[3]}), .b ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, LED_128_Instance_subcells_out[61]}), .c ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, LED_128_Instance_MCS_Instance_0_n37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U52 ( .a ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, LED_128_Instance_mixcolumns_out[34]}), .b ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, LED_128_Instance_mixcolumns_out[18]}), .c ({new_AGEMA_signal_3439, new_AGEMA_signal_3438, LED_128_Instance_MCS_Instance_0_n38}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U51 ( .a ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, LED_128_Instance_MCS_Instance_0_n36}), .b ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, LED_128_Instance_MCS_Instance_0_n35}), .c ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, LED_128_Instance_mixcolumns_out[34]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U50 ( .a ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, LED_128_Instance_subcells_out[62]}), .b ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, LED_128_Instance_MCS_Instance_0_n34}), .c ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, LED_128_Instance_MCS_Instance_0_n36}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U49 ( .a ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, LED_128_Instance_MCS_Instance_0_n33}), .b ({new_AGEMA_signal_3443, new_AGEMA_signal_3442, LED_128_Instance_mixcolumns_out[33]}), .c ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, LED_128_Instance_mixcolumns_out[50]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U48 ( .a ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, LED_128_Instance_mixcolumns_out[2]}), .b ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, LED_128_Instance_MCS_Instance_0_n35}), .c ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, LED_128_Instance_MCS_Instance_0_n33}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U47 ( .a ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, LED_128_Instance_MCS_Instance_0_n32}), .b ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, LED_128_Instance_MCS_Instance_0_n31}), .c ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, LED_128_Instance_mixcolumns_out[49]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U46 ( .a ({new_AGEMA_signal_3625, new_AGEMA_signal_3624, LED_128_Instance_MCS_Instance_0_n30}), .b ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, LED_128_Instance_MCS_Instance_0_n29}), .c ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, LED_128_Instance_MCS_Instance_0_n32}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U45 ( .a ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, LED_128_Instance_subcells_out[63]}), .b ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, LED_128_Instance_mixcolumns_out[1]}), .c ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, LED_128_Instance_MCS_Instance_0_n29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U44 ( .a ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, LED_128_Instance_mixcolumns_out[32]}), .b ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, LED_128_Instance_MCS_Instance_0_n28}), .c ({new_AGEMA_signal_3625, new_AGEMA_signal_3624, LED_128_Instance_MCS_Instance_0_n30}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U43 ( .a ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, LED_128_Instance_MCS_Instance_0_n27}), .b ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, LED_128_Instance_MCS_Instance_0_n26}), .c ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, LED_128_Instance_mixcolumns_out[32]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U42 ( .a ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, LED_128_Instance_subcells_out[42]}), .b ({new_AGEMA_signal_3083, new_AGEMA_signal_3082, LED_128_Instance_mixcolumns_out[3]}), .c ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, LED_128_Instance_MCS_Instance_0_n26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U41 ( .a ({new_AGEMA_signal_6417, new_AGEMA_signal_6415, new_AGEMA_signal_6413}), .b ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, LED_128_Instance_mixcolumns_out[19]}), .c ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, LED_128_Instance_MCS_Instance_0_n27}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U40 ( .a ({new_AGEMA_signal_3627, new_AGEMA_signal_3626, LED_128_Instance_MCS_Instance_0_n25}), .b ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, LED_128_Instance_mixcolumns_out[0]}), .c ({new_AGEMA_signal_3647, new_AGEMA_signal_3646, LED_128_Instance_mixcolumns_out[48]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U39 ( .a ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, LED_128_Instance_mixcolumns_out[19]}), .b ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, LED_128_Instance_MCS_Instance_0_n28}), .c ({new_AGEMA_signal_3627, new_AGEMA_signal_3626, LED_128_Instance_MCS_Instance_0_n25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U38 ( .a ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, LED_128_Instance_subcells_out[62]}), .b ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, LED_128_Instance_mixcolumns_out[35]}), .c ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, LED_128_Instance_MCS_Instance_0_n28}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U37 ( .a ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, LED_128_Instance_MCS_Instance_0_n24}), .b ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, LED_128_Instance_MCS_Instance_0_n23}), .c ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, LED_128_Instance_mixcolumns_out[35]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U36 ( .a ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, LED_128_Instance_subcells_out[63]}), .b ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, LED_128_Instance_subcells_out[41]}), .c ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, LED_128_Instance_MCS_Instance_0_n23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U35 ( .a ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, LED_128_Instance_mixcolumns_out[18]}), .b ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, LED_128_Instance_mixcolumns_out[2]}), .c ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, LED_128_Instance_MCS_Instance_0_n24}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U34 ( .a ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, LED_128_Instance_MCS_Instance_0_n22}), .b ({new_AGEMA_signal_3017, new_AGEMA_signal_3016, LED_128_Instance_MCS_Instance_0_n21}), .c ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, LED_128_Instance_mixcolumns_out[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U33 ( .a ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, LED_128_Instance_MCS_Instance_0_n20}), .b ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, LED_128_Instance_subcells_out[61]}), .c ({new_AGEMA_signal_3017, new_AGEMA_signal_3016, LED_128_Instance_MCS_Instance_0_n21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U32 ( .a ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, LED_128_Instance_mixcolumns_out[1]}), .b ({new_AGEMA_signal_6423, new_AGEMA_signal_6421, new_AGEMA_signal_6419}), .c ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, LED_128_Instance_MCS_Instance_0_n22}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U31 ( .a ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MCS_Instance_0_n19}), .b ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, LED_128_Instance_MCS_Instance_0_n18}), .c ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, LED_128_Instance_mixcolumns_out[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U30 ( .a ({new_AGEMA_signal_6429, new_AGEMA_signal_6427, new_AGEMA_signal_6425}), .b ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, LED_128_Instance_subcells_out[43]}), .c ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, LED_128_Instance_MCS_Instance_0_n18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U29 ( .a ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, LED_128_Instance_MCS_Instance_0_n17}), .b ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, LED_128_Instance_MCS_Instance_0_n34}), .c ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MCS_Instance_0_n19}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U28 ( .a ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, LED_128_Instance_MCS_Instance_0_n16}), .b ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, LED_128_Instance_subcells_out[2]}), .c ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, LED_128_Instance_MCS_Instance_0_n34}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U27 ( .a ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, LED_128_Instance_subcells_out[21]}), .b ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, LED_128_Instance_subcells_out[3]}), .c ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, LED_128_Instance_MCS_Instance_0_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U26 ( .a ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, LED_128_Instance_MCS_Instance_0_n15}), .b ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, LED_128_Instance_MCS_Instance_0_n31}), .c ({new_AGEMA_signal_3443, new_AGEMA_signal_3442, LED_128_Instance_mixcolumns_out[33]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U25 ( .a ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, LED_128_Instance_mixcolumns_out[16]}), .b ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, LED_128_Instance_mixcolumns_out[19]}), .c ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, LED_128_Instance_MCS_Instance_0_n31}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U24 ( .a ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, LED_128_Instance_MCS_Instance_0_n14}), .b ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, LED_128_Instance_MCS_Instance_0_n13}), .c ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, LED_128_Instance_MCS_Instance_0_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U23 ( .a ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, LED_128_Instance_subcells_out[42]}), .b ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, LED_128_Instance_subcells_out[43]}), .c ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, LED_128_Instance_MCS_Instance_0_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U22 ( .a ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, LED_128_Instance_MCS_Instance_0_n12}), .b ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, LED_128_Instance_subcells_out[61]}), .c ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, LED_128_Instance_MCS_Instance_0_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U21 ( .a ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, LED_128_Instance_MCS_Instance_0_n11}), .b ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, LED_128_Instance_MCS_Instance_0_n10}), .c ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, LED_128_Instance_mixcolumns_out[16]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U20 ( .a ({new_AGEMA_signal_3083, new_AGEMA_signal_3082, LED_128_Instance_mixcolumns_out[3]}), .b ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, LED_128_Instance_subcells_out[63]}), .c ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, LED_128_Instance_MCS_Instance_0_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U19 ( .a ({new_AGEMA_signal_6429, new_AGEMA_signal_6427, new_AGEMA_signal_6425}), .b ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, LED_128_Instance_subcells_out[22]}), .c ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, LED_128_Instance_MCS_Instance_0_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U18 ( .a ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, LED_128_Instance_MCS_Instance_0_n9}), .b ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, LED_128_Instance_MCS_Instance_0_n8}), .c ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, LED_128_Instance_mixcolumns_out[19]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U17 ( .a ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, LED_128_Instance_subcells_out[62]}), .b ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, LED_128_Instance_subcells_out[43]}), .c ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, LED_128_Instance_MCS_Instance_0_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U16 ( .a ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, LED_128_Instance_mixcolumns_out[2]}), .b ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, LED_128_Instance_subcells_out[21]}), .c ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, LED_128_Instance_MCS_Instance_0_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U15 ( .a ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, LED_128_Instance_MCS_Instance_0_n7}), .b ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, LED_128_Instance_MCS_Instance_0_n6}), .c ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, LED_128_Instance_mixcolumns_out[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U14 ( .a ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, LED_128_Instance_MCS_Instance_0_n5}), .b ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, LED_128_Instance_subcells_out[3]}), .c ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, LED_128_Instance_MCS_Instance_0_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U13 ( .a ({new_AGEMA_signal_6435, new_AGEMA_signal_6433, new_AGEMA_signal_6431}), .b ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, LED_128_Instance_subcells_out[61]}), .c ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, LED_128_Instance_MCS_Instance_0_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U12 ( .a ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, LED_128_Instance_MCS_Instance_0_n17}), .b ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, LED_128_Instance_MCS_Instance_0_n35}), .c ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, LED_128_Instance_mixcolumns_out[17]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U11 ( .a ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, LED_128_Instance_MCS_Instance_0_n4}), .b ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, LED_128_Instance_MCS_Instance_0_n12}), .c ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, LED_128_Instance_MCS_Instance_0_n35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U10 ( .a ({new_AGEMA_signal_3083, new_AGEMA_signal_3082, LED_128_Instance_mixcolumns_out[3]}), .b ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, LED_128_Instance_mixcolumns_out[0]}), .c ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, LED_128_Instance_MCS_Instance_0_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U9 ( .a ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, LED_128_Instance_subcells_out[23]}), .b ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, LED_128_Instance_MCS_Instance_0_n5}), .c ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, LED_128_Instance_MCS_Instance_0_n4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U8 ( .a ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, LED_128_Instance_subcells_out[22]}), .b ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, LED_128_Instance_subcells_out[41]}), .c ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, LED_128_Instance_MCS_Instance_0_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U7 ( .a ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, LED_128_Instance_subcells_out[63]}), .b ({new_AGEMA_signal_6417, new_AGEMA_signal_6415, new_AGEMA_signal_6413}), .c ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, LED_128_Instance_MCS_Instance_0_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U6 ( .a ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, LED_128_Instance_MCS_Instance_0_n3}), .b ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, LED_128_Instance_MCS_Instance_0_n2}), .c ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, LED_128_Instance_mixcolumns_out[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U5 ( .a ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, LED_128_Instance_subcells_out[63]}), .b ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, LED_128_Instance_subcells_out[43]}), .c ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, LED_128_Instance_MCS_Instance_0_n2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U4 ( .a ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, LED_128_Instance_subcells_out[2]}), .b ({new_AGEMA_signal_6423, new_AGEMA_signal_6421, new_AGEMA_signal_6419}), .c ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, LED_128_Instance_MCS_Instance_0_n3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U3 ( .a ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, LED_128_Instance_MCS_Instance_0_n1}), .b ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, LED_128_Instance_subcells_out[62]}), .c ({new_AGEMA_signal_3083, new_AGEMA_signal_3082, LED_128_Instance_mixcolumns_out[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U2 ( .a ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, LED_128_Instance_MCS_Instance_0_n20}), .b ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, LED_128_Instance_subcells_out[1]}), .c ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, LED_128_Instance_MCS_Instance_0_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U1 ( .a ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, LED_128_Instance_subcells_out[42]}), .b ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, LED_128_Instance_subcells_out[23]}), .c ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, LED_128_Instance_MCS_Instance_0_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U54 ( .a ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, LED_128_Instance_MCS_Instance_1_n38}), .b ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, LED_128_Instance_MCS_Instance_1_n37}), .c ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, LED_128_Instance_mixcolumns_out[55]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U53 ( .a ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, LED_128_Instance_mixcolumns_out[7]}), .b ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, LED_128_Instance_subcells_out[49]}), .c ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, LED_128_Instance_MCS_Instance_1_n37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U52 ( .a ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, LED_128_Instance_mixcolumns_out[38]}), .b ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, LED_128_Instance_mixcolumns_out[22]}), .c ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, LED_128_Instance_MCS_Instance_1_n38}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U51 ( .a ({new_AGEMA_signal_3087, new_AGEMA_signal_3086, LED_128_Instance_MCS_Instance_1_n36}), .b ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, LED_128_Instance_MCS_Instance_1_n35}), .c ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, LED_128_Instance_mixcolumns_out[38]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U50 ( .a ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, LED_128_Instance_subcells_out[50]}), .b ({new_AGEMA_signal_3025, new_AGEMA_signal_3024, LED_128_Instance_MCS_Instance_1_n34}), .c ({new_AGEMA_signal_3087, new_AGEMA_signal_3086, LED_128_Instance_MCS_Instance_1_n36}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U49 ( .a ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, LED_128_Instance_MCS_Instance_1_n33}), .b ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, LED_128_Instance_mixcolumns_out[37]}), .c ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, LED_128_Instance_mixcolumns_out[54]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U48 ( .a ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, LED_128_Instance_mixcolumns_out[6]}), .b ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, LED_128_Instance_MCS_Instance_1_n35}), .c ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, LED_128_Instance_MCS_Instance_1_n33}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U47 ( .a ({new_AGEMA_signal_3649, new_AGEMA_signal_3648, LED_128_Instance_MCS_Instance_1_n32}), .b ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, LED_128_Instance_MCS_Instance_1_n31}), .c ({new_AGEMA_signal_3675, new_AGEMA_signal_3674, LED_128_Instance_mixcolumns_out[53]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U46 ( .a ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, LED_128_Instance_MCS_Instance_1_n30}), .b ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, LED_128_Instance_MCS_Instance_1_n29}), .c ({new_AGEMA_signal_3649, new_AGEMA_signal_3648, LED_128_Instance_MCS_Instance_1_n32}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U45 ( .a ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, LED_128_Instance_subcells_out[51]}), .b ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, LED_128_Instance_mixcolumns_out[5]}), .c ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, LED_128_Instance_MCS_Instance_1_n29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U44 ( .a ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, LED_128_Instance_mixcolumns_out[36]}), .b ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, LED_128_Instance_MCS_Instance_1_n28}), .c ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, LED_128_Instance_MCS_Instance_1_n30}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U43 ( .a ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, LED_128_Instance_MCS_Instance_1_n27}), .b ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, LED_128_Instance_MCS_Instance_1_n26}), .c ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, LED_128_Instance_mixcolumns_out[36]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U42 ( .a ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, LED_128_Instance_subcells_out[46]}), .b ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, LED_128_Instance_mixcolumns_out[7]}), .c ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, LED_128_Instance_MCS_Instance_1_n26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U41 ( .a ({new_AGEMA_signal_6441, new_AGEMA_signal_6439, new_AGEMA_signal_6437}), .b ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, LED_128_Instance_mixcolumns_out[23]}), .c ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, LED_128_Instance_MCS_Instance_1_n27}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U40 ( .a ({new_AGEMA_signal_3631, new_AGEMA_signal_3630, LED_128_Instance_MCS_Instance_1_n25}), .b ({new_AGEMA_signal_3029, new_AGEMA_signal_3028, LED_128_Instance_mixcolumns_out[4]}), .c ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, LED_128_Instance_mixcolumns_out[52]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U39 ( .a ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, LED_128_Instance_mixcolumns_out[23]}), .b ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, LED_128_Instance_MCS_Instance_1_n28}), .c ({new_AGEMA_signal_3631, new_AGEMA_signal_3630, LED_128_Instance_MCS_Instance_1_n25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U38 ( .a ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, LED_128_Instance_subcells_out[50]}), .b ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, LED_128_Instance_mixcolumns_out[39]}), .c ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, LED_128_Instance_MCS_Instance_1_n28}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U37 ( .a ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, LED_128_Instance_MCS_Instance_1_n24}), .b ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, LED_128_Instance_MCS_Instance_1_n23}), .c ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, LED_128_Instance_mixcolumns_out[39]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U36 ( .a ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, LED_128_Instance_subcells_out[51]}), .b ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, LED_128_Instance_subcells_out[45]}), .c ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, LED_128_Instance_MCS_Instance_1_n23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U35 ( .a ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, LED_128_Instance_mixcolumns_out[22]}), .b ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, LED_128_Instance_mixcolumns_out[6]}), .c ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, LED_128_Instance_MCS_Instance_1_n24}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U34 ( .a ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, LED_128_Instance_MCS_Instance_1_n22}), .b ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, LED_128_Instance_MCS_Instance_1_n21}), .c ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, LED_128_Instance_mixcolumns_out[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U33 ( .a ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, LED_128_Instance_MCS_Instance_1_n20}), .b ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, LED_128_Instance_subcells_out[49]}), .c ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, LED_128_Instance_MCS_Instance_1_n21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U32 ( .a ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, LED_128_Instance_mixcolumns_out[5]}), .b ({new_AGEMA_signal_6447, new_AGEMA_signal_6445, new_AGEMA_signal_6443}), .c ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, LED_128_Instance_MCS_Instance_1_n22}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U31 ( .a ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, LED_128_Instance_MCS_Instance_1_n19}), .b ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, LED_128_Instance_MCS_Instance_1_n18}), .c ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, LED_128_Instance_mixcolumns_out[5]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U30 ( .a ({new_AGEMA_signal_6453, new_AGEMA_signal_6451, new_AGEMA_signal_6449}), .b ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, LED_128_Instance_subcells_out[47]}), .c ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, LED_128_Instance_MCS_Instance_1_n18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U29 ( .a ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, LED_128_Instance_MCS_Instance_1_n17}), .b ({new_AGEMA_signal_3025, new_AGEMA_signal_3024, LED_128_Instance_MCS_Instance_1_n34}), .c ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, LED_128_Instance_MCS_Instance_1_n19}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U28 ( .a ({new_AGEMA_signal_2967, new_AGEMA_signal_2966, LED_128_Instance_MCS_Instance_1_n16}), .b ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, LED_128_Instance_subcells_out[6]}), .c ({new_AGEMA_signal_3025, new_AGEMA_signal_3024, LED_128_Instance_MCS_Instance_1_n34}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U27 ( .a ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, LED_128_Instance_subcells_out[25]}), .b ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, LED_128_Instance_subcells_out[7]}), .c ({new_AGEMA_signal_2967, new_AGEMA_signal_2966, LED_128_Instance_MCS_Instance_1_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U26 ( .a ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, LED_128_Instance_MCS_Instance_1_n15}), .b ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, LED_128_Instance_MCS_Instance_1_n31}), .c ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, LED_128_Instance_mixcolumns_out[37]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U25 ( .a ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, LED_128_Instance_mixcolumns_out[20]}), .b ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, LED_128_Instance_mixcolumns_out[23]}), .c ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, LED_128_Instance_MCS_Instance_1_n31}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U24 ( .a ({new_AGEMA_signal_3175, new_AGEMA_signal_3174, LED_128_Instance_MCS_Instance_1_n14}), .b ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, LED_128_Instance_MCS_Instance_1_n13}), .c ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, LED_128_Instance_MCS_Instance_1_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U23 ( .a ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, LED_128_Instance_subcells_out[46]}), .b ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, LED_128_Instance_subcells_out[47]}), .c ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, LED_128_Instance_MCS_Instance_1_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U22 ( .a ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, LED_128_Instance_MCS_Instance_1_n12}), .b ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, LED_128_Instance_subcells_out[49]}), .c ({new_AGEMA_signal_3175, new_AGEMA_signal_3174, LED_128_Instance_MCS_Instance_1_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U21 ( .a ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, LED_128_Instance_MCS_Instance_1_n11}), .b ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, LED_128_Instance_MCS_Instance_1_n10}), .c ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, LED_128_Instance_mixcolumns_out[20]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U20 ( .a ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, LED_128_Instance_mixcolumns_out[7]}), .b ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, LED_128_Instance_subcells_out[51]}), .c ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, LED_128_Instance_MCS_Instance_1_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U19 ( .a ({new_AGEMA_signal_6453, new_AGEMA_signal_6451, new_AGEMA_signal_6449}), .b ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, LED_128_Instance_subcells_out[26]}), .c ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, LED_128_Instance_MCS_Instance_1_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U18 ( .a ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, LED_128_Instance_MCS_Instance_1_n9}), .b ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, LED_128_Instance_MCS_Instance_1_n8}), .c ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, LED_128_Instance_mixcolumns_out[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U17 ( .a ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, LED_128_Instance_subcells_out[50]}), .b ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, LED_128_Instance_subcells_out[47]}), .c ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, LED_128_Instance_MCS_Instance_1_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U16 ( .a ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, LED_128_Instance_mixcolumns_out[6]}), .b ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, LED_128_Instance_subcells_out[25]}), .c ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, LED_128_Instance_MCS_Instance_1_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U15 ( .a ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, LED_128_Instance_MCS_Instance_1_n7}), .b ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, LED_128_Instance_MCS_Instance_1_n6}), .c ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, LED_128_Instance_mixcolumns_out[6]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U14 ( .a ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, LED_128_Instance_MCS_Instance_1_n5}), .b ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, LED_128_Instance_subcells_out[7]}), .c ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, LED_128_Instance_MCS_Instance_1_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U13 ( .a ({new_AGEMA_signal_6459, new_AGEMA_signal_6457, new_AGEMA_signal_6455}), .b ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, LED_128_Instance_subcells_out[49]}), .c ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, LED_128_Instance_MCS_Instance_1_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U12 ( .a ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, LED_128_Instance_MCS_Instance_1_n17}), .b ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, LED_128_Instance_MCS_Instance_1_n35}), .c ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, LED_128_Instance_mixcolumns_out[21]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U11 ( .a ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, LED_128_Instance_MCS_Instance_1_n4}), .b ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, LED_128_Instance_MCS_Instance_1_n12}), .c ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, LED_128_Instance_MCS_Instance_1_n35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U10 ( .a ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, LED_128_Instance_mixcolumns_out[7]}), .b ({new_AGEMA_signal_3029, new_AGEMA_signal_3028, LED_128_Instance_mixcolumns_out[4]}), .c ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, LED_128_Instance_MCS_Instance_1_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U9 ( .a ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, LED_128_Instance_subcells_out[27]}), .b ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, LED_128_Instance_MCS_Instance_1_n5}), .c ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, LED_128_Instance_MCS_Instance_1_n4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U8 ( .a ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, LED_128_Instance_subcells_out[26]}), .b ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, LED_128_Instance_subcells_out[45]}), .c ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, LED_128_Instance_MCS_Instance_1_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U7 ( .a ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, LED_128_Instance_subcells_out[51]}), .b ({new_AGEMA_signal_6441, new_AGEMA_signal_6439, new_AGEMA_signal_6437}), .c ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, LED_128_Instance_MCS_Instance_1_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U6 ( .a ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, LED_128_Instance_MCS_Instance_1_n3}), .b ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, LED_128_Instance_MCS_Instance_1_n2}), .c ({new_AGEMA_signal_3029, new_AGEMA_signal_3028, LED_128_Instance_mixcolumns_out[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U5 ( .a ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, LED_128_Instance_subcells_out[51]}), .b ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, LED_128_Instance_subcells_out[47]}), .c ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, LED_128_Instance_MCS_Instance_1_n2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U4 ( .a ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, LED_128_Instance_subcells_out[6]}), .b ({new_AGEMA_signal_6447, new_AGEMA_signal_6445, new_AGEMA_signal_6443}), .c ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, LED_128_Instance_MCS_Instance_1_n3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U3 ( .a ({new_AGEMA_signal_2975, new_AGEMA_signal_2974, LED_128_Instance_MCS_Instance_1_n1}), .b ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, LED_128_Instance_subcells_out[50]}), .c ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, LED_128_Instance_mixcolumns_out[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U2 ( .a ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, LED_128_Instance_MCS_Instance_1_n20}), .b ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, LED_128_Instance_subcells_out[5]}), .c ({new_AGEMA_signal_2975, new_AGEMA_signal_2974, LED_128_Instance_MCS_Instance_1_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U1 ( .a ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, LED_128_Instance_subcells_out[46]}), .b ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, LED_128_Instance_subcells_out[27]}), .c ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, LED_128_Instance_MCS_Instance_1_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U54 ( .a ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, LED_128_Instance_MCS_Instance_2_n38}), .b ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, LED_128_Instance_MCS_Instance_2_n37}), .c ({new_AGEMA_signal_3451, new_AGEMA_signal_3450, LED_128_Instance_mixcolumns_out[59]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U53 ( .a ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, LED_128_Instance_mixcolumns_out[11]}), .b ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, LED_128_Instance_subcells_out[53]}), .c ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, LED_128_Instance_MCS_Instance_2_n37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U52 ( .a ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, LED_128_Instance_mixcolumns_out[42]}), .b ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, LED_128_Instance_mixcolumns_out[26]}), .c ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, LED_128_Instance_MCS_Instance_2_n38}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U51 ( .a ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MCS_Instance_2_n36}), .b ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, LED_128_Instance_MCS_Instance_2_n35}), .c ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, LED_128_Instance_mixcolumns_out[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U50 ( .a ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, LED_128_Instance_subcells_out[54]}), .b ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, LED_128_Instance_MCS_Instance_2_n34}), .c ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MCS_Instance_2_n36}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U49 ( .a ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, LED_128_Instance_MCS_Instance_2_n33}), .b ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, LED_128_Instance_mixcolumns_out[41]}), .c ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, LED_128_Instance_mixcolumns_out[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U48 ( .a ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, LED_128_Instance_mixcolumns_out[10]}), .b ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, LED_128_Instance_MCS_Instance_2_n35}), .c ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, LED_128_Instance_MCS_Instance_2_n33}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U47 ( .a ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, LED_128_Instance_MCS_Instance_2_n32}), .b ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, LED_128_Instance_MCS_Instance_2_n31}), .c ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, LED_128_Instance_mixcolumns_out[57]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U46 ( .a ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, LED_128_Instance_MCS_Instance_2_n30}), .b ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, LED_128_Instance_MCS_Instance_2_n29}), .c ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, LED_128_Instance_MCS_Instance_2_n32}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U45 ( .a ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, LED_128_Instance_subcells_out[55]}), .b ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, LED_128_Instance_mixcolumns_out[9]}), .c ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, LED_128_Instance_MCS_Instance_2_n29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U44 ( .a ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, LED_128_Instance_mixcolumns_out[40]}), .b ({new_AGEMA_signal_3535, new_AGEMA_signal_3534, LED_128_Instance_MCS_Instance_2_n28}), .c ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, LED_128_Instance_MCS_Instance_2_n30}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U43 ( .a ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, LED_128_Instance_MCS_Instance_2_n27}), .b ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, LED_128_Instance_MCS_Instance_2_n26}), .c ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, LED_128_Instance_mixcolumns_out[40]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U42 ( .a ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, LED_128_Instance_subcells_out[34]}), .b ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, LED_128_Instance_mixcolumns_out[11]}), .c ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, LED_128_Instance_MCS_Instance_2_n26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U41 ( .a ({new_AGEMA_signal_6465, new_AGEMA_signal_6463, new_AGEMA_signal_6461}), .b ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, LED_128_Instance_mixcolumns_out[27]}), .c ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, LED_128_Instance_MCS_Instance_2_n27}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U40 ( .a ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, LED_128_Instance_MCS_Instance_2_n25}), .b ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, LED_128_Instance_mixcolumns_out[8]}), .c ({new_AGEMA_signal_3635, new_AGEMA_signal_3634, LED_128_Instance_mixcolumns_out[56]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U39 ( .a ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, LED_128_Instance_mixcolumns_out[27]}), .b ({new_AGEMA_signal_3535, new_AGEMA_signal_3534, LED_128_Instance_MCS_Instance_2_n28}), .c ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, LED_128_Instance_MCS_Instance_2_n25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U38 ( .a ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, LED_128_Instance_subcells_out[54]}), .b ({new_AGEMA_signal_3455, new_AGEMA_signal_3454, LED_128_Instance_mixcolumns_out[43]}), .c ({new_AGEMA_signal_3535, new_AGEMA_signal_3534, LED_128_Instance_MCS_Instance_2_n28}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U37 ( .a ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, LED_128_Instance_MCS_Instance_2_n24}), .b ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, LED_128_Instance_MCS_Instance_2_n23}), .c ({new_AGEMA_signal_3455, new_AGEMA_signal_3454, LED_128_Instance_mixcolumns_out[43]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U36 ( .a ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, LED_128_Instance_subcells_out[55]}), .b ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, LED_128_Instance_subcells_out[33]}), .c ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, LED_128_Instance_MCS_Instance_2_n23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U35 ( .a ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, LED_128_Instance_mixcolumns_out[26]}), .b ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, LED_128_Instance_mixcolumns_out[10]}), .c ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, LED_128_Instance_MCS_Instance_2_n24}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U34 ( .a ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, LED_128_Instance_MCS_Instance_2_n22}), .b ({new_AGEMA_signal_2979, new_AGEMA_signal_2978, LED_128_Instance_MCS_Instance_2_n21}), .c ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, LED_128_Instance_mixcolumns_out[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U33 ( .a ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, LED_128_Instance_MCS_Instance_2_n20}), .b ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, LED_128_Instance_subcells_out[53]}), .c ({new_AGEMA_signal_2979, new_AGEMA_signal_2978, LED_128_Instance_MCS_Instance_2_n21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U32 ( .a ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, LED_128_Instance_mixcolumns_out[9]}), .b ({new_AGEMA_signal_6471, new_AGEMA_signal_6469, new_AGEMA_signal_6467}), .c ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, LED_128_Instance_MCS_Instance_2_n22}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U31 ( .a ({new_AGEMA_signal_3035, new_AGEMA_signal_3034, LED_128_Instance_MCS_Instance_2_n19}), .b ({new_AGEMA_signal_2981, new_AGEMA_signal_2980, LED_128_Instance_MCS_Instance_2_n18}), .c ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, LED_128_Instance_mixcolumns_out[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U30 ( .a ({new_AGEMA_signal_6477, new_AGEMA_signal_6475, new_AGEMA_signal_6473}), .b ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, LED_128_Instance_subcells_out[35]}), .c ({new_AGEMA_signal_2981, new_AGEMA_signal_2980, LED_128_Instance_MCS_Instance_2_n18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U29 ( .a ({new_AGEMA_signal_2993, new_AGEMA_signal_2992, LED_128_Instance_MCS_Instance_2_n17}), .b ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, LED_128_Instance_MCS_Instance_2_n34}), .c ({new_AGEMA_signal_3035, new_AGEMA_signal_3034, LED_128_Instance_MCS_Instance_2_n19}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U28 ( .a ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, LED_128_Instance_MCS_Instance_2_n16}), .b ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, LED_128_Instance_subcells_out[10]}), .c ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, LED_128_Instance_MCS_Instance_2_n34}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U27 ( .a ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, LED_128_Instance_subcells_out[29]}), .b ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, LED_128_Instance_subcells_out[11]}), .c ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, LED_128_Instance_MCS_Instance_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U26 ( .a ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, LED_128_Instance_MCS_Instance_2_n15}), .b ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, LED_128_Instance_MCS_Instance_2_n31}), .c ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, LED_128_Instance_mixcolumns_out[41]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U25 ( .a ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, LED_128_Instance_mixcolumns_out[24]}), .b ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, LED_128_Instance_mixcolumns_out[27]}), .c ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, LED_128_Instance_MCS_Instance_2_n31}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U24 ( .a ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, LED_128_Instance_MCS_Instance_2_n14}), .b ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, LED_128_Instance_MCS_Instance_2_n13}), .c ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, LED_128_Instance_MCS_Instance_2_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U23 ( .a ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, LED_128_Instance_subcells_out[34]}), .b ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, LED_128_Instance_subcells_out[35]}), .c ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, LED_128_Instance_MCS_Instance_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U22 ( .a ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, LED_128_Instance_MCS_Instance_2_n12}), .b ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, LED_128_Instance_subcells_out[53]}), .c ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, LED_128_Instance_MCS_Instance_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U21 ( .a ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, LED_128_Instance_MCS_Instance_2_n11}), .b ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, LED_128_Instance_MCS_Instance_2_n10}), .c ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, LED_128_Instance_mixcolumns_out[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U20 ( .a ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, LED_128_Instance_mixcolumns_out[11]}), .b ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, LED_128_Instance_subcells_out[55]}), .c ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, LED_128_Instance_MCS_Instance_2_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U19 ( .a ({new_AGEMA_signal_6477, new_AGEMA_signal_6475, new_AGEMA_signal_6473}), .b ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, LED_128_Instance_subcells_out[30]}), .c ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, LED_128_Instance_MCS_Instance_2_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U18 ( .a ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, LED_128_Instance_MCS_Instance_2_n9}), .b ({new_AGEMA_signal_2987, new_AGEMA_signal_2986, LED_128_Instance_MCS_Instance_2_n8}), .c ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, LED_128_Instance_mixcolumns_out[27]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U17 ( .a ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, LED_128_Instance_subcells_out[54]}), .b ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, LED_128_Instance_subcells_out[35]}), .c ({new_AGEMA_signal_2987, new_AGEMA_signal_2986, LED_128_Instance_MCS_Instance_2_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U16 ( .a ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, LED_128_Instance_mixcolumns_out[10]}), .b ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, LED_128_Instance_subcells_out[29]}), .c ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, LED_128_Instance_MCS_Instance_2_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U15 ( .a ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, LED_128_Instance_MCS_Instance_2_n7}), .b ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, LED_128_Instance_MCS_Instance_2_n6}), .c ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, LED_128_Instance_mixcolumns_out[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U14 ( .a ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, LED_128_Instance_MCS_Instance_2_n5}), .b ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, LED_128_Instance_subcells_out[11]}), .c ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, LED_128_Instance_MCS_Instance_2_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U13 ( .a ({new_AGEMA_signal_6483, new_AGEMA_signal_6481, new_AGEMA_signal_6479}), .b ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, LED_128_Instance_subcells_out[53]}), .c ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, LED_128_Instance_MCS_Instance_2_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U12 ( .a ({new_AGEMA_signal_2993, new_AGEMA_signal_2992, LED_128_Instance_MCS_Instance_2_n17}), .b ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, LED_128_Instance_MCS_Instance_2_n35}), .c ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, LED_128_Instance_mixcolumns_out[25]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U11 ( .a ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, LED_128_Instance_MCS_Instance_2_n4}), .b ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, LED_128_Instance_MCS_Instance_2_n12}), .c ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, LED_128_Instance_MCS_Instance_2_n35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U10 ( .a ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, LED_128_Instance_mixcolumns_out[11]}), .b ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, LED_128_Instance_mixcolumns_out[8]}), .c ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, LED_128_Instance_MCS_Instance_2_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U9 ( .a ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, LED_128_Instance_subcells_out[31]}), .b ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, LED_128_Instance_MCS_Instance_2_n5}), .c ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, LED_128_Instance_MCS_Instance_2_n4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U8 ( .a ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, LED_128_Instance_subcells_out[30]}), .b ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, LED_128_Instance_subcells_out[33]}), .c ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, LED_128_Instance_MCS_Instance_2_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U7 ( .a ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, LED_128_Instance_subcells_out[55]}), .b ({new_AGEMA_signal_6465, new_AGEMA_signal_6463, new_AGEMA_signal_6461}), .c ({new_AGEMA_signal_2993, new_AGEMA_signal_2992, LED_128_Instance_MCS_Instance_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U6 ( .a ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, LED_128_Instance_MCS_Instance_2_n3}), .b ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, LED_128_Instance_MCS_Instance_2_n2}), .c ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, LED_128_Instance_mixcolumns_out[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U5 ( .a ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, LED_128_Instance_subcells_out[55]}), .b ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, LED_128_Instance_subcells_out[35]}), .c ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, LED_128_Instance_MCS_Instance_2_n2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U4 ( .a ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, LED_128_Instance_subcells_out[10]}), .b ({new_AGEMA_signal_6471, new_AGEMA_signal_6469, new_AGEMA_signal_6467}), .c ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, LED_128_Instance_MCS_Instance_2_n3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U3 ( .a ({new_AGEMA_signal_2997, new_AGEMA_signal_2996, LED_128_Instance_MCS_Instance_2_n1}), .b ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, LED_128_Instance_subcells_out[54]}), .c ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, LED_128_Instance_mixcolumns_out[11]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U2 ( .a ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, LED_128_Instance_MCS_Instance_2_n20}), .b ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, LED_128_Instance_subcells_out[9]}), .c ({new_AGEMA_signal_2997, new_AGEMA_signal_2996, LED_128_Instance_MCS_Instance_2_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U1 ( .a ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, LED_128_Instance_subcells_out[34]}), .b ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, LED_128_Instance_subcells_out[31]}), .c ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, LED_128_Instance_MCS_Instance_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U54 ( .a ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, LED_128_Instance_MCS_Instance_3_n38}), .b ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, LED_128_Instance_MCS_Instance_3_n37}), .c ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, LED_128_Instance_mixcolumns_out[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U53 ( .a ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, LED_128_Instance_mixcolumns_out[15]}), .b ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, LED_128_Instance_subcells_out[57]}), .c ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, LED_128_Instance_MCS_Instance_3_n37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U52 ( .a ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, LED_128_Instance_mixcolumns_out[46]}), .b ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, LED_128_Instance_mixcolumns_out[30]}), .c ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, LED_128_Instance_MCS_Instance_3_n38}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U51 ( .a ({new_AGEMA_signal_3043, new_AGEMA_signal_3042, LED_128_Instance_MCS_Instance_3_n36}), .b ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, LED_128_Instance_MCS_Instance_3_n35}), .c ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, LED_128_Instance_mixcolumns_out[46]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U50 ( .a ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, LED_128_Instance_subcells_out[58]}), .b ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, LED_128_Instance_MCS_Instance_3_n34}), .c ({new_AGEMA_signal_3043, new_AGEMA_signal_3042, LED_128_Instance_MCS_Instance_3_n36}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U49 ( .a ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, LED_128_Instance_MCS_Instance_3_n33}), .b ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, LED_128_Instance_mixcolumns_out[45]}), .c ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, LED_128_Instance_mixcolumns_out[62]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U48 ( .a ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, LED_128_Instance_mixcolumns_out[14]}), .b ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, LED_128_Instance_MCS_Instance_3_n35}), .c ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, LED_128_Instance_MCS_Instance_3_n33}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U47 ( .a ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, LED_128_Instance_MCS_Instance_3_n32}), .b ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, LED_128_Instance_MCS_Instance_3_n31}), .c ({new_AGEMA_signal_3655, new_AGEMA_signal_3654, LED_128_Instance_mixcolumns_out[61]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U46 ( .a ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, LED_128_Instance_MCS_Instance_3_n30}), .b ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, LED_128_Instance_MCS_Instance_3_n29}), .c ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, LED_128_Instance_MCS_Instance_3_n32}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U45 ( .a ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, LED_128_Instance_subcells_out[59]}), .b ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, LED_128_Instance_mixcolumns_out[13]}), .c ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, LED_128_Instance_MCS_Instance_3_n29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U44 ( .a ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, LED_128_Instance_mixcolumns_out[44]}), .b ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, LED_128_Instance_MCS_Instance_3_n28}), .c ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, LED_128_Instance_MCS_Instance_3_n30}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U43 ( .a ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, LED_128_Instance_MCS_Instance_3_n27}), .b ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, LED_128_Instance_MCS_Instance_3_n26}), .c ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, LED_128_Instance_mixcolumns_out[44]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U42 ( .a ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, LED_128_Instance_subcells_out[38]}), .b ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, LED_128_Instance_mixcolumns_out[15]}), .c ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, LED_128_Instance_MCS_Instance_3_n26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U41 ( .a ({new_AGEMA_signal_6489, new_AGEMA_signal_6487, new_AGEMA_signal_6485}), .b ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, LED_128_Instance_mixcolumns_out[31]}), .c ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, LED_128_Instance_MCS_Instance_3_n27}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U40 ( .a ({new_AGEMA_signal_3595, new_AGEMA_signal_3594, LED_128_Instance_MCS_Instance_3_n25}), .b ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, LED_128_Instance_mixcolumns_out[12]}), .c ({new_AGEMA_signal_3639, new_AGEMA_signal_3638, LED_128_Instance_mixcolumns_out[60]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U39 ( .a ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, LED_128_Instance_mixcolumns_out[31]}), .b ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, LED_128_Instance_MCS_Instance_3_n28}), .c ({new_AGEMA_signal_3595, new_AGEMA_signal_3594, LED_128_Instance_MCS_Instance_3_n25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U38 ( .a ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, LED_128_Instance_subcells_out[58]}), .b ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, LED_128_Instance_mixcolumns_out[47]}), .c ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, LED_128_Instance_MCS_Instance_3_n28}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U37 ( .a ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, LED_128_Instance_MCS_Instance_3_n24}), .b ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, LED_128_Instance_MCS_Instance_3_n23}), .c ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, LED_128_Instance_mixcolumns_out[47]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U36 ( .a ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, LED_128_Instance_subcells_out[59]}), .b ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, LED_128_Instance_subcells_out[37]}), .c ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, LED_128_Instance_MCS_Instance_3_n23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U35 ( .a ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, LED_128_Instance_mixcolumns_out[30]}), .b ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, LED_128_Instance_mixcolumns_out[14]}), .c ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, LED_128_Instance_MCS_Instance_3_n24}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U34 ( .a ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, LED_128_Instance_MCS_Instance_3_n22}), .b ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, LED_128_Instance_MCS_Instance_3_n21}), .c ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, LED_128_Instance_mixcolumns_out[30]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U33 ( .a ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, LED_128_Instance_MCS_Instance_3_n20}), .b ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, LED_128_Instance_subcells_out[57]}), .c ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, LED_128_Instance_MCS_Instance_3_n21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U32 ( .a ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, LED_128_Instance_mixcolumns_out[13]}), .b ({new_AGEMA_signal_6495, new_AGEMA_signal_6493, new_AGEMA_signal_6491}), .c ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, LED_128_Instance_MCS_Instance_3_n22}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U31 ( .a ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, LED_128_Instance_MCS_Instance_3_n19}), .b ({new_AGEMA_signal_2999, new_AGEMA_signal_2998, LED_128_Instance_MCS_Instance_3_n18}), .c ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, LED_128_Instance_mixcolumns_out[13]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U30 ( .a ({new_AGEMA_signal_6501, new_AGEMA_signal_6499, new_AGEMA_signal_6497}), .b ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, LED_128_Instance_subcells_out[39]}), .c ({new_AGEMA_signal_2999, new_AGEMA_signal_2998, LED_128_Instance_MCS_Instance_3_n18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U29 ( .a ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, LED_128_Instance_MCS_Instance_3_n17}), .b ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, LED_128_Instance_MCS_Instance_3_n34}), .c ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, LED_128_Instance_MCS_Instance_3_n19}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U28 ( .a ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, LED_128_Instance_MCS_Instance_3_n16}), .b ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, LED_128_Instance_subcells_out[14]}), .c ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, LED_128_Instance_MCS_Instance_3_n34}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U27 ( .a ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, LED_128_Instance_subcells_out[17]}), .b ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, LED_128_Instance_subcells_out[15]}), .c ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, LED_128_Instance_MCS_Instance_3_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U26 ( .a ({new_AGEMA_signal_3379, new_AGEMA_signal_3378, LED_128_Instance_MCS_Instance_3_n15}), .b ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, LED_128_Instance_MCS_Instance_3_n31}), .c ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, LED_128_Instance_mixcolumns_out[45]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U25 ( .a ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, LED_128_Instance_mixcolumns_out[28]}), .b ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, LED_128_Instance_mixcolumns_out[31]}), .c ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, LED_128_Instance_MCS_Instance_3_n31}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U24 ( .a ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, LED_128_Instance_MCS_Instance_3_n14}), .b ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, LED_128_Instance_MCS_Instance_3_n13}), .c ({new_AGEMA_signal_3379, new_AGEMA_signal_3378, LED_128_Instance_MCS_Instance_3_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U23 ( .a ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, LED_128_Instance_subcells_out[38]}), .b ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, LED_128_Instance_subcells_out[39]}), .c ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, LED_128_Instance_MCS_Instance_3_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U22 ( .a ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, LED_128_Instance_MCS_Instance_3_n12}), .b ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, LED_128_Instance_subcells_out[57]}), .c ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, LED_128_Instance_MCS_Instance_3_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U21 ( .a ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, LED_128_Instance_MCS_Instance_3_n11}), .b ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, LED_128_Instance_MCS_Instance_3_n10}), .c ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, LED_128_Instance_mixcolumns_out[28]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U20 ( .a ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, LED_128_Instance_mixcolumns_out[15]}), .b ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, LED_128_Instance_subcells_out[59]}), .c ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, LED_128_Instance_MCS_Instance_3_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U19 ( .a ({new_AGEMA_signal_6501, new_AGEMA_signal_6499, new_AGEMA_signal_6497}), .b ({new_AGEMA_signal_2827, new_AGEMA_signal_2826, LED_128_Instance_subcells_out[18]}), .c ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, LED_128_Instance_MCS_Instance_3_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U18 ( .a ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, LED_128_Instance_MCS_Instance_3_n9}), .b ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, LED_128_Instance_MCS_Instance_3_n8}), .c ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, LED_128_Instance_mixcolumns_out[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U17 ( .a ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, LED_128_Instance_subcells_out[58]}), .b ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, LED_128_Instance_subcells_out[39]}), .c ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, LED_128_Instance_MCS_Instance_3_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U16 ( .a ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, LED_128_Instance_mixcolumns_out[14]}), .b ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, LED_128_Instance_subcells_out[17]}), .c ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, LED_128_Instance_MCS_Instance_3_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U15 ( .a ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, LED_128_Instance_MCS_Instance_3_n7}), .b ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, LED_128_Instance_MCS_Instance_3_n6}), .c ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, LED_128_Instance_mixcolumns_out[14]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U14 ( .a ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, LED_128_Instance_MCS_Instance_3_n5}), .b ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, LED_128_Instance_subcells_out[15]}), .c ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, LED_128_Instance_MCS_Instance_3_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U13 ( .a ({new_AGEMA_signal_6507, new_AGEMA_signal_6505, new_AGEMA_signal_6503}), .b ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, LED_128_Instance_subcells_out[57]}), .c ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, LED_128_Instance_MCS_Instance_3_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U12 ( .a ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, LED_128_Instance_MCS_Instance_3_n17}), .b ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, LED_128_Instance_MCS_Instance_3_n35}), .c ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, LED_128_Instance_mixcolumns_out[29]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U11 ( .a ({new_AGEMA_signal_3009, new_AGEMA_signal_3008, LED_128_Instance_MCS_Instance_3_n4}), .b ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, LED_128_Instance_MCS_Instance_3_n12}), .c ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, LED_128_Instance_MCS_Instance_3_n35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U10 ( .a ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, LED_128_Instance_mixcolumns_out[15]}), .b ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, LED_128_Instance_mixcolumns_out[12]}), .c ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, LED_128_Instance_MCS_Instance_3_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U9 ( .a ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, LED_128_Instance_subcells_out[19]}), .b ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, LED_128_Instance_MCS_Instance_3_n5}), .c ({new_AGEMA_signal_3009, new_AGEMA_signal_3008, LED_128_Instance_MCS_Instance_3_n4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U8 ( .a ({new_AGEMA_signal_2827, new_AGEMA_signal_2826, LED_128_Instance_subcells_out[18]}), .b ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, LED_128_Instance_subcells_out[37]}), .c ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, LED_128_Instance_MCS_Instance_3_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U7 ( .a ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, LED_128_Instance_subcells_out[59]}), .b ({new_AGEMA_signal_6489, new_AGEMA_signal_6487, new_AGEMA_signal_6485}), .c ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, LED_128_Instance_MCS_Instance_3_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U6 ( .a ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, LED_128_Instance_MCS_Instance_3_n3}), .b ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, LED_128_Instance_MCS_Instance_3_n2}), .c ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, LED_128_Instance_mixcolumns_out[12]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U5 ( .a ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, LED_128_Instance_subcells_out[59]}), .b ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, LED_128_Instance_subcells_out[39]}), .c ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, LED_128_Instance_MCS_Instance_3_n2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U4 ( .a ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, LED_128_Instance_subcells_out[14]}), .b ({new_AGEMA_signal_6495, new_AGEMA_signal_6493, new_AGEMA_signal_6491}), .c ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, LED_128_Instance_MCS_Instance_3_n3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U3 ( .a ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, LED_128_Instance_MCS_Instance_3_n1}), .b ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, LED_128_Instance_subcells_out[58]}), .c ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, LED_128_Instance_mixcolumns_out[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U2 ( .a ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, LED_128_Instance_MCS_Instance_3_n20}), .b ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, LED_128_Instance_subcells_out[13]}), .c ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, LED_128_Instance_MCS_Instance_3_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U1 ( .a ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, LED_128_Instance_subcells_out[38]}), .b ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, LED_128_Instance_subcells_out[19]}), .c ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, LED_128_Instance_MCS_Instance_3_n20}) ) ;
    buf_clk new_AGEMA_reg_buffer_1419 ( .C (CLK), .D (new_AGEMA_signal_4186), .Q (new_AGEMA_signal_4187) ) ;
    buf_clk new_AGEMA_reg_buffer_1423 ( .C (CLK), .D (new_AGEMA_signal_4190), .Q (new_AGEMA_signal_4191) ) ;
    buf_clk new_AGEMA_reg_buffer_1427 ( .C (CLK), .D (new_AGEMA_signal_4194), .Q (new_AGEMA_signal_4195) ) ;
    buf_clk new_AGEMA_reg_buffer_1431 ( .C (CLK), .D (new_AGEMA_signal_4198), .Q (new_AGEMA_signal_4199) ) ;
    buf_clk new_AGEMA_reg_buffer_1435 ( .C (CLK), .D (new_AGEMA_signal_4202), .Q (new_AGEMA_signal_4203) ) ;
    buf_clk new_AGEMA_reg_buffer_1439 ( .C (CLK), .D (new_AGEMA_signal_4206), .Q (new_AGEMA_signal_4207) ) ;
    buf_clk new_AGEMA_reg_buffer_1443 ( .C (CLK), .D (new_AGEMA_signal_4210), .Q (new_AGEMA_signal_4211) ) ;
    buf_clk new_AGEMA_reg_buffer_1447 ( .C (CLK), .D (new_AGEMA_signal_4214), .Q (new_AGEMA_signal_4215) ) ;
    buf_clk new_AGEMA_reg_buffer_1451 ( .C (CLK), .D (new_AGEMA_signal_4218), .Q (new_AGEMA_signal_4219) ) ;
    buf_clk new_AGEMA_reg_buffer_1455 ( .C (CLK), .D (new_AGEMA_signal_4222), .Q (new_AGEMA_signal_4223) ) ;
    buf_clk new_AGEMA_reg_buffer_1459 ( .C (CLK), .D (new_AGEMA_signal_4226), .Q (new_AGEMA_signal_4227) ) ;
    buf_clk new_AGEMA_reg_buffer_1463 ( .C (CLK), .D (new_AGEMA_signal_4230), .Q (new_AGEMA_signal_4231) ) ;
    buf_clk new_AGEMA_reg_buffer_1467 ( .C (CLK), .D (new_AGEMA_signal_4234), .Q (new_AGEMA_signal_4235) ) ;
    buf_clk new_AGEMA_reg_buffer_1471 ( .C (CLK), .D (new_AGEMA_signal_4238), .Q (new_AGEMA_signal_4239) ) ;
    buf_clk new_AGEMA_reg_buffer_1475 ( .C (CLK), .D (new_AGEMA_signal_4242), .Q (new_AGEMA_signal_4243) ) ;
    buf_clk new_AGEMA_reg_buffer_1479 ( .C (CLK), .D (new_AGEMA_signal_4246), .Q (new_AGEMA_signal_4247) ) ;
    buf_clk new_AGEMA_reg_buffer_1483 ( .C (CLK), .D (new_AGEMA_signal_4250), .Q (new_AGEMA_signal_4251) ) ;
    buf_clk new_AGEMA_reg_buffer_1487 ( .C (CLK), .D (new_AGEMA_signal_4254), .Q (new_AGEMA_signal_4255) ) ;
    buf_clk new_AGEMA_reg_buffer_1491 ( .C (CLK), .D (new_AGEMA_signal_4258), .Q (new_AGEMA_signal_4259) ) ;
    buf_clk new_AGEMA_reg_buffer_1495 ( .C (CLK), .D (new_AGEMA_signal_4262), .Q (new_AGEMA_signal_4263) ) ;
    buf_clk new_AGEMA_reg_buffer_1499 ( .C (CLK), .D (new_AGEMA_signal_4266), .Q (new_AGEMA_signal_4267) ) ;
    buf_clk new_AGEMA_reg_buffer_1503 ( .C (CLK), .D (new_AGEMA_signal_4270), .Q (new_AGEMA_signal_4271) ) ;
    buf_clk new_AGEMA_reg_buffer_1507 ( .C (CLK), .D (new_AGEMA_signal_4274), .Q (new_AGEMA_signal_4275) ) ;
    buf_clk new_AGEMA_reg_buffer_1511 ( .C (CLK), .D (new_AGEMA_signal_4278), .Q (new_AGEMA_signal_4279) ) ;
    buf_clk new_AGEMA_reg_buffer_1515 ( .C (CLK), .D (new_AGEMA_signal_4282), .Q (new_AGEMA_signal_4283) ) ;
    buf_clk new_AGEMA_reg_buffer_1519 ( .C (CLK), .D (new_AGEMA_signal_4286), .Q (new_AGEMA_signal_4287) ) ;
    buf_clk new_AGEMA_reg_buffer_1523 ( .C (CLK), .D (new_AGEMA_signal_4290), .Q (new_AGEMA_signal_4291) ) ;
    buf_clk new_AGEMA_reg_buffer_1527 ( .C (CLK), .D (new_AGEMA_signal_4294), .Q (new_AGEMA_signal_4295) ) ;
    buf_clk new_AGEMA_reg_buffer_1531 ( .C (CLK), .D (new_AGEMA_signal_4298), .Q (new_AGEMA_signal_4299) ) ;
    buf_clk new_AGEMA_reg_buffer_1535 ( .C (CLK), .D (new_AGEMA_signal_4302), .Q (new_AGEMA_signal_4303) ) ;
    buf_clk new_AGEMA_reg_buffer_1539 ( .C (CLK), .D (new_AGEMA_signal_4306), .Q (new_AGEMA_signal_4307) ) ;
    buf_clk new_AGEMA_reg_buffer_1543 ( .C (CLK), .D (new_AGEMA_signal_4310), .Q (new_AGEMA_signal_4311) ) ;
    buf_clk new_AGEMA_reg_buffer_1547 ( .C (CLK), .D (new_AGEMA_signal_4314), .Q (new_AGEMA_signal_4315) ) ;
    buf_clk new_AGEMA_reg_buffer_1551 ( .C (CLK), .D (new_AGEMA_signal_4318), .Q (new_AGEMA_signal_4319) ) ;
    buf_clk new_AGEMA_reg_buffer_1555 ( .C (CLK), .D (new_AGEMA_signal_4322), .Q (new_AGEMA_signal_4323) ) ;
    buf_clk new_AGEMA_reg_buffer_1559 ( .C (CLK), .D (new_AGEMA_signal_4326), .Q (new_AGEMA_signal_4327) ) ;
    buf_clk new_AGEMA_reg_buffer_1563 ( .C (CLK), .D (new_AGEMA_signal_4330), .Q (new_AGEMA_signal_4331) ) ;
    buf_clk new_AGEMA_reg_buffer_1567 ( .C (CLK), .D (new_AGEMA_signal_4334), .Q (new_AGEMA_signal_4335) ) ;
    buf_clk new_AGEMA_reg_buffer_1571 ( .C (CLK), .D (new_AGEMA_signal_4338), .Q (new_AGEMA_signal_4339) ) ;
    buf_clk new_AGEMA_reg_buffer_1575 ( .C (CLK), .D (new_AGEMA_signal_4342), .Q (new_AGEMA_signal_4343) ) ;
    buf_clk new_AGEMA_reg_buffer_1579 ( .C (CLK), .D (new_AGEMA_signal_4346), .Q (new_AGEMA_signal_4347) ) ;
    buf_clk new_AGEMA_reg_buffer_1583 ( .C (CLK), .D (new_AGEMA_signal_4350), .Q (new_AGEMA_signal_4351) ) ;
    buf_clk new_AGEMA_reg_buffer_1587 ( .C (CLK), .D (new_AGEMA_signal_4354), .Q (new_AGEMA_signal_4355) ) ;
    buf_clk new_AGEMA_reg_buffer_1591 ( .C (CLK), .D (new_AGEMA_signal_4358), .Q (new_AGEMA_signal_4359) ) ;
    buf_clk new_AGEMA_reg_buffer_1595 ( .C (CLK), .D (new_AGEMA_signal_4362), .Q (new_AGEMA_signal_4363) ) ;
    buf_clk new_AGEMA_reg_buffer_1599 ( .C (CLK), .D (new_AGEMA_signal_4366), .Q (new_AGEMA_signal_4367) ) ;
    buf_clk new_AGEMA_reg_buffer_1603 ( .C (CLK), .D (new_AGEMA_signal_4370), .Q (new_AGEMA_signal_4371) ) ;
    buf_clk new_AGEMA_reg_buffer_1607 ( .C (CLK), .D (new_AGEMA_signal_4374), .Q (new_AGEMA_signal_4375) ) ;
    buf_clk new_AGEMA_reg_buffer_1611 ( .C (CLK), .D (new_AGEMA_signal_4378), .Q (new_AGEMA_signal_4379) ) ;
    buf_clk new_AGEMA_reg_buffer_1615 ( .C (CLK), .D (new_AGEMA_signal_4382), .Q (new_AGEMA_signal_4383) ) ;
    buf_clk new_AGEMA_reg_buffer_1619 ( .C (CLK), .D (new_AGEMA_signal_4386), .Q (new_AGEMA_signal_4387) ) ;
    buf_clk new_AGEMA_reg_buffer_1623 ( .C (CLK), .D (new_AGEMA_signal_4390), .Q (new_AGEMA_signal_4391) ) ;
    buf_clk new_AGEMA_reg_buffer_1627 ( .C (CLK), .D (new_AGEMA_signal_4394), .Q (new_AGEMA_signal_4395) ) ;
    buf_clk new_AGEMA_reg_buffer_1631 ( .C (CLK), .D (new_AGEMA_signal_4398), .Q (new_AGEMA_signal_4399) ) ;
    buf_clk new_AGEMA_reg_buffer_1635 ( .C (CLK), .D (new_AGEMA_signal_4402), .Q (new_AGEMA_signal_4403) ) ;
    buf_clk new_AGEMA_reg_buffer_1639 ( .C (CLK), .D (new_AGEMA_signal_4406), .Q (new_AGEMA_signal_4407) ) ;
    buf_clk new_AGEMA_reg_buffer_1643 ( .C (CLK), .D (new_AGEMA_signal_4410), .Q (new_AGEMA_signal_4411) ) ;
    buf_clk new_AGEMA_reg_buffer_1647 ( .C (CLK), .D (new_AGEMA_signal_4414), .Q (new_AGEMA_signal_4415) ) ;
    buf_clk new_AGEMA_reg_buffer_1651 ( .C (CLK), .D (new_AGEMA_signal_4418), .Q (new_AGEMA_signal_4419) ) ;
    buf_clk new_AGEMA_reg_buffer_1655 ( .C (CLK), .D (new_AGEMA_signal_4422), .Q (new_AGEMA_signal_4423) ) ;
    buf_clk new_AGEMA_reg_buffer_1659 ( .C (CLK), .D (new_AGEMA_signal_4426), .Q (new_AGEMA_signal_4427) ) ;
    buf_clk new_AGEMA_reg_buffer_1663 ( .C (CLK), .D (new_AGEMA_signal_4430), .Q (new_AGEMA_signal_4431) ) ;
    buf_clk new_AGEMA_reg_buffer_1667 ( .C (CLK), .D (new_AGEMA_signal_4434), .Q (new_AGEMA_signal_4435) ) ;
    buf_clk new_AGEMA_reg_buffer_1671 ( .C (CLK), .D (new_AGEMA_signal_4438), .Q (new_AGEMA_signal_4439) ) ;
    buf_clk new_AGEMA_reg_buffer_1675 ( .C (CLK), .D (new_AGEMA_signal_4442), .Q (new_AGEMA_signal_4443) ) ;
    buf_clk new_AGEMA_reg_buffer_1679 ( .C (CLK), .D (new_AGEMA_signal_4446), .Q (new_AGEMA_signal_4447) ) ;
    buf_clk new_AGEMA_reg_buffer_1683 ( .C (CLK), .D (new_AGEMA_signal_4450), .Q (new_AGEMA_signal_4451) ) ;
    buf_clk new_AGEMA_reg_buffer_1687 ( .C (CLK), .D (new_AGEMA_signal_4454), .Q (new_AGEMA_signal_4455) ) ;
    buf_clk new_AGEMA_reg_buffer_1691 ( .C (CLK), .D (new_AGEMA_signal_4458), .Q (new_AGEMA_signal_4459) ) ;
    buf_clk new_AGEMA_reg_buffer_1695 ( .C (CLK), .D (new_AGEMA_signal_4462), .Q (new_AGEMA_signal_4463) ) ;
    buf_clk new_AGEMA_reg_buffer_1699 ( .C (CLK), .D (new_AGEMA_signal_4466), .Q (new_AGEMA_signal_4467) ) ;
    buf_clk new_AGEMA_reg_buffer_1703 ( .C (CLK), .D (new_AGEMA_signal_4470), .Q (new_AGEMA_signal_4471) ) ;
    buf_clk new_AGEMA_reg_buffer_1707 ( .C (CLK), .D (new_AGEMA_signal_4474), .Q (new_AGEMA_signal_4475) ) ;
    buf_clk new_AGEMA_reg_buffer_1711 ( .C (CLK), .D (new_AGEMA_signal_4478), .Q (new_AGEMA_signal_4479) ) ;
    buf_clk new_AGEMA_reg_buffer_1715 ( .C (CLK), .D (new_AGEMA_signal_4482), .Q (new_AGEMA_signal_4483) ) ;
    buf_clk new_AGEMA_reg_buffer_1719 ( .C (CLK), .D (new_AGEMA_signal_4486), .Q (new_AGEMA_signal_4487) ) ;
    buf_clk new_AGEMA_reg_buffer_1723 ( .C (CLK), .D (new_AGEMA_signal_4490), .Q (new_AGEMA_signal_4491) ) ;
    buf_clk new_AGEMA_reg_buffer_1727 ( .C (CLK), .D (new_AGEMA_signal_4494), .Q (new_AGEMA_signal_4495) ) ;
    buf_clk new_AGEMA_reg_buffer_1731 ( .C (CLK), .D (new_AGEMA_signal_4498), .Q (new_AGEMA_signal_4499) ) ;
    buf_clk new_AGEMA_reg_buffer_1735 ( .C (CLK), .D (new_AGEMA_signal_4502), .Q (new_AGEMA_signal_4503) ) ;
    buf_clk new_AGEMA_reg_buffer_1739 ( .C (CLK), .D (new_AGEMA_signal_4506), .Q (new_AGEMA_signal_4507) ) ;
    buf_clk new_AGEMA_reg_buffer_1743 ( .C (CLK), .D (new_AGEMA_signal_4510), .Q (new_AGEMA_signal_4511) ) ;
    buf_clk new_AGEMA_reg_buffer_1747 ( .C (CLK), .D (new_AGEMA_signal_4514), .Q (new_AGEMA_signal_4515) ) ;
    buf_clk new_AGEMA_reg_buffer_1751 ( .C (CLK), .D (new_AGEMA_signal_4518), .Q (new_AGEMA_signal_4519) ) ;
    buf_clk new_AGEMA_reg_buffer_1755 ( .C (CLK), .D (new_AGEMA_signal_4522), .Q (new_AGEMA_signal_4523) ) ;
    buf_clk new_AGEMA_reg_buffer_1759 ( .C (CLK), .D (new_AGEMA_signal_4526), .Q (new_AGEMA_signal_4527) ) ;
    buf_clk new_AGEMA_reg_buffer_1763 ( .C (CLK), .D (new_AGEMA_signal_4530), .Q (new_AGEMA_signal_4531) ) ;
    buf_clk new_AGEMA_reg_buffer_1767 ( .C (CLK), .D (new_AGEMA_signal_4534), .Q (new_AGEMA_signal_4535) ) ;
    buf_clk new_AGEMA_reg_buffer_1771 ( .C (CLK), .D (new_AGEMA_signal_4538), .Q (new_AGEMA_signal_4539) ) ;
    buf_clk new_AGEMA_reg_buffer_1775 ( .C (CLK), .D (new_AGEMA_signal_4542), .Q (new_AGEMA_signal_4543) ) ;
    buf_clk new_AGEMA_reg_buffer_1779 ( .C (CLK), .D (new_AGEMA_signal_4546), .Q (new_AGEMA_signal_4547) ) ;
    buf_clk new_AGEMA_reg_buffer_1783 ( .C (CLK), .D (new_AGEMA_signal_4550), .Q (new_AGEMA_signal_4551) ) ;
    buf_clk new_AGEMA_reg_buffer_1787 ( .C (CLK), .D (new_AGEMA_signal_4554), .Q (new_AGEMA_signal_4555) ) ;
    buf_clk new_AGEMA_reg_buffer_1791 ( .C (CLK), .D (new_AGEMA_signal_4558), .Q (new_AGEMA_signal_4559) ) ;
    buf_clk new_AGEMA_reg_buffer_1795 ( .C (CLK), .D (new_AGEMA_signal_4562), .Q (new_AGEMA_signal_4563) ) ;
    buf_clk new_AGEMA_reg_buffer_1799 ( .C (CLK), .D (new_AGEMA_signal_4566), .Q (new_AGEMA_signal_4567) ) ;
    buf_clk new_AGEMA_reg_buffer_1803 ( .C (CLK), .D (new_AGEMA_signal_4570), .Q (new_AGEMA_signal_4571) ) ;
    buf_clk new_AGEMA_reg_buffer_1807 ( .C (CLK), .D (new_AGEMA_signal_4574), .Q (new_AGEMA_signal_4575) ) ;
    buf_clk new_AGEMA_reg_buffer_1811 ( .C (CLK), .D (new_AGEMA_signal_4578), .Q (new_AGEMA_signal_4579) ) ;
    buf_clk new_AGEMA_reg_buffer_1815 ( .C (CLK), .D (new_AGEMA_signal_4582), .Q (new_AGEMA_signal_4583) ) ;
    buf_clk new_AGEMA_reg_buffer_1819 ( .C (CLK), .D (new_AGEMA_signal_4586), .Q (new_AGEMA_signal_4587) ) ;
    buf_clk new_AGEMA_reg_buffer_1823 ( .C (CLK), .D (new_AGEMA_signal_4590), .Q (new_AGEMA_signal_4591) ) ;
    buf_clk new_AGEMA_reg_buffer_1827 ( .C (CLK), .D (new_AGEMA_signal_4594), .Q (new_AGEMA_signal_4595) ) ;
    buf_clk new_AGEMA_reg_buffer_1831 ( .C (CLK), .D (new_AGEMA_signal_4598), .Q (new_AGEMA_signal_4599) ) ;
    buf_clk new_AGEMA_reg_buffer_1835 ( .C (CLK), .D (new_AGEMA_signal_4602), .Q (new_AGEMA_signal_4603) ) ;
    buf_clk new_AGEMA_reg_buffer_1839 ( .C (CLK), .D (new_AGEMA_signal_4606), .Q (new_AGEMA_signal_4607) ) ;
    buf_clk new_AGEMA_reg_buffer_1843 ( .C (CLK), .D (new_AGEMA_signal_4610), .Q (new_AGEMA_signal_4611) ) ;
    buf_clk new_AGEMA_reg_buffer_1847 ( .C (CLK), .D (new_AGEMA_signal_4614), .Q (new_AGEMA_signal_4615) ) ;
    buf_clk new_AGEMA_reg_buffer_1851 ( .C (CLK), .D (new_AGEMA_signal_4618), .Q (new_AGEMA_signal_4619) ) ;
    buf_clk new_AGEMA_reg_buffer_1855 ( .C (CLK), .D (new_AGEMA_signal_4622), .Q (new_AGEMA_signal_4623) ) ;
    buf_clk new_AGEMA_reg_buffer_1859 ( .C (CLK), .D (new_AGEMA_signal_4626), .Q (new_AGEMA_signal_4627) ) ;
    buf_clk new_AGEMA_reg_buffer_1863 ( .C (CLK), .D (new_AGEMA_signal_4630), .Q (new_AGEMA_signal_4631) ) ;
    buf_clk new_AGEMA_reg_buffer_1867 ( .C (CLK), .D (new_AGEMA_signal_4634), .Q (new_AGEMA_signal_4635) ) ;
    buf_clk new_AGEMA_reg_buffer_1871 ( .C (CLK), .D (new_AGEMA_signal_4638), .Q (new_AGEMA_signal_4639) ) ;
    buf_clk new_AGEMA_reg_buffer_1875 ( .C (CLK), .D (new_AGEMA_signal_4642), .Q (new_AGEMA_signal_4643) ) ;
    buf_clk new_AGEMA_reg_buffer_1879 ( .C (CLK), .D (new_AGEMA_signal_4646), .Q (new_AGEMA_signal_4647) ) ;
    buf_clk new_AGEMA_reg_buffer_1883 ( .C (CLK), .D (new_AGEMA_signal_4650), .Q (new_AGEMA_signal_4651) ) ;
    buf_clk new_AGEMA_reg_buffer_1887 ( .C (CLK), .D (new_AGEMA_signal_4654), .Q (new_AGEMA_signal_4655) ) ;
    buf_clk new_AGEMA_reg_buffer_1891 ( .C (CLK), .D (new_AGEMA_signal_4658), .Q (new_AGEMA_signal_4659) ) ;
    buf_clk new_AGEMA_reg_buffer_1895 ( .C (CLK), .D (new_AGEMA_signal_4662), .Q (new_AGEMA_signal_4663) ) ;
    buf_clk new_AGEMA_reg_buffer_1899 ( .C (CLK), .D (new_AGEMA_signal_4666), .Q (new_AGEMA_signal_4667) ) ;
    buf_clk new_AGEMA_reg_buffer_1903 ( .C (CLK), .D (new_AGEMA_signal_4670), .Q (new_AGEMA_signal_4671) ) ;
    buf_clk new_AGEMA_reg_buffer_1907 ( .C (CLK), .D (new_AGEMA_signal_4674), .Q (new_AGEMA_signal_4675) ) ;
    buf_clk new_AGEMA_reg_buffer_1911 ( .C (CLK), .D (new_AGEMA_signal_4678), .Q (new_AGEMA_signal_4679) ) ;
    buf_clk new_AGEMA_reg_buffer_1915 ( .C (CLK), .D (new_AGEMA_signal_4682), .Q (new_AGEMA_signal_4683) ) ;
    buf_clk new_AGEMA_reg_buffer_1919 ( .C (CLK), .D (new_AGEMA_signal_4686), .Q (new_AGEMA_signal_4687) ) ;
    buf_clk new_AGEMA_reg_buffer_1923 ( .C (CLK), .D (new_AGEMA_signal_4690), .Q (new_AGEMA_signal_4691) ) ;
    buf_clk new_AGEMA_reg_buffer_1927 ( .C (CLK), .D (new_AGEMA_signal_4694), .Q (new_AGEMA_signal_4695) ) ;
    buf_clk new_AGEMA_reg_buffer_1931 ( .C (CLK), .D (new_AGEMA_signal_4698), .Q (new_AGEMA_signal_4699) ) ;
    buf_clk new_AGEMA_reg_buffer_1935 ( .C (CLK), .D (new_AGEMA_signal_4702), .Q (new_AGEMA_signal_4703) ) ;
    buf_clk new_AGEMA_reg_buffer_1939 ( .C (CLK), .D (new_AGEMA_signal_4706), .Q (new_AGEMA_signal_4707) ) ;
    buf_clk new_AGEMA_reg_buffer_1943 ( .C (CLK), .D (new_AGEMA_signal_4710), .Q (new_AGEMA_signal_4711) ) ;
    buf_clk new_AGEMA_reg_buffer_1947 ( .C (CLK), .D (new_AGEMA_signal_4714), .Q (new_AGEMA_signal_4715) ) ;
    buf_clk new_AGEMA_reg_buffer_1951 ( .C (CLK), .D (new_AGEMA_signal_4718), .Q (new_AGEMA_signal_4719) ) ;
    buf_clk new_AGEMA_reg_buffer_1955 ( .C (CLK), .D (new_AGEMA_signal_4722), .Q (new_AGEMA_signal_4723) ) ;
    buf_clk new_AGEMA_reg_buffer_1959 ( .C (CLK), .D (new_AGEMA_signal_4726), .Q (new_AGEMA_signal_4727) ) ;
    buf_clk new_AGEMA_reg_buffer_1963 ( .C (CLK), .D (new_AGEMA_signal_4730), .Q (new_AGEMA_signal_4731) ) ;
    buf_clk new_AGEMA_reg_buffer_1967 ( .C (CLK), .D (new_AGEMA_signal_4734), .Q (new_AGEMA_signal_4735) ) ;
    buf_clk new_AGEMA_reg_buffer_1971 ( .C (CLK), .D (new_AGEMA_signal_4738), .Q (new_AGEMA_signal_4739) ) ;
    buf_clk new_AGEMA_reg_buffer_1975 ( .C (CLK), .D (new_AGEMA_signal_4742), .Q (new_AGEMA_signal_4743) ) ;
    buf_clk new_AGEMA_reg_buffer_1979 ( .C (CLK), .D (new_AGEMA_signal_4746), .Q (new_AGEMA_signal_4747) ) ;
    buf_clk new_AGEMA_reg_buffer_1983 ( .C (CLK), .D (new_AGEMA_signal_4750), .Q (new_AGEMA_signal_4751) ) ;
    buf_clk new_AGEMA_reg_buffer_1987 ( .C (CLK), .D (new_AGEMA_signal_4754), .Q (new_AGEMA_signal_4755) ) ;
    buf_clk new_AGEMA_reg_buffer_1991 ( .C (CLK), .D (new_AGEMA_signal_4758), .Q (new_AGEMA_signal_4759) ) ;
    buf_clk new_AGEMA_reg_buffer_1995 ( .C (CLK), .D (new_AGEMA_signal_4762), .Q (new_AGEMA_signal_4763) ) ;
    buf_clk new_AGEMA_reg_buffer_1999 ( .C (CLK), .D (new_AGEMA_signal_4766), .Q (new_AGEMA_signal_4767) ) ;
    buf_clk new_AGEMA_reg_buffer_2003 ( .C (CLK), .D (new_AGEMA_signal_4770), .Q (new_AGEMA_signal_4771) ) ;
    buf_clk new_AGEMA_reg_buffer_2007 ( .C (CLK), .D (new_AGEMA_signal_4774), .Q (new_AGEMA_signal_4775) ) ;
    buf_clk new_AGEMA_reg_buffer_2011 ( .C (CLK), .D (new_AGEMA_signal_4778), .Q (new_AGEMA_signal_4779) ) ;
    buf_clk new_AGEMA_reg_buffer_2015 ( .C (CLK), .D (new_AGEMA_signal_4782), .Q (new_AGEMA_signal_4783) ) ;
    buf_clk new_AGEMA_reg_buffer_2019 ( .C (CLK), .D (new_AGEMA_signal_4786), .Q (new_AGEMA_signal_4787) ) ;
    buf_clk new_AGEMA_reg_buffer_2023 ( .C (CLK), .D (new_AGEMA_signal_4790), .Q (new_AGEMA_signal_4791) ) ;
    buf_clk new_AGEMA_reg_buffer_2027 ( .C (CLK), .D (new_AGEMA_signal_4794), .Q (new_AGEMA_signal_4795) ) ;
    buf_clk new_AGEMA_reg_buffer_2031 ( .C (CLK), .D (new_AGEMA_signal_4798), .Q (new_AGEMA_signal_4799) ) ;
    buf_clk new_AGEMA_reg_buffer_2035 ( .C (CLK), .D (new_AGEMA_signal_4802), .Q (new_AGEMA_signal_4803) ) ;
    buf_clk new_AGEMA_reg_buffer_2039 ( .C (CLK), .D (new_AGEMA_signal_4806), .Q (new_AGEMA_signal_4807) ) ;
    buf_clk new_AGEMA_reg_buffer_2043 ( .C (CLK), .D (new_AGEMA_signal_4810), .Q (new_AGEMA_signal_4811) ) ;
    buf_clk new_AGEMA_reg_buffer_2047 ( .C (CLK), .D (new_AGEMA_signal_4814), .Q (new_AGEMA_signal_4815) ) ;
    buf_clk new_AGEMA_reg_buffer_2051 ( .C (CLK), .D (new_AGEMA_signal_4818), .Q (new_AGEMA_signal_4819) ) ;
    buf_clk new_AGEMA_reg_buffer_2055 ( .C (CLK), .D (new_AGEMA_signal_4822), .Q (new_AGEMA_signal_4823) ) ;
    buf_clk new_AGEMA_reg_buffer_2059 ( .C (CLK), .D (new_AGEMA_signal_4826), .Q (new_AGEMA_signal_4827) ) ;
    buf_clk new_AGEMA_reg_buffer_2063 ( .C (CLK), .D (new_AGEMA_signal_4830), .Q (new_AGEMA_signal_4831) ) ;
    buf_clk new_AGEMA_reg_buffer_2067 ( .C (CLK), .D (new_AGEMA_signal_4834), .Q (new_AGEMA_signal_4835) ) ;
    buf_clk new_AGEMA_reg_buffer_2071 ( .C (CLK), .D (new_AGEMA_signal_4838), .Q (new_AGEMA_signal_4839) ) ;
    buf_clk new_AGEMA_reg_buffer_2075 ( .C (CLK), .D (new_AGEMA_signal_4842), .Q (new_AGEMA_signal_4843) ) ;
    buf_clk new_AGEMA_reg_buffer_2079 ( .C (CLK), .D (new_AGEMA_signal_4846), .Q (new_AGEMA_signal_4847) ) ;
    buf_clk new_AGEMA_reg_buffer_2083 ( .C (CLK), .D (new_AGEMA_signal_4850), .Q (new_AGEMA_signal_4851) ) ;
    buf_clk new_AGEMA_reg_buffer_2087 ( .C (CLK), .D (new_AGEMA_signal_4854), .Q (new_AGEMA_signal_4855) ) ;
    buf_clk new_AGEMA_reg_buffer_2091 ( .C (CLK), .D (new_AGEMA_signal_4858), .Q (new_AGEMA_signal_4859) ) ;
    buf_clk new_AGEMA_reg_buffer_2095 ( .C (CLK), .D (new_AGEMA_signal_4862), .Q (new_AGEMA_signal_4863) ) ;
    buf_clk new_AGEMA_reg_buffer_2099 ( .C (CLK), .D (new_AGEMA_signal_4866), .Q (new_AGEMA_signal_4867) ) ;
    buf_clk new_AGEMA_reg_buffer_2103 ( .C (CLK), .D (new_AGEMA_signal_4870), .Q (new_AGEMA_signal_4871) ) ;
    buf_clk new_AGEMA_reg_buffer_2107 ( .C (CLK), .D (new_AGEMA_signal_4874), .Q (new_AGEMA_signal_4875) ) ;
    buf_clk new_AGEMA_reg_buffer_2111 ( .C (CLK), .D (new_AGEMA_signal_4878), .Q (new_AGEMA_signal_4879) ) ;
    buf_clk new_AGEMA_reg_buffer_2115 ( .C (CLK), .D (new_AGEMA_signal_4882), .Q (new_AGEMA_signal_4883) ) ;
    buf_clk new_AGEMA_reg_buffer_2119 ( .C (CLK), .D (new_AGEMA_signal_4886), .Q (new_AGEMA_signal_4887) ) ;
    buf_clk new_AGEMA_reg_buffer_2123 ( .C (CLK), .D (new_AGEMA_signal_4890), .Q (new_AGEMA_signal_4891) ) ;
    buf_clk new_AGEMA_reg_buffer_2127 ( .C (CLK), .D (new_AGEMA_signal_4894), .Q (new_AGEMA_signal_4895) ) ;
    buf_clk new_AGEMA_reg_buffer_2131 ( .C (CLK), .D (new_AGEMA_signal_4898), .Q (new_AGEMA_signal_4899) ) ;
    buf_clk new_AGEMA_reg_buffer_2135 ( .C (CLK), .D (new_AGEMA_signal_4902), .Q (new_AGEMA_signal_4903) ) ;
    buf_clk new_AGEMA_reg_buffer_2139 ( .C (CLK), .D (new_AGEMA_signal_4906), .Q (new_AGEMA_signal_4907) ) ;
    buf_clk new_AGEMA_reg_buffer_2143 ( .C (CLK), .D (new_AGEMA_signal_4910), .Q (new_AGEMA_signal_4911) ) ;
    buf_clk new_AGEMA_reg_buffer_2147 ( .C (CLK), .D (new_AGEMA_signal_4914), .Q (new_AGEMA_signal_4915) ) ;
    buf_clk new_AGEMA_reg_buffer_2151 ( .C (CLK), .D (new_AGEMA_signal_4918), .Q (new_AGEMA_signal_4919) ) ;
    buf_clk new_AGEMA_reg_buffer_2155 ( .C (CLK), .D (new_AGEMA_signal_4922), .Q (new_AGEMA_signal_4923) ) ;
    buf_clk new_AGEMA_reg_buffer_2159 ( .C (CLK), .D (new_AGEMA_signal_4926), .Q (new_AGEMA_signal_4927) ) ;
    buf_clk new_AGEMA_reg_buffer_2163 ( .C (CLK), .D (new_AGEMA_signal_4930), .Q (new_AGEMA_signal_4931) ) ;
    buf_clk new_AGEMA_reg_buffer_2167 ( .C (CLK), .D (new_AGEMA_signal_4934), .Q (new_AGEMA_signal_4935) ) ;
    buf_clk new_AGEMA_reg_buffer_2171 ( .C (CLK), .D (new_AGEMA_signal_4938), .Q (new_AGEMA_signal_4939) ) ;
    buf_clk new_AGEMA_reg_buffer_2175 ( .C (CLK), .D (new_AGEMA_signal_4942), .Q (new_AGEMA_signal_4943) ) ;
    buf_clk new_AGEMA_reg_buffer_2179 ( .C (CLK), .D (new_AGEMA_signal_4946), .Q (new_AGEMA_signal_4947) ) ;
    buf_clk new_AGEMA_reg_buffer_2183 ( .C (CLK), .D (new_AGEMA_signal_4950), .Q (new_AGEMA_signal_4951) ) ;
    buf_clk new_AGEMA_reg_buffer_2187 ( .C (CLK), .D (new_AGEMA_signal_4954), .Q (new_AGEMA_signal_4955) ) ;
    buf_clk new_AGEMA_reg_buffer_2191 ( .C (CLK), .D (new_AGEMA_signal_4958), .Q (new_AGEMA_signal_4959) ) ;
    buf_clk new_AGEMA_reg_buffer_2195 ( .C (CLK), .D (new_AGEMA_signal_4962), .Q (new_AGEMA_signal_4963) ) ;
    buf_clk new_AGEMA_reg_buffer_2199 ( .C (CLK), .D (new_AGEMA_signal_4966), .Q (new_AGEMA_signal_4967) ) ;
    buf_clk new_AGEMA_reg_buffer_2203 ( .C (CLK), .D (new_AGEMA_signal_4970), .Q (new_AGEMA_signal_4971) ) ;
    buf_clk new_AGEMA_reg_buffer_2207 ( .C (CLK), .D (new_AGEMA_signal_4974), .Q (new_AGEMA_signal_4975) ) ;
    buf_clk new_AGEMA_reg_buffer_2211 ( .C (CLK), .D (new_AGEMA_signal_4978), .Q (new_AGEMA_signal_4979) ) ;
    buf_clk new_AGEMA_reg_buffer_2215 ( .C (CLK), .D (new_AGEMA_signal_4982), .Q (new_AGEMA_signal_4983) ) ;
    buf_clk new_AGEMA_reg_buffer_2219 ( .C (CLK), .D (new_AGEMA_signal_4986), .Q (new_AGEMA_signal_4987) ) ;
    buf_clk new_AGEMA_reg_buffer_2223 ( .C (CLK), .D (new_AGEMA_signal_4990), .Q (new_AGEMA_signal_4991) ) ;
    buf_clk new_AGEMA_reg_buffer_2227 ( .C (CLK), .D (new_AGEMA_signal_4994), .Q (new_AGEMA_signal_4995) ) ;
    buf_clk new_AGEMA_reg_buffer_2231 ( .C (CLK), .D (new_AGEMA_signal_4998), .Q (new_AGEMA_signal_4999) ) ;
    buf_clk new_AGEMA_reg_buffer_2235 ( .C (CLK), .D (new_AGEMA_signal_5002), .Q (new_AGEMA_signal_5003) ) ;
    buf_clk new_AGEMA_reg_buffer_2239 ( .C (CLK), .D (new_AGEMA_signal_5006), .Q (new_AGEMA_signal_5007) ) ;
    buf_clk new_AGEMA_reg_buffer_2243 ( .C (CLK), .D (new_AGEMA_signal_5010), .Q (new_AGEMA_signal_5011) ) ;
    buf_clk new_AGEMA_reg_buffer_2247 ( .C (CLK), .D (new_AGEMA_signal_5014), .Q (new_AGEMA_signal_5015) ) ;
    buf_clk new_AGEMA_reg_buffer_2251 ( .C (CLK), .D (new_AGEMA_signal_5018), .Q (new_AGEMA_signal_5019) ) ;
    buf_clk new_AGEMA_reg_buffer_2255 ( .C (CLK), .D (new_AGEMA_signal_5022), .Q (new_AGEMA_signal_5023) ) ;
    buf_clk new_AGEMA_reg_buffer_2259 ( .C (CLK), .D (new_AGEMA_signal_5026), .Q (new_AGEMA_signal_5027) ) ;
    buf_clk new_AGEMA_reg_buffer_2263 ( .C (CLK), .D (new_AGEMA_signal_5030), .Q (new_AGEMA_signal_5031) ) ;
    buf_clk new_AGEMA_reg_buffer_2267 ( .C (CLK), .D (new_AGEMA_signal_5034), .Q (new_AGEMA_signal_5035) ) ;
    buf_clk new_AGEMA_reg_buffer_2271 ( .C (CLK), .D (new_AGEMA_signal_5038), .Q (new_AGEMA_signal_5039) ) ;
    buf_clk new_AGEMA_reg_buffer_2275 ( .C (CLK), .D (new_AGEMA_signal_5042), .Q (new_AGEMA_signal_5043) ) ;
    buf_clk new_AGEMA_reg_buffer_2279 ( .C (CLK), .D (new_AGEMA_signal_5046), .Q (new_AGEMA_signal_5047) ) ;
    buf_clk new_AGEMA_reg_buffer_2283 ( .C (CLK), .D (new_AGEMA_signal_5050), .Q (new_AGEMA_signal_5051) ) ;
    buf_clk new_AGEMA_reg_buffer_2287 ( .C (CLK), .D (new_AGEMA_signal_5054), .Q (new_AGEMA_signal_5055) ) ;
    buf_clk new_AGEMA_reg_buffer_2291 ( .C (CLK), .D (new_AGEMA_signal_5058), .Q (new_AGEMA_signal_5059) ) ;
    buf_clk new_AGEMA_reg_buffer_2295 ( .C (CLK), .D (new_AGEMA_signal_5062), .Q (new_AGEMA_signal_5063) ) ;
    buf_clk new_AGEMA_reg_buffer_2299 ( .C (CLK), .D (new_AGEMA_signal_5066), .Q (new_AGEMA_signal_5067) ) ;
    buf_clk new_AGEMA_reg_buffer_2303 ( .C (CLK), .D (new_AGEMA_signal_5070), .Q (new_AGEMA_signal_5071) ) ;
    buf_clk new_AGEMA_reg_buffer_2307 ( .C (CLK), .D (new_AGEMA_signal_5074), .Q (new_AGEMA_signal_5075) ) ;
    buf_clk new_AGEMA_reg_buffer_2311 ( .C (CLK), .D (new_AGEMA_signal_5078), .Q (new_AGEMA_signal_5079) ) ;
    buf_clk new_AGEMA_reg_buffer_2315 ( .C (CLK), .D (new_AGEMA_signal_5082), .Q (new_AGEMA_signal_5083) ) ;
    buf_clk new_AGEMA_reg_buffer_2319 ( .C (CLK), .D (new_AGEMA_signal_5086), .Q (new_AGEMA_signal_5087) ) ;
    buf_clk new_AGEMA_reg_buffer_2323 ( .C (CLK), .D (new_AGEMA_signal_5090), .Q (new_AGEMA_signal_5091) ) ;
    buf_clk new_AGEMA_reg_buffer_2327 ( .C (CLK), .D (new_AGEMA_signal_5094), .Q (new_AGEMA_signal_5095) ) ;
    buf_clk new_AGEMA_reg_buffer_2331 ( .C (CLK), .D (new_AGEMA_signal_5098), .Q (new_AGEMA_signal_5099) ) ;
    buf_clk new_AGEMA_reg_buffer_2335 ( .C (CLK), .D (new_AGEMA_signal_5102), .Q (new_AGEMA_signal_5103) ) ;
    buf_clk new_AGEMA_reg_buffer_2339 ( .C (CLK), .D (new_AGEMA_signal_5106), .Q (new_AGEMA_signal_5107) ) ;
    buf_clk new_AGEMA_reg_buffer_2343 ( .C (CLK), .D (new_AGEMA_signal_5110), .Q (new_AGEMA_signal_5111) ) ;
    buf_clk new_AGEMA_reg_buffer_2347 ( .C (CLK), .D (new_AGEMA_signal_5114), .Q (new_AGEMA_signal_5115) ) ;
    buf_clk new_AGEMA_reg_buffer_2351 ( .C (CLK), .D (new_AGEMA_signal_5118), .Q (new_AGEMA_signal_5119) ) ;
    buf_clk new_AGEMA_reg_buffer_2355 ( .C (CLK), .D (new_AGEMA_signal_5122), .Q (new_AGEMA_signal_5123) ) ;
    buf_clk new_AGEMA_reg_buffer_2359 ( .C (CLK), .D (new_AGEMA_signal_5126), .Q (new_AGEMA_signal_5127) ) ;
    buf_clk new_AGEMA_reg_buffer_2363 ( .C (CLK), .D (new_AGEMA_signal_5130), .Q (new_AGEMA_signal_5131) ) ;
    buf_clk new_AGEMA_reg_buffer_2367 ( .C (CLK), .D (new_AGEMA_signal_5134), .Q (new_AGEMA_signal_5135) ) ;
    buf_clk new_AGEMA_reg_buffer_2371 ( .C (CLK), .D (new_AGEMA_signal_5138), .Q (new_AGEMA_signal_5139) ) ;
    buf_clk new_AGEMA_reg_buffer_2375 ( .C (CLK), .D (new_AGEMA_signal_5142), .Q (new_AGEMA_signal_5143) ) ;
    buf_clk new_AGEMA_reg_buffer_2379 ( .C (CLK), .D (new_AGEMA_signal_5146), .Q (new_AGEMA_signal_5147) ) ;
    buf_clk new_AGEMA_reg_buffer_2383 ( .C (CLK), .D (new_AGEMA_signal_5150), .Q (new_AGEMA_signal_5151) ) ;
    buf_clk new_AGEMA_reg_buffer_2387 ( .C (CLK), .D (new_AGEMA_signal_5154), .Q (new_AGEMA_signal_5155) ) ;
    buf_clk new_AGEMA_reg_buffer_2391 ( .C (CLK), .D (new_AGEMA_signal_5158), .Q (new_AGEMA_signal_5159) ) ;
    buf_clk new_AGEMA_reg_buffer_2395 ( .C (CLK), .D (new_AGEMA_signal_5162), .Q (new_AGEMA_signal_5163) ) ;
    buf_clk new_AGEMA_reg_buffer_2399 ( .C (CLK), .D (new_AGEMA_signal_5166), .Q (new_AGEMA_signal_5167) ) ;
    buf_clk new_AGEMA_reg_buffer_2403 ( .C (CLK), .D (new_AGEMA_signal_5170), .Q (new_AGEMA_signal_5171) ) ;
    buf_clk new_AGEMA_reg_buffer_2407 ( .C (CLK), .D (new_AGEMA_signal_5174), .Q (new_AGEMA_signal_5175) ) ;
    buf_clk new_AGEMA_reg_buffer_2411 ( .C (CLK), .D (new_AGEMA_signal_5178), .Q (new_AGEMA_signal_5179) ) ;
    buf_clk new_AGEMA_reg_buffer_2415 ( .C (CLK), .D (new_AGEMA_signal_5182), .Q (new_AGEMA_signal_5183) ) ;
    buf_clk new_AGEMA_reg_buffer_2419 ( .C (CLK), .D (new_AGEMA_signal_5186), .Q (new_AGEMA_signal_5187) ) ;
    buf_clk new_AGEMA_reg_buffer_2423 ( .C (CLK), .D (new_AGEMA_signal_5190), .Q (new_AGEMA_signal_5191) ) ;
    buf_clk new_AGEMA_reg_buffer_2427 ( .C (CLK), .D (new_AGEMA_signal_5194), .Q (new_AGEMA_signal_5195) ) ;
    buf_clk new_AGEMA_reg_buffer_2431 ( .C (CLK), .D (new_AGEMA_signal_5198), .Q (new_AGEMA_signal_5199) ) ;
    buf_clk new_AGEMA_reg_buffer_2435 ( .C (CLK), .D (new_AGEMA_signal_5202), .Q (new_AGEMA_signal_5203) ) ;
    buf_clk new_AGEMA_reg_buffer_2439 ( .C (CLK), .D (new_AGEMA_signal_5206), .Q (new_AGEMA_signal_5207) ) ;
    buf_clk new_AGEMA_reg_buffer_2443 ( .C (CLK), .D (new_AGEMA_signal_5210), .Q (new_AGEMA_signal_5211) ) ;
    buf_clk new_AGEMA_reg_buffer_2447 ( .C (CLK), .D (new_AGEMA_signal_5214), .Q (new_AGEMA_signal_5215) ) ;
    buf_clk new_AGEMA_reg_buffer_2451 ( .C (CLK), .D (new_AGEMA_signal_5218), .Q (new_AGEMA_signal_5219) ) ;
    buf_clk new_AGEMA_reg_buffer_2455 ( .C (CLK), .D (new_AGEMA_signal_5222), .Q (new_AGEMA_signal_5223) ) ;
    buf_clk new_AGEMA_reg_buffer_2459 ( .C (CLK), .D (new_AGEMA_signal_5226), .Q (new_AGEMA_signal_5227) ) ;
    buf_clk new_AGEMA_reg_buffer_2463 ( .C (CLK), .D (new_AGEMA_signal_5230), .Q (new_AGEMA_signal_5231) ) ;
    buf_clk new_AGEMA_reg_buffer_2467 ( .C (CLK), .D (new_AGEMA_signal_5234), .Q (new_AGEMA_signal_5235) ) ;
    buf_clk new_AGEMA_reg_buffer_2471 ( .C (CLK), .D (new_AGEMA_signal_5238), .Q (new_AGEMA_signal_5239) ) ;
    buf_clk new_AGEMA_reg_buffer_2475 ( .C (CLK), .D (new_AGEMA_signal_5242), .Q (new_AGEMA_signal_5243) ) ;
    buf_clk new_AGEMA_reg_buffer_2479 ( .C (CLK), .D (new_AGEMA_signal_5246), .Q (new_AGEMA_signal_5247) ) ;
    buf_clk new_AGEMA_reg_buffer_2483 ( .C (CLK), .D (new_AGEMA_signal_5250), .Q (new_AGEMA_signal_5251) ) ;
    buf_clk new_AGEMA_reg_buffer_2487 ( .C (CLK), .D (new_AGEMA_signal_5254), .Q (new_AGEMA_signal_5255) ) ;
    buf_clk new_AGEMA_reg_buffer_2491 ( .C (CLK), .D (new_AGEMA_signal_5258), .Q (new_AGEMA_signal_5259) ) ;
    buf_clk new_AGEMA_reg_buffer_2495 ( .C (CLK), .D (new_AGEMA_signal_5262), .Q (new_AGEMA_signal_5263) ) ;
    buf_clk new_AGEMA_reg_buffer_2499 ( .C (CLK), .D (new_AGEMA_signal_5266), .Q (new_AGEMA_signal_5267) ) ;
    buf_clk new_AGEMA_reg_buffer_2503 ( .C (CLK), .D (new_AGEMA_signal_5270), .Q (new_AGEMA_signal_5271) ) ;
    buf_clk new_AGEMA_reg_buffer_2507 ( .C (CLK), .D (new_AGEMA_signal_5274), .Q (new_AGEMA_signal_5275) ) ;
    buf_clk new_AGEMA_reg_buffer_2511 ( .C (CLK), .D (new_AGEMA_signal_5278), .Q (new_AGEMA_signal_5279) ) ;
    buf_clk new_AGEMA_reg_buffer_2515 ( .C (CLK), .D (new_AGEMA_signal_5282), .Q (new_AGEMA_signal_5283) ) ;
    buf_clk new_AGEMA_reg_buffer_2519 ( .C (CLK), .D (new_AGEMA_signal_5286), .Q (new_AGEMA_signal_5287) ) ;
    buf_clk new_AGEMA_reg_buffer_2523 ( .C (CLK), .D (new_AGEMA_signal_5290), .Q (new_AGEMA_signal_5291) ) ;
    buf_clk new_AGEMA_reg_buffer_2527 ( .C (CLK), .D (new_AGEMA_signal_5294), .Q (new_AGEMA_signal_5295) ) ;
    buf_clk new_AGEMA_reg_buffer_2531 ( .C (CLK), .D (new_AGEMA_signal_5298), .Q (new_AGEMA_signal_5299) ) ;
    buf_clk new_AGEMA_reg_buffer_2535 ( .C (CLK), .D (new_AGEMA_signal_5302), .Q (new_AGEMA_signal_5303) ) ;
    buf_clk new_AGEMA_reg_buffer_2539 ( .C (CLK), .D (new_AGEMA_signal_5306), .Q (new_AGEMA_signal_5307) ) ;
    buf_clk new_AGEMA_reg_buffer_2543 ( .C (CLK), .D (new_AGEMA_signal_5310), .Q (new_AGEMA_signal_5311) ) ;
    buf_clk new_AGEMA_reg_buffer_2547 ( .C (CLK), .D (new_AGEMA_signal_5314), .Q (new_AGEMA_signal_5315) ) ;
    buf_clk new_AGEMA_reg_buffer_2551 ( .C (CLK), .D (new_AGEMA_signal_5318), .Q (new_AGEMA_signal_5319) ) ;
    buf_clk new_AGEMA_reg_buffer_2555 ( .C (CLK), .D (new_AGEMA_signal_5322), .Q (new_AGEMA_signal_5323) ) ;
    buf_clk new_AGEMA_reg_buffer_2559 ( .C (CLK), .D (new_AGEMA_signal_5326), .Q (new_AGEMA_signal_5327) ) ;
    buf_clk new_AGEMA_reg_buffer_2563 ( .C (CLK), .D (new_AGEMA_signal_5330), .Q (new_AGEMA_signal_5331) ) ;
    buf_clk new_AGEMA_reg_buffer_2567 ( .C (CLK), .D (new_AGEMA_signal_5334), .Q (new_AGEMA_signal_5335) ) ;
    buf_clk new_AGEMA_reg_buffer_2571 ( .C (CLK), .D (new_AGEMA_signal_5338), .Q (new_AGEMA_signal_5339) ) ;
    buf_clk new_AGEMA_reg_buffer_2575 ( .C (CLK), .D (new_AGEMA_signal_5342), .Q (new_AGEMA_signal_5343) ) ;
    buf_clk new_AGEMA_reg_buffer_2579 ( .C (CLK), .D (new_AGEMA_signal_5346), .Q (new_AGEMA_signal_5347) ) ;
    buf_clk new_AGEMA_reg_buffer_2583 ( .C (CLK), .D (new_AGEMA_signal_5350), .Q (new_AGEMA_signal_5351) ) ;
    buf_clk new_AGEMA_reg_buffer_2587 ( .C (CLK), .D (new_AGEMA_signal_5354), .Q (new_AGEMA_signal_5355) ) ;
    buf_clk new_AGEMA_reg_buffer_2591 ( .C (CLK), .D (new_AGEMA_signal_5358), .Q (new_AGEMA_signal_5359) ) ;
    buf_clk new_AGEMA_reg_buffer_2595 ( .C (CLK), .D (new_AGEMA_signal_5362), .Q (new_AGEMA_signal_5363) ) ;
    buf_clk new_AGEMA_reg_buffer_2599 ( .C (CLK), .D (new_AGEMA_signal_5366), .Q (new_AGEMA_signal_5367) ) ;
    buf_clk new_AGEMA_reg_buffer_2603 ( .C (CLK), .D (new_AGEMA_signal_5370), .Q (new_AGEMA_signal_5371) ) ;
    buf_clk new_AGEMA_reg_buffer_2607 ( .C (CLK), .D (new_AGEMA_signal_5374), .Q (new_AGEMA_signal_5375) ) ;
    buf_clk new_AGEMA_reg_buffer_2611 ( .C (CLK), .D (new_AGEMA_signal_5378), .Q (new_AGEMA_signal_5379) ) ;
    buf_clk new_AGEMA_reg_buffer_2615 ( .C (CLK), .D (new_AGEMA_signal_5382), .Q (new_AGEMA_signal_5383) ) ;
    buf_clk new_AGEMA_reg_buffer_2619 ( .C (CLK), .D (new_AGEMA_signal_5386), .Q (new_AGEMA_signal_5387) ) ;
    buf_clk new_AGEMA_reg_buffer_2623 ( .C (CLK), .D (new_AGEMA_signal_5390), .Q (new_AGEMA_signal_5391) ) ;
    buf_clk new_AGEMA_reg_buffer_2627 ( .C (CLK), .D (new_AGEMA_signal_5394), .Q (new_AGEMA_signal_5395) ) ;
    buf_clk new_AGEMA_reg_buffer_2631 ( .C (CLK), .D (new_AGEMA_signal_5398), .Q (new_AGEMA_signal_5399) ) ;
    buf_clk new_AGEMA_reg_buffer_2635 ( .C (CLK), .D (new_AGEMA_signal_5402), .Q (new_AGEMA_signal_5403) ) ;
    buf_clk new_AGEMA_reg_buffer_2639 ( .C (CLK), .D (new_AGEMA_signal_5406), .Q (new_AGEMA_signal_5407) ) ;
    buf_clk new_AGEMA_reg_buffer_2643 ( .C (CLK), .D (new_AGEMA_signal_5410), .Q (new_AGEMA_signal_5411) ) ;
    buf_clk new_AGEMA_reg_buffer_2647 ( .C (CLK), .D (new_AGEMA_signal_5414), .Q (new_AGEMA_signal_5415) ) ;
    buf_clk new_AGEMA_reg_buffer_2651 ( .C (CLK), .D (new_AGEMA_signal_5418), .Q (new_AGEMA_signal_5419) ) ;
    buf_clk new_AGEMA_reg_buffer_2655 ( .C (CLK), .D (new_AGEMA_signal_5422), .Q (new_AGEMA_signal_5423) ) ;
    buf_clk new_AGEMA_reg_buffer_2659 ( .C (CLK), .D (new_AGEMA_signal_5426), .Q (new_AGEMA_signal_5427) ) ;
    buf_clk new_AGEMA_reg_buffer_2663 ( .C (CLK), .D (new_AGEMA_signal_5430), .Q (new_AGEMA_signal_5431) ) ;
    buf_clk new_AGEMA_reg_buffer_2667 ( .C (CLK), .D (new_AGEMA_signal_5434), .Q (new_AGEMA_signal_5435) ) ;
    buf_clk new_AGEMA_reg_buffer_2671 ( .C (CLK), .D (new_AGEMA_signal_5438), .Q (new_AGEMA_signal_5439) ) ;
    buf_clk new_AGEMA_reg_buffer_2675 ( .C (CLK), .D (new_AGEMA_signal_5442), .Q (new_AGEMA_signal_5443) ) ;
    buf_clk new_AGEMA_reg_buffer_2679 ( .C (CLK), .D (new_AGEMA_signal_5446), .Q (new_AGEMA_signal_5447) ) ;
    buf_clk new_AGEMA_reg_buffer_2683 ( .C (CLK), .D (new_AGEMA_signal_5450), .Q (new_AGEMA_signal_5451) ) ;
    buf_clk new_AGEMA_reg_buffer_2687 ( .C (CLK), .D (new_AGEMA_signal_5454), .Q (new_AGEMA_signal_5455) ) ;
    buf_clk new_AGEMA_reg_buffer_2691 ( .C (CLK), .D (new_AGEMA_signal_5458), .Q (new_AGEMA_signal_5459) ) ;
    buf_clk new_AGEMA_reg_buffer_2695 ( .C (CLK), .D (new_AGEMA_signal_5462), .Q (new_AGEMA_signal_5463) ) ;
    buf_clk new_AGEMA_reg_buffer_2699 ( .C (CLK), .D (new_AGEMA_signal_5466), .Q (new_AGEMA_signal_5467) ) ;
    buf_clk new_AGEMA_reg_buffer_2703 ( .C (CLK), .D (new_AGEMA_signal_5470), .Q (new_AGEMA_signal_5471) ) ;
    buf_clk new_AGEMA_reg_buffer_2707 ( .C (CLK), .D (new_AGEMA_signal_5474), .Q (new_AGEMA_signal_5475) ) ;
    buf_clk new_AGEMA_reg_buffer_2711 ( .C (CLK), .D (new_AGEMA_signal_5478), .Q (new_AGEMA_signal_5479) ) ;
    buf_clk new_AGEMA_reg_buffer_2715 ( .C (CLK), .D (new_AGEMA_signal_5482), .Q (new_AGEMA_signal_5483) ) ;
    buf_clk new_AGEMA_reg_buffer_2719 ( .C (CLK), .D (new_AGEMA_signal_5486), .Q (new_AGEMA_signal_5487) ) ;
    buf_clk new_AGEMA_reg_buffer_2723 ( .C (CLK), .D (new_AGEMA_signal_5490), .Q (new_AGEMA_signal_5491) ) ;
    buf_clk new_AGEMA_reg_buffer_2727 ( .C (CLK), .D (new_AGEMA_signal_5494), .Q (new_AGEMA_signal_5495) ) ;
    buf_clk new_AGEMA_reg_buffer_2731 ( .C (CLK), .D (new_AGEMA_signal_5498), .Q (new_AGEMA_signal_5499) ) ;
    buf_clk new_AGEMA_reg_buffer_2735 ( .C (CLK), .D (new_AGEMA_signal_5502), .Q (new_AGEMA_signal_5503) ) ;
    buf_clk new_AGEMA_reg_buffer_2739 ( .C (CLK), .D (new_AGEMA_signal_5506), .Q (new_AGEMA_signal_5507) ) ;
    buf_clk new_AGEMA_reg_buffer_2743 ( .C (CLK), .D (new_AGEMA_signal_5510), .Q (new_AGEMA_signal_5511) ) ;
    buf_clk new_AGEMA_reg_buffer_2747 ( .C (CLK), .D (new_AGEMA_signal_5514), .Q (new_AGEMA_signal_5515) ) ;
    buf_clk new_AGEMA_reg_buffer_2751 ( .C (CLK), .D (new_AGEMA_signal_5518), .Q (new_AGEMA_signal_5519) ) ;
    buf_clk new_AGEMA_reg_buffer_2755 ( .C (CLK), .D (new_AGEMA_signal_5522), .Q (new_AGEMA_signal_5523) ) ;
    buf_clk new_AGEMA_reg_buffer_2759 ( .C (CLK), .D (new_AGEMA_signal_5526), .Q (new_AGEMA_signal_5527) ) ;
    buf_clk new_AGEMA_reg_buffer_2763 ( .C (CLK), .D (new_AGEMA_signal_5530), .Q (new_AGEMA_signal_5531) ) ;
    buf_clk new_AGEMA_reg_buffer_2767 ( .C (CLK), .D (new_AGEMA_signal_5534), .Q (new_AGEMA_signal_5535) ) ;
    buf_clk new_AGEMA_reg_buffer_2771 ( .C (CLK), .D (new_AGEMA_signal_5538), .Q (new_AGEMA_signal_5539) ) ;
    buf_clk new_AGEMA_reg_buffer_2775 ( .C (CLK), .D (new_AGEMA_signal_5542), .Q (new_AGEMA_signal_5543) ) ;
    buf_clk new_AGEMA_reg_buffer_2779 ( .C (CLK), .D (new_AGEMA_signal_5546), .Q (new_AGEMA_signal_5547) ) ;
    buf_clk new_AGEMA_reg_buffer_2783 ( .C (CLK), .D (new_AGEMA_signal_5550), .Q (new_AGEMA_signal_5551) ) ;
    buf_clk new_AGEMA_reg_buffer_2787 ( .C (CLK), .D (new_AGEMA_signal_5554), .Q (new_AGEMA_signal_5555) ) ;
    buf_clk new_AGEMA_reg_buffer_2791 ( .C (CLK), .D (new_AGEMA_signal_5558), .Q (new_AGEMA_signal_5559) ) ;
    buf_clk new_AGEMA_reg_buffer_2795 ( .C (CLK), .D (new_AGEMA_signal_5562), .Q (new_AGEMA_signal_5563) ) ;
    buf_clk new_AGEMA_reg_buffer_2799 ( .C (CLK), .D (new_AGEMA_signal_5566), .Q (new_AGEMA_signal_5567) ) ;
    buf_clk new_AGEMA_reg_buffer_2803 ( .C (CLK), .D (new_AGEMA_signal_5570), .Q (new_AGEMA_signal_5571) ) ;
    buf_clk new_AGEMA_reg_buffer_2807 ( .C (CLK), .D (new_AGEMA_signal_5574), .Q (new_AGEMA_signal_5575) ) ;
    buf_clk new_AGEMA_reg_buffer_2811 ( .C (CLK), .D (new_AGEMA_signal_5578), .Q (new_AGEMA_signal_5579) ) ;
    buf_clk new_AGEMA_reg_buffer_2815 ( .C (CLK), .D (new_AGEMA_signal_5582), .Q (new_AGEMA_signal_5583) ) ;
    buf_clk new_AGEMA_reg_buffer_2819 ( .C (CLK), .D (new_AGEMA_signal_5586), .Q (new_AGEMA_signal_5587) ) ;
    buf_clk new_AGEMA_reg_buffer_2823 ( .C (CLK), .D (new_AGEMA_signal_5590), .Q (new_AGEMA_signal_5591) ) ;
    buf_clk new_AGEMA_reg_buffer_2827 ( .C (CLK), .D (new_AGEMA_signal_5594), .Q (new_AGEMA_signal_5595) ) ;
    buf_clk new_AGEMA_reg_buffer_2831 ( .C (CLK), .D (new_AGEMA_signal_5598), .Q (new_AGEMA_signal_5599) ) ;
    buf_clk new_AGEMA_reg_buffer_2835 ( .C (CLK), .D (new_AGEMA_signal_5602), .Q (new_AGEMA_signal_5603) ) ;
    buf_clk new_AGEMA_reg_buffer_2839 ( .C (CLK), .D (new_AGEMA_signal_5606), .Q (new_AGEMA_signal_5607) ) ;
    buf_clk new_AGEMA_reg_buffer_2843 ( .C (CLK), .D (new_AGEMA_signal_5610), .Q (new_AGEMA_signal_5611) ) ;
    buf_clk new_AGEMA_reg_buffer_2847 ( .C (CLK), .D (new_AGEMA_signal_5614), .Q (new_AGEMA_signal_5615) ) ;
    buf_clk new_AGEMA_reg_buffer_2851 ( .C (CLK), .D (new_AGEMA_signal_5618), .Q (new_AGEMA_signal_5619) ) ;
    buf_clk new_AGEMA_reg_buffer_2855 ( .C (CLK), .D (new_AGEMA_signal_5622), .Q (new_AGEMA_signal_5623) ) ;
    buf_clk new_AGEMA_reg_buffer_2859 ( .C (CLK), .D (new_AGEMA_signal_5626), .Q (new_AGEMA_signal_5627) ) ;
    buf_clk new_AGEMA_reg_buffer_2863 ( .C (CLK), .D (new_AGEMA_signal_5630), .Q (new_AGEMA_signal_5631) ) ;
    buf_clk new_AGEMA_reg_buffer_2867 ( .C (CLK), .D (new_AGEMA_signal_5634), .Q (new_AGEMA_signal_5635) ) ;
    buf_clk new_AGEMA_reg_buffer_2871 ( .C (CLK), .D (new_AGEMA_signal_5638), .Q (new_AGEMA_signal_5639) ) ;
    buf_clk new_AGEMA_reg_buffer_2875 ( .C (CLK), .D (new_AGEMA_signal_5642), .Q (new_AGEMA_signal_5643) ) ;
    buf_clk new_AGEMA_reg_buffer_2879 ( .C (CLK), .D (new_AGEMA_signal_5646), .Q (new_AGEMA_signal_5647) ) ;
    buf_clk new_AGEMA_reg_buffer_2883 ( .C (CLK), .D (new_AGEMA_signal_5650), .Q (new_AGEMA_signal_5651) ) ;
    buf_clk new_AGEMA_reg_buffer_2887 ( .C (CLK), .D (new_AGEMA_signal_5654), .Q (new_AGEMA_signal_5655) ) ;
    buf_clk new_AGEMA_reg_buffer_2891 ( .C (CLK), .D (new_AGEMA_signal_5658), .Q (new_AGEMA_signal_5659) ) ;
    buf_clk new_AGEMA_reg_buffer_2895 ( .C (CLK), .D (new_AGEMA_signal_5662), .Q (new_AGEMA_signal_5663) ) ;
    buf_clk new_AGEMA_reg_buffer_2899 ( .C (CLK), .D (new_AGEMA_signal_5666), .Q (new_AGEMA_signal_5667) ) ;
    buf_clk new_AGEMA_reg_buffer_2903 ( .C (CLK), .D (new_AGEMA_signal_5670), .Q (new_AGEMA_signal_5671) ) ;
    buf_clk new_AGEMA_reg_buffer_2907 ( .C (CLK), .D (new_AGEMA_signal_5674), .Q (new_AGEMA_signal_5675) ) ;
    buf_clk new_AGEMA_reg_buffer_2911 ( .C (CLK), .D (new_AGEMA_signal_5678), .Q (new_AGEMA_signal_5679) ) ;
    buf_clk new_AGEMA_reg_buffer_2915 ( .C (CLK), .D (new_AGEMA_signal_5682), .Q (new_AGEMA_signal_5683) ) ;
    buf_clk new_AGEMA_reg_buffer_2919 ( .C (CLK), .D (new_AGEMA_signal_5686), .Q (new_AGEMA_signal_5687) ) ;
    buf_clk new_AGEMA_reg_buffer_2923 ( .C (CLK), .D (new_AGEMA_signal_5690), .Q (new_AGEMA_signal_5691) ) ;
    buf_clk new_AGEMA_reg_buffer_2927 ( .C (CLK), .D (new_AGEMA_signal_5694), .Q (new_AGEMA_signal_5695) ) ;
    buf_clk new_AGEMA_reg_buffer_2931 ( .C (CLK), .D (new_AGEMA_signal_5698), .Q (new_AGEMA_signal_5699) ) ;
    buf_clk new_AGEMA_reg_buffer_2935 ( .C (CLK), .D (new_AGEMA_signal_5702), .Q (new_AGEMA_signal_5703) ) ;
    buf_clk new_AGEMA_reg_buffer_2939 ( .C (CLK), .D (new_AGEMA_signal_5706), .Q (new_AGEMA_signal_5707) ) ;
    buf_clk new_AGEMA_reg_buffer_2943 ( .C (CLK), .D (new_AGEMA_signal_5710), .Q (new_AGEMA_signal_5711) ) ;
    buf_clk new_AGEMA_reg_buffer_2947 ( .C (CLK), .D (new_AGEMA_signal_5714), .Q (new_AGEMA_signal_5715) ) ;
    buf_clk new_AGEMA_reg_buffer_2951 ( .C (CLK), .D (new_AGEMA_signal_5718), .Q (new_AGEMA_signal_5719) ) ;
    buf_clk new_AGEMA_reg_buffer_2955 ( .C (CLK), .D (new_AGEMA_signal_5722), .Q (new_AGEMA_signal_5723) ) ;
    buf_clk new_AGEMA_reg_buffer_2959 ( .C (CLK), .D (new_AGEMA_signal_5726), .Q (new_AGEMA_signal_5727) ) ;
    buf_clk new_AGEMA_reg_buffer_2963 ( .C (CLK), .D (new_AGEMA_signal_5730), .Q (new_AGEMA_signal_5731) ) ;
    buf_clk new_AGEMA_reg_buffer_2967 ( .C (CLK), .D (new_AGEMA_signal_5734), .Q (new_AGEMA_signal_5735) ) ;
    buf_clk new_AGEMA_reg_buffer_2971 ( .C (CLK), .D (new_AGEMA_signal_5738), .Q (new_AGEMA_signal_5739) ) ;
    buf_clk new_AGEMA_reg_buffer_2985 ( .C (CLK), .D (new_AGEMA_signal_5752), .Q (new_AGEMA_signal_5753) ) ;
    buf_clk new_AGEMA_reg_buffer_2987 ( .C (CLK), .D (new_AGEMA_signal_5754), .Q (new_AGEMA_signal_5755) ) ;
    buf_clk new_AGEMA_reg_buffer_2989 ( .C (CLK), .D (new_AGEMA_signal_5756), .Q (new_AGEMA_signal_5757) ) ;
    buf_clk new_AGEMA_reg_buffer_2993 ( .C (CLK), .D (new_AGEMA_signal_5760), .Q (new_AGEMA_signal_5761) ) ;
    buf_clk new_AGEMA_reg_buffer_2997 ( .C (CLK), .D (new_AGEMA_signal_5764), .Q (new_AGEMA_signal_5765) ) ;
    buf_clk new_AGEMA_reg_buffer_3001 ( .C (CLK), .D (new_AGEMA_signal_5768), .Q (new_AGEMA_signal_5769) ) ;
    buf_clk new_AGEMA_reg_buffer_3005 ( .C (CLK), .D (new_AGEMA_signal_5772), .Q (new_AGEMA_signal_5773) ) ;
    buf_clk new_AGEMA_reg_buffer_3009 ( .C (CLK), .D (new_AGEMA_signal_5776), .Q (new_AGEMA_signal_5777) ) ;
    buf_clk new_AGEMA_reg_buffer_3013 ( .C (CLK), .D (new_AGEMA_signal_5780), .Q (new_AGEMA_signal_5781) ) ;
    buf_clk new_AGEMA_reg_buffer_3015 ( .C (CLK), .D (new_AGEMA_signal_5782), .Q (new_AGEMA_signal_5783) ) ;
    buf_clk new_AGEMA_reg_buffer_3017 ( .C (CLK), .D (new_AGEMA_signal_5784), .Q (new_AGEMA_signal_5785) ) ;
    buf_clk new_AGEMA_reg_buffer_3019 ( .C (CLK), .D (new_AGEMA_signal_5786), .Q (new_AGEMA_signal_5787) ) ;
    buf_clk new_AGEMA_reg_buffer_3033 ( .C (CLK), .D (new_AGEMA_signal_5800), .Q (new_AGEMA_signal_5801) ) ;
    buf_clk new_AGEMA_reg_buffer_3035 ( .C (CLK), .D (new_AGEMA_signal_5802), .Q (new_AGEMA_signal_5803) ) ;
    buf_clk new_AGEMA_reg_buffer_3037 ( .C (CLK), .D (new_AGEMA_signal_5804), .Q (new_AGEMA_signal_5805) ) ;
    buf_clk new_AGEMA_reg_buffer_3041 ( .C (CLK), .D (new_AGEMA_signal_5808), .Q (new_AGEMA_signal_5809) ) ;
    buf_clk new_AGEMA_reg_buffer_3045 ( .C (CLK), .D (new_AGEMA_signal_5812), .Q (new_AGEMA_signal_5813) ) ;
    buf_clk new_AGEMA_reg_buffer_3049 ( .C (CLK), .D (new_AGEMA_signal_5816), .Q (new_AGEMA_signal_5817) ) ;
    buf_clk new_AGEMA_reg_buffer_3053 ( .C (CLK), .D (new_AGEMA_signal_5820), .Q (new_AGEMA_signal_5821) ) ;
    buf_clk new_AGEMA_reg_buffer_3057 ( .C (CLK), .D (new_AGEMA_signal_5824), .Q (new_AGEMA_signal_5825) ) ;
    buf_clk new_AGEMA_reg_buffer_3061 ( .C (CLK), .D (new_AGEMA_signal_5828), .Q (new_AGEMA_signal_5829) ) ;
    buf_clk new_AGEMA_reg_buffer_3063 ( .C (CLK), .D (new_AGEMA_signal_5830), .Q (new_AGEMA_signal_5831) ) ;
    buf_clk new_AGEMA_reg_buffer_3065 ( .C (CLK), .D (new_AGEMA_signal_5832), .Q (new_AGEMA_signal_5833) ) ;
    buf_clk new_AGEMA_reg_buffer_3067 ( .C (CLK), .D (new_AGEMA_signal_5834), .Q (new_AGEMA_signal_5835) ) ;
    buf_clk new_AGEMA_reg_buffer_3081 ( .C (CLK), .D (new_AGEMA_signal_5848), .Q (new_AGEMA_signal_5849) ) ;
    buf_clk new_AGEMA_reg_buffer_3083 ( .C (CLK), .D (new_AGEMA_signal_5850), .Q (new_AGEMA_signal_5851) ) ;
    buf_clk new_AGEMA_reg_buffer_3085 ( .C (CLK), .D (new_AGEMA_signal_5852), .Q (new_AGEMA_signal_5853) ) ;
    buf_clk new_AGEMA_reg_buffer_3089 ( .C (CLK), .D (new_AGEMA_signal_5856), .Q (new_AGEMA_signal_5857) ) ;
    buf_clk new_AGEMA_reg_buffer_3093 ( .C (CLK), .D (new_AGEMA_signal_5860), .Q (new_AGEMA_signal_5861) ) ;
    buf_clk new_AGEMA_reg_buffer_3097 ( .C (CLK), .D (new_AGEMA_signal_5864), .Q (new_AGEMA_signal_5865) ) ;
    buf_clk new_AGEMA_reg_buffer_3099 ( .C (CLK), .D (new_AGEMA_signal_5866), .Q (new_AGEMA_signal_5867) ) ;
    buf_clk new_AGEMA_reg_buffer_3101 ( .C (CLK), .D (new_AGEMA_signal_5868), .Q (new_AGEMA_signal_5869) ) ;
    buf_clk new_AGEMA_reg_buffer_3103 ( .C (CLK), .D (new_AGEMA_signal_5870), .Q (new_AGEMA_signal_5871) ) ;
    buf_clk new_AGEMA_reg_buffer_3117 ( .C (CLK), .D (new_AGEMA_signal_5884), .Q (new_AGEMA_signal_5885) ) ;
    buf_clk new_AGEMA_reg_buffer_3119 ( .C (CLK), .D (new_AGEMA_signal_5886), .Q (new_AGEMA_signal_5887) ) ;
    buf_clk new_AGEMA_reg_buffer_3121 ( .C (CLK), .D (new_AGEMA_signal_5888), .Q (new_AGEMA_signal_5889) ) ;
    buf_clk new_AGEMA_reg_buffer_3125 ( .C (CLK), .D (new_AGEMA_signal_5892), .Q (new_AGEMA_signal_5893) ) ;
    buf_clk new_AGEMA_reg_buffer_3129 ( .C (CLK), .D (new_AGEMA_signal_5896), .Q (new_AGEMA_signal_5897) ) ;
    buf_clk new_AGEMA_reg_buffer_3133 ( .C (CLK), .D (new_AGEMA_signal_5900), .Q (new_AGEMA_signal_5901) ) ;
    buf_clk new_AGEMA_reg_buffer_3135 ( .C (CLK), .D (new_AGEMA_signal_5902), .Q (new_AGEMA_signal_5903) ) ;
    buf_clk new_AGEMA_reg_buffer_3137 ( .C (CLK), .D (new_AGEMA_signal_5904), .Q (new_AGEMA_signal_5905) ) ;
    buf_clk new_AGEMA_reg_buffer_3139 ( .C (CLK), .D (new_AGEMA_signal_5906), .Q (new_AGEMA_signal_5907) ) ;
    buf_clk new_AGEMA_reg_buffer_3153 ( .C (CLK), .D (new_AGEMA_signal_5920), .Q (new_AGEMA_signal_5921) ) ;
    buf_clk new_AGEMA_reg_buffer_3155 ( .C (CLK), .D (new_AGEMA_signal_5922), .Q (new_AGEMA_signal_5923) ) ;
    buf_clk new_AGEMA_reg_buffer_3157 ( .C (CLK), .D (new_AGEMA_signal_5924), .Q (new_AGEMA_signal_5925) ) ;
    buf_clk new_AGEMA_reg_buffer_3161 ( .C (CLK), .D (new_AGEMA_signal_5928), .Q (new_AGEMA_signal_5929) ) ;
    buf_clk new_AGEMA_reg_buffer_3165 ( .C (CLK), .D (new_AGEMA_signal_5932), .Q (new_AGEMA_signal_5933) ) ;
    buf_clk new_AGEMA_reg_buffer_3169 ( .C (CLK), .D (new_AGEMA_signal_5936), .Q (new_AGEMA_signal_5937) ) ;
    buf_clk new_AGEMA_reg_buffer_3173 ( .C (CLK), .D (new_AGEMA_signal_5940), .Q (new_AGEMA_signal_5941) ) ;
    buf_clk new_AGEMA_reg_buffer_3177 ( .C (CLK), .D (new_AGEMA_signal_5944), .Q (new_AGEMA_signal_5945) ) ;
    buf_clk new_AGEMA_reg_buffer_3181 ( .C (CLK), .D (new_AGEMA_signal_5948), .Q (new_AGEMA_signal_5949) ) ;
    buf_clk new_AGEMA_reg_buffer_3183 ( .C (CLK), .D (new_AGEMA_signal_5950), .Q (new_AGEMA_signal_5951) ) ;
    buf_clk new_AGEMA_reg_buffer_3185 ( .C (CLK), .D (new_AGEMA_signal_5952), .Q (new_AGEMA_signal_5953) ) ;
    buf_clk new_AGEMA_reg_buffer_3187 ( .C (CLK), .D (new_AGEMA_signal_5954), .Q (new_AGEMA_signal_5955) ) ;
    buf_clk new_AGEMA_reg_buffer_3201 ( .C (CLK), .D (new_AGEMA_signal_5968), .Q (new_AGEMA_signal_5969) ) ;
    buf_clk new_AGEMA_reg_buffer_3203 ( .C (CLK), .D (new_AGEMA_signal_5970), .Q (new_AGEMA_signal_5971) ) ;
    buf_clk new_AGEMA_reg_buffer_3205 ( .C (CLK), .D (new_AGEMA_signal_5972), .Q (new_AGEMA_signal_5973) ) ;
    buf_clk new_AGEMA_reg_buffer_3209 ( .C (CLK), .D (new_AGEMA_signal_5976), .Q (new_AGEMA_signal_5977) ) ;
    buf_clk new_AGEMA_reg_buffer_3213 ( .C (CLK), .D (new_AGEMA_signal_5980), .Q (new_AGEMA_signal_5981) ) ;
    buf_clk new_AGEMA_reg_buffer_3217 ( .C (CLK), .D (new_AGEMA_signal_5984), .Q (new_AGEMA_signal_5985) ) ;
    buf_clk new_AGEMA_reg_buffer_3221 ( .C (CLK), .D (new_AGEMA_signal_5988), .Q (new_AGEMA_signal_5989) ) ;
    buf_clk new_AGEMA_reg_buffer_3225 ( .C (CLK), .D (new_AGEMA_signal_5992), .Q (new_AGEMA_signal_5993) ) ;
    buf_clk new_AGEMA_reg_buffer_3229 ( .C (CLK), .D (new_AGEMA_signal_5996), .Q (new_AGEMA_signal_5997) ) ;
    buf_clk new_AGEMA_reg_buffer_3231 ( .C (CLK), .D (new_AGEMA_signal_5998), .Q (new_AGEMA_signal_5999) ) ;
    buf_clk new_AGEMA_reg_buffer_3233 ( .C (CLK), .D (new_AGEMA_signal_6000), .Q (new_AGEMA_signal_6001) ) ;
    buf_clk new_AGEMA_reg_buffer_3235 ( .C (CLK), .D (new_AGEMA_signal_6002), .Q (new_AGEMA_signal_6003) ) ;
    buf_clk new_AGEMA_reg_buffer_3249 ( .C (CLK), .D (new_AGEMA_signal_6016), .Q (new_AGEMA_signal_6017) ) ;
    buf_clk new_AGEMA_reg_buffer_3251 ( .C (CLK), .D (new_AGEMA_signal_6018), .Q (new_AGEMA_signal_6019) ) ;
    buf_clk new_AGEMA_reg_buffer_3253 ( .C (CLK), .D (new_AGEMA_signal_6020), .Q (new_AGEMA_signal_6021) ) ;
    buf_clk new_AGEMA_reg_buffer_3257 ( .C (CLK), .D (new_AGEMA_signal_6024), .Q (new_AGEMA_signal_6025) ) ;
    buf_clk new_AGEMA_reg_buffer_3261 ( .C (CLK), .D (new_AGEMA_signal_6028), .Q (new_AGEMA_signal_6029) ) ;
    buf_clk new_AGEMA_reg_buffer_3265 ( .C (CLK), .D (new_AGEMA_signal_6032), .Q (new_AGEMA_signal_6033) ) ;
    buf_clk new_AGEMA_reg_buffer_3267 ( .C (CLK), .D (new_AGEMA_signal_6034), .Q (new_AGEMA_signal_6035) ) ;
    buf_clk new_AGEMA_reg_buffer_3269 ( .C (CLK), .D (new_AGEMA_signal_6036), .Q (new_AGEMA_signal_6037) ) ;
    buf_clk new_AGEMA_reg_buffer_3271 ( .C (CLK), .D (new_AGEMA_signal_6038), .Q (new_AGEMA_signal_6039) ) ;
    buf_clk new_AGEMA_reg_buffer_3285 ( .C (CLK), .D (new_AGEMA_signal_6052), .Q (new_AGEMA_signal_6053) ) ;
    buf_clk new_AGEMA_reg_buffer_3287 ( .C (CLK), .D (new_AGEMA_signal_6054), .Q (new_AGEMA_signal_6055) ) ;
    buf_clk new_AGEMA_reg_buffer_3289 ( .C (CLK), .D (new_AGEMA_signal_6056), .Q (new_AGEMA_signal_6057) ) ;
    buf_clk new_AGEMA_reg_buffer_3293 ( .C (CLK), .D (new_AGEMA_signal_6060), .Q (new_AGEMA_signal_6061) ) ;
    buf_clk new_AGEMA_reg_buffer_3297 ( .C (CLK), .D (new_AGEMA_signal_6064), .Q (new_AGEMA_signal_6065) ) ;
    buf_clk new_AGEMA_reg_buffer_3301 ( .C (CLK), .D (new_AGEMA_signal_6068), .Q (new_AGEMA_signal_6069) ) ;
    buf_clk new_AGEMA_reg_buffer_3303 ( .C (CLK), .D (new_AGEMA_signal_6070), .Q (new_AGEMA_signal_6071) ) ;
    buf_clk new_AGEMA_reg_buffer_3305 ( .C (CLK), .D (new_AGEMA_signal_6072), .Q (new_AGEMA_signal_6073) ) ;
    buf_clk new_AGEMA_reg_buffer_3307 ( .C (CLK), .D (new_AGEMA_signal_6074), .Q (new_AGEMA_signal_6075) ) ;
    buf_clk new_AGEMA_reg_buffer_3321 ( .C (CLK), .D (new_AGEMA_signal_6088), .Q (new_AGEMA_signal_6089) ) ;
    buf_clk new_AGEMA_reg_buffer_3323 ( .C (CLK), .D (new_AGEMA_signal_6090), .Q (new_AGEMA_signal_6091) ) ;
    buf_clk new_AGEMA_reg_buffer_3325 ( .C (CLK), .D (new_AGEMA_signal_6092), .Q (new_AGEMA_signal_6093) ) ;
    buf_clk new_AGEMA_reg_buffer_3329 ( .C (CLK), .D (new_AGEMA_signal_6096), .Q (new_AGEMA_signal_6097) ) ;
    buf_clk new_AGEMA_reg_buffer_3333 ( .C (CLK), .D (new_AGEMA_signal_6100), .Q (new_AGEMA_signal_6101) ) ;
    buf_clk new_AGEMA_reg_buffer_3337 ( .C (CLK), .D (new_AGEMA_signal_6104), .Q (new_AGEMA_signal_6105) ) ;
    buf_clk new_AGEMA_reg_buffer_3341 ( .C (CLK), .D (new_AGEMA_signal_6108), .Q (new_AGEMA_signal_6109) ) ;
    buf_clk new_AGEMA_reg_buffer_3345 ( .C (CLK), .D (new_AGEMA_signal_6112), .Q (new_AGEMA_signal_6113) ) ;
    buf_clk new_AGEMA_reg_buffer_3349 ( .C (CLK), .D (new_AGEMA_signal_6116), .Q (new_AGEMA_signal_6117) ) ;
    buf_clk new_AGEMA_reg_buffer_3351 ( .C (CLK), .D (new_AGEMA_signal_6118), .Q (new_AGEMA_signal_6119) ) ;
    buf_clk new_AGEMA_reg_buffer_3353 ( .C (CLK), .D (new_AGEMA_signal_6120), .Q (new_AGEMA_signal_6121) ) ;
    buf_clk new_AGEMA_reg_buffer_3355 ( .C (CLK), .D (new_AGEMA_signal_6122), .Q (new_AGEMA_signal_6123) ) ;
    buf_clk new_AGEMA_reg_buffer_3369 ( .C (CLK), .D (new_AGEMA_signal_6136), .Q (new_AGEMA_signal_6137) ) ;
    buf_clk new_AGEMA_reg_buffer_3371 ( .C (CLK), .D (new_AGEMA_signal_6138), .Q (new_AGEMA_signal_6139) ) ;
    buf_clk new_AGEMA_reg_buffer_3373 ( .C (CLK), .D (new_AGEMA_signal_6140), .Q (new_AGEMA_signal_6141) ) ;
    buf_clk new_AGEMA_reg_buffer_3377 ( .C (CLK), .D (new_AGEMA_signal_6144), .Q (new_AGEMA_signal_6145) ) ;
    buf_clk new_AGEMA_reg_buffer_3381 ( .C (CLK), .D (new_AGEMA_signal_6148), .Q (new_AGEMA_signal_6149) ) ;
    buf_clk new_AGEMA_reg_buffer_3385 ( .C (CLK), .D (new_AGEMA_signal_6152), .Q (new_AGEMA_signal_6153) ) ;
    buf_clk new_AGEMA_reg_buffer_3389 ( .C (CLK), .D (new_AGEMA_signal_6156), .Q (new_AGEMA_signal_6157) ) ;
    buf_clk new_AGEMA_reg_buffer_3393 ( .C (CLK), .D (new_AGEMA_signal_6160), .Q (new_AGEMA_signal_6161) ) ;
    buf_clk new_AGEMA_reg_buffer_3397 ( .C (CLK), .D (new_AGEMA_signal_6164), .Q (new_AGEMA_signal_6165) ) ;
    buf_clk new_AGEMA_reg_buffer_3399 ( .C (CLK), .D (new_AGEMA_signal_6166), .Q (new_AGEMA_signal_6167) ) ;
    buf_clk new_AGEMA_reg_buffer_3401 ( .C (CLK), .D (new_AGEMA_signal_6168), .Q (new_AGEMA_signal_6169) ) ;
    buf_clk new_AGEMA_reg_buffer_3403 ( .C (CLK), .D (new_AGEMA_signal_6170), .Q (new_AGEMA_signal_6171) ) ;
    buf_clk new_AGEMA_reg_buffer_3417 ( .C (CLK), .D (new_AGEMA_signal_6184), .Q (new_AGEMA_signal_6185) ) ;
    buf_clk new_AGEMA_reg_buffer_3419 ( .C (CLK), .D (new_AGEMA_signal_6186), .Q (new_AGEMA_signal_6187) ) ;
    buf_clk new_AGEMA_reg_buffer_3421 ( .C (CLK), .D (new_AGEMA_signal_6188), .Q (new_AGEMA_signal_6189) ) ;
    buf_clk new_AGEMA_reg_buffer_3425 ( .C (CLK), .D (new_AGEMA_signal_6192), .Q (new_AGEMA_signal_6193) ) ;
    buf_clk new_AGEMA_reg_buffer_3429 ( .C (CLK), .D (new_AGEMA_signal_6196), .Q (new_AGEMA_signal_6197) ) ;
    buf_clk new_AGEMA_reg_buffer_3433 ( .C (CLK), .D (new_AGEMA_signal_6200), .Q (new_AGEMA_signal_6201) ) ;
    buf_clk new_AGEMA_reg_buffer_3435 ( .C (CLK), .D (new_AGEMA_signal_6202), .Q (new_AGEMA_signal_6203) ) ;
    buf_clk new_AGEMA_reg_buffer_3437 ( .C (CLK), .D (new_AGEMA_signal_6204), .Q (new_AGEMA_signal_6205) ) ;
    buf_clk new_AGEMA_reg_buffer_3439 ( .C (CLK), .D (new_AGEMA_signal_6206), .Q (new_AGEMA_signal_6207) ) ;
    buf_clk new_AGEMA_reg_buffer_3453 ( .C (CLK), .D (new_AGEMA_signal_6220), .Q (new_AGEMA_signal_6221) ) ;
    buf_clk new_AGEMA_reg_buffer_3455 ( .C (CLK), .D (new_AGEMA_signal_6222), .Q (new_AGEMA_signal_6223) ) ;
    buf_clk new_AGEMA_reg_buffer_3457 ( .C (CLK), .D (new_AGEMA_signal_6224), .Q (new_AGEMA_signal_6225) ) ;
    buf_clk new_AGEMA_reg_buffer_3461 ( .C (CLK), .D (new_AGEMA_signal_6228), .Q (new_AGEMA_signal_6229) ) ;
    buf_clk new_AGEMA_reg_buffer_3465 ( .C (CLK), .D (new_AGEMA_signal_6232), .Q (new_AGEMA_signal_6233) ) ;
    buf_clk new_AGEMA_reg_buffer_3469 ( .C (CLK), .D (new_AGEMA_signal_6236), .Q (new_AGEMA_signal_6237) ) ;
    buf_clk new_AGEMA_reg_buffer_3471 ( .C (CLK), .D (new_AGEMA_signal_6238), .Q (new_AGEMA_signal_6239) ) ;
    buf_clk new_AGEMA_reg_buffer_3473 ( .C (CLK), .D (new_AGEMA_signal_6240), .Q (new_AGEMA_signal_6241) ) ;
    buf_clk new_AGEMA_reg_buffer_3475 ( .C (CLK), .D (new_AGEMA_signal_6242), .Q (new_AGEMA_signal_6243) ) ;
    buf_clk new_AGEMA_reg_buffer_3489 ( .C (CLK), .D (new_AGEMA_signal_6256), .Q (new_AGEMA_signal_6257) ) ;
    buf_clk new_AGEMA_reg_buffer_3491 ( .C (CLK), .D (new_AGEMA_signal_6258), .Q (new_AGEMA_signal_6259) ) ;
    buf_clk new_AGEMA_reg_buffer_3493 ( .C (CLK), .D (new_AGEMA_signal_6260), .Q (new_AGEMA_signal_6261) ) ;
    buf_clk new_AGEMA_reg_buffer_3497 ( .C (CLK), .D (new_AGEMA_signal_6264), .Q (new_AGEMA_signal_6265) ) ;
    buf_clk new_AGEMA_reg_buffer_3501 ( .C (CLK), .D (new_AGEMA_signal_6268), .Q (new_AGEMA_signal_6269) ) ;
    buf_clk new_AGEMA_reg_buffer_3505 ( .C (CLK), .D (new_AGEMA_signal_6272), .Q (new_AGEMA_signal_6273) ) ;
    buf_clk new_AGEMA_reg_buffer_3509 ( .C (CLK), .D (new_AGEMA_signal_6276), .Q (new_AGEMA_signal_6277) ) ;
    buf_clk new_AGEMA_reg_buffer_3513 ( .C (CLK), .D (new_AGEMA_signal_6280), .Q (new_AGEMA_signal_6281) ) ;
    buf_clk new_AGEMA_reg_buffer_3517 ( .C (CLK), .D (new_AGEMA_signal_6284), .Q (new_AGEMA_signal_6285) ) ;
    buf_clk new_AGEMA_reg_buffer_3519 ( .C (CLK), .D (new_AGEMA_signal_6286), .Q (new_AGEMA_signal_6287) ) ;
    buf_clk new_AGEMA_reg_buffer_3521 ( .C (CLK), .D (new_AGEMA_signal_6288), .Q (new_AGEMA_signal_6289) ) ;
    buf_clk new_AGEMA_reg_buffer_3523 ( .C (CLK), .D (new_AGEMA_signal_6290), .Q (new_AGEMA_signal_6291) ) ;
    buf_clk new_AGEMA_reg_buffer_3537 ( .C (CLK), .D (new_AGEMA_signal_6304), .Q (new_AGEMA_signal_6305) ) ;
    buf_clk new_AGEMA_reg_buffer_3539 ( .C (CLK), .D (new_AGEMA_signal_6306), .Q (new_AGEMA_signal_6307) ) ;
    buf_clk new_AGEMA_reg_buffer_3541 ( .C (CLK), .D (new_AGEMA_signal_6308), .Q (new_AGEMA_signal_6309) ) ;
    buf_clk new_AGEMA_reg_buffer_3545 ( .C (CLK), .D (new_AGEMA_signal_6312), .Q (new_AGEMA_signal_6313) ) ;
    buf_clk new_AGEMA_reg_buffer_3549 ( .C (CLK), .D (new_AGEMA_signal_6316), .Q (new_AGEMA_signal_6317) ) ;
    buf_clk new_AGEMA_reg_buffer_3553 ( .C (CLK), .D (new_AGEMA_signal_6320), .Q (new_AGEMA_signal_6321) ) ;
    buf_clk new_AGEMA_reg_buffer_3557 ( .C (CLK), .D (new_AGEMA_signal_6324), .Q (new_AGEMA_signal_6325) ) ;
    buf_clk new_AGEMA_reg_buffer_3561 ( .C (CLK), .D (new_AGEMA_signal_6328), .Q (new_AGEMA_signal_6329) ) ;
    buf_clk new_AGEMA_reg_buffer_3565 ( .C (CLK), .D (new_AGEMA_signal_6332), .Q (new_AGEMA_signal_6333) ) ;
    buf_clk new_AGEMA_reg_buffer_3567 ( .C (CLK), .D (new_AGEMA_signal_6334), .Q (new_AGEMA_signal_6335) ) ;
    buf_clk new_AGEMA_reg_buffer_3569 ( .C (CLK), .D (new_AGEMA_signal_6336), .Q (new_AGEMA_signal_6337) ) ;
    buf_clk new_AGEMA_reg_buffer_3571 ( .C (CLK), .D (new_AGEMA_signal_6338), .Q (new_AGEMA_signal_6339) ) ;
    buf_clk new_AGEMA_reg_buffer_3585 ( .C (CLK), .D (new_AGEMA_signal_6352), .Q (new_AGEMA_signal_6353) ) ;
    buf_clk new_AGEMA_reg_buffer_3587 ( .C (CLK), .D (new_AGEMA_signal_6354), .Q (new_AGEMA_signal_6355) ) ;
    buf_clk new_AGEMA_reg_buffer_3589 ( .C (CLK), .D (new_AGEMA_signal_6356), .Q (new_AGEMA_signal_6357) ) ;
    buf_clk new_AGEMA_reg_buffer_3593 ( .C (CLK), .D (new_AGEMA_signal_6360), .Q (new_AGEMA_signal_6361) ) ;
    buf_clk new_AGEMA_reg_buffer_3597 ( .C (CLK), .D (new_AGEMA_signal_6364), .Q (new_AGEMA_signal_6365) ) ;
    buf_clk new_AGEMA_reg_buffer_3601 ( .C (CLK), .D (new_AGEMA_signal_6368), .Q (new_AGEMA_signal_6369) ) ;
    buf_clk new_AGEMA_reg_buffer_3603 ( .C (CLK), .D (new_AGEMA_signal_6370), .Q (new_AGEMA_signal_6371) ) ;
    buf_clk new_AGEMA_reg_buffer_3605 ( .C (CLK), .D (new_AGEMA_signal_6372), .Q (new_AGEMA_signal_6373) ) ;
    buf_clk new_AGEMA_reg_buffer_3607 ( .C (CLK), .D (new_AGEMA_signal_6374), .Q (new_AGEMA_signal_6375) ) ;
    buf_clk new_AGEMA_reg_buffer_3621 ( .C (CLK), .D (new_AGEMA_signal_6388), .Q (new_AGEMA_signal_6389) ) ;
    buf_clk new_AGEMA_reg_buffer_3623 ( .C (CLK), .D (new_AGEMA_signal_6390), .Q (new_AGEMA_signal_6391) ) ;
    buf_clk new_AGEMA_reg_buffer_3625 ( .C (CLK), .D (new_AGEMA_signal_6392), .Q (new_AGEMA_signal_6393) ) ;
    buf_clk new_AGEMA_reg_buffer_3629 ( .C (CLK), .D (new_AGEMA_signal_6396), .Q (new_AGEMA_signal_6397) ) ;
    buf_clk new_AGEMA_reg_buffer_3633 ( .C (CLK), .D (new_AGEMA_signal_6400), .Q (new_AGEMA_signal_6401) ) ;
    buf_clk new_AGEMA_reg_buffer_3637 ( .C (CLK), .D (new_AGEMA_signal_6404), .Q (new_AGEMA_signal_6405) ) ;
    buf_clk new_AGEMA_reg_buffer_3639 ( .C (CLK), .D (new_AGEMA_signal_6406), .Q (new_AGEMA_signal_6407) ) ;
    buf_clk new_AGEMA_reg_buffer_3641 ( .C (CLK), .D (new_AGEMA_signal_6408), .Q (new_AGEMA_signal_6409) ) ;
    buf_clk new_AGEMA_reg_buffer_3643 ( .C (CLK), .D (new_AGEMA_signal_6410), .Q (new_AGEMA_signal_6411) ) ;
    buf_clk new_AGEMA_reg_buffer_3645 ( .C (CLK), .D (new_AGEMA_signal_6412), .Q (new_AGEMA_signal_6413) ) ;
    buf_clk new_AGEMA_reg_buffer_3647 ( .C (CLK), .D (new_AGEMA_signal_6414), .Q (new_AGEMA_signal_6415) ) ;
    buf_clk new_AGEMA_reg_buffer_3649 ( .C (CLK), .D (new_AGEMA_signal_6416), .Q (new_AGEMA_signal_6417) ) ;
    buf_clk new_AGEMA_reg_buffer_3651 ( .C (CLK), .D (new_AGEMA_signal_6418), .Q (new_AGEMA_signal_6419) ) ;
    buf_clk new_AGEMA_reg_buffer_3653 ( .C (CLK), .D (new_AGEMA_signal_6420), .Q (new_AGEMA_signal_6421) ) ;
    buf_clk new_AGEMA_reg_buffer_3655 ( .C (CLK), .D (new_AGEMA_signal_6422), .Q (new_AGEMA_signal_6423) ) ;
    buf_clk new_AGEMA_reg_buffer_3657 ( .C (CLK), .D (new_AGEMA_signal_6424), .Q (new_AGEMA_signal_6425) ) ;
    buf_clk new_AGEMA_reg_buffer_3659 ( .C (CLK), .D (new_AGEMA_signal_6426), .Q (new_AGEMA_signal_6427) ) ;
    buf_clk new_AGEMA_reg_buffer_3661 ( .C (CLK), .D (new_AGEMA_signal_6428), .Q (new_AGEMA_signal_6429) ) ;
    buf_clk new_AGEMA_reg_buffer_3663 ( .C (CLK), .D (new_AGEMA_signal_6430), .Q (new_AGEMA_signal_6431) ) ;
    buf_clk new_AGEMA_reg_buffer_3665 ( .C (CLK), .D (new_AGEMA_signal_6432), .Q (new_AGEMA_signal_6433) ) ;
    buf_clk new_AGEMA_reg_buffer_3667 ( .C (CLK), .D (new_AGEMA_signal_6434), .Q (new_AGEMA_signal_6435) ) ;
    buf_clk new_AGEMA_reg_buffer_3669 ( .C (CLK), .D (new_AGEMA_signal_6436), .Q (new_AGEMA_signal_6437) ) ;
    buf_clk new_AGEMA_reg_buffer_3671 ( .C (CLK), .D (new_AGEMA_signal_6438), .Q (new_AGEMA_signal_6439) ) ;
    buf_clk new_AGEMA_reg_buffer_3673 ( .C (CLK), .D (new_AGEMA_signal_6440), .Q (new_AGEMA_signal_6441) ) ;
    buf_clk new_AGEMA_reg_buffer_3675 ( .C (CLK), .D (new_AGEMA_signal_6442), .Q (new_AGEMA_signal_6443) ) ;
    buf_clk new_AGEMA_reg_buffer_3677 ( .C (CLK), .D (new_AGEMA_signal_6444), .Q (new_AGEMA_signal_6445) ) ;
    buf_clk new_AGEMA_reg_buffer_3679 ( .C (CLK), .D (new_AGEMA_signal_6446), .Q (new_AGEMA_signal_6447) ) ;
    buf_clk new_AGEMA_reg_buffer_3681 ( .C (CLK), .D (new_AGEMA_signal_6448), .Q (new_AGEMA_signal_6449) ) ;
    buf_clk new_AGEMA_reg_buffer_3683 ( .C (CLK), .D (new_AGEMA_signal_6450), .Q (new_AGEMA_signal_6451) ) ;
    buf_clk new_AGEMA_reg_buffer_3685 ( .C (CLK), .D (new_AGEMA_signal_6452), .Q (new_AGEMA_signal_6453) ) ;
    buf_clk new_AGEMA_reg_buffer_3687 ( .C (CLK), .D (new_AGEMA_signal_6454), .Q (new_AGEMA_signal_6455) ) ;
    buf_clk new_AGEMA_reg_buffer_3689 ( .C (CLK), .D (new_AGEMA_signal_6456), .Q (new_AGEMA_signal_6457) ) ;
    buf_clk new_AGEMA_reg_buffer_3691 ( .C (CLK), .D (new_AGEMA_signal_6458), .Q (new_AGEMA_signal_6459) ) ;
    buf_clk new_AGEMA_reg_buffer_3693 ( .C (CLK), .D (new_AGEMA_signal_6460), .Q (new_AGEMA_signal_6461) ) ;
    buf_clk new_AGEMA_reg_buffer_3695 ( .C (CLK), .D (new_AGEMA_signal_6462), .Q (new_AGEMA_signal_6463) ) ;
    buf_clk new_AGEMA_reg_buffer_3697 ( .C (CLK), .D (new_AGEMA_signal_6464), .Q (new_AGEMA_signal_6465) ) ;
    buf_clk new_AGEMA_reg_buffer_3699 ( .C (CLK), .D (new_AGEMA_signal_6466), .Q (new_AGEMA_signal_6467) ) ;
    buf_clk new_AGEMA_reg_buffer_3701 ( .C (CLK), .D (new_AGEMA_signal_6468), .Q (new_AGEMA_signal_6469) ) ;
    buf_clk new_AGEMA_reg_buffer_3703 ( .C (CLK), .D (new_AGEMA_signal_6470), .Q (new_AGEMA_signal_6471) ) ;
    buf_clk new_AGEMA_reg_buffer_3705 ( .C (CLK), .D (new_AGEMA_signal_6472), .Q (new_AGEMA_signal_6473) ) ;
    buf_clk new_AGEMA_reg_buffer_3707 ( .C (CLK), .D (new_AGEMA_signal_6474), .Q (new_AGEMA_signal_6475) ) ;
    buf_clk new_AGEMA_reg_buffer_3709 ( .C (CLK), .D (new_AGEMA_signal_6476), .Q (new_AGEMA_signal_6477) ) ;
    buf_clk new_AGEMA_reg_buffer_3711 ( .C (CLK), .D (new_AGEMA_signal_6478), .Q (new_AGEMA_signal_6479) ) ;
    buf_clk new_AGEMA_reg_buffer_3713 ( .C (CLK), .D (new_AGEMA_signal_6480), .Q (new_AGEMA_signal_6481) ) ;
    buf_clk new_AGEMA_reg_buffer_3715 ( .C (CLK), .D (new_AGEMA_signal_6482), .Q (new_AGEMA_signal_6483) ) ;
    buf_clk new_AGEMA_reg_buffer_3717 ( .C (CLK), .D (new_AGEMA_signal_6484), .Q (new_AGEMA_signal_6485) ) ;
    buf_clk new_AGEMA_reg_buffer_3719 ( .C (CLK), .D (new_AGEMA_signal_6486), .Q (new_AGEMA_signal_6487) ) ;
    buf_clk new_AGEMA_reg_buffer_3721 ( .C (CLK), .D (new_AGEMA_signal_6488), .Q (new_AGEMA_signal_6489) ) ;
    buf_clk new_AGEMA_reg_buffer_3723 ( .C (CLK), .D (new_AGEMA_signal_6490), .Q (new_AGEMA_signal_6491) ) ;
    buf_clk new_AGEMA_reg_buffer_3725 ( .C (CLK), .D (new_AGEMA_signal_6492), .Q (new_AGEMA_signal_6493) ) ;
    buf_clk new_AGEMA_reg_buffer_3727 ( .C (CLK), .D (new_AGEMA_signal_6494), .Q (new_AGEMA_signal_6495) ) ;
    buf_clk new_AGEMA_reg_buffer_3729 ( .C (CLK), .D (new_AGEMA_signal_6496), .Q (new_AGEMA_signal_6497) ) ;
    buf_clk new_AGEMA_reg_buffer_3731 ( .C (CLK), .D (new_AGEMA_signal_6498), .Q (new_AGEMA_signal_6499) ) ;
    buf_clk new_AGEMA_reg_buffer_3733 ( .C (CLK), .D (new_AGEMA_signal_6500), .Q (new_AGEMA_signal_6501) ) ;
    buf_clk new_AGEMA_reg_buffer_3735 ( .C (CLK), .D (new_AGEMA_signal_6502), .Q (new_AGEMA_signal_6503) ) ;
    buf_clk new_AGEMA_reg_buffer_3737 ( .C (CLK), .D (new_AGEMA_signal_6504), .Q (new_AGEMA_signal_6505) ) ;
    buf_clk new_AGEMA_reg_buffer_3739 ( .C (CLK), .D (new_AGEMA_signal_6506), .Q (new_AGEMA_signal_6507) ) ;
    buf_clk new_AGEMA_reg_buffer_3743 ( .C (CLK), .D (new_AGEMA_signal_6510), .Q (new_AGEMA_signal_6511) ) ;
    buf_clk new_AGEMA_reg_buffer_3747 ( .C (CLK), .D (new_AGEMA_signal_6514), .Q (new_AGEMA_signal_6515) ) ;
    buf_clk new_AGEMA_reg_buffer_3751 ( .C (CLK), .D (new_AGEMA_signal_6518), .Q (new_AGEMA_signal_6519) ) ;
    buf_clk new_AGEMA_reg_buffer_3755 ( .C (CLK), .D (new_AGEMA_signal_6522), .Q (new_AGEMA_signal_6523) ) ;
    buf_clk new_AGEMA_reg_buffer_3759 ( .C (CLK), .D (new_AGEMA_signal_6526), .Q (new_AGEMA_signal_6527) ) ;
    buf_clk new_AGEMA_reg_buffer_3763 ( .C (CLK), .D (new_AGEMA_signal_6530), .Q (new_AGEMA_signal_6531) ) ;
    buf_clk new_AGEMA_reg_buffer_3767 ( .C (CLK), .D (new_AGEMA_signal_6534), .Q (new_AGEMA_signal_6535) ) ;
    buf_clk new_AGEMA_reg_buffer_3771 ( .C (CLK), .D (new_AGEMA_signal_6538), .Q (new_AGEMA_signal_6539) ) ;
    buf_clk new_AGEMA_reg_buffer_3775 ( .C (CLK), .D (new_AGEMA_signal_6542), .Q (new_AGEMA_signal_6543) ) ;
    buf_clk new_AGEMA_reg_buffer_3779 ( .C (CLK), .D (new_AGEMA_signal_6546), .Q (new_AGEMA_signal_6547) ) ;
    buf_clk new_AGEMA_reg_buffer_3783 ( .C (CLK), .D (new_AGEMA_signal_6550), .Q (new_AGEMA_signal_6551) ) ;

    /* register cells */
    DFF_X1 LED_128_Instance_ks_reg_0__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_6511), .Q (LED_128_Instance_ks_reg_0__Q), .QN () ) ;
    DFF_X1 LED_128_Instance_ks_reg_1__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_6515), .Q (LED_128_Instance_n26), .QN () ) ;
    DFF_X1 LED_128_Instance_ks_reg_2__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_6519), .Q (LED_128_Instance_n25), .QN () ) ;
    DFF_X1 LED_128_Instance_ks_reg_3__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_6523), .Q (LED_128_Instance_n2), .QN () ) ;
    DFF_X1 LED_128_Instance_roundconstant_reg_0__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_6527), .Q (roundconstant[0]), .QN () ) ;
    DFF_X1 LED_128_Instance_roundconstant_reg_1__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_6531), .Q (roundconstant[1]), .QN () ) ;
    DFF_X1 LED_128_Instance_roundconstant_reg_2__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_6535), .Q (roundconstant[2]), .QN () ) ;
    DFF_X1 LED_128_Instance_roundconstant_reg_3__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_6539), .Q (roundconstant[3]), .QN () ) ;
    DFF_X1 LED_128_Instance_roundconstant_reg_4__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_6543), .Q (roundconstant[4]), .QN () ) ;
    DFF_X1 LED_128_Instance_roundconstant_reg_5__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_6547), .Q (roundconstant[5]), .QN () ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_0__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_state1[0]}), .Q ({OUT_ciphertext_s2[0], OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_1__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, LED_128_Instance_state1[1]}), .Q ({OUT_ciphertext_s2[1], OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_2__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, LED_128_Instance_state1[2]}), .Q ({OUT_ciphertext_s2[2], OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_3__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, LED_128_Instance_state1[3]}), .Q ({OUT_ciphertext_s2[3], OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_4__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, LED_128_Instance_state1[4]}), .Q ({OUT_ciphertext_s2[4], OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_5__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, LED_128_Instance_state1[5]}), .Q ({OUT_ciphertext_s2[5], OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_6__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, LED_128_Instance_state1[6]}), .Q ({OUT_ciphertext_s2[6], OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_7__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, LED_128_Instance_state1[7]}), .Q ({OUT_ciphertext_s2[7], OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_8__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, LED_128_Instance_state1[8]}), .Q ({OUT_ciphertext_s2[8], OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_9__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, LED_128_Instance_state1[9]}), .Q ({OUT_ciphertext_s2[9], OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_10__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, LED_128_Instance_state1[10]}), .Q ({OUT_ciphertext_s2[10], OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_11__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3151, new_AGEMA_signal_3150, LED_128_Instance_state1[11]}), .Q ({OUT_ciphertext_s2[11], OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_12__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, LED_128_Instance_state1[12]}), .Q ({OUT_ciphertext_s2[12], OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_13__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, LED_128_Instance_state1[13]}), .Q ({OUT_ciphertext_s2[13], OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_14__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, LED_128_Instance_state1[14]}), .Q ({OUT_ciphertext_s2[14], OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_15__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, LED_128_Instance_state1[15]}), .Q ({OUT_ciphertext_s2[15], OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_16__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, LED_128_Instance_state1[16]}), .Q ({OUT_ciphertext_s2[16], OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_17__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, LED_128_Instance_state1[17]}), .Q ({OUT_ciphertext_s2[17], OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_18__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3483, new_AGEMA_signal_3482, LED_128_Instance_state1[18]}), .Q ({OUT_ciphertext_s2[18], OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_19__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, LED_128_Instance_state1[19]}), .Q ({OUT_ciphertext_s2[19], OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_20__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, LED_128_Instance_state1[20]}), .Q ({OUT_ciphertext_s2[20], OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_21__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, LED_128_Instance_state1[21]}), .Q ({OUT_ciphertext_s2[21], OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_22__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3487, new_AGEMA_signal_3486, LED_128_Instance_state1[22]}), .Q ({OUT_ciphertext_s2[22], OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_23__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, LED_128_Instance_state1[23]}), .Q ({OUT_ciphertext_s2[23], OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_24__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, LED_128_Instance_state1[24]}), .Q ({OUT_ciphertext_s2[24], OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_25__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, LED_128_Instance_state1[25]}), .Q ({OUT_ciphertext_s2[25], OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_26__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, LED_128_Instance_state1[26]}), .Q ({OUT_ciphertext_s2[26], OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_27__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, LED_128_Instance_state1[27]}), .Q ({OUT_ciphertext_s2[27], OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_28__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, LED_128_Instance_state1[28]}), .Q ({OUT_ciphertext_s2[28], OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_29__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, LED_128_Instance_state1[29]}), .Q ({OUT_ciphertext_s2[29], OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_30__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, LED_128_Instance_state1[30]}), .Q ({OUT_ciphertext_s2[30], OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_31__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, LED_128_Instance_state1[31]}), .Q ({OUT_ciphertext_s2[31], OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_32__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, LED_128_Instance_state1[32]}), .Q ({OUT_ciphertext_s2[32], OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_33__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3559, new_AGEMA_signal_3558, LED_128_Instance_state1[33]}), .Q ({OUT_ciphertext_s2[33], OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_34__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3499, new_AGEMA_signal_3498, LED_128_Instance_state1[34]}), .Q ({OUT_ciphertext_s2[34], OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_35__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, LED_128_Instance_state1[35]}), .Q ({OUT_ciphertext_s2[35], OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_36__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, LED_128_Instance_state1[36]}), .Q ({OUT_ciphertext_s2[36], OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_37__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, LED_128_Instance_state1[37]}), .Q ({OUT_ciphertext_s2[37], OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_38__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, LED_128_Instance_state1[38]}), .Q ({OUT_ciphertext_s2[38], OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_39__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, LED_128_Instance_state1[39]}), .Q ({OUT_ciphertext_s2[39], OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_40__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3511, new_AGEMA_signal_3510, LED_128_Instance_state1[40]}), .Q ({OUT_ciphertext_s2[40], OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_41__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, LED_128_Instance_state1[41]}), .Q ({OUT_ciphertext_s2[41], OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_42__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, LED_128_Instance_state1[42]}), .Q ({OUT_ciphertext_s2[42], OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_43__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, LED_128_Instance_state1[43]}), .Q ({OUT_ciphertext_s2[43], OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_44__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3519, new_AGEMA_signal_3518, LED_128_Instance_state1[44]}), .Q ({OUT_ciphertext_s2[44], OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_45__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, LED_128_Instance_state1[45]}), .Q ({OUT_ciphertext_s2[45], OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_46__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3523, new_AGEMA_signal_3522, LED_128_Instance_state1[46]}), .Q ({OUT_ciphertext_s2[46], OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_47__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3571, new_AGEMA_signal_3570, LED_128_Instance_state1[47]}), .Q ({OUT_ciphertext_s2[47], OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_48__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3683, new_AGEMA_signal_3682, LED_128_Instance_state1[48]}), .Q ({OUT_ciphertext_s2[48], OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_49__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3699, new_AGEMA_signal_3698, LED_128_Instance_state1[49]}), .Q ({OUT_ciphertext_s2[49], OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_50__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3607, new_AGEMA_signal_3606, LED_128_Instance_state1[50]}), .Q ({OUT_ciphertext_s2[50], OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_51__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, LED_128_Instance_state1[51]}), .Q ({OUT_ciphertext_s2[51], OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_52__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3687, new_AGEMA_signal_3686, LED_128_Instance_state1[52]}), .Q ({OUT_ciphertext_s2[52], OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_53__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3703, new_AGEMA_signal_3702, LED_128_Instance_state1[53]}), .Q ({OUT_ciphertext_s2[53], OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_54__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, LED_128_Instance_state1[54]}), .Q ({OUT_ciphertext_s2[54], OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_55__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, LED_128_Instance_state1[55]}), .Q ({OUT_ciphertext_s2[55], OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_56__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3667, new_AGEMA_signal_3666, LED_128_Instance_state1[56]}), .Q ({OUT_ciphertext_s2[56], OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_57__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3691, new_AGEMA_signal_3690, LED_128_Instance_state1[57]}), .Q ({OUT_ciphertext_s2[57], OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_58__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, LED_128_Instance_state1[58]}), .Q ({OUT_ciphertext_s2[58], OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_59__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, LED_128_Instance_state1[59]}), .Q ({OUT_ciphertext_s2[59], OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_60__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3671, new_AGEMA_signal_3670, LED_128_Instance_state1[60]}), .Q ({OUT_ciphertext_s2[60], OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_61__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, LED_128_Instance_state1[61]}), .Q ({OUT_ciphertext_s2[61], OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_62__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3619, new_AGEMA_signal_3618, LED_128_Instance_state1[62]}), .Q ({OUT_ciphertext_s2[62], OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) LED_128_Instance_cipherstate_reg_63__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_3623, new_AGEMA_signal_3622, LED_128_Instance_state1[63]}), .Q ({OUT_ciphertext_s2[63], OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}) ) ;
    DFF_X1 internal_done_reg_FF_FF ( .CK (CLK), .D (new_AGEMA_signal_6551), .Q (OUT_done), .QN () ) ;
endmodule
