////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module CRAFT in file /AGEMA/Designs/CRAFT_round-based/AGEMA/CRAFT.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module CRAFT_HPC2_Pipeline_d2 (plaintext_s0, key_s0, clk, rst, key_s1, key_s2, plaintext_s1, plaintext_s2, Fresh, ciphertext_s0, done, ciphertext_s1, ciphertext_s2);
    input [63:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input rst ;
    input [127:0] key_s1 ;
    input [127:0] key_s2 ;
    input [63:0] plaintext_s1 ;
    input [63:0] plaintext_s2 ;
    input [767:0] Fresh ;
    output [63:0] ciphertext_s0 ;
    output done ;
    output [63:0] ciphertext_s1 ;
    output [63:0] ciphertext_s2 ;
    wire RoundConstant_4_ ;
    wire RoundConstant_0 ;
    wire done_internal ;
    wire MCInst_XOR_r0_Inst_0_n2 ;
    wire MCInst_XOR_r0_Inst_0_n1 ;
    wire MCInst_XOR_r1_Inst_0_n1 ;
    wire MCInst_XOR_r0_Inst_1_n2 ;
    wire MCInst_XOR_r0_Inst_1_n1 ;
    wire MCInst_XOR_r1_Inst_1_n1 ;
    wire MCInst_XOR_r0_Inst_2_n2 ;
    wire MCInst_XOR_r0_Inst_2_n1 ;
    wire MCInst_XOR_r1_Inst_2_n1 ;
    wire MCInst_XOR_r0_Inst_3_n2 ;
    wire MCInst_XOR_r0_Inst_3_n1 ;
    wire MCInst_XOR_r1_Inst_3_n1 ;
    wire MCInst_XOR_r0_Inst_4_n2 ;
    wire MCInst_XOR_r0_Inst_4_n1 ;
    wire MCInst_XOR_r1_Inst_4_n1 ;
    wire MCInst_XOR_r0_Inst_5_n2 ;
    wire MCInst_XOR_r0_Inst_5_n1 ;
    wire MCInst_XOR_r1_Inst_5_n1 ;
    wire MCInst_XOR_r0_Inst_6_n2 ;
    wire MCInst_XOR_r0_Inst_6_n1 ;
    wire MCInst_XOR_r1_Inst_6_n1 ;
    wire MCInst_XOR_r0_Inst_7_n2 ;
    wire MCInst_XOR_r0_Inst_7_n1 ;
    wire MCInst_XOR_r1_Inst_7_n1 ;
    wire MCInst_XOR_r0_Inst_8_n2 ;
    wire MCInst_XOR_r0_Inst_8_n1 ;
    wire MCInst_XOR_r1_Inst_8_n1 ;
    wire MCInst_XOR_r0_Inst_9_n2 ;
    wire MCInst_XOR_r0_Inst_9_n1 ;
    wire MCInst_XOR_r1_Inst_9_n1 ;
    wire MCInst_XOR_r0_Inst_10_n2 ;
    wire MCInst_XOR_r0_Inst_10_n1 ;
    wire MCInst_XOR_r1_Inst_10_n1 ;
    wire MCInst_XOR_r0_Inst_11_n2 ;
    wire MCInst_XOR_r0_Inst_11_n1 ;
    wire MCInst_XOR_r1_Inst_11_n1 ;
    wire MCInst_XOR_r0_Inst_12_n2 ;
    wire MCInst_XOR_r0_Inst_12_n1 ;
    wire MCInst_XOR_r1_Inst_12_n1 ;
    wire MCInst_XOR_r0_Inst_13_n2 ;
    wire MCInst_XOR_r0_Inst_13_n1 ;
    wire MCInst_XOR_r1_Inst_13_n1 ;
    wire MCInst_XOR_r0_Inst_14_n2 ;
    wire MCInst_XOR_r0_Inst_14_n1 ;
    wire MCInst_XOR_r1_Inst_14_n1 ;
    wire MCInst_XOR_r0_Inst_15_n2 ;
    wire MCInst_XOR_r0_Inst_15_n1 ;
    wire MCInst_XOR_r1_Inst_15_n1 ;
    wire AddKeyXOR1_XORInst_0_0_n1 ;
    wire AddKeyXOR1_XORInst_0_1_n1 ;
    wire AddKeyXOR1_XORInst_0_2_n1 ;
    wire AddKeyXOR1_XORInst_0_3_n1 ;
    wire AddKeyXOR1_XORInst_1_0_n1 ;
    wire AddKeyXOR1_XORInst_1_1_n1 ;
    wire AddKeyXOR1_XORInst_1_2_n1 ;
    wire AddKeyXOR1_XORInst_1_3_n1 ;
    wire AddKeyXOR1_XORInst_2_0_n1 ;
    wire AddKeyXOR1_XORInst_2_1_n1 ;
    wire AddKeyXOR1_XORInst_2_2_n1 ;
    wire AddKeyXOR1_XORInst_2_3_n1 ;
    wire AddKeyXOR1_XORInst_3_0_n1 ;
    wire AddKeyXOR1_XORInst_3_1_n1 ;
    wire AddKeyXOR1_XORInst_3_2_n1 ;
    wire AddKeyXOR1_XORInst_3_3_n1 ;
    wire AddKeyConstXOR_XORInst_0_0_n2 ;
    wire AddKeyConstXOR_XORInst_0_0_n1 ;
    wire AddKeyConstXOR_XORInst_0_1_n2 ;
    wire AddKeyConstXOR_XORInst_0_1_n1 ;
    wire AddKeyConstXOR_XORInst_0_2_n2 ;
    wire AddKeyConstXOR_XORInst_0_2_n1 ;
    wire AddKeyConstXOR_XORInst_0_3_n2 ;
    wire AddKeyConstXOR_XORInst_0_3_n1 ;
    wire AddKeyConstXOR_XORInst_1_0_n2 ;
    wire AddKeyConstXOR_XORInst_1_0_n1 ;
    wire AddKeyConstXOR_XORInst_1_1_n2 ;
    wire AddKeyConstXOR_XORInst_1_1_n1 ;
    wire AddKeyConstXOR_XORInst_1_2_n2 ;
    wire AddKeyConstXOR_XORInst_1_2_n1 ;
    wire AddKeyConstXOR_XORInst_1_3_n2 ;
    wire AddKeyConstXOR_XORInst_1_3_n1 ;
    wire AddKeyXOR2_XORInst_0_0_n1 ;
    wire AddKeyXOR2_XORInst_0_1_n1 ;
    wire AddKeyXOR2_XORInst_0_2_n1 ;
    wire AddKeyXOR2_XORInst_0_3_n1 ;
    wire AddKeyXOR2_XORInst_1_0_n1 ;
    wire AddKeyXOR2_XORInst_1_1_n1 ;
    wire AddKeyXOR2_XORInst_1_2_n1 ;
    wire AddKeyXOR2_XORInst_1_3_n1 ;
    wire AddKeyXOR2_XORInst_2_0_n1 ;
    wire AddKeyXOR2_XORInst_2_1_n1 ;
    wire AddKeyXOR2_XORInst_2_2_n1 ;
    wire AddKeyXOR2_XORInst_2_3_n1 ;
    wire AddKeyXOR2_XORInst_3_0_n1 ;
    wire AddKeyXOR2_XORInst_3_1_n1 ;
    wire AddKeyXOR2_XORInst_3_2_n1 ;
    wire AddKeyXOR2_XORInst_3_3_n1 ;
    wire AddKeyXOR2_XORInst_4_0_n1 ;
    wire AddKeyXOR2_XORInst_4_1_n1 ;
    wire AddKeyXOR2_XORInst_4_2_n1 ;
    wire AddKeyXOR2_XORInst_4_3_n1 ;
    wire AddKeyXOR2_XORInst_5_0_n1 ;
    wire AddKeyXOR2_XORInst_5_1_n1 ;
    wire AddKeyXOR2_XORInst_5_2_n1 ;
    wire AddKeyXOR2_XORInst_5_3_n1 ;
    wire AddKeyXOR2_XORInst_6_0_n1 ;
    wire AddKeyXOR2_XORInst_6_1_n1 ;
    wire AddKeyXOR2_XORInst_6_2_n1 ;
    wire AddKeyXOR2_XORInst_6_3_n1 ;
    wire AddKeyXOR2_XORInst_7_0_n1 ;
    wire AddKeyXOR2_XORInst_7_1_n1 ;
    wire AddKeyXOR2_XORInst_7_2_n1 ;
    wire AddKeyXOR2_XORInst_7_3_n1 ;
    wire AddKeyXOR2_XORInst_8_0_n1 ;
    wire AddKeyXOR2_XORInst_8_1_n1 ;
    wire AddKeyXOR2_XORInst_8_2_n1 ;
    wire AddKeyXOR2_XORInst_8_3_n1 ;
    wire AddKeyXOR2_XORInst_9_0_n1 ;
    wire AddKeyXOR2_XORInst_9_1_n1 ;
    wire AddKeyXOR2_XORInst_9_2_n1 ;
    wire AddKeyXOR2_XORInst_9_3_n1 ;
    wire SubCellInst_SboxInst_0_n15 ;
    wire SubCellInst_SboxInst_0_n14 ;
    wire SubCellInst_SboxInst_0_n13 ;
    wire SubCellInst_SboxInst_0_n12 ;
    wire SubCellInst_SboxInst_0_n11 ;
    wire SubCellInst_SboxInst_0_n10 ;
    wire SubCellInst_SboxInst_0_n9 ;
    wire SubCellInst_SboxInst_0_n8 ;
    wire SubCellInst_SboxInst_0_n7 ;
    wire SubCellInst_SboxInst_0_n6 ;
    wire SubCellInst_SboxInst_0_n5 ;
    wire SubCellInst_SboxInst_0_n4 ;
    wire SubCellInst_SboxInst_0_n3 ;
    wire SubCellInst_SboxInst_0_n2 ;
    wire SubCellInst_SboxInst_0_n1 ;
    wire SubCellInst_SboxInst_1_n15 ;
    wire SubCellInst_SboxInst_1_n14 ;
    wire SubCellInst_SboxInst_1_n13 ;
    wire SubCellInst_SboxInst_1_n12 ;
    wire SubCellInst_SboxInst_1_n11 ;
    wire SubCellInst_SboxInst_1_n10 ;
    wire SubCellInst_SboxInst_1_n9 ;
    wire SubCellInst_SboxInst_1_n8 ;
    wire SubCellInst_SboxInst_1_n7 ;
    wire SubCellInst_SboxInst_1_n6 ;
    wire SubCellInst_SboxInst_1_n5 ;
    wire SubCellInst_SboxInst_1_n4 ;
    wire SubCellInst_SboxInst_1_n3 ;
    wire SubCellInst_SboxInst_1_n2 ;
    wire SubCellInst_SboxInst_1_n1 ;
    wire SubCellInst_SboxInst_2_n15 ;
    wire SubCellInst_SboxInst_2_n14 ;
    wire SubCellInst_SboxInst_2_n13 ;
    wire SubCellInst_SboxInst_2_n12 ;
    wire SubCellInst_SboxInst_2_n11 ;
    wire SubCellInst_SboxInst_2_n10 ;
    wire SubCellInst_SboxInst_2_n9 ;
    wire SubCellInst_SboxInst_2_n8 ;
    wire SubCellInst_SboxInst_2_n7 ;
    wire SubCellInst_SboxInst_2_n6 ;
    wire SubCellInst_SboxInst_2_n5 ;
    wire SubCellInst_SboxInst_2_n4 ;
    wire SubCellInst_SboxInst_2_n3 ;
    wire SubCellInst_SboxInst_2_n2 ;
    wire SubCellInst_SboxInst_2_n1 ;
    wire SubCellInst_SboxInst_3_n15 ;
    wire SubCellInst_SboxInst_3_n14 ;
    wire SubCellInst_SboxInst_3_n13 ;
    wire SubCellInst_SboxInst_3_n12 ;
    wire SubCellInst_SboxInst_3_n11 ;
    wire SubCellInst_SboxInst_3_n10 ;
    wire SubCellInst_SboxInst_3_n9 ;
    wire SubCellInst_SboxInst_3_n8 ;
    wire SubCellInst_SboxInst_3_n7 ;
    wire SubCellInst_SboxInst_3_n6 ;
    wire SubCellInst_SboxInst_3_n5 ;
    wire SubCellInst_SboxInst_3_n4 ;
    wire SubCellInst_SboxInst_3_n3 ;
    wire SubCellInst_SboxInst_3_n2 ;
    wire SubCellInst_SboxInst_3_n1 ;
    wire SubCellInst_SboxInst_4_n15 ;
    wire SubCellInst_SboxInst_4_n14 ;
    wire SubCellInst_SboxInst_4_n13 ;
    wire SubCellInst_SboxInst_4_n12 ;
    wire SubCellInst_SboxInst_4_n11 ;
    wire SubCellInst_SboxInst_4_n10 ;
    wire SubCellInst_SboxInst_4_n9 ;
    wire SubCellInst_SboxInst_4_n8 ;
    wire SubCellInst_SboxInst_4_n7 ;
    wire SubCellInst_SboxInst_4_n6 ;
    wire SubCellInst_SboxInst_4_n5 ;
    wire SubCellInst_SboxInst_4_n4 ;
    wire SubCellInst_SboxInst_4_n3 ;
    wire SubCellInst_SboxInst_4_n2 ;
    wire SubCellInst_SboxInst_4_n1 ;
    wire SubCellInst_SboxInst_5_n15 ;
    wire SubCellInst_SboxInst_5_n14 ;
    wire SubCellInst_SboxInst_5_n13 ;
    wire SubCellInst_SboxInst_5_n12 ;
    wire SubCellInst_SboxInst_5_n11 ;
    wire SubCellInst_SboxInst_5_n10 ;
    wire SubCellInst_SboxInst_5_n9 ;
    wire SubCellInst_SboxInst_5_n8 ;
    wire SubCellInst_SboxInst_5_n7 ;
    wire SubCellInst_SboxInst_5_n6 ;
    wire SubCellInst_SboxInst_5_n5 ;
    wire SubCellInst_SboxInst_5_n4 ;
    wire SubCellInst_SboxInst_5_n3 ;
    wire SubCellInst_SboxInst_5_n2 ;
    wire SubCellInst_SboxInst_5_n1 ;
    wire SubCellInst_SboxInst_6_n15 ;
    wire SubCellInst_SboxInst_6_n14 ;
    wire SubCellInst_SboxInst_6_n13 ;
    wire SubCellInst_SboxInst_6_n12 ;
    wire SubCellInst_SboxInst_6_n11 ;
    wire SubCellInst_SboxInst_6_n10 ;
    wire SubCellInst_SboxInst_6_n9 ;
    wire SubCellInst_SboxInst_6_n8 ;
    wire SubCellInst_SboxInst_6_n7 ;
    wire SubCellInst_SboxInst_6_n6 ;
    wire SubCellInst_SboxInst_6_n5 ;
    wire SubCellInst_SboxInst_6_n4 ;
    wire SubCellInst_SboxInst_6_n3 ;
    wire SubCellInst_SboxInst_6_n2 ;
    wire SubCellInst_SboxInst_6_n1 ;
    wire SubCellInst_SboxInst_7_n15 ;
    wire SubCellInst_SboxInst_7_n14 ;
    wire SubCellInst_SboxInst_7_n13 ;
    wire SubCellInst_SboxInst_7_n12 ;
    wire SubCellInst_SboxInst_7_n11 ;
    wire SubCellInst_SboxInst_7_n10 ;
    wire SubCellInst_SboxInst_7_n9 ;
    wire SubCellInst_SboxInst_7_n8 ;
    wire SubCellInst_SboxInst_7_n7 ;
    wire SubCellInst_SboxInst_7_n6 ;
    wire SubCellInst_SboxInst_7_n5 ;
    wire SubCellInst_SboxInst_7_n4 ;
    wire SubCellInst_SboxInst_7_n3 ;
    wire SubCellInst_SboxInst_7_n2 ;
    wire SubCellInst_SboxInst_7_n1 ;
    wire SubCellInst_SboxInst_8_n15 ;
    wire SubCellInst_SboxInst_8_n14 ;
    wire SubCellInst_SboxInst_8_n13 ;
    wire SubCellInst_SboxInst_8_n12 ;
    wire SubCellInst_SboxInst_8_n11 ;
    wire SubCellInst_SboxInst_8_n10 ;
    wire SubCellInst_SboxInst_8_n9 ;
    wire SubCellInst_SboxInst_8_n8 ;
    wire SubCellInst_SboxInst_8_n7 ;
    wire SubCellInst_SboxInst_8_n6 ;
    wire SubCellInst_SboxInst_8_n5 ;
    wire SubCellInst_SboxInst_8_n4 ;
    wire SubCellInst_SboxInst_8_n3 ;
    wire SubCellInst_SboxInst_8_n2 ;
    wire SubCellInst_SboxInst_8_n1 ;
    wire SubCellInst_SboxInst_9_n15 ;
    wire SubCellInst_SboxInst_9_n14 ;
    wire SubCellInst_SboxInst_9_n13 ;
    wire SubCellInst_SboxInst_9_n12 ;
    wire SubCellInst_SboxInst_9_n11 ;
    wire SubCellInst_SboxInst_9_n10 ;
    wire SubCellInst_SboxInst_9_n9 ;
    wire SubCellInst_SboxInst_9_n8 ;
    wire SubCellInst_SboxInst_9_n7 ;
    wire SubCellInst_SboxInst_9_n6 ;
    wire SubCellInst_SboxInst_9_n5 ;
    wire SubCellInst_SboxInst_9_n4 ;
    wire SubCellInst_SboxInst_9_n3 ;
    wire SubCellInst_SboxInst_9_n2 ;
    wire SubCellInst_SboxInst_9_n1 ;
    wire SubCellInst_SboxInst_10_n15 ;
    wire SubCellInst_SboxInst_10_n14 ;
    wire SubCellInst_SboxInst_10_n13 ;
    wire SubCellInst_SboxInst_10_n12 ;
    wire SubCellInst_SboxInst_10_n11 ;
    wire SubCellInst_SboxInst_10_n10 ;
    wire SubCellInst_SboxInst_10_n9 ;
    wire SubCellInst_SboxInst_10_n8 ;
    wire SubCellInst_SboxInst_10_n7 ;
    wire SubCellInst_SboxInst_10_n6 ;
    wire SubCellInst_SboxInst_10_n5 ;
    wire SubCellInst_SboxInst_10_n4 ;
    wire SubCellInst_SboxInst_10_n3 ;
    wire SubCellInst_SboxInst_10_n2 ;
    wire SubCellInst_SboxInst_10_n1 ;
    wire SubCellInst_SboxInst_11_n15 ;
    wire SubCellInst_SboxInst_11_n14 ;
    wire SubCellInst_SboxInst_11_n13 ;
    wire SubCellInst_SboxInst_11_n12 ;
    wire SubCellInst_SboxInst_11_n11 ;
    wire SubCellInst_SboxInst_11_n10 ;
    wire SubCellInst_SboxInst_11_n9 ;
    wire SubCellInst_SboxInst_11_n8 ;
    wire SubCellInst_SboxInst_11_n7 ;
    wire SubCellInst_SboxInst_11_n6 ;
    wire SubCellInst_SboxInst_11_n5 ;
    wire SubCellInst_SboxInst_11_n4 ;
    wire SubCellInst_SboxInst_11_n3 ;
    wire SubCellInst_SboxInst_11_n2 ;
    wire SubCellInst_SboxInst_11_n1 ;
    wire SubCellInst_SboxInst_12_n15 ;
    wire SubCellInst_SboxInst_12_n14 ;
    wire SubCellInst_SboxInst_12_n13 ;
    wire SubCellInst_SboxInst_12_n12 ;
    wire SubCellInst_SboxInst_12_n11 ;
    wire SubCellInst_SboxInst_12_n10 ;
    wire SubCellInst_SboxInst_12_n9 ;
    wire SubCellInst_SboxInst_12_n8 ;
    wire SubCellInst_SboxInst_12_n7 ;
    wire SubCellInst_SboxInst_12_n6 ;
    wire SubCellInst_SboxInst_12_n5 ;
    wire SubCellInst_SboxInst_12_n4 ;
    wire SubCellInst_SboxInst_12_n3 ;
    wire SubCellInst_SboxInst_12_n2 ;
    wire SubCellInst_SboxInst_12_n1 ;
    wire SubCellInst_SboxInst_13_n15 ;
    wire SubCellInst_SboxInst_13_n14 ;
    wire SubCellInst_SboxInst_13_n13 ;
    wire SubCellInst_SboxInst_13_n12 ;
    wire SubCellInst_SboxInst_13_n11 ;
    wire SubCellInst_SboxInst_13_n10 ;
    wire SubCellInst_SboxInst_13_n9 ;
    wire SubCellInst_SboxInst_13_n8 ;
    wire SubCellInst_SboxInst_13_n7 ;
    wire SubCellInst_SboxInst_13_n6 ;
    wire SubCellInst_SboxInst_13_n5 ;
    wire SubCellInst_SboxInst_13_n4 ;
    wire SubCellInst_SboxInst_13_n3 ;
    wire SubCellInst_SboxInst_13_n2 ;
    wire SubCellInst_SboxInst_13_n1 ;
    wire SubCellInst_SboxInst_14_n15 ;
    wire SubCellInst_SboxInst_14_n14 ;
    wire SubCellInst_SboxInst_14_n13 ;
    wire SubCellInst_SboxInst_14_n12 ;
    wire SubCellInst_SboxInst_14_n11 ;
    wire SubCellInst_SboxInst_14_n10 ;
    wire SubCellInst_SboxInst_14_n9 ;
    wire SubCellInst_SboxInst_14_n8 ;
    wire SubCellInst_SboxInst_14_n7 ;
    wire SubCellInst_SboxInst_14_n6 ;
    wire SubCellInst_SboxInst_14_n5 ;
    wire SubCellInst_SboxInst_14_n4 ;
    wire SubCellInst_SboxInst_14_n3 ;
    wire SubCellInst_SboxInst_14_n2 ;
    wire SubCellInst_SboxInst_14_n1 ;
    wire SubCellInst_SboxInst_15_n15 ;
    wire SubCellInst_SboxInst_15_n14 ;
    wire SubCellInst_SboxInst_15_n13 ;
    wire SubCellInst_SboxInst_15_n12 ;
    wire SubCellInst_SboxInst_15_n11 ;
    wire SubCellInst_SboxInst_15_n10 ;
    wire SubCellInst_SboxInst_15_n9 ;
    wire SubCellInst_SboxInst_15_n8 ;
    wire SubCellInst_SboxInst_15_n7 ;
    wire SubCellInst_SboxInst_15_n6 ;
    wire SubCellInst_SboxInst_15_n5 ;
    wire SubCellInst_SboxInst_15_n4 ;
    wire SubCellInst_SboxInst_15_n3 ;
    wire SubCellInst_SboxInst_15_n2 ;
    wire SubCellInst_SboxInst_15_n1 ;
    wire KeyMUX_n9 ;
    wire KeyMUX_n8 ;
    wire KeyMUX_n7 ;
    wire FSMSignalsInst_n5 ;
    wire FSMSignalsInst_n4 ;
    wire FSMSignalsInst_n3 ;
    wire FSMSignalsInst_n2 ;
    wire FSMSignalsInst_n1 ;
    wire selectsUpdateInst_n3 ;
    wire [63:0] Feedback ;
    wire [63:32] MCInput ;
    wire [63:0] MCOutput ;
    wire [63:0] SelectedKey ;
    wire [63:0] AddRoundKeyOutput ;
    wire [1:0] selects ;
    wire [6:0] FSMReg ;
    wire [6:0] FSMUpdate ;
    wire [1:0] selectsReg ;
    wire [1:0] selectsNext ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4235 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4282 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4290 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4308 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4318 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4325 ;
    wire new_AGEMA_signal_4326 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4336 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4354 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4361 ;
    wire new_AGEMA_signal_4362 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4372 ;
    wire new_AGEMA_signal_4373 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4378 ;
    wire new_AGEMA_signal_4379 ;
    wire new_AGEMA_signal_4380 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4382 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4497 ;
    wire new_AGEMA_signal_4498 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5195 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5202 ;
    wire new_AGEMA_signal_5203 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5207 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5213 ;
    wire new_AGEMA_signal_5214 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5219 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5226 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5231 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5238 ;
    wire new_AGEMA_signal_5239 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5249 ;
    wire new_AGEMA_signal_5250 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5255 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5262 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5273 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5291 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5303 ;
    wire new_AGEMA_signal_5304 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5309 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6654 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;
    wire new_AGEMA_signal_6672 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6677 ;
    wire new_AGEMA_signal_6678 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6682 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6688 ;
    wire new_AGEMA_signal_6689 ;
    wire new_AGEMA_signal_6690 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6695 ;
    wire new_AGEMA_signal_6696 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6700 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6706 ;
    wire new_AGEMA_signal_6707 ;
    wire new_AGEMA_signal_6708 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6713 ;
    wire new_AGEMA_signal_6714 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6718 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6724 ;
    wire new_AGEMA_signal_6725 ;
    wire new_AGEMA_signal_6726 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7036 ;
    wire new_AGEMA_signal_7037 ;
    wire new_AGEMA_signal_7038 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7042 ;
    wire new_AGEMA_signal_7043 ;
    wire new_AGEMA_signal_7044 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7048 ;
    wire new_AGEMA_signal_7049 ;
    wire new_AGEMA_signal_7050 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7054 ;
    wire new_AGEMA_signal_7055 ;
    wire new_AGEMA_signal_7056 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7060 ;
    wire new_AGEMA_signal_7061 ;
    wire new_AGEMA_signal_7062 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7066 ;
    wire new_AGEMA_signal_7067 ;
    wire new_AGEMA_signal_7068 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7072 ;
    wire new_AGEMA_signal_7073 ;
    wire new_AGEMA_signal_7074 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7078 ;
    wire new_AGEMA_signal_7079 ;
    wire new_AGEMA_signal_7080 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7084 ;
    wire new_AGEMA_signal_7085 ;
    wire new_AGEMA_signal_7086 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7090 ;
    wire new_AGEMA_signal_7091 ;
    wire new_AGEMA_signal_7092 ;
    wire new_AGEMA_signal_7093 ;
    wire new_AGEMA_signal_7094 ;
    wire new_AGEMA_signal_7095 ;
    wire new_AGEMA_signal_7096 ;
    wire new_AGEMA_signal_7097 ;
    wire new_AGEMA_signal_7098 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7102 ;
    wire new_AGEMA_signal_7103 ;
    wire new_AGEMA_signal_7104 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7108 ;
    wire new_AGEMA_signal_7109 ;
    wire new_AGEMA_signal_7110 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7114 ;
    wire new_AGEMA_signal_7115 ;
    wire new_AGEMA_signal_7116 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7120 ;
    wire new_AGEMA_signal_7121 ;
    wire new_AGEMA_signal_7122 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7126 ;
    wire new_AGEMA_signal_7127 ;
    wire new_AGEMA_signal_7128 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7132 ;
    wire new_AGEMA_signal_7133 ;
    wire new_AGEMA_signal_7134 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7138 ;
    wire new_AGEMA_signal_7139 ;
    wire new_AGEMA_signal_7140 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7144 ;
    wire new_AGEMA_signal_7145 ;
    wire new_AGEMA_signal_7146 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7150 ;
    wire new_AGEMA_signal_7151 ;
    wire new_AGEMA_signal_7152 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7156 ;
    wire new_AGEMA_signal_7157 ;
    wire new_AGEMA_signal_7158 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7162 ;
    wire new_AGEMA_signal_7163 ;
    wire new_AGEMA_signal_7164 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7168 ;
    wire new_AGEMA_signal_7169 ;
    wire new_AGEMA_signal_7170 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7174 ;
    wire new_AGEMA_signal_7175 ;
    wire new_AGEMA_signal_7176 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7180 ;
    wire new_AGEMA_signal_7181 ;
    wire new_AGEMA_signal_7182 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7186 ;
    wire new_AGEMA_signal_7187 ;
    wire new_AGEMA_signal_7188 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7192 ;
    wire new_AGEMA_signal_7193 ;
    wire new_AGEMA_signal_7194 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7198 ;
    wire new_AGEMA_signal_7199 ;
    wire new_AGEMA_signal_7200 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7204 ;
    wire new_AGEMA_signal_7205 ;
    wire new_AGEMA_signal_7206 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7489 ;
    wire new_AGEMA_signal_7490 ;
    wire new_AGEMA_signal_7491 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7495 ;
    wire new_AGEMA_signal_7496 ;
    wire new_AGEMA_signal_7497 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7499 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7501 ;
    wire new_AGEMA_signal_7502 ;
    wire new_AGEMA_signal_7503 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7507 ;
    wire new_AGEMA_signal_7508 ;
    wire new_AGEMA_signal_7509 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7513 ;
    wire new_AGEMA_signal_7514 ;
    wire new_AGEMA_signal_7515 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7519 ;
    wire new_AGEMA_signal_7520 ;
    wire new_AGEMA_signal_7521 ;
    wire new_AGEMA_signal_7522 ;

    /* cells in depth 0 */
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2030, new_AGEMA_signal_2029, SelectedKey[40]}), .b ({1'b0, 1'b0, RoundConstant_0}), .c ({new_AGEMA_signal_2396, new_AGEMA_signal_2395, AddKeyConstXOR_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2036, new_AGEMA_signal_2035, SelectedKey[41]}), .b ({1'b0, 1'b0, FSMUpdate[0]}), .c ({new_AGEMA_signal_2398, new_AGEMA_signal_2397, AddKeyConstXOR_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2042, new_AGEMA_signal_2041, SelectedKey[42]}), .b ({1'b0, 1'b0, FSMUpdate[1]}), .c ({new_AGEMA_signal_2400, new_AGEMA_signal_2399, AddKeyConstXOR_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2048, new_AGEMA_signal_2047, SelectedKey[43]}), .b ({1'b0, 1'b0, 1'b0}), .c ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, AddKeyConstXOR_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, SelectedKey[44]}), .b ({1'b0, 1'b0, RoundConstant_4_}), .c ({new_AGEMA_signal_2404, new_AGEMA_signal_2403, AddKeyConstXOR_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2060, new_AGEMA_signal_2059, SelectedKey[45]}), .b ({1'b0, 1'b0, FSMUpdate[3]}), .c ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, AddKeyConstXOR_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2066, new_AGEMA_signal_2065, SelectedKey[46]}), .b ({1'b0, 1'b0, FSMUpdate[4]}), .c ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, AddKeyConstXOR_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, SelectedKey[47]}), .b ({1'b0, 1'b0, FSMUpdate[5]}), .c ({new_AGEMA_signal_2410, new_AGEMA_signal_2409, AddKeyConstXOR_XORInst_1_3_n1}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U4 ( .a ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_1030, new_AGEMA_signal_1029, SubCellInst_SboxInst_0_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U2 ( .a ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_1032, new_AGEMA_signal_1031, SubCellInst_SboxInst_0_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U1 ( .a ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, SubCellInst_SboxInst_0_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U4 ( .a ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, SubCellInst_SboxInst_1_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U2 ( .a ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .b ({new_AGEMA_signal_1048, new_AGEMA_signal_1047, SubCellInst_SboxInst_1_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U1 ( .a ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .b ({new_AGEMA_signal_1050, new_AGEMA_signal_1049, SubCellInst_SboxInst_1_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U4 ( .a ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .b ({new_AGEMA_signal_1062, new_AGEMA_signal_1061, SubCellInst_SboxInst_2_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U2 ( .a ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, SubCellInst_SboxInst_2_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U1 ( .a ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({new_AGEMA_signal_1066, new_AGEMA_signal_1065, SubCellInst_SboxInst_2_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U4 ( .a ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_1078, new_AGEMA_signal_1077, SubCellInst_SboxInst_3_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U2 ( .a ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_1080, new_AGEMA_signal_1079, SubCellInst_SboxInst_3_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U1 ( .a ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .b ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, SubCellInst_SboxInst_3_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U4 ( .a ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, SubCellInst_SboxInst_4_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U2 ( .a ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .b ({new_AGEMA_signal_1096, new_AGEMA_signal_1095, SubCellInst_SboxInst_4_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U1 ( .a ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .b ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, SubCellInst_SboxInst_4_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U4 ( .a ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .b ({new_AGEMA_signal_1110, new_AGEMA_signal_1109, SubCellInst_SboxInst_5_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U2 ( .a ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, SubCellInst_SboxInst_5_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U1 ( .a ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, SubCellInst_SboxInst_5_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U4 ( .a ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_1126, new_AGEMA_signal_1125, SubCellInst_SboxInst_6_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U2 ( .a ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .b ({new_AGEMA_signal_1128, new_AGEMA_signal_1127, SubCellInst_SboxInst_6_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U1 ( .a ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .b ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, SubCellInst_SboxInst_6_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U4 ( .a ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .b ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, SubCellInst_SboxInst_7_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U2 ( .a ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, SubCellInst_SboxInst_7_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U1 ( .a ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({new_AGEMA_signal_1146, new_AGEMA_signal_1145, SubCellInst_SboxInst_7_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U4 ( .a ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, SubCellInst_SboxInst_8_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U2 ( .a ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .b ({new_AGEMA_signal_1160, new_AGEMA_signal_1159, SubCellInst_SboxInst_8_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U1 ( .a ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .b ({new_AGEMA_signal_1162, new_AGEMA_signal_1161, SubCellInst_SboxInst_8_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U4 ( .a ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_1174, new_AGEMA_signal_1173, SubCellInst_SboxInst_9_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U2 ( .a ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_1176, new_AGEMA_signal_1175, SubCellInst_SboxInst_9_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U1 ( .a ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, SubCellInst_SboxInst_9_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U4 ( .a ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, SubCellInst_SboxInst_10_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U2 ( .a ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_1192, new_AGEMA_signal_1191, SubCellInst_SboxInst_10_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U1 ( .a ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .b ({new_AGEMA_signal_1194, new_AGEMA_signal_1193, SubCellInst_SboxInst_10_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U4 ( .a ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .b ({new_AGEMA_signal_1206, new_AGEMA_signal_1205, SubCellInst_SboxInst_11_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U2 ( .a ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, SubCellInst_SboxInst_11_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U1 ( .a ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({new_AGEMA_signal_1210, new_AGEMA_signal_1209, SubCellInst_SboxInst_11_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U4 ( .a ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .b ({new_AGEMA_signal_1222, new_AGEMA_signal_1221, SubCellInst_SboxInst_12_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U2 ( .a ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({new_AGEMA_signal_1224, new_AGEMA_signal_1223, SubCellInst_SboxInst_12_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U1 ( .a ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({new_AGEMA_signal_1226, new_AGEMA_signal_1225, SubCellInst_SboxInst_12_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U4 ( .a ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, SubCellInst_SboxInst_13_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U2 ( .a ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .b ({new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_13_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U1 ( .a ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .b ({new_AGEMA_signal_1242, new_AGEMA_signal_1241, SubCellInst_SboxInst_13_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U4 ( .a ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .b ({new_AGEMA_signal_1254, new_AGEMA_signal_1253, SubCellInst_SboxInst_14_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U2 ( .a ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, SubCellInst_SboxInst_14_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U1 ( .a ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_14_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U4 ( .a ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_1270, new_AGEMA_signal_1269, SubCellInst_SboxInst_15_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U2 ( .a ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .b ({new_AGEMA_signal_1272, new_AGEMA_signal_1271, SubCellInst_SboxInst_15_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U1 ( .a ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .b ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, SubCellInst_SboxInst_15_n9}) ) ;
    INV_X1 KeyMUX_U3 ( .A (selects[0]), .ZN (KeyMUX_n9) ) ;
    INV_X1 KeyMUX_U2 ( .A (KeyMUX_n9), .ZN (KeyMUX_n8) ) ;
    INV_X1 KeyMUX_U1 ( .A (KeyMUX_n9), .ZN (KeyMUX_n7) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_0_U1 ( .s (selects[0]), .b ({key_s2[64], key_s1[64], key_s0[64]}), .a ({key_s2[0], key_s1[0], key_s0[0]}), .c ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, SelectedKey[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_1_U1 ( .s (KeyMUX_n8), .b ({key_s2[65], key_s1[65], key_s0[65]}), .a ({key_s2[1], key_s1[1], key_s0[1]}), .c ({new_AGEMA_signal_1856, new_AGEMA_signal_1855, SelectedKey[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_2_U1 ( .s (selects[0]), .b ({key_s2[66], key_s1[66], key_s0[66]}), .a ({key_s2[2], key_s1[2], key_s0[2]}), .c ({new_AGEMA_signal_1478, new_AGEMA_signal_1477, SelectedKey[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_3_U1 ( .s (KeyMUX_n8), .b ({key_s2[67], key_s1[67], key_s0[67]}), .a ({key_s2[3], key_s1[3], key_s0[3]}), .c ({new_AGEMA_signal_1862, new_AGEMA_signal_1861, SelectedKey[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_4_U1 ( .s (KeyMUX_n8), .b ({key_s2[68], key_s1[68], key_s0[68]}), .a ({key_s2[4], key_s1[4], key_s0[4]}), .c ({new_AGEMA_signal_1868, new_AGEMA_signal_1867, SelectedKey[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_5_U1 ( .s (KeyMUX_n8), .b ({key_s2[69], key_s1[69], key_s0[69]}), .a ({key_s2[5], key_s1[5], key_s0[5]}), .c ({new_AGEMA_signal_1874, new_AGEMA_signal_1873, SelectedKey[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_6_U1 ( .s (KeyMUX_n8), .b ({key_s2[70], key_s1[70], key_s0[70]}), .a ({key_s2[6], key_s1[6], key_s0[6]}), .c ({new_AGEMA_signal_1880, new_AGEMA_signal_1879, SelectedKey[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_7_U1 ( .s (KeyMUX_n8), .b ({key_s2[71], key_s1[71], key_s0[71]}), .a ({key_s2[7], key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_1886, new_AGEMA_signal_1885, SelectedKey[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_8_U1 ( .s (KeyMUX_n8), .b ({key_s2[72], key_s1[72], key_s0[72]}), .a ({key_s2[8], key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_1892, new_AGEMA_signal_1891, SelectedKey[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_9_U1 ( .s (KeyMUX_n8), .b ({key_s2[73], key_s1[73], key_s0[73]}), .a ({key_s2[9], key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_1898, new_AGEMA_signal_1897, SelectedKey[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_10_U1 ( .s (KeyMUX_n8), .b ({key_s2[74], key_s1[74], key_s0[74]}), .a ({key_s2[10], key_s1[10], key_s0[10]}), .c ({new_AGEMA_signal_1904, new_AGEMA_signal_1903, SelectedKey[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_11_U1 ( .s (KeyMUX_n8), .b ({key_s2[75], key_s1[75], key_s0[75]}), .a ({key_s2[11], key_s1[11], key_s0[11]}), .c ({new_AGEMA_signal_1910, new_AGEMA_signal_1909, SelectedKey[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_12_U1 ( .s (KeyMUX_n8), .b ({key_s2[76], key_s1[76], key_s0[76]}), .a ({key_s2[12], key_s1[12], key_s0[12]}), .c ({new_AGEMA_signal_1916, new_AGEMA_signal_1915, SelectedKey[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_13_U1 ( .s (KeyMUX_n8), .b ({key_s2[77], key_s1[77], key_s0[77]}), .a ({key_s2[13], key_s1[13], key_s0[13]}), .c ({new_AGEMA_signal_1922, new_AGEMA_signal_1921, SelectedKey[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_14_U1 ( .s (KeyMUX_n8), .b ({key_s2[78], key_s1[78], key_s0[78]}), .a ({key_s2[14], key_s1[14], key_s0[14]}), .c ({new_AGEMA_signal_1928, new_AGEMA_signal_1927, SelectedKey[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_15_U1 ( .s (KeyMUX_n8), .b ({key_s2[79], key_s1[79], key_s0[79]}), .a ({key_s2[15], key_s1[15], key_s0[15]}), .c ({new_AGEMA_signal_1934, new_AGEMA_signal_1933, SelectedKey[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_16_U1 ( .s (KeyMUX_n8), .b ({key_s2[80], key_s1[80], key_s0[80]}), .a ({key_s2[16], key_s1[16], key_s0[16]}), .c ({new_AGEMA_signal_1940, new_AGEMA_signal_1939, SelectedKey[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_17_U1 ( .s (KeyMUX_n8), .b ({key_s2[81], key_s1[81], key_s0[81]}), .a ({key_s2[17], key_s1[17], key_s0[17]}), .c ({new_AGEMA_signal_1946, new_AGEMA_signal_1945, SelectedKey[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_18_U1 ( .s (KeyMUX_n8), .b ({key_s2[82], key_s1[82], key_s0[82]}), .a ({key_s2[18], key_s1[18], key_s0[18]}), .c ({new_AGEMA_signal_1952, new_AGEMA_signal_1951, SelectedKey[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_19_U1 ( .s (KeyMUX_n8), .b ({key_s2[83], key_s1[83], key_s0[83]}), .a ({key_s2[19], key_s1[19], key_s0[19]}), .c ({new_AGEMA_signal_1958, new_AGEMA_signal_1957, SelectedKey[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_20_U1 ( .s (KeyMUX_n8), .b ({key_s2[84], key_s1[84], key_s0[84]}), .a ({key_s2[20], key_s1[20], key_s0[20]}), .c ({new_AGEMA_signal_1964, new_AGEMA_signal_1963, SelectedKey[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_21_U1 ( .s (KeyMUX_n8), .b ({key_s2[85], key_s1[85], key_s0[85]}), .a ({key_s2[21], key_s1[21], key_s0[21]}), .c ({new_AGEMA_signal_1970, new_AGEMA_signal_1969, SelectedKey[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_22_U1 ( .s (selects[0]), .b ({key_s2[86], key_s1[86], key_s0[86]}), .a ({key_s2[22], key_s1[22], key_s0[22]}), .c ({new_AGEMA_signal_1484, new_AGEMA_signal_1483, SelectedKey[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_23_U1 ( .s (selects[0]), .b ({key_s2[87], key_s1[87], key_s0[87]}), .a ({key_s2[23], key_s1[23], key_s0[23]}), .c ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, SelectedKey[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_24_U1 ( .s (selects[0]), .b ({key_s2[88], key_s1[88], key_s0[88]}), .a ({key_s2[24], key_s1[24], key_s0[24]}), .c ({new_AGEMA_signal_1496, new_AGEMA_signal_1495, SelectedKey[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_25_U1 ( .s (selects[0]), .b ({key_s2[89], key_s1[89], key_s0[89]}), .a ({key_s2[25], key_s1[25], key_s0[25]}), .c ({new_AGEMA_signal_1502, new_AGEMA_signal_1501, SelectedKey[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_26_U1 ( .s (selects[0]), .b ({key_s2[90], key_s1[90], key_s0[90]}), .a ({key_s2[26], key_s1[26], key_s0[26]}), .c ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, SelectedKey[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_27_U1 ( .s (selects[0]), .b ({key_s2[91], key_s1[91], key_s0[91]}), .a ({key_s2[27], key_s1[27], key_s0[27]}), .c ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, SelectedKey[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_28_U1 ( .s (KeyMUX_n7), .b ({key_s2[92], key_s1[92], key_s0[92]}), .a ({key_s2[28], key_s1[28], key_s0[28]}), .c ({new_AGEMA_signal_1976, new_AGEMA_signal_1975, SelectedKey[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_29_U1 ( .s (KeyMUX_n7), .b ({key_s2[93], key_s1[93], key_s0[93]}), .a ({key_s2[29], key_s1[29], key_s0[29]}), .c ({new_AGEMA_signal_1982, new_AGEMA_signal_1981, SelectedKey[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_30_U1 ( .s (KeyMUX_n7), .b ({key_s2[94], key_s1[94], key_s0[94]}), .a ({key_s2[30], key_s1[30], key_s0[30]}), .c ({new_AGEMA_signal_1988, new_AGEMA_signal_1987, SelectedKey[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_31_U1 ( .s (KeyMUX_n7), .b ({key_s2[95], key_s1[95], key_s0[95]}), .a ({key_s2[31], key_s1[31], key_s0[31]}), .c ({new_AGEMA_signal_1994, new_AGEMA_signal_1993, SelectedKey[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_32_U1 ( .s (KeyMUX_n7), .b ({key_s2[96], key_s1[96], key_s0[96]}), .a ({key_s2[32], key_s1[32], key_s0[32]}), .c ({new_AGEMA_signal_2000, new_AGEMA_signal_1999, SelectedKey[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_33_U1 ( .s (selects[0]), .b ({key_s2[97], key_s1[97], key_s0[97]}), .a ({key_s2[33], key_s1[33], key_s0[33]}), .c ({new_AGEMA_signal_1520, new_AGEMA_signal_1519, SelectedKey[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_34_U1 ( .s (KeyMUX_n7), .b ({key_s2[98], key_s1[98], key_s0[98]}), .a ({key_s2[34], key_s1[34], key_s0[34]}), .c ({new_AGEMA_signal_2006, new_AGEMA_signal_2005, SelectedKey[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_35_U1 ( .s (KeyMUX_n7), .b ({key_s2[99], key_s1[99], key_s0[99]}), .a ({key_s2[35], key_s1[35], key_s0[35]}), .c ({new_AGEMA_signal_2012, new_AGEMA_signal_2011, SelectedKey[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_36_U1 ( .s (selects[0]), .b ({key_s2[100], key_s1[100], key_s0[100]}), .a ({key_s2[36], key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, SelectedKey[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_37_U1 ( .s (KeyMUX_n7), .b ({key_s2[101], key_s1[101], key_s0[101]}), .a ({key_s2[37], key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_2018, new_AGEMA_signal_2017, SelectedKey[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_38_U1 ( .s (KeyMUX_n7), .b ({key_s2[102], key_s1[102], key_s0[102]}), .a ({key_s2[38], key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_2024, new_AGEMA_signal_2023, SelectedKey[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_39_U1 ( .s (selects[0]), .b ({key_s2[103], key_s1[103], key_s0[103]}), .a ({key_s2[39], key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_1532, new_AGEMA_signal_1531, SelectedKey[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_40_U1 ( .s (KeyMUX_n7), .b ({key_s2[104], key_s1[104], key_s0[104]}), .a ({key_s2[40], key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_2030, new_AGEMA_signal_2029, SelectedKey[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_41_U1 ( .s (KeyMUX_n7), .b ({key_s2[105], key_s1[105], key_s0[105]}), .a ({key_s2[41], key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_2036, new_AGEMA_signal_2035, SelectedKey[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_42_U1 ( .s (KeyMUX_n7), .b ({key_s2[106], key_s1[106], key_s0[106]}), .a ({key_s2[42], key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_2042, new_AGEMA_signal_2041, SelectedKey[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_43_U1 ( .s (KeyMUX_n7), .b ({key_s2[107], key_s1[107], key_s0[107]}), .a ({key_s2[43], key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_2048, new_AGEMA_signal_2047, SelectedKey[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_44_U1 ( .s (KeyMUX_n7), .b ({key_s2[108], key_s1[108], key_s0[108]}), .a ({key_s2[44], key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, SelectedKey[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_45_U1 ( .s (KeyMUX_n7), .b ({key_s2[109], key_s1[109], key_s0[109]}), .a ({key_s2[45], key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_2060, new_AGEMA_signal_2059, SelectedKey[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_46_U1 ( .s (KeyMUX_n7), .b ({key_s2[110], key_s1[110], key_s0[110]}), .a ({key_s2[46], key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_2066, new_AGEMA_signal_2065, SelectedKey[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_47_U1 ( .s (KeyMUX_n7), .b ({key_s2[111], key_s1[111], key_s0[111]}), .a ({key_s2[47], key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, SelectedKey[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_48_U1 ( .s (KeyMUX_n7), .b ({key_s2[112], key_s1[112], key_s0[112]}), .a ({key_s2[48], key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, SelectedKey[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_49_U1 ( .s (KeyMUX_n7), .b ({key_s2[113], key_s1[113], key_s0[113]}), .a ({key_s2[49], key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_2084, new_AGEMA_signal_2083, SelectedKey[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_50_U1 ( .s (KeyMUX_n7), .b ({key_s2[114], key_s1[114], key_s0[114]}), .a ({key_s2[50], key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, SelectedKey[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_51_U1 ( .s (KeyMUX_n7), .b ({key_s2[115], key_s1[115], key_s0[115]}), .a ({key_s2[51], key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_2096, new_AGEMA_signal_2095, SelectedKey[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_52_U1 ( .s (KeyMUX_n7), .b ({key_s2[116], key_s1[116], key_s0[116]}), .a ({key_s2[52], key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_2102, new_AGEMA_signal_2101, SelectedKey[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_53_U1 ( .s (selects[0]), .b ({key_s2[117], key_s1[117], key_s0[117]}), .a ({key_s2[53], key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_1538, new_AGEMA_signal_1537, SelectedKey[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_54_U1 ( .s (selects[0]), .b ({key_s2[118], key_s1[118], key_s0[118]}), .a ({key_s2[54], key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, SelectedKey[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_55_U1 ( .s (KeyMUX_n7), .b ({key_s2[119], key_s1[119], key_s0[119]}), .a ({key_s2[55], key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_2108, new_AGEMA_signal_2107, SelectedKey[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_56_U1 ( .s (selects[0]), .b ({key_s2[120], key_s1[120], key_s0[120]}), .a ({key_s2[56], key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, SelectedKey[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_57_U1 ( .s (KeyMUX_n7), .b ({key_s2[121], key_s1[121], key_s0[121]}), .a ({key_s2[57], key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, SelectedKey[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_58_U1 ( .s (KeyMUX_n7), .b ({key_s2[122], key_s1[122], key_s0[122]}), .a ({key_s2[58], key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_2120, new_AGEMA_signal_2119, SelectedKey[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_59_U1 ( .s (selects[0]), .b ({key_s2[123], key_s1[123], key_s0[123]}), .a ({key_s2[59], key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, SelectedKey[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_60_U1 ( .s (KeyMUX_n7), .b ({key_s2[124], key_s1[124], key_s0[124]}), .a ({key_s2[60], key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, SelectedKey[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_61_U1 ( .s (KeyMUX_n7), .b ({key_s2[125], key_s1[125], key_s0[125]}), .a ({key_s2[61], key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_2132, new_AGEMA_signal_2131, SelectedKey[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_62_U1 ( .s (selects[0]), .b ({key_s2[126], key_s1[126], key_s0[126]}), .a ({key_s2[62], key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, SelectedKey[62]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyMUX_MUXInst_63_U1 ( .s (KeyMUX_n7), .b ({key_s2[127], key_s1[127], key_s0[127]}), .a ({key_s2[63], key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_2138, new_AGEMA_signal_2137, SelectedKey[63]}) ) ;
    MUX2_X1 FSMMUX_MUXInst_0_U1 ( .S (rst), .A (FSMReg[0]), .B (1'b1), .Z (RoundConstant_0) ) ;
    MUX2_X1 FSMMUX_MUXInst_1_U1 ( .S (rst), .A (FSMReg[1]), .B (1'b0), .Z (FSMUpdate[0]) ) ;
    MUX2_X1 FSMMUX_MUXInst_2_U1 ( .S (rst), .A (FSMReg[2]), .B (1'b0), .Z (FSMUpdate[1]) ) ;
    MUX2_X1 FSMMUX_MUXInst_3_U1 ( .S (rst), .A (FSMReg[3]), .B (1'b1), .Z (RoundConstant_4_) ) ;
    MUX2_X1 FSMMUX_MUXInst_4_U1 ( .S (rst), .A (FSMReg[4]), .B (1'b0), .Z (FSMUpdate[3]) ) ;
    MUX2_X1 FSMMUX_MUXInst_5_U1 ( .S (rst), .A (FSMReg[5]), .B (1'b0), .Z (FSMUpdate[4]) ) ;
    MUX2_X1 FSMMUX_MUXInst_6_U1 ( .S (rst), .A (FSMReg[6]), .B (1'b0), .Z (FSMUpdate[5]) ) ;
    XOR2_X1 FSMUpdateInst_U2 ( .A (RoundConstant_4_), .B (FSMUpdate[3]), .Z (FSMUpdate[6]) ) ;
    XOR2_X1 FSMUpdateInst_U1 ( .A (FSMUpdate[0]), .B (RoundConstant_0), .Z (FSMUpdate[2]) ) ;
    AND2_X1 FSMSignalsInst_U6 ( .A1 (FSMUpdate[5]), .A2 (FSMSignalsInst_n5), .ZN (done_internal) ) ;
    NOR2_X1 FSMSignalsInst_U5 ( .A1 (FSMSignalsInst_n4), .A2 (FSMSignalsInst_n3), .ZN (FSMSignalsInst_n5) ) ;
    NAND2_X1 FSMSignalsInst_U4 ( .A1 (FSMSignalsInst_n2), .A2 (FSMSignalsInst_n1), .ZN (FSMSignalsInst_n3) ) ;
    NOR2_X1 FSMSignalsInst_U3 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdate[4]), .ZN (FSMSignalsInst_n1) ) ;
    NOR2_X1 FSMSignalsInst_U2 ( .A1 (FSMUpdate[0]), .A2 (RoundConstant_4_), .ZN (FSMSignalsInst_n2) ) ;
    NAND2_X1 FSMSignalsInst_U1 ( .A1 (RoundConstant_0), .A2 (FSMUpdate[1]), .ZN (FSMSignalsInst_n4) ) ;
    MUX2_X1 selectsMUX_MUXInst_0_U1 ( .S (rst), .A (selectsReg[0]), .B (1'b0), .Z (selects[0]) ) ;
    MUX2_X1 selectsMUX_MUXInst_1_U1 ( .S (rst), .A (selectsReg[1]), .B (1'b0), .Z (selects[1]) ) ;
    XNOR2_X1 selectsUpdateInst_U3 ( .A (selectsUpdateInst_n3), .B (selects[1]), .ZN (selectsNext[1]) ) ;
    XNOR2_X1 selectsUpdateInst_U2 ( .A (selects[0]), .B (1'b0), .ZN (selectsUpdateInst_n3) ) ;
    INV_X1 selectsUpdateInst_U1 ( .A (selects[0]), .ZN (selectsNext[0]) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_819 ( .C (clk), .D (ciphertext_s0[61]), .Q (new_AGEMA_signal_3595) ) ;
    buf_clk new_AGEMA_reg_buffer_821 ( .C (clk), .D (ciphertext_s1[61]), .Q (new_AGEMA_signal_3597) ) ;
    buf_clk new_AGEMA_reg_buffer_823 ( .C (clk), .D (ciphertext_s2[61]), .Q (new_AGEMA_signal_3599) ) ;
    buf_clk new_AGEMA_reg_buffer_825 ( .C (clk), .D (SubCellInst_SboxInst_0_n9), .Q (new_AGEMA_signal_3601) ) ;
    buf_clk new_AGEMA_reg_buffer_827 ( .C (clk), .D (new_AGEMA_signal_1033), .Q (new_AGEMA_signal_3603) ) ;
    buf_clk new_AGEMA_reg_buffer_829 ( .C (clk), .D (new_AGEMA_signal_1034), .Q (new_AGEMA_signal_3605) ) ;
    buf_clk new_AGEMA_reg_buffer_831 ( .C (clk), .D (ciphertext_s0[60]), .Q (new_AGEMA_signal_3607) ) ;
    buf_clk new_AGEMA_reg_buffer_833 ( .C (clk), .D (ciphertext_s1[60]), .Q (new_AGEMA_signal_3609) ) ;
    buf_clk new_AGEMA_reg_buffer_835 ( .C (clk), .D (ciphertext_s2[60]), .Q (new_AGEMA_signal_3611) ) ;
    buf_clk new_AGEMA_reg_buffer_837 ( .C (clk), .D (SubCellInst_SboxInst_0_n7), .Q (new_AGEMA_signal_3613) ) ;
    buf_clk new_AGEMA_reg_buffer_839 ( .C (clk), .D (new_AGEMA_signal_1029), .Q (new_AGEMA_signal_3615) ) ;
    buf_clk new_AGEMA_reg_buffer_841 ( .C (clk), .D (new_AGEMA_signal_1030), .Q (new_AGEMA_signal_3617) ) ;
    buf_clk new_AGEMA_reg_buffer_843 ( .C (clk), .D (ciphertext_s0[49]), .Q (new_AGEMA_signal_3619) ) ;
    buf_clk new_AGEMA_reg_buffer_845 ( .C (clk), .D (ciphertext_s1[49]), .Q (new_AGEMA_signal_3621) ) ;
    buf_clk new_AGEMA_reg_buffer_847 ( .C (clk), .D (ciphertext_s2[49]), .Q (new_AGEMA_signal_3623) ) ;
    buf_clk new_AGEMA_reg_buffer_849 ( .C (clk), .D (SubCellInst_SboxInst_1_n9), .Q (new_AGEMA_signal_3625) ) ;
    buf_clk new_AGEMA_reg_buffer_851 ( .C (clk), .D (new_AGEMA_signal_1049), .Q (new_AGEMA_signal_3627) ) ;
    buf_clk new_AGEMA_reg_buffer_853 ( .C (clk), .D (new_AGEMA_signal_1050), .Q (new_AGEMA_signal_3629) ) ;
    buf_clk new_AGEMA_reg_buffer_855 ( .C (clk), .D (ciphertext_s0[48]), .Q (new_AGEMA_signal_3631) ) ;
    buf_clk new_AGEMA_reg_buffer_857 ( .C (clk), .D (ciphertext_s1[48]), .Q (new_AGEMA_signal_3633) ) ;
    buf_clk new_AGEMA_reg_buffer_859 ( .C (clk), .D (ciphertext_s2[48]), .Q (new_AGEMA_signal_3635) ) ;
    buf_clk new_AGEMA_reg_buffer_861 ( .C (clk), .D (SubCellInst_SboxInst_1_n7), .Q (new_AGEMA_signal_3637) ) ;
    buf_clk new_AGEMA_reg_buffer_863 ( .C (clk), .D (new_AGEMA_signal_1045), .Q (new_AGEMA_signal_3639) ) ;
    buf_clk new_AGEMA_reg_buffer_865 ( .C (clk), .D (new_AGEMA_signal_1046), .Q (new_AGEMA_signal_3641) ) ;
    buf_clk new_AGEMA_reg_buffer_867 ( .C (clk), .D (ciphertext_s0[53]), .Q (new_AGEMA_signal_3643) ) ;
    buf_clk new_AGEMA_reg_buffer_869 ( .C (clk), .D (ciphertext_s1[53]), .Q (new_AGEMA_signal_3645) ) ;
    buf_clk new_AGEMA_reg_buffer_871 ( .C (clk), .D (ciphertext_s2[53]), .Q (new_AGEMA_signal_3647) ) ;
    buf_clk new_AGEMA_reg_buffer_873 ( .C (clk), .D (SubCellInst_SboxInst_2_n9), .Q (new_AGEMA_signal_3649) ) ;
    buf_clk new_AGEMA_reg_buffer_875 ( .C (clk), .D (new_AGEMA_signal_1065), .Q (new_AGEMA_signal_3651) ) ;
    buf_clk new_AGEMA_reg_buffer_877 ( .C (clk), .D (new_AGEMA_signal_1066), .Q (new_AGEMA_signal_3653) ) ;
    buf_clk new_AGEMA_reg_buffer_879 ( .C (clk), .D (ciphertext_s0[52]), .Q (new_AGEMA_signal_3655) ) ;
    buf_clk new_AGEMA_reg_buffer_881 ( .C (clk), .D (ciphertext_s1[52]), .Q (new_AGEMA_signal_3657) ) ;
    buf_clk new_AGEMA_reg_buffer_883 ( .C (clk), .D (ciphertext_s2[52]), .Q (new_AGEMA_signal_3659) ) ;
    buf_clk new_AGEMA_reg_buffer_885 ( .C (clk), .D (SubCellInst_SboxInst_2_n7), .Q (new_AGEMA_signal_3661) ) ;
    buf_clk new_AGEMA_reg_buffer_887 ( .C (clk), .D (new_AGEMA_signal_1061), .Q (new_AGEMA_signal_3663) ) ;
    buf_clk new_AGEMA_reg_buffer_889 ( .C (clk), .D (new_AGEMA_signal_1062), .Q (new_AGEMA_signal_3665) ) ;
    buf_clk new_AGEMA_reg_buffer_891 ( .C (clk), .D (ciphertext_s0[57]), .Q (new_AGEMA_signal_3667) ) ;
    buf_clk new_AGEMA_reg_buffer_893 ( .C (clk), .D (ciphertext_s1[57]), .Q (new_AGEMA_signal_3669) ) ;
    buf_clk new_AGEMA_reg_buffer_895 ( .C (clk), .D (ciphertext_s2[57]), .Q (new_AGEMA_signal_3671) ) ;
    buf_clk new_AGEMA_reg_buffer_897 ( .C (clk), .D (SubCellInst_SboxInst_3_n9), .Q (new_AGEMA_signal_3673) ) ;
    buf_clk new_AGEMA_reg_buffer_899 ( .C (clk), .D (new_AGEMA_signal_1081), .Q (new_AGEMA_signal_3675) ) ;
    buf_clk new_AGEMA_reg_buffer_901 ( .C (clk), .D (new_AGEMA_signal_1082), .Q (new_AGEMA_signal_3677) ) ;
    buf_clk new_AGEMA_reg_buffer_903 ( .C (clk), .D (ciphertext_s0[56]), .Q (new_AGEMA_signal_3679) ) ;
    buf_clk new_AGEMA_reg_buffer_905 ( .C (clk), .D (ciphertext_s1[56]), .Q (new_AGEMA_signal_3681) ) ;
    buf_clk new_AGEMA_reg_buffer_907 ( .C (clk), .D (ciphertext_s2[56]), .Q (new_AGEMA_signal_3683) ) ;
    buf_clk new_AGEMA_reg_buffer_909 ( .C (clk), .D (SubCellInst_SboxInst_3_n7), .Q (new_AGEMA_signal_3685) ) ;
    buf_clk new_AGEMA_reg_buffer_911 ( .C (clk), .D (new_AGEMA_signal_1077), .Q (new_AGEMA_signal_3687) ) ;
    buf_clk new_AGEMA_reg_buffer_913 ( .C (clk), .D (new_AGEMA_signal_1078), .Q (new_AGEMA_signal_3689) ) ;
    buf_clk new_AGEMA_reg_buffer_915 ( .C (clk), .D (ciphertext_s0[33]), .Q (new_AGEMA_signal_3691) ) ;
    buf_clk new_AGEMA_reg_buffer_917 ( .C (clk), .D (ciphertext_s1[33]), .Q (new_AGEMA_signal_3693) ) ;
    buf_clk new_AGEMA_reg_buffer_919 ( .C (clk), .D (ciphertext_s2[33]), .Q (new_AGEMA_signal_3695) ) ;
    buf_clk new_AGEMA_reg_buffer_921 ( .C (clk), .D (SubCellInst_SboxInst_4_n9), .Q (new_AGEMA_signal_3697) ) ;
    buf_clk new_AGEMA_reg_buffer_923 ( .C (clk), .D (new_AGEMA_signal_1097), .Q (new_AGEMA_signal_3699) ) ;
    buf_clk new_AGEMA_reg_buffer_925 ( .C (clk), .D (new_AGEMA_signal_1098), .Q (new_AGEMA_signal_3701) ) ;
    buf_clk new_AGEMA_reg_buffer_927 ( .C (clk), .D (ciphertext_s0[32]), .Q (new_AGEMA_signal_3703) ) ;
    buf_clk new_AGEMA_reg_buffer_929 ( .C (clk), .D (ciphertext_s1[32]), .Q (new_AGEMA_signal_3705) ) ;
    buf_clk new_AGEMA_reg_buffer_931 ( .C (clk), .D (ciphertext_s2[32]), .Q (new_AGEMA_signal_3707) ) ;
    buf_clk new_AGEMA_reg_buffer_933 ( .C (clk), .D (SubCellInst_SboxInst_4_n7), .Q (new_AGEMA_signal_3709) ) ;
    buf_clk new_AGEMA_reg_buffer_935 ( .C (clk), .D (new_AGEMA_signal_1093), .Q (new_AGEMA_signal_3711) ) ;
    buf_clk new_AGEMA_reg_buffer_937 ( .C (clk), .D (new_AGEMA_signal_1094), .Q (new_AGEMA_signal_3713) ) ;
    buf_clk new_AGEMA_reg_buffer_939 ( .C (clk), .D (ciphertext_s0[45]), .Q (new_AGEMA_signal_3715) ) ;
    buf_clk new_AGEMA_reg_buffer_941 ( .C (clk), .D (ciphertext_s1[45]), .Q (new_AGEMA_signal_3717) ) ;
    buf_clk new_AGEMA_reg_buffer_943 ( .C (clk), .D (ciphertext_s2[45]), .Q (new_AGEMA_signal_3719) ) ;
    buf_clk new_AGEMA_reg_buffer_945 ( .C (clk), .D (SubCellInst_SboxInst_5_n9), .Q (new_AGEMA_signal_3721) ) ;
    buf_clk new_AGEMA_reg_buffer_947 ( .C (clk), .D (new_AGEMA_signal_1113), .Q (new_AGEMA_signal_3723) ) ;
    buf_clk new_AGEMA_reg_buffer_949 ( .C (clk), .D (new_AGEMA_signal_1114), .Q (new_AGEMA_signal_3725) ) ;
    buf_clk new_AGEMA_reg_buffer_951 ( .C (clk), .D (ciphertext_s0[44]), .Q (new_AGEMA_signal_3727) ) ;
    buf_clk new_AGEMA_reg_buffer_953 ( .C (clk), .D (ciphertext_s1[44]), .Q (new_AGEMA_signal_3729) ) ;
    buf_clk new_AGEMA_reg_buffer_955 ( .C (clk), .D (ciphertext_s2[44]), .Q (new_AGEMA_signal_3731) ) ;
    buf_clk new_AGEMA_reg_buffer_957 ( .C (clk), .D (SubCellInst_SboxInst_5_n7), .Q (new_AGEMA_signal_3733) ) ;
    buf_clk new_AGEMA_reg_buffer_959 ( .C (clk), .D (new_AGEMA_signal_1109), .Q (new_AGEMA_signal_3735) ) ;
    buf_clk new_AGEMA_reg_buffer_961 ( .C (clk), .D (new_AGEMA_signal_1110), .Q (new_AGEMA_signal_3737) ) ;
    buf_clk new_AGEMA_reg_buffer_963 ( .C (clk), .D (ciphertext_s0[41]), .Q (new_AGEMA_signal_3739) ) ;
    buf_clk new_AGEMA_reg_buffer_965 ( .C (clk), .D (ciphertext_s1[41]), .Q (new_AGEMA_signal_3741) ) ;
    buf_clk new_AGEMA_reg_buffer_967 ( .C (clk), .D (ciphertext_s2[41]), .Q (new_AGEMA_signal_3743) ) ;
    buf_clk new_AGEMA_reg_buffer_969 ( .C (clk), .D (SubCellInst_SboxInst_6_n9), .Q (new_AGEMA_signal_3745) ) ;
    buf_clk new_AGEMA_reg_buffer_971 ( .C (clk), .D (new_AGEMA_signal_1129), .Q (new_AGEMA_signal_3747) ) ;
    buf_clk new_AGEMA_reg_buffer_973 ( .C (clk), .D (new_AGEMA_signal_1130), .Q (new_AGEMA_signal_3749) ) ;
    buf_clk new_AGEMA_reg_buffer_975 ( .C (clk), .D (ciphertext_s0[40]), .Q (new_AGEMA_signal_3751) ) ;
    buf_clk new_AGEMA_reg_buffer_977 ( .C (clk), .D (ciphertext_s1[40]), .Q (new_AGEMA_signal_3753) ) ;
    buf_clk new_AGEMA_reg_buffer_979 ( .C (clk), .D (ciphertext_s2[40]), .Q (new_AGEMA_signal_3755) ) ;
    buf_clk new_AGEMA_reg_buffer_981 ( .C (clk), .D (SubCellInst_SboxInst_6_n7), .Q (new_AGEMA_signal_3757) ) ;
    buf_clk new_AGEMA_reg_buffer_983 ( .C (clk), .D (new_AGEMA_signal_1125), .Q (new_AGEMA_signal_3759) ) ;
    buf_clk new_AGEMA_reg_buffer_985 ( .C (clk), .D (new_AGEMA_signal_1126), .Q (new_AGEMA_signal_3761) ) ;
    buf_clk new_AGEMA_reg_buffer_987 ( .C (clk), .D (ciphertext_s0[37]), .Q (new_AGEMA_signal_3763) ) ;
    buf_clk new_AGEMA_reg_buffer_989 ( .C (clk), .D (ciphertext_s1[37]), .Q (new_AGEMA_signal_3765) ) ;
    buf_clk new_AGEMA_reg_buffer_991 ( .C (clk), .D (ciphertext_s2[37]), .Q (new_AGEMA_signal_3767) ) ;
    buf_clk new_AGEMA_reg_buffer_993 ( .C (clk), .D (SubCellInst_SboxInst_7_n9), .Q (new_AGEMA_signal_3769) ) ;
    buf_clk new_AGEMA_reg_buffer_995 ( .C (clk), .D (new_AGEMA_signal_1145), .Q (new_AGEMA_signal_3771) ) ;
    buf_clk new_AGEMA_reg_buffer_997 ( .C (clk), .D (new_AGEMA_signal_1146), .Q (new_AGEMA_signal_3773) ) ;
    buf_clk new_AGEMA_reg_buffer_999 ( .C (clk), .D (ciphertext_s0[36]), .Q (new_AGEMA_signal_3775) ) ;
    buf_clk new_AGEMA_reg_buffer_1001 ( .C (clk), .D (ciphertext_s1[36]), .Q (new_AGEMA_signal_3777) ) ;
    buf_clk new_AGEMA_reg_buffer_1003 ( .C (clk), .D (ciphertext_s2[36]), .Q (new_AGEMA_signal_3779) ) ;
    buf_clk new_AGEMA_reg_buffer_1005 ( .C (clk), .D (SubCellInst_SboxInst_7_n7), .Q (new_AGEMA_signal_3781) ) ;
    buf_clk new_AGEMA_reg_buffer_1007 ( .C (clk), .D (new_AGEMA_signal_1141), .Q (new_AGEMA_signal_3783) ) ;
    buf_clk new_AGEMA_reg_buffer_1009 ( .C (clk), .D (new_AGEMA_signal_1142), .Q (new_AGEMA_signal_3785) ) ;
    buf_clk new_AGEMA_reg_buffer_1011 ( .C (clk), .D (ciphertext_s0[17]), .Q (new_AGEMA_signal_3787) ) ;
    buf_clk new_AGEMA_reg_buffer_1013 ( .C (clk), .D (ciphertext_s1[17]), .Q (new_AGEMA_signal_3789) ) ;
    buf_clk new_AGEMA_reg_buffer_1015 ( .C (clk), .D (ciphertext_s2[17]), .Q (new_AGEMA_signal_3791) ) ;
    buf_clk new_AGEMA_reg_buffer_1017 ( .C (clk), .D (SubCellInst_SboxInst_8_n9), .Q (new_AGEMA_signal_3793) ) ;
    buf_clk new_AGEMA_reg_buffer_1019 ( .C (clk), .D (new_AGEMA_signal_1161), .Q (new_AGEMA_signal_3795) ) ;
    buf_clk new_AGEMA_reg_buffer_1021 ( .C (clk), .D (new_AGEMA_signal_1162), .Q (new_AGEMA_signal_3797) ) ;
    buf_clk new_AGEMA_reg_buffer_1023 ( .C (clk), .D (ciphertext_s0[16]), .Q (new_AGEMA_signal_3799) ) ;
    buf_clk new_AGEMA_reg_buffer_1025 ( .C (clk), .D (ciphertext_s1[16]), .Q (new_AGEMA_signal_3801) ) ;
    buf_clk new_AGEMA_reg_buffer_1027 ( .C (clk), .D (ciphertext_s2[16]), .Q (new_AGEMA_signal_3803) ) ;
    buf_clk new_AGEMA_reg_buffer_1029 ( .C (clk), .D (SubCellInst_SboxInst_8_n7), .Q (new_AGEMA_signal_3805) ) ;
    buf_clk new_AGEMA_reg_buffer_1031 ( .C (clk), .D (new_AGEMA_signal_1157), .Q (new_AGEMA_signal_3807) ) ;
    buf_clk new_AGEMA_reg_buffer_1033 ( .C (clk), .D (new_AGEMA_signal_1158), .Q (new_AGEMA_signal_3809) ) ;
    buf_clk new_AGEMA_reg_buffer_1035 ( .C (clk), .D (ciphertext_s0[29]), .Q (new_AGEMA_signal_3811) ) ;
    buf_clk new_AGEMA_reg_buffer_1037 ( .C (clk), .D (ciphertext_s1[29]), .Q (new_AGEMA_signal_3813) ) ;
    buf_clk new_AGEMA_reg_buffer_1039 ( .C (clk), .D (ciphertext_s2[29]), .Q (new_AGEMA_signal_3815) ) ;
    buf_clk new_AGEMA_reg_buffer_1041 ( .C (clk), .D (SubCellInst_SboxInst_9_n9), .Q (new_AGEMA_signal_3817) ) ;
    buf_clk new_AGEMA_reg_buffer_1043 ( .C (clk), .D (new_AGEMA_signal_1177), .Q (new_AGEMA_signal_3819) ) ;
    buf_clk new_AGEMA_reg_buffer_1045 ( .C (clk), .D (new_AGEMA_signal_1178), .Q (new_AGEMA_signal_3821) ) ;
    buf_clk new_AGEMA_reg_buffer_1047 ( .C (clk), .D (ciphertext_s0[28]), .Q (new_AGEMA_signal_3823) ) ;
    buf_clk new_AGEMA_reg_buffer_1049 ( .C (clk), .D (ciphertext_s1[28]), .Q (new_AGEMA_signal_3825) ) ;
    buf_clk new_AGEMA_reg_buffer_1051 ( .C (clk), .D (ciphertext_s2[28]), .Q (new_AGEMA_signal_3827) ) ;
    buf_clk new_AGEMA_reg_buffer_1053 ( .C (clk), .D (SubCellInst_SboxInst_9_n7), .Q (new_AGEMA_signal_3829) ) ;
    buf_clk new_AGEMA_reg_buffer_1055 ( .C (clk), .D (new_AGEMA_signal_1173), .Q (new_AGEMA_signal_3831) ) ;
    buf_clk new_AGEMA_reg_buffer_1057 ( .C (clk), .D (new_AGEMA_signal_1174), .Q (new_AGEMA_signal_3833) ) ;
    buf_clk new_AGEMA_reg_buffer_1059 ( .C (clk), .D (ciphertext_s0[25]), .Q (new_AGEMA_signal_3835) ) ;
    buf_clk new_AGEMA_reg_buffer_1061 ( .C (clk), .D (ciphertext_s1[25]), .Q (new_AGEMA_signal_3837) ) ;
    buf_clk new_AGEMA_reg_buffer_1063 ( .C (clk), .D (ciphertext_s2[25]), .Q (new_AGEMA_signal_3839) ) ;
    buf_clk new_AGEMA_reg_buffer_1065 ( .C (clk), .D (SubCellInst_SboxInst_10_n9), .Q (new_AGEMA_signal_3841) ) ;
    buf_clk new_AGEMA_reg_buffer_1067 ( .C (clk), .D (new_AGEMA_signal_1193), .Q (new_AGEMA_signal_3843) ) ;
    buf_clk new_AGEMA_reg_buffer_1069 ( .C (clk), .D (new_AGEMA_signal_1194), .Q (new_AGEMA_signal_3845) ) ;
    buf_clk new_AGEMA_reg_buffer_1071 ( .C (clk), .D (ciphertext_s0[24]), .Q (new_AGEMA_signal_3847) ) ;
    buf_clk new_AGEMA_reg_buffer_1073 ( .C (clk), .D (ciphertext_s1[24]), .Q (new_AGEMA_signal_3849) ) ;
    buf_clk new_AGEMA_reg_buffer_1075 ( .C (clk), .D (ciphertext_s2[24]), .Q (new_AGEMA_signal_3851) ) ;
    buf_clk new_AGEMA_reg_buffer_1077 ( .C (clk), .D (SubCellInst_SboxInst_10_n7), .Q (new_AGEMA_signal_3853) ) ;
    buf_clk new_AGEMA_reg_buffer_1079 ( .C (clk), .D (new_AGEMA_signal_1189), .Q (new_AGEMA_signal_3855) ) ;
    buf_clk new_AGEMA_reg_buffer_1081 ( .C (clk), .D (new_AGEMA_signal_1190), .Q (new_AGEMA_signal_3857) ) ;
    buf_clk new_AGEMA_reg_buffer_1083 ( .C (clk), .D (ciphertext_s0[21]), .Q (new_AGEMA_signal_3859) ) ;
    buf_clk new_AGEMA_reg_buffer_1085 ( .C (clk), .D (ciphertext_s1[21]), .Q (new_AGEMA_signal_3861) ) ;
    buf_clk new_AGEMA_reg_buffer_1087 ( .C (clk), .D (ciphertext_s2[21]), .Q (new_AGEMA_signal_3863) ) ;
    buf_clk new_AGEMA_reg_buffer_1089 ( .C (clk), .D (SubCellInst_SboxInst_11_n9), .Q (new_AGEMA_signal_3865) ) ;
    buf_clk new_AGEMA_reg_buffer_1091 ( .C (clk), .D (new_AGEMA_signal_1209), .Q (new_AGEMA_signal_3867) ) ;
    buf_clk new_AGEMA_reg_buffer_1093 ( .C (clk), .D (new_AGEMA_signal_1210), .Q (new_AGEMA_signal_3869) ) ;
    buf_clk new_AGEMA_reg_buffer_1095 ( .C (clk), .D (ciphertext_s0[20]), .Q (new_AGEMA_signal_3871) ) ;
    buf_clk new_AGEMA_reg_buffer_1097 ( .C (clk), .D (ciphertext_s1[20]), .Q (new_AGEMA_signal_3873) ) ;
    buf_clk new_AGEMA_reg_buffer_1099 ( .C (clk), .D (ciphertext_s2[20]), .Q (new_AGEMA_signal_3875) ) ;
    buf_clk new_AGEMA_reg_buffer_1101 ( .C (clk), .D (SubCellInst_SboxInst_11_n7), .Q (new_AGEMA_signal_3877) ) ;
    buf_clk new_AGEMA_reg_buffer_1103 ( .C (clk), .D (new_AGEMA_signal_1205), .Q (new_AGEMA_signal_3879) ) ;
    buf_clk new_AGEMA_reg_buffer_1105 ( .C (clk), .D (new_AGEMA_signal_1206), .Q (new_AGEMA_signal_3881) ) ;
    buf_clk new_AGEMA_reg_buffer_1107 ( .C (clk), .D (ciphertext_s0[5]), .Q (new_AGEMA_signal_3883) ) ;
    buf_clk new_AGEMA_reg_buffer_1109 ( .C (clk), .D (ciphertext_s1[5]), .Q (new_AGEMA_signal_3885) ) ;
    buf_clk new_AGEMA_reg_buffer_1111 ( .C (clk), .D (ciphertext_s2[5]), .Q (new_AGEMA_signal_3887) ) ;
    buf_clk new_AGEMA_reg_buffer_1113 ( .C (clk), .D (SubCellInst_SboxInst_12_n9), .Q (new_AGEMA_signal_3889) ) ;
    buf_clk new_AGEMA_reg_buffer_1115 ( .C (clk), .D (new_AGEMA_signal_1225), .Q (new_AGEMA_signal_3891) ) ;
    buf_clk new_AGEMA_reg_buffer_1117 ( .C (clk), .D (new_AGEMA_signal_1226), .Q (new_AGEMA_signal_3893) ) ;
    buf_clk new_AGEMA_reg_buffer_1119 ( .C (clk), .D (ciphertext_s0[4]), .Q (new_AGEMA_signal_3895) ) ;
    buf_clk new_AGEMA_reg_buffer_1121 ( .C (clk), .D (ciphertext_s1[4]), .Q (new_AGEMA_signal_3897) ) ;
    buf_clk new_AGEMA_reg_buffer_1123 ( .C (clk), .D (ciphertext_s2[4]), .Q (new_AGEMA_signal_3899) ) ;
    buf_clk new_AGEMA_reg_buffer_1125 ( .C (clk), .D (SubCellInst_SboxInst_12_n7), .Q (new_AGEMA_signal_3901) ) ;
    buf_clk new_AGEMA_reg_buffer_1127 ( .C (clk), .D (new_AGEMA_signal_1221), .Q (new_AGEMA_signal_3903) ) ;
    buf_clk new_AGEMA_reg_buffer_1129 ( .C (clk), .D (new_AGEMA_signal_1222), .Q (new_AGEMA_signal_3905) ) ;
    buf_clk new_AGEMA_reg_buffer_1131 ( .C (clk), .D (ciphertext_s0[9]), .Q (new_AGEMA_signal_3907) ) ;
    buf_clk new_AGEMA_reg_buffer_1133 ( .C (clk), .D (ciphertext_s1[9]), .Q (new_AGEMA_signal_3909) ) ;
    buf_clk new_AGEMA_reg_buffer_1135 ( .C (clk), .D (ciphertext_s2[9]), .Q (new_AGEMA_signal_3911) ) ;
    buf_clk new_AGEMA_reg_buffer_1137 ( .C (clk), .D (SubCellInst_SboxInst_13_n9), .Q (new_AGEMA_signal_3913) ) ;
    buf_clk new_AGEMA_reg_buffer_1139 ( .C (clk), .D (new_AGEMA_signal_1241), .Q (new_AGEMA_signal_3915) ) ;
    buf_clk new_AGEMA_reg_buffer_1141 ( .C (clk), .D (new_AGEMA_signal_1242), .Q (new_AGEMA_signal_3917) ) ;
    buf_clk new_AGEMA_reg_buffer_1143 ( .C (clk), .D (ciphertext_s0[8]), .Q (new_AGEMA_signal_3919) ) ;
    buf_clk new_AGEMA_reg_buffer_1145 ( .C (clk), .D (ciphertext_s1[8]), .Q (new_AGEMA_signal_3921) ) ;
    buf_clk new_AGEMA_reg_buffer_1147 ( .C (clk), .D (ciphertext_s2[8]), .Q (new_AGEMA_signal_3923) ) ;
    buf_clk new_AGEMA_reg_buffer_1149 ( .C (clk), .D (SubCellInst_SboxInst_13_n7), .Q (new_AGEMA_signal_3925) ) ;
    buf_clk new_AGEMA_reg_buffer_1151 ( .C (clk), .D (new_AGEMA_signal_1237), .Q (new_AGEMA_signal_3927) ) ;
    buf_clk new_AGEMA_reg_buffer_1153 ( .C (clk), .D (new_AGEMA_signal_1238), .Q (new_AGEMA_signal_3929) ) ;
    buf_clk new_AGEMA_reg_buffer_1155 ( .C (clk), .D (ciphertext_s0[13]), .Q (new_AGEMA_signal_3931) ) ;
    buf_clk new_AGEMA_reg_buffer_1157 ( .C (clk), .D (ciphertext_s1[13]), .Q (new_AGEMA_signal_3933) ) ;
    buf_clk new_AGEMA_reg_buffer_1159 ( .C (clk), .D (ciphertext_s2[13]), .Q (new_AGEMA_signal_3935) ) ;
    buf_clk new_AGEMA_reg_buffer_1161 ( .C (clk), .D (SubCellInst_SboxInst_14_n9), .Q (new_AGEMA_signal_3937) ) ;
    buf_clk new_AGEMA_reg_buffer_1163 ( .C (clk), .D (new_AGEMA_signal_1257), .Q (new_AGEMA_signal_3939) ) ;
    buf_clk new_AGEMA_reg_buffer_1165 ( .C (clk), .D (new_AGEMA_signal_1258), .Q (new_AGEMA_signal_3941) ) ;
    buf_clk new_AGEMA_reg_buffer_1167 ( .C (clk), .D (ciphertext_s0[12]), .Q (new_AGEMA_signal_3943) ) ;
    buf_clk new_AGEMA_reg_buffer_1169 ( .C (clk), .D (ciphertext_s1[12]), .Q (new_AGEMA_signal_3945) ) ;
    buf_clk new_AGEMA_reg_buffer_1171 ( .C (clk), .D (ciphertext_s2[12]), .Q (new_AGEMA_signal_3947) ) ;
    buf_clk new_AGEMA_reg_buffer_1173 ( .C (clk), .D (SubCellInst_SboxInst_14_n7), .Q (new_AGEMA_signal_3949) ) ;
    buf_clk new_AGEMA_reg_buffer_1175 ( .C (clk), .D (new_AGEMA_signal_1253), .Q (new_AGEMA_signal_3951) ) ;
    buf_clk new_AGEMA_reg_buffer_1177 ( .C (clk), .D (new_AGEMA_signal_1254), .Q (new_AGEMA_signal_3953) ) ;
    buf_clk new_AGEMA_reg_buffer_1179 ( .C (clk), .D (ciphertext_s0[1]), .Q (new_AGEMA_signal_3955) ) ;
    buf_clk new_AGEMA_reg_buffer_1181 ( .C (clk), .D (ciphertext_s1[1]), .Q (new_AGEMA_signal_3957) ) ;
    buf_clk new_AGEMA_reg_buffer_1183 ( .C (clk), .D (ciphertext_s2[1]), .Q (new_AGEMA_signal_3959) ) ;
    buf_clk new_AGEMA_reg_buffer_1185 ( .C (clk), .D (SubCellInst_SboxInst_15_n9), .Q (new_AGEMA_signal_3961) ) ;
    buf_clk new_AGEMA_reg_buffer_1187 ( .C (clk), .D (new_AGEMA_signal_1273), .Q (new_AGEMA_signal_3963) ) ;
    buf_clk new_AGEMA_reg_buffer_1189 ( .C (clk), .D (new_AGEMA_signal_1274), .Q (new_AGEMA_signal_3965) ) ;
    buf_clk new_AGEMA_reg_buffer_1191 ( .C (clk), .D (ciphertext_s0[0]), .Q (new_AGEMA_signal_3967) ) ;
    buf_clk new_AGEMA_reg_buffer_1193 ( .C (clk), .D (ciphertext_s1[0]), .Q (new_AGEMA_signal_3969) ) ;
    buf_clk new_AGEMA_reg_buffer_1195 ( .C (clk), .D (ciphertext_s2[0]), .Q (new_AGEMA_signal_3971) ) ;
    buf_clk new_AGEMA_reg_buffer_1197 ( .C (clk), .D (SubCellInst_SboxInst_15_n7), .Q (new_AGEMA_signal_3973) ) ;
    buf_clk new_AGEMA_reg_buffer_1199 ( .C (clk), .D (new_AGEMA_signal_1269), .Q (new_AGEMA_signal_3975) ) ;
    buf_clk new_AGEMA_reg_buffer_1201 ( .C (clk), .D (new_AGEMA_signal_1270), .Q (new_AGEMA_signal_3977) ) ;
    buf_clk new_AGEMA_reg_buffer_1203 ( .C (clk), .D (rst), .Q (new_AGEMA_signal_3979) ) ;
    buf_clk new_AGEMA_reg_buffer_1209 ( .C (clk), .D (plaintext_s0[1]), .Q (new_AGEMA_signal_3985) ) ;
    buf_clk new_AGEMA_reg_buffer_1215 ( .C (clk), .D (plaintext_s1[1]), .Q (new_AGEMA_signal_3991) ) ;
    buf_clk new_AGEMA_reg_buffer_1221 ( .C (clk), .D (plaintext_s2[1]), .Q (new_AGEMA_signal_3997) ) ;
    buf_clk new_AGEMA_reg_buffer_1227 ( .C (clk), .D (plaintext_s0[3]), .Q (new_AGEMA_signal_4003) ) ;
    buf_clk new_AGEMA_reg_buffer_1233 ( .C (clk), .D (plaintext_s1[3]), .Q (new_AGEMA_signal_4009) ) ;
    buf_clk new_AGEMA_reg_buffer_1239 ( .C (clk), .D (plaintext_s2[3]), .Q (new_AGEMA_signal_4015) ) ;
    buf_clk new_AGEMA_reg_buffer_1245 ( .C (clk), .D (plaintext_s0[5]), .Q (new_AGEMA_signal_4021) ) ;
    buf_clk new_AGEMA_reg_buffer_1251 ( .C (clk), .D (plaintext_s1[5]), .Q (new_AGEMA_signal_4027) ) ;
    buf_clk new_AGEMA_reg_buffer_1257 ( .C (clk), .D (plaintext_s2[5]), .Q (new_AGEMA_signal_4033) ) ;
    buf_clk new_AGEMA_reg_buffer_1263 ( .C (clk), .D (plaintext_s0[7]), .Q (new_AGEMA_signal_4039) ) ;
    buf_clk new_AGEMA_reg_buffer_1269 ( .C (clk), .D (plaintext_s1[7]), .Q (new_AGEMA_signal_4045) ) ;
    buf_clk new_AGEMA_reg_buffer_1275 ( .C (clk), .D (plaintext_s2[7]), .Q (new_AGEMA_signal_4051) ) ;
    buf_clk new_AGEMA_reg_buffer_1281 ( .C (clk), .D (plaintext_s0[9]), .Q (new_AGEMA_signal_4057) ) ;
    buf_clk new_AGEMA_reg_buffer_1287 ( .C (clk), .D (plaintext_s1[9]), .Q (new_AGEMA_signal_4063) ) ;
    buf_clk new_AGEMA_reg_buffer_1293 ( .C (clk), .D (plaintext_s2[9]), .Q (new_AGEMA_signal_4069) ) ;
    buf_clk new_AGEMA_reg_buffer_1299 ( .C (clk), .D (plaintext_s0[11]), .Q (new_AGEMA_signal_4075) ) ;
    buf_clk new_AGEMA_reg_buffer_1305 ( .C (clk), .D (plaintext_s1[11]), .Q (new_AGEMA_signal_4081) ) ;
    buf_clk new_AGEMA_reg_buffer_1311 ( .C (clk), .D (plaintext_s2[11]), .Q (new_AGEMA_signal_4087) ) ;
    buf_clk new_AGEMA_reg_buffer_1317 ( .C (clk), .D (plaintext_s0[13]), .Q (new_AGEMA_signal_4093) ) ;
    buf_clk new_AGEMA_reg_buffer_1323 ( .C (clk), .D (plaintext_s1[13]), .Q (new_AGEMA_signal_4099) ) ;
    buf_clk new_AGEMA_reg_buffer_1329 ( .C (clk), .D (plaintext_s2[13]), .Q (new_AGEMA_signal_4105) ) ;
    buf_clk new_AGEMA_reg_buffer_1335 ( .C (clk), .D (plaintext_s0[15]), .Q (new_AGEMA_signal_4111) ) ;
    buf_clk new_AGEMA_reg_buffer_1341 ( .C (clk), .D (plaintext_s1[15]), .Q (new_AGEMA_signal_4117) ) ;
    buf_clk new_AGEMA_reg_buffer_1347 ( .C (clk), .D (plaintext_s2[15]), .Q (new_AGEMA_signal_4123) ) ;
    buf_clk new_AGEMA_reg_buffer_1353 ( .C (clk), .D (plaintext_s0[17]), .Q (new_AGEMA_signal_4129) ) ;
    buf_clk new_AGEMA_reg_buffer_1359 ( .C (clk), .D (plaintext_s1[17]), .Q (new_AGEMA_signal_4135) ) ;
    buf_clk new_AGEMA_reg_buffer_1365 ( .C (clk), .D (plaintext_s2[17]), .Q (new_AGEMA_signal_4141) ) ;
    buf_clk new_AGEMA_reg_buffer_1371 ( .C (clk), .D (plaintext_s0[19]), .Q (new_AGEMA_signal_4147) ) ;
    buf_clk new_AGEMA_reg_buffer_1377 ( .C (clk), .D (plaintext_s1[19]), .Q (new_AGEMA_signal_4153) ) ;
    buf_clk new_AGEMA_reg_buffer_1383 ( .C (clk), .D (plaintext_s2[19]), .Q (new_AGEMA_signal_4159) ) ;
    buf_clk new_AGEMA_reg_buffer_1389 ( .C (clk), .D (plaintext_s0[21]), .Q (new_AGEMA_signal_4165) ) ;
    buf_clk new_AGEMA_reg_buffer_1395 ( .C (clk), .D (plaintext_s1[21]), .Q (new_AGEMA_signal_4171) ) ;
    buf_clk new_AGEMA_reg_buffer_1401 ( .C (clk), .D (plaintext_s2[21]), .Q (new_AGEMA_signal_4177) ) ;
    buf_clk new_AGEMA_reg_buffer_1407 ( .C (clk), .D (plaintext_s0[23]), .Q (new_AGEMA_signal_4183) ) ;
    buf_clk new_AGEMA_reg_buffer_1413 ( .C (clk), .D (plaintext_s1[23]), .Q (new_AGEMA_signal_4189) ) ;
    buf_clk new_AGEMA_reg_buffer_1419 ( .C (clk), .D (plaintext_s2[23]), .Q (new_AGEMA_signal_4195) ) ;
    buf_clk new_AGEMA_reg_buffer_1425 ( .C (clk), .D (plaintext_s0[25]), .Q (new_AGEMA_signal_4201) ) ;
    buf_clk new_AGEMA_reg_buffer_1431 ( .C (clk), .D (plaintext_s1[25]), .Q (new_AGEMA_signal_4207) ) ;
    buf_clk new_AGEMA_reg_buffer_1437 ( .C (clk), .D (plaintext_s2[25]), .Q (new_AGEMA_signal_4213) ) ;
    buf_clk new_AGEMA_reg_buffer_1443 ( .C (clk), .D (plaintext_s0[27]), .Q (new_AGEMA_signal_4219) ) ;
    buf_clk new_AGEMA_reg_buffer_1449 ( .C (clk), .D (plaintext_s1[27]), .Q (new_AGEMA_signal_4225) ) ;
    buf_clk new_AGEMA_reg_buffer_1455 ( .C (clk), .D (plaintext_s2[27]), .Q (new_AGEMA_signal_4231) ) ;
    buf_clk new_AGEMA_reg_buffer_1461 ( .C (clk), .D (plaintext_s0[29]), .Q (new_AGEMA_signal_4237) ) ;
    buf_clk new_AGEMA_reg_buffer_1467 ( .C (clk), .D (plaintext_s1[29]), .Q (new_AGEMA_signal_4243) ) ;
    buf_clk new_AGEMA_reg_buffer_1473 ( .C (clk), .D (plaintext_s2[29]), .Q (new_AGEMA_signal_4249) ) ;
    buf_clk new_AGEMA_reg_buffer_1479 ( .C (clk), .D (plaintext_s0[31]), .Q (new_AGEMA_signal_4255) ) ;
    buf_clk new_AGEMA_reg_buffer_1485 ( .C (clk), .D (plaintext_s1[31]), .Q (new_AGEMA_signal_4261) ) ;
    buf_clk new_AGEMA_reg_buffer_1491 ( .C (clk), .D (plaintext_s2[31]), .Q (new_AGEMA_signal_4267) ) ;
    buf_clk new_AGEMA_reg_buffer_1497 ( .C (clk), .D (plaintext_s0[33]), .Q (new_AGEMA_signal_4273) ) ;
    buf_clk new_AGEMA_reg_buffer_1503 ( .C (clk), .D (plaintext_s1[33]), .Q (new_AGEMA_signal_4279) ) ;
    buf_clk new_AGEMA_reg_buffer_1509 ( .C (clk), .D (plaintext_s2[33]), .Q (new_AGEMA_signal_4285) ) ;
    buf_clk new_AGEMA_reg_buffer_1515 ( .C (clk), .D (plaintext_s0[35]), .Q (new_AGEMA_signal_4291) ) ;
    buf_clk new_AGEMA_reg_buffer_1521 ( .C (clk), .D (plaintext_s1[35]), .Q (new_AGEMA_signal_4297) ) ;
    buf_clk new_AGEMA_reg_buffer_1527 ( .C (clk), .D (plaintext_s2[35]), .Q (new_AGEMA_signal_4303) ) ;
    buf_clk new_AGEMA_reg_buffer_1533 ( .C (clk), .D (plaintext_s0[37]), .Q (new_AGEMA_signal_4309) ) ;
    buf_clk new_AGEMA_reg_buffer_1539 ( .C (clk), .D (plaintext_s1[37]), .Q (new_AGEMA_signal_4315) ) ;
    buf_clk new_AGEMA_reg_buffer_1545 ( .C (clk), .D (plaintext_s2[37]), .Q (new_AGEMA_signal_4321) ) ;
    buf_clk new_AGEMA_reg_buffer_1551 ( .C (clk), .D (plaintext_s0[39]), .Q (new_AGEMA_signal_4327) ) ;
    buf_clk new_AGEMA_reg_buffer_1557 ( .C (clk), .D (plaintext_s1[39]), .Q (new_AGEMA_signal_4333) ) ;
    buf_clk new_AGEMA_reg_buffer_1563 ( .C (clk), .D (plaintext_s2[39]), .Q (new_AGEMA_signal_4339) ) ;
    buf_clk new_AGEMA_reg_buffer_1569 ( .C (clk), .D (plaintext_s0[41]), .Q (new_AGEMA_signal_4345) ) ;
    buf_clk new_AGEMA_reg_buffer_1575 ( .C (clk), .D (plaintext_s1[41]), .Q (new_AGEMA_signal_4351) ) ;
    buf_clk new_AGEMA_reg_buffer_1581 ( .C (clk), .D (plaintext_s2[41]), .Q (new_AGEMA_signal_4357) ) ;
    buf_clk new_AGEMA_reg_buffer_1587 ( .C (clk), .D (plaintext_s0[43]), .Q (new_AGEMA_signal_4363) ) ;
    buf_clk new_AGEMA_reg_buffer_1593 ( .C (clk), .D (plaintext_s1[43]), .Q (new_AGEMA_signal_4369) ) ;
    buf_clk new_AGEMA_reg_buffer_1599 ( .C (clk), .D (plaintext_s2[43]), .Q (new_AGEMA_signal_4375) ) ;
    buf_clk new_AGEMA_reg_buffer_1605 ( .C (clk), .D (plaintext_s0[45]), .Q (new_AGEMA_signal_4381) ) ;
    buf_clk new_AGEMA_reg_buffer_1611 ( .C (clk), .D (plaintext_s1[45]), .Q (new_AGEMA_signal_4387) ) ;
    buf_clk new_AGEMA_reg_buffer_1617 ( .C (clk), .D (plaintext_s2[45]), .Q (new_AGEMA_signal_4393) ) ;
    buf_clk new_AGEMA_reg_buffer_1623 ( .C (clk), .D (plaintext_s0[47]), .Q (new_AGEMA_signal_4399) ) ;
    buf_clk new_AGEMA_reg_buffer_1629 ( .C (clk), .D (plaintext_s1[47]), .Q (new_AGEMA_signal_4405) ) ;
    buf_clk new_AGEMA_reg_buffer_1635 ( .C (clk), .D (plaintext_s2[47]), .Q (new_AGEMA_signal_4411) ) ;
    buf_clk new_AGEMA_reg_buffer_1641 ( .C (clk), .D (plaintext_s0[49]), .Q (new_AGEMA_signal_4417) ) ;
    buf_clk new_AGEMA_reg_buffer_1647 ( .C (clk), .D (plaintext_s1[49]), .Q (new_AGEMA_signal_4423) ) ;
    buf_clk new_AGEMA_reg_buffer_1653 ( .C (clk), .D (plaintext_s2[49]), .Q (new_AGEMA_signal_4429) ) ;
    buf_clk new_AGEMA_reg_buffer_1659 ( .C (clk), .D (plaintext_s0[51]), .Q (new_AGEMA_signal_4435) ) ;
    buf_clk new_AGEMA_reg_buffer_1665 ( .C (clk), .D (plaintext_s1[51]), .Q (new_AGEMA_signal_4441) ) ;
    buf_clk new_AGEMA_reg_buffer_1671 ( .C (clk), .D (plaintext_s2[51]), .Q (new_AGEMA_signal_4447) ) ;
    buf_clk new_AGEMA_reg_buffer_1677 ( .C (clk), .D (plaintext_s0[53]), .Q (new_AGEMA_signal_4453) ) ;
    buf_clk new_AGEMA_reg_buffer_1683 ( .C (clk), .D (plaintext_s1[53]), .Q (new_AGEMA_signal_4459) ) ;
    buf_clk new_AGEMA_reg_buffer_1689 ( .C (clk), .D (plaintext_s2[53]), .Q (new_AGEMA_signal_4465) ) ;
    buf_clk new_AGEMA_reg_buffer_1695 ( .C (clk), .D (plaintext_s0[55]), .Q (new_AGEMA_signal_4471) ) ;
    buf_clk new_AGEMA_reg_buffer_1701 ( .C (clk), .D (plaintext_s1[55]), .Q (new_AGEMA_signal_4477) ) ;
    buf_clk new_AGEMA_reg_buffer_1707 ( .C (clk), .D (plaintext_s2[55]), .Q (new_AGEMA_signal_4483) ) ;
    buf_clk new_AGEMA_reg_buffer_1713 ( .C (clk), .D (plaintext_s0[57]), .Q (new_AGEMA_signal_4489) ) ;
    buf_clk new_AGEMA_reg_buffer_1719 ( .C (clk), .D (plaintext_s1[57]), .Q (new_AGEMA_signal_4495) ) ;
    buf_clk new_AGEMA_reg_buffer_1725 ( .C (clk), .D (plaintext_s2[57]), .Q (new_AGEMA_signal_4501) ) ;
    buf_clk new_AGEMA_reg_buffer_1731 ( .C (clk), .D (plaintext_s0[59]), .Q (new_AGEMA_signal_4507) ) ;
    buf_clk new_AGEMA_reg_buffer_1737 ( .C (clk), .D (plaintext_s1[59]), .Q (new_AGEMA_signal_4513) ) ;
    buf_clk new_AGEMA_reg_buffer_1743 ( .C (clk), .D (plaintext_s2[59]), .Q (new_AGEMA_signal_4519) ) ;
    buf_clk new_AGEMA_reg_buffer_1749 ( .C (clk), .D (plaintext_s0[61]), .Q (new_AGEMA_signal_4525) ) ;
    buf_clk new_AGEMA_reg_buffer_1755 ( .C (clk), .D (plaintext_s1[61]), .Q (new_AGEMA_signal_4531) ) ;
    buf_clk new_AGEMA_reg_buffer_1761 ( .C (clk), .D (plaintext_s2[61]), .Q (new_AGEMA_signal_4537) ) ;
    buf_clk new_AGEMA_reg_buffer_1767 ( .C (clk), .D (plaintext_s0[63]), .Q (new_AGEMA_signal_4543) ) ;
    buf_clk new_AGEMA_reg_buffer_1773 ( .C (clk), .D (plaintext_s1[63]), .Q (new_AGEMA_signal_4549) ) ;
    buf_clk new_AGEMA_reg_buffer_1779 ( .C (clk), .D (plaintext_s2[63]), .Q (new_AGEMA_signal_4555) ) ;
    buf_clk new_AGEMA_reg_buffer_1785 ( .C (clk), .D (SelectedKey[49]), .Q (new_AGEMA_signal_4561) ) ;
    buf_clk new_AGEMA_reg_buffer_1791 ( .C (clk), .D (new_AGEMA_signal_2083), .Q (new_AGEMA_signal_4567) ) ;
    buf_clk new_AGEMA_reg_buffer_1797 ( .C (clk), .D (new_AGEMA_signal_2084), .Q (new_AGEMA_signal_4573) ) ;
    buf_clk new_AGEMA_reg_buffer_1803 ( .C (clk), .D (SelectedKey[51]), .Q (new_AGEMA_signal_4579) ) ;
    buf_clk new_AGEMA_reg_buffer_1809 ( .C (clk), .D (new_AGEMA_signal_2095), .Q (new_AGEMA_signal_4585) ) ;
    buf_clk new_AGEMA_reg_buffer_1815 ( .C (clk), .D (new_AGEMA_signal_2096), .Q (new_AGEMA_signal_4591) ) ;
    buf_clk new_AGEMA_reg_buffer_1821 ( .C (clk), .D (SelectedKey[53]), .Q (new_AGEMA_signal_4597) ) ;
    buf_clk new_AGEMA_reg_buffer_1827 ( .C (clk), .D (new_AGEMA_signal_1537), .Q (new_AGEMA_signal_4603) ) ;
    buf_clk new_AGEMA_reg_buffer_1833 ( .C (clk), .D (new_AGEMA_signal_1538), .Q (new_AGEMA_signal_4609) ) ;
    buf_clk new_AGEMA_reg_buffer_1839 ( .C (clk), .D (SelectedKey[55]), .Q (new_AGEMA_signal_4615) ) ;
    buf_clk new_AGEMA_reg_buffer_1845 ( .C (clk), .D (new_AGEMA_signal_2107), .Q (new_AGEMA_signal_4621) ) ;
    buf_clk new_AGEMA_reg_buffer_1851 ( .C (clk), .D (new_AGEMA_signal_2108), .Q (new_AGEMA_signal_4627) ) ;
    buf_clk new_AGEMA_reg_buffer_1857 ( .C (clk), .D (SelectedKey[57]), .Q (new_AGEMA_signal_4633) ) ;
    buf_clk new_AGEMA_reg_buffer_1863 ( .C (clk), .D (new_AGEMA_signal_2113), .Q (new_AGEMA_signal_4639) ) ;
    buf_clk new_AGEMA_reg_buffer_1869 ( .C (clk), .D (new_AGEMA_signal_2114), .Q (new_AGEMA_signal_4645) ) ;
    buf_clk new_AGEMA_reg_buffer_1875 ( .C (clk), .D (SelectedKey[59]), .Q (new_AGEMA_signal_4651) ) ;
    buf_clk new_AGEMA_reg_buffer_1881 ( .C (clk), .D (new_AGEMA_signal_1555), .Q (new_AGEMA_signal_4657) ) ;
    buf_clk new_AGEMA_reg_buffer_1887 ( .C (clk), .D (new_AGEMA_signal_1556), .Q (new_AGEMA_signal_4663) ) ;
    buf_clk new_AGEMA_reg_buffer_1893 ( .C (clk), .D (SelectedKey[61]), .Q (new_AGEMA_signal_4669) ) ;
    buf_clk new_AGEMA_reg_buffer_1899 ( .C (clk), .D (new_AGEMA_signal_2131), .Q (new_AGEMA_signal_4675) ) ;
    buf_clk new_AGEMA_reg_buffer_1905 ( .C (clk), .D (new_AGEMA_signal_2132), .Q (new_AGEMA_signal_4681) ) ;
    buf_clk new_AGEMA_reg_buffer_1911 ( .C (clk), .D (SelectedKey[63]), .Q (new_AGEMA_signal_4687) ) ;
    buf_clk new_AGEMA_reg_buffer_1917 ( .C (clk), .D (new_AGEMA_signal_2137), .Q (new_AGEMA_signal_4693) ) ;
    buf_clk new_AGEMA_reg_buffer_1923 ( .C (clk), .D (new_AGEMA_signal_2138), .Q (new_AGEMA_signal_4699) ) ;
    buf_clk new_AGEMA_reg_buffer_1929 ( .C (clk), .D (AddKeyConstXOR_XORInst_0_1_n1), .Q (new_AGEMA_signal_4705) ) ;
    buf_clk new_AGEMA_reg_buffer_1935 ( .C (clk), .D (new_AGEMA_signal_2397), .Q (new_AGEMA_signal_4711) ) ;
    buf_clk new_AGEMA_reg_buffer_1941 ( .C (clk), .D (new_AGEMA_signal_2398), .Q (new_AGEMA_signal_4717) ) ;
    buf_clk new_AGEMA_reg_buffer_1947 ( .C (clk), .D (AddKeyConstXOR_XORInst_0_3_n1), .Q (new_AGEMA_signal_4723) ) ;
    buf_clk new_AGEMA_reg_buffer_1953 ( .C (clk), .D (new_AGEMA_signal_2401), .Q (new_AGEMA_signal_4729) ) ;
    buf_clk new_AGEMA_reg_buffer_1959 ( .C (clk), .D (new_AGEMA_signal_2402), .Q (new_AGEMA_signal_4735) ) ;
    buf_clk new_AGEMA_reg_buffer_1965 ( .C (clk), .D (AddKeyConstXOR_XORInst_1_1_n1), .Q (new_AGEMA_signal_4741) ) ;
    buf_clk new_AGEMA_reg_buffer_1971 ( .C (clk), .D (new_AGEMA_signal_2405), .Q (new_AGEMA_signal_4747) ) ;
    buf_clk new_AGEMA_reg_buffer_1977 ( .C (clk), .D (new_AGEMA_signal_2406), .Q (new_AGEMA_signal_4753) ) ;
    buf_clk new_AGEMA_reg_buffer_1983 ( .C (clk), .D (AddKeyConstXOR_XORInst_1_3_n1), .Q (new_AGEMA_signal_4759) ) ;
    buf_clk new_AGEMA_reg_buffer_1989 ( .C (clk), .D (new_AGEMA_signal_2409), .Q (new_AGEMA_signal_4765) ) ;
    buf_clk new_AGEMA_reg_buffer_1995 ( .C (clk), .D (new_AGEMA_signal_2410), .Q (new_AGEMA_signal_4771) ) ;
    buf_clk new_AGEMA_reg_buffer_2001 ( .C (clk), .D (SelectedKey[1]), .Q (new_AGEMA_signal_4777) ) ;
    buf_clk new_AGEMA_reg_buffer_2007 ( .C (clk), .D (new_AGEMA_signal_1855), .Q (new_AGEMA_signal_4783) ) ;
    buf_clk new_AGEMA_reg_buffer_2013 ( .C (clk), .D (new_AGEMA_signal_1856), .Q (new_AGEMA_signal_4789) ) ;
    buf_clk new_AGEMA_reg_buffer_2019 ( .C (clk), .D (SelectedKey[3]), .Q (new_AGEMA_signal_4795) ) ;
    buf_clk new_AGEMA_reg_buffer_2025 ( .C (clk), .D (new_AGEMA_signal_1861), .Q (new_AGEMA_signal_4801) ) ;
    buf_clk new_AGEMA_reg_buffer_2031 ( .C (clk), .D (new_AGEMA_signal_1862), .Q (new_AGEMA_signal_4807) ) ;
    buf_clk new_AGEMA_reg_buffer_2037 ( .C (clk), .D (SelectedKey[5]), .Q (new_AGEMA_signal_4813) ) ;
    buf_clk new_AGEMA_reg_buffer_2043 ( .C (clk), .D (new_AGEMA_signal_1873), .Q (new_AGEMA_signal_4819) ) ;
    buf_clk new_AGEMA_reg_buffer_2049 ( .C (clk), .D (new_AGEMA_signal_1874), .Q (new_AGEMA_signal_4825) ) ;
    buf_clk new_AGEMA_reg_buffer_2055 ( .C (clk), .D (SelectedKey[7]), .Q (new_AGEMA_signal_4831) ) ;
    buf_clk new_AGEMA_reg_buffer_2061 ( .C (clk), .D (new_AGEMA_signal_1885), .Q (new_AGEMA_signal_4837) ) ;
    buf_clk new_AGEMA_reg_buffer_2067 ( .C (clk), .D (new_AGEMA_signal_1886), .Q (new_AGEMA_signal_4843) ) ;
    buf_clk new_AGEMA_reg_buffer_2073 ( .C (clk), .D (SelectedKey[9]), .Q (new_AGEMA_signal_4849) ) ;
    buf_clk new_AGEMA_reg_buffer_2079 ( .C (clk), .D (new_AGEMA_signal_1897), .Q (new_AGEMA_signal_4855) ) ;
    buf_clk new_AGEMA_reg_buffer_2085 ( .C (clk), .D (new_AGEMA_signal_1898), .Q (new_AGEMA_signal_4861) ) ;
    buf_clk new_AGEMA_reg_buffer_2091 ( .C (clk), .D (SelectedKey[11]), .Q (new_AGEMA_signal_4867) ) ;
    buf_clk new_AGEMA_reg_buffer_2097 ( .C (clk), .D (new_AGEMA_signal_1909), .Q (new_AGEMA_signal_4873) ) ;
    buf_clk new_AGEMA_reg_buffer_2103 ( .C (clk), .D (new_AGEMA_signal_1910), .Q (new_AGEMA_signal_4879) ) ;
    buf_clk new_AGEMA_reg_buffer_2109 ( .C (clk), .D (SelectedKey[13]), .Q (new_AGEMA_signal_4885) ) ;
    buf_clk new_AGEMA_reg_buffer_2115 ( .C (clk), .D (new_AGEMA_signal_1921), .Q (new_AGEMA_signal_4891) ) ;
    buf_clk new_AGEMA_reg_buffer_2121 ( .C (clk), .D (new_AGEMA_signal_1922), .Q (new_AGEMA_signal_4897) ) ;
    buf_clk new_AGEMA_reg_buffer_2127 ( .C (clk), .D (SelectedKey[15]), .Q (new_AGEMA_signal_4903) ) ;
    buf_clk new_AGEMA_reg_buffer_2133 ( .C (clk), .D (new_AGEMA_signal_1933), .Q (new_AGEMA_signal_4909) ) ;
    buf_clk new_AGEMA_reg_buffer_2139 ( .C (clk), .D (new_AGEMA_signal_1934), .Q (new_AGEMA_signal_4915) ) ;
    buf_clk new_AGEMA_reg_buffer_2145 ( .C (clk), .D (SelectedKey[17]), .Q (new_AGEMA_signal_4921) ) ;
    buf_clk new_AGEMA_reg_buffer_2151 ( .C (clk), .D (new_AGEMA_signal_1945), .Q (new_AGEMA_signal_4927) ) ;
    buf_clk new_AGEMA_reg_buffer_2157 ( .C (clk), .D (new_AGEMA_signal_1946), .Q (new_AGEMA_signal_4933) ) ;
    buf_clk new_AGEMA_reg_buffer_2163 ( .C (clk), .D (SelectedKey[19]), .Q (new_AGEMA_signal_4939) ) ;
    buf_clk new_AGEMA_reg_buffer_2169 ( .C (clk), .D (new_AGEMA_signal_1957), .Q (new_AGEMA_signal_4945) ) ;
    buf_clk new_AGEMA_reg_buffer_2175 ( .C (clk), .D (new_AGEMA_signal_1958), .Q (new_AGEMA_signal_4951) ) ;
    buf_clk new_AGEMA_reg_buffer_2181 ( .C (clk), .D (SelectedKey[21]), .Q (new_AGEMA_signal_4957) ) ;
    buf_clk new_AGEMA_reg_buffer_2187 ( .C (clk), .D (new_AGEMA_signal_1969), .Q (new_AGEMA_signal_4963) ) ;
    buf_clk new_AGEMA_reg_buffer_2193 ( .C (clk), .D (new_AGEMA_signal_1970), .Q (new_AGEMA_signal_4969) ) ;
    buf_clk new_AGEMA_reg_buffer_2199 ( .C (clk), .D (SelectedKey[23]), .Q (new_AGEMA_signal_4975) ) ;
    buf_clk new_AGEMA_reg_buffer_2205 ( .C (clk), .D (new_AGEMA_signal_1489), .Q (new_AGEMA_signal_4981) ) ;
    buf_clk new_AGEMA_reg_buffer_2211 ( .C (clk), .D (new_AGEMA_signal_1490), .Q (new_AGEMA_signal_4987) ) ;
    buf_clk new_AGEMA_reg_buffer_2217 ( .C (clk), .D (SelectedKey[25]), .Q (new_AGEMA_signal_4993) ) ;
    buf_clk new_AGEMA_reg_buffer_2223 ( .C (clk), .D (new_AGEMA_signal_1501), .Q (new_AGEMA_signal_4999) ) ;
    buf_clk new_AGEMA_reg_buffer_2229 ( .C (clk), .D (new_AGEMA_signal_1502), .Q (new_AGEMA_signal_5005) ) ;
    buf_clk new_AGEMA_reg_buffer_2235 ( .C (clk), .D (SelectedKey[27]), .Q (new_AGEMA_signal_5011) ) ;
    buf_clk new_AGEMA_reg_buffer_2241 ( .C (clk), .D (new_AGEMA_signal_1513), .Q (new_AGEMA_signal_5017) ) ;
    buf_clk new_AGEMA_reg_buffer_2247 ( .C (clk), .D (new_AGEMA_signal_1514), .Q (new_AGEMA_signal_5023) ) ;
    buf_clk new_AGEMA_reg_buffer_2253 ( .C (clk), .D (SelectedKey[29]), .Q (new_AGEMA_signal_5029) ) ;
    buf_clk new_AGEMA_reg_buffer_2259 ( .C (clk), .D (new_AGEMA_signal_1981), .Q (new_AGEMA_signal_5035) ) ;
    buf_clk new_AGEMA_reg_buffer_2265 ( .C (clk), .D (new_AGEMA_signal_1982), .Q (new_AGEMA_signal_5041) ) ;
    buf_clk new_AGEMA_reg_buffer_2271 ( .C (clk), .D (SelectedKey[31]), .Q (new_AGEMA_signal_5047) ) ;
    buf_clk new_AGEMA_reg_buffer_2277 ( .C (clk), .D (new_AGEMA_signal_1993), .Q (new_AGEMA_signal_5053) ) ;
    buf_clk new_AGEMA_reg_buffer_2283 ( .C (clk), .D (new_AGEMA_signal_1994), .Q (new_AGEMA_signal_5059) ) ;
    buf_clk new_AGEMA_reg_buffer_2289 ( .C (clk), .D (SelectedKey[33]), .Q (new_AGEMA_signal_5065) ) ;
    buf_clk new_AGEMA_reg_buffer_2295 ( .C (clk), .D (new_AGEMA_signal_1519), .Q (new_AGEMA_signal_5071) ) ;
    buf_clk new_AGEMA_reg_buffer_2301 ( .C (clk), .D (new_AGEMA_signal_1520), .Q (new_AGEMA_signal_5077) ) ;
    buf_clk new_AGEMA_reg_buffer_2307 ( .C (clk), .D (SelectedKey[35]), .Q (new_AGEMA_signal_5083) ) ;
    buf_clk new_AGEMA_reg_buffer_2313 ( .C (clk), .D (new_AGEMA_signal_2011), .Q (new_AGEMA_signal_5089) ) ;
    buf_clk new_AGEMA_reg_buffer_2319 ( .C (clk), .D (new_AGEMA_signal_2012), .Q (new_AGEMA_signal_5095) ) ;
    buf_clk new_AGEMA_reg_buffer_2325 ( .C (clk), .D (SelectedKey[37]), .Q (new_AGEMA_signal_5101) ) ;
    buf_clk new_AGEMA_reg_buffer_2331 ( .C (clk), .D (new_AGEMA_signal_2017), .Q (new_AGEMA_signal_5107) ) ;
    buf_clk new_AGEMA_reg_buffer_2337 ( .C (clk), .D (new_AGEMA_signal_2018), .Q (new_AGEMA_signal_5113) ) ;
    buf_clk new_AGEMA_reg_buffer_2343 ( .C (clk), .D (SelectedKey[39]), .Q (new_AGEMA_signal_5119) ) ;
    buf_clk new_AGEMA_reg_buffer_2349 ( .C (clk), .D (new_AGEMA_signal_1531), .Q (new_AGEMA_signal_5125) ) ;
    buf_clk new_AGEMA_reg_buffer_2355 ( .C (clk), .D (new_AGEMA_signal_1532), .Q (new_AGEMA_signal_5131) ) ;
    buf_clk new_AGEMA_reg_buffer_2651 ( .C (clk), .D (plaintext_s0[0]), .Q (new_AGEMA_signal_5427) ) ;
    buf_clk new_AGEMA_reg_buffer_2659 ( .C (clk), .D (plaintext_s1[0]), .Q (new_AGEMA_signal_5435) ) ;
    buf_clk new_AGEMA_reg_buffer_2667 ( .C (clk), .D (plaintext_s2[0]), .Q (new_AGEMA_signal_5443) ) ;
    buf_clk new_AGEMA_reg_buffer_2675 ( .C (clk), .D (plaintext_s0[2]), .Q (new_AGEMA_signal_5451) ) ;
    buf_clk new_AGEMA_reg_buffer_2683 ( .C (clk), .D (plaintext_s1[2]), .Q (new_AGEMA_signal_5459) ) ;
    buf_clk new_AGEMA_reg_buffer_2691 ( .C (clk), .D (plaintext_s2[2]), .Q (new_AGEMA_signal_5467) ) ;
    buf_clk new_AGEMA_reg_buffer_2699 ( .C (clk), .D (plaintext_s0[4]), .Q (new_AGEMA_signal_5475) ) ;
    buf_clk new_AGEMA_reg_buffer_2707 ( .C (clk), .D (plaintext_s1[4]), .Q (new_AGEMA_signal_5483) ) ;
    buf_clk new_AGEMA_reg_buffer_2715 ( .C (clk), .D (plaintext_s2[4]), .Q (new_AGEMA_signal_5491) ) ;
    buf_clk new_AGEMA_reg_buffer_2723 ( .C (clk), .D (plaintext_s0[6]), .Q (new_AGEMA_signal_5499) ) ;
    buf_clk new_AGEMA_reg_buffer_2731 ( .C (clk), .D (plaintext_s1[6]), .Q (new_AGEMA_signal_5507) ) ;
    buf_clk new_AGEMA_reg_buffer_2739 ( .C (clk), .D (plaintext_s2[6]), .Q (new_AGEMA_signal_5515) ) ;
    buf_clk new_AGEMA_reg_buffer_2747 ( .C (clk), .D (plaintext_s0[8]), .Q (new_AGEMA_signal_5523) ) ;
    buf_clk new_AGEMA_reg_buffer_2755 ( .C (clk), .D (plaintext_s1[8]), .Q (new_AGEMA_signal_5531) ) ;
    buf_clk new_AGEMA_reg_buffer_2763 ( .C (clk), .D (plaintext_s2[8]), .Q (new_AGEMA_signal_5539) ) ;
    buf_clk new_AGEMA_reg_buffer_2771 ( .C (clk), .D (plaintext_s0[10]), .Q (new_AGEMA_signal_5547) ) ;
    buf_clk new_AGEMA_reg_buffer_2779 ( .C (clk), .D (plaintext_s1[10]), .Q (new_AGEMA_signal_5555) ) ;
    buf_clk new_AGEMA_reg_buffer_2787 ( .C (clk), .D (plaintext_s2[10]), .Q (new_AGEMA_signal_5563) ) ;
    buf_clk new_AGEMA_reg_buffer_2795 ( .C (clk), .D (plaintext_s0[12]), .Q (new_AGEMA_signal_5571) ) ;
    buf_clk new_AGEMA_reg_buffer_2803 ( .C (clk), .D (plaintext_s1[12]), .Q (new_AGEMA_signal_5579) ) ;
    buf_clk new_AGEMA_reg_buffer_2811 ( .C (clk), .D (plaintext_s2[12]), .Q (new_AGEMA_signal_5587) ) ;
    buf_clk new_AGEMA_reg_buffer_2819 ( .C (clk), .D (plaintext_s0[14]), .Q (new_AGEMA_signal_5595) ) ;
    buf_clk new_AGEMA_reg_buffer_2827 ( .C (clk), .D (plaintext_s1[14]), .Q (new_AGEMA_signal_5603) ) ;
    buf_clk new_AGEMA_reg_buffer_2835 ( .C (clk), .D (plaintext_s2[14]), .Q (new_AGEMA_signal_5611) ) ;
    buf_clk new_AGEMA_reg_buffer_2843 ( .C (clk), .D (plaintext_s0[16]), .Q (new_AGEMA_signal_5619) ) ;
    buf_clk new_AGEMA_reg_buffer_2851 ( .C (clk), .D (plaintext_s1[16]), .Q (new_AGEMA_signal_5627) ) ;
    buf_clk new_AGEMA_reg_buffer_2859 ( .C (clk), .D (plaintext_s2[16]), .Q (new_AGEMA_signal_5635) ) ;
    buf_clk new_AGEMA_reg_buffer_2867 ( .C (clk), .D (plaintext_s0[18]), .Q (new_AGEMA_signal_5643) ) ;
    buf_clk new_AGEMA_reg_buffer_2875 ( .C (clk), .D (plaintext_s1[18]), .Q (new_AGEMA_signal_5651) ) ;
    buf_clk new_AGEMA_reg_buffer_2883 ( .C (clk), .D (plaintext_s2[18]), .Q (new_AGEMA_signal_5659) ) ;
    buf_clk new_AGEMA_reg_buffer_2891 ( .C (clk), .D (plaintext_s0[20]), .Q (new_AGEMA_signal_5667) ) ;
    buf_clk new_AGEMA_reg_buffer_2899 ( .C (clk), .D (plaintext_s1[20]), .Q (new_AGEMA_signal_5675) ) ;
    buf_clk new_AGEMA_reg_buffer_2907 ( .C (clk), .D (plaintext_s2[20]), .Q (new_AGEMA_signal_5683) ) ;
    buf_clk new_AGEMA_reg_buffer_2915 ( .C (clk), .D (plaintext_s0[22]), .Q (new_AGEMA_signal_5691) ) ;
    buf_clk new_AGEMA_reg_buffer_2923 ( .C (clk), .D (plaintext_s1[22]), .Q (new_AGEMA_signal_5699) ) ;
    buf_clk new_AGEMA_reg_buffer_2931 ( .C (clk), .D (plaintext_s2[22]), .Q (new_AGEMA_signal_5707) ) ;
    buf_clk new_AGEMA_reg_buffer_2939 ( .C (clk), .D (plaintext_s0[24]), .Q (new_AGEMA_signal_5715) ) ;
    buf_clk new_AGEMA_reg_buffer_2947 ( .C (clk), .D (plaintext_s1[24]), .Q (new_AGEMA_signal_5723) ) ;
    buf_clk new_AGEMA_reg_buffer_2955 ( .C (clk), .D (plaintext_s2[24]), .Q (new_AGEMA_signal_5731) ) ;
    buf_clk new_AGEMA_reg_buffer_2963 ( .C (clk), .D (plaintext_s0[26]), .Q (new_AGEMA_signal_5739) ) ;
    buf_clk new_AGEMA_reg_buffer_2971 ( .C (clk), .D (plaintext_s1[26]), .Q (new_AGEMA_signal_5747) ) ;
    buf_clk new_AGEMA_reg_buffer_2979 ( .C (clk), .D (plaintext_s2[26]), .Q (new_AGEMA_signal_5755) ) ;
    buf_clk new_AGEMA_reg_buffer_2987 ( .C (clk), .D (plaintext_s0[28]), .Q (new_AGEMA_signal_5763) ) ;
    buf_clk new_AGEMA_reg_buffer_2995 ( .C (clk), .D (plaintext_s1[28]), .Q (new_AGEMA_signal_5771) ) ;
    buf_clk new_AGEMA_reg_buffer_3003 ( .C (clk), .D (plaintext_s2[28]), .Q (new_AGEMA_signal_5779) ) ;
    buf_clk new_AGEMA_reg_buffer_3011 ( .C (clk), .D (plaintext_s0[30]), .Q (new_AGEMA_signal_5787) ) ;
    buf_clk new_AGEMA_reg_buffer_3019 ( .C (clk), .D (plaintext_s1[30]), .Q (new_AGEMA_signal_5795) ) ;
    buf_clk new_AGEMA_reg_buffer_3027 ( .C (clk), .D (plaintext_s2[30]), .Q (new_AGEMA_signal_5803) ) ;
    buf_clk new_AGEMA_reg_buffer_3035 ( .C (clk), .D (plaintext_s0[32]), .Q (new_AGEMA_signal_5811) ) ;
    buf_clk new_AGEMA_reg_buffer_3043 ( .C (clk), .D (plaintext_s1[32]), .Q (new_AGEMA_signal_5819) ) ;
    buf_clk new_AGEMA_reg_buffer_3051 ( .C (clk), .D (plaintext_s2[32]), .Q (new_AGEMA_signal_5827) ) ;
    buf_clk new_AGEMA_reg_buffer_3059 ( .C (clk), .D (plaintext_s0[34]), .Q (new_AGEMA_signal_5835) ) ;
    buf_clk new_AGEMA_reg_buffer_3067 ( .C (clk), .D (plaintext_s1[34]), .Q (new_AGEMA_signal_5843) ) ;
    buf_clk new_AGEMA_reg_buffer_3075 ( .C (clk), .D (plaintext_s2[34]), .Q (new_AGEMA_signal_5851) ) ;
    buf_clk new_AGEMA_reg_buffer_3083 ( .C (clk), .D (plaintext_s0[36]), .Q (new_AGEMA_signal_5859) ) ;
    buf_clk new_AGEMA_reg_buffer_3091 ( .C (clk), .D (plaintext_s1[36]), .Q (new_AGEMA_signal_5867) ) ;
    buf_clk new_AGEMA_reg_buffer_3099 ( .C (clk), .D (plaintext_s2[36]), .Q (new_AGEMA_signal_5875) ) ;
    buf_clk new_AGEMA_reg_buffer_3107 ( .C (clk), .D (plaintext_s0[38]), .Q (new_AGEMA_signal_5883) ) ;
    buf_clk new_AGEMA_reg_buffer_3115 ( .C (clk), .D (plaintext_s1[38]), .Q (new_AGEMA_signal_5891) ) ;
    buf_clk new_AGEMA_reg_buffer_3123 ( .C (clk), .D (plaintext_s2[38]), .Q (new_AGEMA_signal_5899) ) ;
    buf_clk new_AGEMA_reg_buffer_3131 ( .C (clk), .D (plaintext_s0[40]), .Q (new_AGEMA_signal_5907) ) ;
    buf_clk new_AGEMA_reg_buffer_3139 ( .C (clk), .D (plaintext_s1[40]), .Q (new_AGEMA_signal_5915) ) ;
    buf_clk new_AGEMA_reg_buffer_3147 ( .C (clk), .D (plaintext_s2[40]), .Q (new_AGEMA_signal_5923) ) ;
    buf_clk new_AGEMA_reg_buffer_3155 ( .C (clk), .D (plaintext_s0[42]), .Q (new_AGEMA_signal_5931) ) ;
    buf_clk new_AGEMA_reg_buffer_3163 ( .C (clk), .D (plaintext_s1[42]), .Q (new_AGEMA_signal_5939) ) ;
    buf_clk new_AGEMA_reg_buffer_3171 ( .C (clk), .D (plaintext_s2[42]), .Q (new_AGEMA_signal_5947) ) ;
    buf_clk new_AGEMA_reg_buffer_3179 ( .C (clk), .D (plaintext_s0[44]), .Q (new_AGEMA_signal_5955) ) ;
    buf_clk new_AGEMA_reg_buffer_3187 ( .C (clk), .D (plaintext_s1[44]), .Q (new_AGEMA_signal_5963) ) ;
    buf_clk new_AGEMA_reg_buffer_3195 ( .C (clk), .D (plaintext_s2[44]), .Q (new_AGEMA_signal_5971) ) ;
    buf_clk new_AGEMA_reg_buffer_3203 ( .C (clk), .D (plaintext_s0[46]), .Q (new_AGEMA_signal_5979) ) ;
    buf_clk new_AGEMA_reg_buffer_3211 ( .C (clk), .D (plaintext_s1[46]), .Q (new_AGEMA_signal_5987) ) ;
    buf_clk new_AGEMA_reg_buffer_3219 ( .C (clk), .D (plaintext_s2[46]), .Q (new_AGEMA_signal_5995) ) ;
    buf_clk new_AGEMA_reg_buffer_3227 ( .C (clk), .D (plaintext_s0[48]), .Q (new_AGEMA_signal_6003) ) ;
    buf_clk new_AGEMA_reg_buffer_3235 ( .C (clk), .D (plaintext_s1[48]), .Q (new_AGEMA_signal_6011) ) ;
    buf_clk new_AGEMA_reg_buffer_3243 ( .C (clk), .D (plaintext_s2[48]), .Q (new_AGEMA_signal_6019) ) ;
    buf_clk new_AGEMA_reg_buffer_3251 ( .C (clk), .D (plaintext_s0[50]), .Q (new_AGEMA_signal_6027) ) ;
    buf_clk new_AGEMA_reg_buffer_3259 ( .C (clk), .D (plaintext_s1[50]), .Q (new_AGEMA_signal_6035) ) ;
    buf_clk new_AGEMA_reg_buffer_3267 ( .C (clk), .D (plaintext_s2[50]), .Q (new_AGEMA_signal_6043) ) ;
    buf_clk new_AGEMA_reg_buffer_3275 ( .C (clk), .D (plaintext_s0[52]), .Q (new_AGEMA_signal_6051) ) ;
    buf_clk new_AGEMA_reg_buffer_3283 ( .C (clk), .D (plaintext_s1[52]), .Q (new_AGEMA_signal_6059) ) ;
    buf_clk new_AGEMA_reg_buffer_3291 ( .C (clk), .D (plaintext_s2[52]), .Q (new_AGEMA_signal_6067) ) ;
    buf_clk new_AGEMA_reg_buffer_3299 ( .C (clk), .D (plaintext_s0[54]), .Q (new_AGEMA_signal_6075) ) ;
    buf_clk new_AGEMA_reg_buffer_3307 ( .C (clk), .D (plaintext_s1[54]), .Q (new_AGEMA_signal_6083) ) ;
    buf_clk new_AGEMA_reg_buffer_3315 ( .C (clk), .D (plaintext_s2[54]), .Q (new_AGEMA_signal_6091) ) ;
    buf_clk new_AGEMA_reg_buffer_3323 ( .C (clk), .D (plaintext_s0[56]), .Q (new_AGEMA_signal_6099) ) ;
    buf_clk new_AGEMA_reg_buffer_3331 ( .C (clk), .D (plaintext_s1[56]), .Q (new_AGEMA_signal_6107) ) ;
    buf_clk new_AGEMA_reg_buffer_3339 ( .C (clk), .D (plaintext_s2[56]), .Q (new_AGEMA_signal_6115) ) ;
    buf_clk new_AGEMA_reg_buffer_3347 ( .C (clk), .D (plaintext_s0[58]), .Q (new_AGEMA_signal_6123) ) ;
    buf_clk new_AGEMA_reg_buffer_3355 ( .C (clk), .D (plaintext_s1[58]), .Q (new_AGEMA_signal_6131) ) ;
    buf_clk new_AGEMA_reg_buffer_3363 ( .C (clk), .D (plaintext_s2[58]), .Q (new_AGEMA_signal_6139) ) ;
    buf_clk new_AGEMA_reg_buffer_3371 ( .C (clk), .D (plaintext_s0[60]), .Q (new_AGEMA_signal_6147) ) ;
    buf_clk new_AGEMA_reg_buffer_3379 ( .C (clk), .D (plaintext_s1[60]), .Q (new_AGEMA_signal_6155) ) ;
    buf_clk new_AGEMA_reg_buffer_3387 ( .C (clk), .D (plaintext_s2[60]), .Q (new_AGEMA_signal_6163) ) ;
    buf_clk new_AGEMA_reg_buffer_3395 ( .C (clk), .D (plaintext_s0[62]), .Q (new_AGEMA_signal_6171) ) ;
    buf_clk new_AGEMA_reg_buffer_3403 ( .C (clk), .D (plaintext_s1[62]), .Q (new_AGEMA_signal_6179) ) ;
    buf_clk new_AGEMA_reg_buffer_3411 ( .C (clk), .D (plaintext_s2[62]), .Q (new_AGEMA_signal_6187) ) ;
    buf_clk new_AGEMA_reg_buffer_3419 ( .C (clk), .D (SelectedKey[48]), .Q (new_AGEMA_signal_6195) ) ;
    buf_clk new_AGEMA_reg_buffer_3427 ( .C (clk), .D (new_AGEMA_signal_2077), .Q (new_AGEMA_signal_6203) ) ;
    buf_clk new_AGEMA_reg_buffer_3435 ( .C (clk), .D (new_AGEMA_signal_2078), .Q (new_AGEMA_signal_6211) ) ;
    buf_clk new_AGEMA_reg_buffer_3443 ( .C (clk), .D (SelectedKey[50]), .Q (new_AGEMA_signal_6219) ) ;
    buf_clk new_AGEMA_reg_buffer_3451 ( .C (clk), .D (new_AGEMA_signal_2089), .Q (new_AGEMA_signal_6227) ) ;
    buf_clk new_AGEMA_reg_buffer_3459 ( .C (clk), .D (new_AGEMA_signal_2090), .Q (new_AGEMA_signal_6235) ) ;
    buf_clk new_AGEMA_reg_buffer_3467 ( .C (clk), .D (SelectedKey[52]), .Q (new_AGEMA_signal_6243) ) ;
    buf_clk new_AGEMA_reg_buffer_3475 ( .C (clk), .D (new_AGEMA_signal_2101), .Q (new_AGEMA_signal_6251) ) ;
    buf_clk new_AGEMA_reg_buffer_3483 ( .C (clk), .D (new_AGEMA_signal_2102), .Q (new_AGEMA_signal_6259) ) ;
    buf_clk new_AGEMA_reg_buffer_3491 ( .C (clk), .D (SelectedKey[54]), .Q (new_AGEMA_signal_6267) ) ;
    buf_clk new_AGEMA_reg_buffer_3499 ( .C (clk), .D (new_AGEMA_signal_1543), .Q (new_AGEMA_signal_6275) ) ;
    buf_clk new_AGEMA_reg_buffer_3507 ( .C (clk), .D (new_AGEMA_signal_1544), .Q (new_AGEMA_signal_6283) ) ;
    buf_clk new_AGEMA_reg_buffer_3515 ( .C (clk), .D (SelectedKey[56]), .Q (new_AGEMA_signal_6291) ) ;
    buf_clk new_AGEMA_reg_buffer_3523 ( .C (clk), .D (new_AGEMA_signal_1549), .Q (new_AGEMA_signal_6299) ) ;
    buf_clk new_AGEMA_reg_buffer_3531 ( .C (clk), .D (new_AGEMA_signal_1550), .Q (new_AGEMA_signal_6307) ) ;
    buf_clk new_AGEMA_reg_buffer_3539 ( .C (clk), .D (SelectedKey[58]), .Q (new_AGEMA_signal_6315) ) ;
    buf_clk new_AGEMA_reg_buffer_3547 ( .C (clk), .D (new_AGEMA_signal_2119), .Q (new_AGEMA_signal_6323) ) ;
    buf_clk new_AGEMA_reg_buffer_3555 ( .C (clk), .D (new_AGEMA_signal_2120), .Q (new_AGEMA_signal_6331) ) ;
    buf_clk new_AGEMA_reg_buffer_3563 ( .C (clk), .D (SelectedKey[60]), .Q (new_AGEMA_signal_6339) ) ;
    buf_clk new_AGEMA_reg_buffer_3571 ( .C (clk), .D (new_AGEMA_signal_2125), .Q (new_AGEMA_signal_6347) ) ;
    buf_clk new_AGEMA_reg_buffer_3579 ( .C (clk), .D (new_AGEMA_signal_2126), .Q (new_AGEMA_signal_6355) ) ;
    buf_clk new_AGEMA_reg_buffer_3587 ( .C (clk), .D (SelectedKey[62]), .Q (new_AGEMA_signal_6363) ) ;
    buf_clk new_AGEMA_reg_buffer_3595 ( .C (clk), .D (new_AGEMA_signal_1561), .Q (new_AGEMA_signal_6371) ) ;
    buf_clk new_AGEMA_reg_buffer_3603 ( .C (clk), .D (new_AGEMA_signal_1562), .Q (new_AGEMA_signal_6379) ) ;
    buf_clk new_AGEMA_reg_buffer_3611 ( .C (clk), .D (AddKeyConstXOR_XORInst_0_0_n1), .Q (new_AGEMA_signal_6387) ) ;
    buf_clk new_AGEMA_reg_buffer_3619 ( .C (clk), .D (new_AGEMA_signal_2395), .Q (new_AGEMA_signal_6395) ) ;
    buf_clk new_AGEMA_reg_buffer_3627 ( .C (clk), .D (new_AGEMA_signal_2396), .Q (new_AGEMA_signal_6403) ) ;
    buf_clk new_AGEMA_reg_buffer_3635 ( .C (clk), .D (AddKeyConstXOR_XORInst_0_2_n1), .Q (new_AGEMA_signal_6411) ) ;
    buf_clk new_AGEMA_reg_buffer_3643 ( .C (clk), .D (new_AGEMA_signal_2399), .Q (new_AGEMA_signal_6419) ) ;
    buf_clk new_AGEMA_reg_buffer_3651 ( .C (clk), .D (new_AGEMA_signal_2400), .Q (new_AGEMA_signal_6427) ) ;
    buf_clk new_AGEMA_reg_buffer_3659 ( .C (clk), .D (AddKeyConstXOR_XORInst_1_0_n1), .Q (new_AGEMA_signal_6435) ) ;
    buf_clk new_AGEMA_reg_buffer_3667 ( .C (clk), .D (new_AGEMA_signal_2403), .Q (new_AGEMA_signal_6443) ) ;
    buf_clk new_AGEMA_reg_buffer_3675 ( .C (clk), .D (new_AGEMA_signal_2404), .Q (new_AGEMA_signal_6451) ) ;
    buf_clk new_AGEMA_reg_buffer_3683 ( .C (clk), .D (AddKeyConstXOR_XORInst_1_2_n1), .Q (new_AGEMA_signal_6459) ) ;
    buf_clk new_AGEMA_reg_buffer_3691 ( .C (clk), .D (new_AGEMA_signal_2407), .Q (new_AGEMA_signal_6467) ) ;
    buf_clk new_AGEMA_reg_buffer_3699 ( .C (clk), .D (new_AGEMA_signal_2408), .Q (new_AGEMA_signal_6475) ) ;
    buf_clk new_AGEMA_reg_buffer_3707 ( .C (clk), .D (SelectedKey[0]), .Q (new_AGEMA_signal_6483) ) ;
    buf_clk new_AGEMA_reg_buffer_3715 ( .C (clk), .D (new_AGEMA_signal_1471), .Q (new_AGEMA_signal_6491) ) ;
    buf_clk new_AGEMA_reg_buffer_3723 ( .C (clk), .D (new_AGEMA_signal_1472), .Q (new_AGEMA_signal_6499) ) ;
    buf_clk new_AGEMA_reg_buffer_3731 ( .C (clk), .D (SelectedKey[2]), .Q (new_AGEMA_signal_6507) ) ;
    buf_clk new_AGEMA_reg_buffer_3739 ( .C (clk), .D (new_AGEMA_signal_1477), .Q (new_AGEMA_signal_6515) ) ;
    buf_clk new_AGEMA_reg_buffer_3747 ( .C (clk), .D (new_AGEMA_signal_1478), .Q (new_AGEMA_signal_6523) ) ;
    buf_clk new_AGEMA_reg_buffer_3755 ( .C (clk), .D (SelectedKey[4]), .Q (new_AGEMA_signal_6531) ) ;
    buf_clk new_AGEMA_reg_buffer_3763 ( .C (clk), .D (new_AGEMA_signal_1867), .Q (new_AGEMA_signal_6539) ) ;
    buf_clk new_AGEMA_reg_buffer_3771 ( .C (clk), .D (new_AGEMA_signal_1868), .Q (new_AGEMA_signal_6547) ) ;
    buf_clk new_AGEMA_reg_buffer_3779 ( .C (clk), .D (SelectedKey[6]), .Q (new_AGEMA_signal_6555) ) ;
    buf_clk new_AGEMA_reg_buffer_3787 ( .C (clk), .D (new_AGEMA_signal_1879), .Q (new_AGEMA_signal_6563) ) ;
    buf_clk new_AGEMA_reg_buffer_3795 ( .C (clk), .D (new_AGEMA_signal_1880), .Q (new_AGEMA_signal_6571) ) ;
    buf_clk new_AGEMA_reg_buffer_3803 ( .C (clk), .D (SelectedKey[8]), .Q (new_AGEMA_signal_6579) ) ;
    buf_clk new_AGEMA_reg_buffer_3811 ( .C (clk), .D (new_AGEMA_signal_1891), .Q (new_AGEMA_signal_6587) ) ;
    buf_clk new_AGEMA_reg_buffer_3819 ( .C (clk), .D (new_AGEMA_signal_1892), .Q (new_AGEMA_signal_6595) ) ;
    buf_clk new_AGEMA_reg_buffer_3827 ( .C (clk), .D (SelectedKey[10]), .Q (new_AGEMA_signal_6603) ) ;
    buf_clk new_AGEMA_reg_buffer_3835 ( .C (clk), .D (new_AGEMA_signal_1903), .Q (new_AGEMA_signal_6611) ) ;
    buf_clk new_AGEMA_reg_buffer_3843 ( .C (clk), .D (new_AGEMA_signal_1904), .Q (new_AGEMA_signal_6619) ) ;
    buf_clk new_AGEMA_reg_buffer_3851 ( .C (clk), .D (SelectedKey[12]), .Q (new_AGEMA_signal_6627) ) ;
    buf_clk new_AGEMA_reg_buffer_3859 ( .C (clk), .D (new_AGEMA_signal_1915), .Q (new_AGEMA_signal_6635) ) ;
    buf_clk new_AGEMA_reg_buffer_3867 ( .C (clk), .D (new_AGEMA_signal_1916), .Q (new_AGEMA_signal_6643) ) ;
    buf_clk new_AGEMA_reg_buffer_3875 ( .C (clk), .D (SelectedKey[14]), .Q (new_AGEMA_signal_6651) ) ;
    buf_clk new_AGEMA_reg_buffer_3883 ( .C (clk), .D (new_AGEMA_signal_1927), .Q (new_AGEMA_signal_6659) ) ;
    buf_clk new_AGEMA_reg_buffer_3891 ( .C (clk), .D (new_AGEMA_signal_1928), .Q (new_AGEMA_signal_6667) ) ;
    buf_clk new_AGEMA_reg_buffer_3899 ( .C (clk), .D (SelectedKey[16]), .Q (new_AGEMA_signal_6675) ) ;
    buf_clk new_AGEMA_reg_buffer_3907 ( .C (clk), .D (new_AGEMA_signal_1939), .Q (new_AGEMA_signal_6683) ) ;
    buf_clk new_AGEMA_reg_buffer_3915 ( .C (clk), .D (new_AGEMA_signal_1940), .Q (new_AGEMA_signal_6691) ) ;
    buf_clk new_AGEMA_reg_buffer_3923 ( .C (clk), .D (SelectedKey[18]), .Q (new_AGEMA_signal_6699) ) ;
    buf_clk new_AGEMA_reg_buffer_3931 ( .C (clk), .D (new_AGEMA_signal_1951), .Q (new_AGEMA_signal_6707) ) ;
    buf_clk new_AGEMA_reg_buffer_3939 ( .C (clk), .D (new_AGEMA_signal_1952), .Q (new_AGEMA_signal_6715) ) ;
    buf_clk new_AGEMA_reg_buffer_3947 ( .C (clk), .D (SelectedKey[20]), .Q (new_AGEMA_signal_6723) ) ;
    buf_clk new_AGEMA_reg_buffer_3955 ( .C (clk), .D (new_AGEMA_signal_1963), .Q (new_AGEMA_signal_6731) ) ;
    buf_clk new_AGEMA_reg_buffer_3963 ( .C (clk), .D (new_AGEMA_signal_1964), .Q (new_AGEMA_signal_6739) ) ;
    buf_clk new_AGEMA_reg_buffer_3971 ( .C (clk), .D (SelectedKey[22]), .Q (new_AGEMA_signal_6747) ) ;
    buf_clk new_AGEMA_reg_buffer_3979 ( .C (clk), .D (new_AGEMA_signal_1483), .Q (new_AGEMA_signal_6755) ) ;
    buf_clk new_AGEMA_reg_buffer_3987 ( .C (clk), .D (new_AGEMA_signal_1484), .Q (new_AGEMA_signal_6763) ) ;
    buf_clk new_AGEMA_reg_buffer_3995 ( .C (clk), .D (SelectedKey[24]), .Q (new_AGEMA_signal_6771) ) ;
    buf_clk new_AGEMA_reg_buffer_4003 ( .C (clk), .D (new_AGEMA_signal_1495), .Q (new_AGEMA_signal_6779) ) ;
    buf_clk new_AGEMA_reg_buffer_4011 ( .C (clk), .D (new_AGEMA_signal_1496), .Q (new_AGEMA_signal_6787) ) ;
    buf_clk new_AGEMA_reg_buffer_4019 ( .C (clk), .D (SelectedKey[26]), .Q (new_AGEMA_signal_6795) ) ;
    buf_clk new_AGEMA_reg_buffer_4027 ( .C (clk), .D (new_AGEMA_signal_1507), .Q (new_AGEMA_signal_6803) ) ;
    buf_clk new_AGEMA_reg_buffer_4035 ( .C (clk), .D (new_AGEMA_signal_1508), .Q (new_AGEMA_signal_6811) ) ;
    buf_clk new_AGEMA_reg_buffer_4043 ( .C (clk), .D (SelectedKey[28]), .Q (new_AGEMA_signal_6819) ) ;
    buf_clk new_AGEMA_reg_buffer_4051 ( .C (clk), .D (new_AGEMA_signal_1975), .Q (new_AGEMA_signal_6827) ) ;
    buf_clk new_AGEMA_reg_buffer_4059 ( .C (clk), .D (new_AGEMA_signal_1976), .Q (new_AGEMA_signal_6835) ) ;
    buf_clk new_AGEMA_reg_buffer_4067 ( .C (clk), .D (SelectedKey[30]), .Q (new_AGEMA_signal_6843) ) ;
    buf_clk new_AGEMA_reg_buffer_4075 ( .C (clk), .D (new_AGEMA_signal_1987), .Q (new_AGEMA_signal_6851) ) ;
    buf_clk new_AGEMA_reg_buffer_4083 ( .C (clk), .D (new_AGEMA_signal_1988), .Q (new_AGEMA_signal_6859) ) ;
    buf_clk new_AGEMA_reg_buffer_4091 ( .C (clk), .D (SelectedKey[32]), .Q (new_AGEMA_signal_6867) ) ;
    buf_clk new_AGEMA_reg_buffer_4099 ( .C (clk), .D (new_AGEMA_signal_1999), .Q (new_AGEMA_signal_6875) ) ;
    buf_clk new_AGEMA_reg_buffer_4107 ( .C (clk), .D (new_AGEMA_signal_2000), .Q (new_AGEMA_signal_6883) ) ;
    buf_clk new_AGEMA_reg_buffer_4115 ( .C (clk), .D (SelectedKey[34]), .Q (new_AGEMA_signal_6891) ) ;
    buf_clk new_AGEMA_reg_buffer_4123 ( .C (clk), .D (new_AGEMA_signal_2005), .Q (new_AGEMA_signal_6899) ) ;
    buf_clk new_AGEMA_reg_buffer_4131 ( .C (clk), .D (new_AGEMA_signal_2006), .Q (new_AGEMA_signal_6907) ) ;
    buf_clk new_AGEMA_reg_buffer_4139 ( .C (clk), .D (SelectedKey[36]), .Q (new_AGEMA_signal_6915) ) ;
    buf_clk new_AGEMA_reg_buffer_4147 ( .C (clk), .D (new_AGEMA_signal_1525), .Q (new_AGEMA_signal_6923) ) ;
    buf_clk new_AGEMA_reg_buffer_4155 ( .C (clk), .D (new_AGEMA_signal_1526), .Q (new_AGEMA_signal_6931) ) ;
    buf_clk new_AGEMA_reg_buffer_4163 ( .C (clk), .D (SelectedKey[38]), .Q (new_AGEMA_signal_6939) ) ;
    buf_clk new_AGEMA_reg_buffer_4171 ( .C (clk), .D (new_AGEMA_signal_2023), .Q (new_AGEMA_signal_6947) ) ;
    buf_clk new_AGEMA_reg_buffer_4179 ( .C (clk), .D (new_AGEMA_signal_2024), .Q (new_AGEMA_signal_6955) ) ;
    buf_clk new_AGEMA_reg_buffer_4667 ( .C (clk), .D (FSMUpdate[6]), .Q (new_AGEMA_signal_7443) ) ;
    buf_clk new_AGEMA_reg_buffer_4675 ( .C (clk), .D (FSMUpdate[5]), .Q (new_AGEMA_signal_7451) ) ;
    buf_clk new_AGEMA_reg_buffer_4683 ( .C (clk), .D (FSMUpdate[4]), .Q (new_AGEMA_signal_7459) ) ;
    buf_clk new_AGEMA_reg_buffer_4691 ( .C (clk), .D (FSMUpdate[3]), .Q (new_AGEMA_signal_7467) ) ;
    buf_clk new_AGEMA_reg_buffer_4699 ( .C (clk), .D (FSMUpdate[2]), .Q (new_AGEMA_signal_7475) ) ;
    buf_clk new_AGEMA_reg_buffer_4707 ( .C (clk), .D (FSMUpdate[1]), .Q (new_AGEMA_signal_7483) ) ;
    buf_clk new_AGEMA_reg_buffer_4715 ( .C (clk), .D (FSMUpdate[0]), .Q (new_AGEMA_signal_7491) ) ;
    buf_clk new_AGEMA_reg_buffer_4723 ( .C (clk), .D (selectsNext[1]), .Q (new_AGEMA_signal_7499) ) ;
    buf_clk new_AGEMA_reg_buffer_4731 ( .C (clk), .D (selectsNext[0]), .Q (new_AGEMA_signal_7507) ) ;
    buf_clk new_AGEMA_reg_buffer_4739 ( .C (clk), .D (done_internal), .Q (new_AGEMA_signal_7515) ) ;

    /* cells in depth 2 */
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U14 ( .a ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_1024, new_AGEMA_signal_1023, SubCellInst_SboxInst_0_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U13 ( .a ({new_AGEMA_signal_1032, new_AGEMA_signal_1031, SubCellInst_SboxInst_0_n8}), .b ({new_AGEMA_signal_1030, new_AGEMA_signal_1029, SubCellInst_SboxInst_0_n7}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, SubCellInst_SboxInst_0_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U10 ( .a ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, SubCellInst_SboxInst_0_n9}), .clk (clk), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, SubCellInst_SboxInst_0_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U9 ( .a ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_1032, new_AGEMA_signal_1031, SubCellInst_SboxInst_0_n8}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({new_AGEMA_signal_1282, new_AGEMA_signal_1281, SubCellInst_SboxInst_0_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U5 ( .a ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, SubCellInst_SboxInst_0_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U3 ( .a ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, SubCellInst_SboxInst_0_n9}), .b ({new_AGEMA_signal_1032, new_AGEMA_signal_1031, SubCellInst_SboxInst_0_n8}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, SubCellInst_SboxInst_0_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U14 ( .a ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .b ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .clk (clk), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_1040, new_AGEMA_signal_1039, SubCellInst_SboxInst_1_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U13 ( .a ({new_AGEMA_signal_1048, new_AGEMA_signal_1047, SubCellInst_SboxInst_1_n8}), .b ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, SubCellInst_SboxInst_1_n7}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({new_AGEMA_signal_1290, new_AGEMA_signal_1289, SubCellInst_SboxInst_1_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U10 ( .a ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .b ({new_AGEMA_signal_1050, new_AGEMA_signal_1049, SubCellInst_SboxInst_1_n9}), .clk (clk), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, SubCellInst_SboxInst_1_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U9 ( .a ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .b ({new_AGEMA_signal_1048, new_AGEMA_signal_1047, SubCellInst_SboxInst_1_n8}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({new_AGEMA_signal_1294, new_AGEMA_signal_1293, SubCellInst_SboxInst_1_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U5 ( .a ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .b ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .clk (clk), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_1044, new_AGEMA_signal_1043, SubCellInst_SboxInst_1_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U3 ( .a ({new_AGEMA_signal_1050, new_AGEMA_signal_1049, SubCellInst_SboxInst_1_n9}), .b ({new_AGEMA_signal_1048, new_AGEMA_signal_1047, SubCellInst_SboxInst_1_n8}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({new_AGEMA_signal_1298, new_AGEMA_signal_1297, SubCellInst_SboxInst_1_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U14 ( .a ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_1056, new_AGEMA_signal_1055, SubCellInst_SboxInst_2_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U13 ( .a ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, SubCellInst_SboxInst_2_n8}), .b ({new_AGEMA_signal_1062, new_AGEMA_signal_1061, SubCellInst_SboxInst_2_n7}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({new_AGEMA_signal_1302, new_AGEMA_signal_1301, SubCellInst_SboxInst_2_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U10 ( .a ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({new_AGEMA_signal_1066, new_AGEMA_signal_1065, SubCellInst_SboxInst_2_n9}), .clk (clk), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, SubCellInst_SboxInst_2_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U9 ( .a ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, SubCellInst_SboxInst_2_n8}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({new_AGEMA_signal_1306, new_AGEMA_signal_1305, SubCellInst_SboxInst_2_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U5 ( .a ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_1060, new_AGEMA_signal_1059, SubCellInst_SboxInst_2_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U3 ( .a ({new_AGEMA_signal_1066, new_AGEMA_signal_1065, SubCellInst_SboxInst_2_n9}), .b ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, SubCellInst_SboxInst_2_n8}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({new_AGEMA_signal_1310, new_AGEMA_signal_1309, SubCellInst_SboxInst_2_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U14 ( .a ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .clk (clk), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_1072, new_AGEMA_signal_1071, SubCellInst_SboxInst_3_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U13 ( .a ({new_AGEMA_signal_1080, new_AGEMA_signal_1079, SubCellInst_SboxInst_3_n8}), .b ({new_AGEMA_signal_1078, new_AGEMA_signal_1077, SubCellInst_SboxInst_3_n7}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({new_AGEMA_signal_1314, new_AGEMA_signal_1313, SubCellInst_SboxInst_3_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U10 ( .a ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, SubCellInst_SboxInst_3_n9}), .clk (clk), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, SubCellInst_SboxInst_3_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U9 ( .a ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .b ({new_AGEMA_signal_1080, new_AGEMA_signal_1079, SubCellInst_SboxInst_3_n8}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({new_AGEMA_signal_1318, new_AGEMA_signal_1317, SubCellInst_SboxInst_3_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U5 ( .a ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .clk (clk), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, SubCellInst_SboxInst_3_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U3 ( .a ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, SubCellInst_SboxInst_3_n9}), .b ({new_AGEMA_signal_1080, new_AGEMA_signal_1079, SubCellInst_SboxInst_3_n8}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, SubCellInst_SboxInst_3_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U14 ( .a ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .b ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .clk (clk), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, SubCellInst_SboxInst_4_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U13 ( .a ({new_AGEMA_signal_1096, new_AGEMA_signal_1095, SubCellInst_SboxInst_4_n8}), .b ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, SubCellInst_SboxInst_4_n7}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({new_AGEMA_signal_1326, new_AGEMA_signal_1325, SubCellInst_SboxInst_4_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U10 ( .a ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .b ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, SubCellInst_SboxInst_4_n9}), .clk (clk), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, SubCellInst_SboxInst_4_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U9 ( .a ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .b ({new_AGEMA_signal_1096, new_AGEMA_signal_1095, SubCellInst_SboxInst_4_n8}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({new_AGEMA_signal_1330, new_AGEMA_signal_1329, SubCellInst_SboxInst_4_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U5 ( .a ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .b ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .clk (clk), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_1092, new_AGEMA_signal_1091, SubCellInst_SboxInst_4_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U3 ( .a ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, SubCellInst_SboxInst_4_n9}), .b ({new_AGEMA_signal_1096, new_AGEMA_signal_1095, SubCellInst_SboxInst_4_n8}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({new_AGEMA_signal_1334, new_AGEMA_signal_1333, SubCellInst_SboxInst_4_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U14 ( .a ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_1104, new_AGEMA_signal_1103, SubCellInst_SboxInst_5_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U13 ( .a ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, SubCellInst_SboxInst_5_n8}), .b ({new_AGEMA_signal_1110, new_AGEMA_signal_1109, SubCellInst_SboxInst_5_n7}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({new_AGEMA_signal_1338, new_AGEMA_signal_1337, SubCellInst_SboxInst_5_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U10 ( .a ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, SubCellInst_SboxInst_5_n9}), .clk (clk), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, SubCellInst_SboxInst_5_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U9 ( .a ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, SubCellInst_SboxInst_5_n8}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({new_AGEMA_signal_1342, new_AGEMA_signal_1341, SubCellInst_SboxInst_5_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U5 ( .a ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r ({Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_1108, new_AGEMA_signal_1107, SubCellInst_SboxInst_5_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U3 ( .a ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, SubCellInst_SboxInst_5_n9}), .b ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, SubCellInst_SboxInst_5_n8}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105]}), .c ({new_AGEMA_signal_1346, new_AGEMA_signal_1345, SubCellInst_SboxInst_5_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U14 ( .a ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .b ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .clk (clk), .r ({Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_1120, new_AGEMA_signal_1119, SubCellInst_SboxInst_6_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U13 ( .a ({new_AGEMA_signal_1128, new_AGEMA_signal_1127, SubCellInst_SboxInst_6_n8}), .b ({new_AGEMA_signal_1126, new_AGEMA_signal_1125, SubCellInst_SboxInst_6_n7}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111]}), .c ({new_AGEMA_signal_1350, new_AGEMA_signal_1349, SubCellInst_SboxInst_6_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U10 ( .a ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .b ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, SubCellInst_SboxInst_6_n9}), .clk (clk), .r ({Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_1352, new_AGEMA_signal_1351, SubCellInst_SboxInst_6_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U9 ( .a ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .b ({new_AGEMA_signal_1128, new_AGEMA_signal_1127, SubCellInst_SboxInst_6_n8}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117]}), .c ({new_AGEMA_signal_1354, new_AGEMA_signal_1353, SubCellInst_SboxInst_6_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U5 ( .a ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .b ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .clk (clk), .r ({Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, SubCellInst_SboxInst_6_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U3 ( .a ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, SubCellInst_SboxInst_6_n9}), .b ({new_AGEMA_signal_1128, new_AGEMA_signal_1127, SubCellInst_SboxInst_6_n8}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123]}), .c ({new_AGEMA_signal_1358, new_AGEMA_signal_1357, SubCellInst_SboxInst_6_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U14 ( .a ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r ({Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, SubCellInst_SboxInst_7_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U13 ( .a ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, SubCellInst_SboxInst_7_n8}), .b ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, SubCellInst_SboxInst_7_n7}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129]}), .c ({new_AGEMA_signal_1362, new_AGEMA_signal_1361, SubCellInst_SboxInst_7_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U10 ( .a ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({new_AGEMA_signal_1146, new_AGEMA_signal_1145, SubCellInst_SboxInst_7_n9}), .clk (clk), .r ({Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_1364, new_AGEMA_signal_1363, SubCellInst_SboxInst_7_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U9 ( .a ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, SubCellInst_SboxInst_7_n8}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135]}), .c ({new_AGEMA_signal_1366, new_AGEMA_signal_1365, SubCellInst_SboxInst_7_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U5 ( .a ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r ({Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_1140, new_AGEMA_signal_1139, SubCellInst_SboxInst_7_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U3 ( .a ({new_AGEMA_signal_1146, new_AGEMA_signal_1145, SubCellInst_SboxInst_7_n9}), .b ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, SubCellInst_SboxInst_7_n8}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141]}), .c ({new_AGEMA_signal_1370, new_AGEMA_signal_1369, SubCellInst_SboxInst_7_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U14 ( .a ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .b ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .clk (clk), .r ({Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_1152, new_AGEMA_signal_1151, SubCellInst_SboxInst_8_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U13 ( .a ({new_AGEMA_signal_1160, new_AGEMA_signal_1159, SubCellInst_SboxInst_8_n8}), .b ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, SubCellInst_SboxInst_8_n7}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147]}), .c ({new_AGEMA_signal_1374, new_AGEMA_signal_1373, SubCellInst_SboxInst_8_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U10 ( .a ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .b ({new_AGEMA_signal_1162, new_AGEMA_signal_1161, SubCellInst_SboxInst_8_n9}), .clk (clk), .r ({Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_1376, new_AGEMA_signal_1375, SubCellInst_SboxInst_8_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U9 ( .a ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .b ({new_AGEMA_signal_1160, new_AGEMA_signal_1159, SubCellInst_SboxInst_8_n8}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153]}), .c ({new_AGEMA_signal_1378, new_AGEMA_signal_1377, SubCellInst_SboxInst_8_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U5 ( .a ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .b ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .clk (clk), .r ({Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_1156, new_AGEMA_signal_1155, SubCellInst_SboxInst_8_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U3 ( .a ({new_AGEMA_signal_1162, new_AGEMA_signal_1161, SubCellInst_SboxInst_8_n9}), .b ({new_AGEMA_signal_1160, new_AGEMA_signal_1159, SubCellInst_SboxInst_8_n8}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159]}), .c ({new_AGEMA_signal_1382, new_AGEMA_signal_1381, SubCellInst_SboxInst_8_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U14 ( .a ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r ({Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_1168, new_AGEMA_signal_1167, SubCellInst_SboxInst_9_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U13 ( .a ({new_AGEMA_signal_1176, new_AGEMA_signal_1175, SubCellInst_SboxInst_9_n8}), .b ({new_AGEMA_signal_1174, new_AGEMA_signal_1173, SubCellInst_SboxInst_9_n7}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165]}), .c ({new_AGEMA_signal_1386, new_AGEMA_signal_1385, SubCellInst_SboxInst_9_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U10 ( .a ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, SubCellInst_SboxInst_9_n9}), .clk (clk), .r ({Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_1388, new_AGEMA_signal_1387, SubCellInst_SboxInst_9_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U9 ( .a ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_1176, new_AGEMA_signal_1175, SubCellInst_SboxInst_9_n8}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171]}), .c ({new_AGEMA_signal_1390, new_AGEMA_signal_1389, SubCellInst_SboxInst_9_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U5 ( .a ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r ({Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_1172, new_AGEMA_signal_1171, SubCellInst_SboxInst_9_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U3 ( .a ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, SubCellInst_SboxInst_9_n9}), .b ({new_AGEMA_signal_1176, new_AGEMA_signal_1175, SubCellInst_SboxInst_9_n8}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177]}), .c ({new_AGEMA_signal_1394, new_AGEMA_signal_1393, SubCellInst_SboxInst_9_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U14 ( .a ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .clk (clk), .r ({Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_1184, new_AGEMA_signal_1183, SubCellInst_SboxInst_10_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U13 ( .a ({new_AGEMA_signal_1192, new_AGEMA_signal_1191, SubCellInst_SboxInst_10_n8}), .b ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, SubCellInst_SboxInst_10_n7}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183]}), .c ({new_AGEMA_signal_1398, new_AGEMA_signal_1397, SubCellInst_SboxInst_10_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U10 ( .a ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_1194, new_AGEMA_signal_1193, SubCellInst_SboxInst_10_n9}), .clk (clk), .r ({Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_1400, new_AGEMA_signal_1399, SubCellInst_SboxInst_10_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U9 ( .a ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .b ({new_AGEMA_signal_1192, new_AGEMA_signal_1191, SubCellInst_SboxInst_10_n8}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189]}), .c ({new_AGEMA_signal_1402, new_AGEMA_signal_1401, SubCellInst_SboxInst_10_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U5 ( .a ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .clk (clk), .r ({Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_1188, new_AGEMA_signal_1187, SubCellInst_SboxInst_10_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U3 ( .a ({new_AGEMA_signal_1194, new_AGEMA_signal_1193, SubCellInst_SboxInst_10_n9}), .b ({new_AGEMA_signal_1192, new_AGEMA_signal_1191, SubCellInst_SboxInst_10_n8}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195]}), .c ({new_AGEMA_signal_1406, new_AGEMA_signal_1405, SubCellInst_SboxInst_10_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U14 ( .a ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r ({Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_1200, new_AGEMA_signal_1199, SubCellInst_SboxInst_11_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U13 ( .a ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, SubCellInst_SboxInst_11_n8}), .b ({new_AGEMA_signal_1206, new_AGEMA_signal_1205, SubCellInst_SboxInst_11_n7}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201]}), .c ({new_AGEMA_signal_1410, new_AGEMA_signal_1409, SubCellInst_SboxInst_11_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U10 ( .a ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({new_AGEMA_signal_1210, new_AGEMA_signal_1209, SubCellInst_SboxInst_11_n9}), .clk (clk), .r ({Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_1412, new_AGEMA_signal_1411, SubCellInst_SboxInst_11_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U9 ( .a ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, SubCellInst_SboxInst_11_n8}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207]}), .c ({new_AGEMA_signal_1414, new_AGEMA_signal_1413, SubCellInst_SboxInst_11_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U5 ( .a ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r ({Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_1204, new_AGEMA_signal_1203, SubCellInst_SboxInst_11_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U3 ( .a ({new_AGEMA_signal_1210, new_AGEMA_signal_1209, SubCellInst_SboxInst_11_n9}), .b ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, SubCellInst_SboxInst_11_n8}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213]}), .c ({new_AGEMA_signal_1418, new_AGEMA_signal_1417, SubCellInst_SboxInst_11_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U14 ( .a ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r ({Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_1216, new_AGEMA_signal_1215, SubCellInst_SboxInst_12_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U13 ( .a ({new_AGEMA_signal_1224, new_AGEMA_signal_1223, SubCellInst_SboxInst_12_n8}), .b ({new_AGEMA_signal_1222, new_AGEMA_signal_1221, SubCellInst_SboxInst_12_n7}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219]}), .c ({new_AGEMA_signal_1422, new_AGEMA_signal_1421, SubCellInst_SboxInst_12_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U10 ( .a ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({new_AGEMA_signal_1226, new_AGEMA_signal_1225, SubCellInst_SboxInst_12_n9}), .clk (clk), .r ({Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_1424, new_AGEMA_signal_1423, SubCellInst_SboxInst_12_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U9 ( .a ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({new_AGEMA_signal_1224, new_AGEMA_signal_1223, SubCellInst_SboxInst_12_n8}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225]}), .c ({new_AGEMA_signal_1426, new_AGEMA_signal_1425, SubCellInst_SboxInst_12_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U5 ( .a ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r ({Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, SubCellInst_SboxInst_12_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U3 ( .a ({new_AGEMA_signal_1226, new_AGEMA_signal_1225, SubCellInst_SboxInst_12_n9}), .b ({new_AGEMA_signal_1224, new_AGEMA_signal_1223, SubCellInst_SboxInst_12_n8}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231]}), .c ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, SubCellInst_SboxInst_12_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U14 ( .a ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .b ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .clk (clk), .r ({Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, SubCellInst_SboxInst_13_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U13 ( .a ({new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_13_n8}), .b ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, SubCellInst_SboxInst_13_n7}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237]}), .c ({new_AGEMA_signal_1434, new_AGEMA_signal_1433, SubCellInst_SboxInst_13_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U10 ( .a ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .b ({new_AGEMA_signal_1242, new_AGEMA_signal_1241, SubCellInst_SboxInst_13_n9}), .clk (clk), .r ({Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_1436, new_AGEMA_signal_1435, SubCellInst_SboxInst_13_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U9 ( .a ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .b ({new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_13_n8}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243]}), .c ({new_AGEMA_signal_1438, new_AGEMA_signal_1437, SubCellInst_SboxInst_13_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U5 ( .a ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .b ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .clk (clk), .r ({Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_1236, new_AGEMA_signal_1235, SubCellInst_SboxInst_13_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U3 ( .a ({new_AGEMA_signal_1242, new_AGEMA_signal_1241, SubCellInst_SboxInst_13_n9}), .b ({new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_13_n8}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249]}), .c ({new_AGEMA_signal_1442, new_AGEMA_signal_1441, SubCellInst_SboxInst_13_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U14 ( .a ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r ({Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_1248, new_AGEMA_signal_1247, SubCellInst_SboxInst_14_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U13 ( .a ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, SubCellInst_SboxInst_14_n8}), .b ({new_AGEMA_signal_1254, new_AGEMA_signal_1253, SubCellInst_SboxInst_14_n7}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255]}), .c ({new_AGEMA_signal_1446, new_AGEMA_signal_1445, SubCellInst_SboxInst_14_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U10 ( .a ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_14_n9}), .clk (clk), .r ({Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_1448, new_AGEMA_signal_1447, SubCellInst_SboxInst_14_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U9 ( .a ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, SubCellInst_SboxInst_14_n8}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261]}), .c ({new_AGEMA_signal_1450, new_AGEMA_signal_1449, SubCellInst_SboxInst_14_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U5 ( .a ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r ({Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_1252, new_AGEMA_signal_1251, SubCellInst_SboxInst_14_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U3 ( .a ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_14_n9}), .b ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, SubCellInst_SboxInst_14_n8}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267]}), .c ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, SubCellInst_SboxInst_14_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U14 ( .a ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .b ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .clk (clk), .r ({Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_1264, new_AGEMA_signal_1263, SubCellInst_SboxInst_15_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U13 ( .a ({new_AGEMA_signal_1272, new_AGEMA_signal_1271, SubCellInst_SboxInst_15_n8}), .b ({new_AGEMA_signal_1270, new_AGEMA_signal_1269, SubCellInst_SboxInst_15_n7}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273]}), .c ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, SubCellInst_SboxInst_15_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U10 ( .a ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .b ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, SubCellInst_SboxInst_15_n9}), .clk (clk), .r ({Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_1460, new_AGEMA_signal_1459, SubCellInst_SboxInst_15_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U9 ( .a ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .b ({new_AGEMA_signal_1272, new_AGEMA_signal_1271, SubCellInst_SboxInst_15_n8}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279]}), .c ({new_AGEMA_signal_1462, new_AGEMA_signal_1461, SubCellInst_SboxInst_15_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U5 ( .a ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .b ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .clk (clk), .r ({Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, SubCellInst_SboxInst_15_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U3 ( .a ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, SubCellInst_SboxInst_15_n9}), .b ({new_AGEMA_signal_1272, new_AGEMA_signal_1271, SubCellInst_SboxInst_15_n8}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285]}), .c ({new_AGEMA_signal_1466, new_AGEMA_signal_1465, SubCellInst_SboxInst_15_n13}) ) ;
    buf_clk new_AGEMA_reg_buffer_820 ( .C (clk), .D (new_AGEMA_signal_3595), .Q (new_AGEMA_signal_3596) ) ;
    buf_clk new_AGEMA_reg_buffer_822 ( .C (clk), .D (new_AGEMA_signal_3597), .Q (new_AGEMA_signal_3598) ) ;
    buf_clk new_AGEMA_reg_buffer_824 ( .C (clk), .D (new_AGEMA_signal_3599), .Q (new_AGEMA_signal_3600) ) ;
    buf_clk new_AGEMA_reg_buffer_826 ( .C (clk), .D (new_AGEMA_signal_3601), .Q (new_AGEMA_signal_3602) ) ;
    buf_clk new_AGEMA_reg_buffer_828 ( .C (clk), .D (new_AGEMA_signal_3603), .Q (new_AGEMA_signal_3604) ) ;
    buf_clk new_AGEMA_reg_buffer_830 ( .C (clk), .D (new_AGEMA_signal_3605), .Q (new_AGEMA_signal_3606) ) ;
    buf_clk new_AGEMA_reg_buffer_832 ( .C (clk), .D (new_AGEMA_signal_3607), .Q (new_AGEMA_signal_3608) ) ;
    buf_clk new_AGEMA_reg_buffer_834 ( .C (clk), .D (new_AGEMA_signal_3609), .Q (new_AGEMA_signal_3610) ) ;
    buf_clk new_AGEMA_reg_buffer_836 ( .C (clk), .D (new_AGEMA_signal_3611), .Q (new_AGEMA_signal_3612) ) ;
    buf_clk new_AGEMA_reg_buffer_838 ( .C (clk), .D (new_AGEMA_signal_3613), .Q (new_AGEMA_signal_3614) ) ;
    buf_clk new_AGEMA_reg_buffer_840 ( .C (clk), .D (new_AGEMA_signal_3615), .Q (new_AGEMA_signal_3616) ) ;
    buf_clk new_AGEMA_reg_buffer_842 ( .C (clk), .D (new_AGEMA_signal_3617), .Q (new_AGEMA_signal_3618) ) ;
    buf_clk new_AGEMA_reg_buffer_844 ( .C (clk), .D (new_AGEMA_signal_3619), .Q (new_AGEMA_signal_3620) ) ;
    buf_clk new_AGEMA_reg_buffer_846 ( .C (clk), .D (new_AGEMA_signal_3621), .Q (new_AGEMA_signal_3622) ) ;
    buf_clk new_AGEMA_reg_buffer_848 ( .C (clk), .D (new_AGEMA_signal_3623), .Q (new_AGEMA_signal_3624) ) ;
    buf_clk new_AGEMA_reg_buffer_850 ( .C (clk), .D (new_AGEMA_signal_3625), .Q (new_AGEMA_signal_3626) ) ;
    buf_clk new_AGEMA_reg_buffer_852 ( .C (clk), .D (new_AGEMA_signal_3627), .Q (new_AGEMA_signal_3628) ) ;
    buf_clk new_AGEMA_reg_buffer_854 ( .C (clk), .D (new_AGEMA_signal_3629), .Q (new_AGEMA_signal_3630) ) ;
    buf_clk new_AGEMA_reg_buffer_856 ( .C (clk), .D (new_AGEMA_signal_3631), .Q (new_AGEMA_signal_3632) ) ;
    buf_clk new_AGEMA_reg_buffer_858 ( .C (clk), .D (new_AGEMA_signal_3633), .Q (new_AGEMA_signal_3634) ) ;
    buf_clk new_AGEMA_reg_buffer_860 ( .C (clk), .D (new_AGEMA_signal_3635), .Q (new_AGEMA_signal_3636) ) ;
    buf_clk new_AGEMA_reg_buffer_862 ( .C (clk), .D (new_AGEMA_signal_3637), .Q (new_AGEMA_signal_3638) ) ;
    buf_clk new_AGEMA_reg_buffer_864 ( .C (clk), .D (new_AGEMA_signal_3639), .Q (new_AGEMA_signal_3640) ) ;
    buf_clk new_AGEMA_reg_buffer_866 ( .C (clk), .D (new_AGEMA_signal_3641), .Q (new_AGEMA_signal_3642) ) ;
    buf_clk new_AGEMA_reg_buffer_868 ( .C (clk), .D (new_AGEMA_signal_3643), .Q (new_AGEMA_signal_3644) ) ;
    buf_clk new_AGEMA_reg_buffer_870 ( .C (clk), .D (new_AGEMA_signal_3645), .Q (new_AGEMA_signal_3646) ) ;
    buf_clk new_AGEMA_reg_buffer_872 ( .C (clk), .D (new_AGEMA_signal_3647), .Q (new_AGEMA_signal_3648) ) ;
    buf_clk new_AGEMA_reg_buffer_874 ( .C (clk), .D (new_AGEMA_signal_3649), .Q (new_AGEMA_signal_3650) ) ;
    buf_clk new_AGEMA_reg_buffer_876 ( .C (clk), .D (new_AGEMA_signal_3651), .Q (new_AGEMA_signal_3652) ) ;
    buf_clk new_AGEMA_reg_buffer_878 ( .C (clk), .D (new_AGEMA_signal_3653), .Q (new_AGEMA_signal_3654) ) ;
    buf_clk new_AGEMA_reg_buffer_880 ( .C (clk), .D (new_AGEMA_signal_3655), .Q (new_AGEMA_signal_3656) ) ;
    buf_clk new_AGEMA_reg_buffer_882 ( .C (clk), .D (new_AGEMA_signal_3657), .Q (new_AGEMA_signal_3658) ) ;
    buf_clk new_AGEMA_reg_buffer_884 ( .C (clk), .D (new_AGEMA_signal_3659), .Q (new_AGEMA_signal_3660) ) ;
    buf_clk new_AGEMA_reg_buffer_886 ( .C (clk), .D (new_AGEMA_signal_3661), .Q (new_AGEMA_signal_3662) ) ;
    buf_clk new_AGEMA_reg_buffer_888 ( .C (clk), .D (new_AGEMA_signal_3663), .Q (new_AGEMA_signal_3664) ) ;
    buf_clk new_AGEMA_reg_buffer_890 ( .C (clk), .D (new_AGEMA_signal_3665), .Q (new_AGEMA_signal_3666) ) ;
    buf_clk new_AGEMA_reg_buffer_892 ( .C (clk), .D (new_AGEMA_signal_3667), .Q (new_AGEMA_signal_3668) ) ;
    buf_clk new_AGEMA_reg_buffer_894 ( .C (clk), .D (new_AGEMA_signal_3669), .Q (new_AGEMA_signal_3670) ) ;
    buf_clk new_AGEMA_reg_buffer_896 ( .C (clk), .D (new_AGEMA_signal_3671), .Q (new_AGEMA_signal_3672) ) ;
    buf_clk new_AGEMA_reg_buffer_898 ( .C (clk), .D (new_AGEMA_signal_3673), .Q (new_AGEMA_signal_3674) ) ;
    buf_clk new_AGEMA_reg_buffer_900 ( .C (clk), .D (new_AGEMA_signal_3675), .Q (new_AGEMA_signal_3676) ) ;
    buf_clk new_AGEMA_reg_buffer_902 ( .C (clk), .D (new_AGEMA_signal_3677), .Q (new_AGEMA_signal_3678) ) ;
    buf_clk new_AGEMA_reg_buffer_904 ( .C (clk), .D (new_AGEMA_signal_3679), .Q (new_AGEMA_signal_3680) ) ;
    buf_clk new_AGEMA_reg_buffer_906 ( .C (clk), .D (new_AGEMA_signal_3681), .Q (new_AGEMA_signal_3682) ) ;
    buf_clk new_AGEMA_reg_buffer_908 ( .C (clk), .D (new_AGEMA_signal_3683), .Q (new_AGEMA_signal_3684) ) ;
    buf_clk new_AGEMA_reg_buffer_910 ( .C (clk), .D (new_AGEMA_signal_3685), .Q (new_AGEMA_signal_3686) ) ;
    buf_clk new_AGEMA_reg_buffer_912 ( .C (clk), .D (new_AGEMA_signal_3687), .Q (new_AGEMA_signal_3688) ) ;
    buf_clk new_AGEMA_reg_buffer_914 ( .C (clk), .D (new_AGEMA_signal_3689), .Q (new_AGEMA_signal_3690) ) ;
    buf_clk new_AGEMA_reg_buffer_916 ( .C (clk), .D (new_AGEMA_signal_3691), .Q (new_AGEMA_signal_3692) ) ;
    buf_clk new_AGEMA_reg_buffer_918 ( .C (clk), .D (new_AGEMA_signal_3693), .Q (new_AGEMA_signal_3694) ) ;
    buf_clk new_AGEMA_reg_buffer_920 ( .C (clk), .D (new_AGEMA_signal_3695), .Q (new_AGEMA_signal_3696) ) ;
    buf_clk new_AGEMA_reg_buffer_922 ( .C (clk), .D (new_AGEMA_signal_3697), .Q (new_AGEMA_signal_3698) ) ;
    buf_clk new_AGEMA_reg_buffer_924 ( .C (clk), .D (new_AGEMA_signal_3699), .Q (new_AGEMA_signal_3700) ) ;
    buf_clk new_AGEMA_reg_buffer_926 ( .C (clk), .D (new_AGEMA_signal_3701), .Q (new_AGEMA_signal_3702) ) ;
    buf_clk new_AGEMA_reg_buffer_928 ( .C (clk), .D (new_AGEMA_signal_3703), .Q (new_AGEMA_signal_3704) ) ;
    buf_clk new_AGEMA_reg_buffer_930 ( .C (clk), .D (new_AGEMA_signal_3705), .Q (new_AGEMA_signal_3706) ) ;
    buf_clk new_AGEMA_reg_buffer_932 ( .C (clk), .D (new_AGEMA_signal_3707), .Q (new_AGEMA_signal_3708) ) ;
    buf_clk new_AGEMA_reg_buffer_934 ( .C (clk), .D (new_AGEMA_signal_3709), .Q (new_AGEMA_signal_3710) ) ;
    buf_clk new_AGEMA_reg_buffer_936 ( .C (clk), .D (new_AGEMA_signal_3711), .Q (new_AGEMA_signal_3712) ) ;
    buf_clk new_AGEMA_reg_buffer_938 ( .C (clk), .D (new_AGEMA_signal_3713), .Q (new_AGEMA_signal_3714) ) ;
    buf_clk new_AGEMA_reg_buffer_940 ( .C (clk), .D (new_AGEMA_signal_3715), .Q (new_AGEMA_signal_3716) ) ;
    buf_clk new_AGEMA_reg_buffer_942 ( .C (clk), .D (new_AGEMA_signal_3717), .Q (new_AGEMA_signal_3718) ) ;
    buf_clk new_AGEMA_reg_buffer_944 ( .C (clk), .D (new_AGEMA_signal_3719), .Q (new_AGEMA_signal_3720) ) ;
    buf_clk new_AGEMA_reg_buffer_946 ( .C (clk), .D (new_AGEMA_signal_3721), .Q (new_AGEMA_signal_3722) ) ;
    buf_clk new_AGEMA_reg_buffer_948 ( .C (clk), .D (new_AGEMA_signal_3723), .Q (new_AGEMA_signal_3724) ) ;
    buf_clk new_AGEMA_reg_buffer_950 ( .C (clk), .D (new_AGEMA_signal_3725), .Q (new_AGEMA_signal_3726) ) ;
    buf_clk new_AGEMA_reg_buffer_952 ( .C (clk), .D (new_AGEMA_signal_3727), .Q (new_AGEMA_signal_3728) ) ;
    buf_clk new_AGEMA_reg_buffer_954 ( .C (clk), .D (new_AGEMA_signal_3729), .Q (new_AGEMA_signal_3730) ) ;
    buf_clk new_AGEMA_reg_buffer_956 ( .C (clk), .D (new_AGEMA_signal_3731), .Q (new_AGEMA_signal_3732) ) ;
    buf_clk new_AGEMA_reg_buffer_958 ( .C (clk), .D (new_AGEMA_signal_3733), .Q (new_AGEMA_signal_3734) ) ;
    buf_clk new_AGEMA_reg_buffer_960 ( .C (clk), .D (new_AGEMA_signal_3735), .Q (new_AGEMA_signal_3736) ) ;
    buf_clk new_AGEMA_reg_buffer_962 ( .C (clk), .D (new_AGEMA_signal_3737), .Q (new_AGEMA_signal_3738) ) ;
    buf_clk new_AGEMA_reg_buffer_964 ( .C (clk), .D (new_AGEMA_signal_3739), .Q (new_AGEMA_signal_3740) ) ;
    buf_clk new_AGEMA_reg_buffer_966 ( .C (clk), .D (new_AGEMA_signal_3741), .Q (new_AGEMA_signal_3742) ) ;
    buf_clk new_AGEMA_reg_buffer_968 ( .C (clk), .D (new_AGEMA_signal_3743), .Q (new_AGEMA_signal_3744) ) ;
    buf_clk new_AGEMA_reg_buffer_970 ( .C (clk), .D (new_AGEMA_signal_3745), .Q (new_AGEMA_signal_3746) ) ;
    buf_clk new_AGEMA_reg_buffer_972 ( .C (clk), .D (new_AGEMA_signal_3747), .Q (new_AGEMA_signal_3748) ) ;
    buf_clk new_AGEMA_reg_buffer_974 ( .C (clk), .D (new_AGEMA_signal_3749), .Q (new_AGEMA_signal_3750) ) ;
    buf_clk new_AGEMA_reg_buffer_976 ( .C (clk), .D (new_AGEMA_signal_3751), .Q (new_AGEMA_signal_3752) ) ;
    buf_clk new_AGEMA_reg_buffer_978 ( .C (clk), .D (new_AGEMA_signal_3753), .Q (new_AGEMA_signal_3754) ) ;
    buf_clk new_AGEMA_reg_buffer_980 ( .C (clk), .D (new_AGEMA_signal_3755), .Q (new_AGEMA_signal_3756) ) ;
    buf_clk new_AGEMA_reg_buffer_982 ( .C (clk), .D (new_AGEMA_signal_3757), .Q (new_AGEMA_signal_3758) ) ;
    buf_clk new_AGEMA_reg_buffer_984 ( .C (clk), .D (new_AGEMA_signal_3759), .Q (new_AGEMA_signal_3760) ) ;
    buf_clk new_AGEMA_reg_buffer_986 ( .C (clk), .D (new_AGEMA_signal_3761), .Q (new_AGEMA_signal_3762) ) ;
    buf_clk new_AGEMA_reg_buffer_988 ( .C (clk), .D (new_AGEMA_signal_3763), .Q (new_AGEMA_signal_3764) ) ;
    buf_clk new_AGEMA_reg_buffer_990 ( .C (clk), .D (new_AGEMA_signal_3765), .Q (new_AGEMA_signal_3766) ) ;
    buf_clk new_AGEMA_reg_buffer_992 ( .C (clk), .D (new_AGEMA_signal_3767), .Q (new_AGEMA_signal_3768) ) ;
    buf_clk new_AGEMA_reg_buffer_994 ( .C (clk), .D (new_AGEMA_signal_3769), .Q (new_AGEMA_signal_3770) ) ;
    buf_clk new_AGEMA_reg_buffer_996 ( .C (clk), .D (new_AGEMA_signal_3771), .Q (new_AGEMA_signal_3772) ) ;
    buf_clk new_AGEMA_reg_buffer_998 ( .C (clk), .D (new_AGEMA_signal_3773), .Q (new_AGEMA_signal_3774) ) ;
    buf_clk new_AGEMA_reg_buffer_1000 ( .C (clk), .D (new_AGEMA_signal_3775), .Q (new_AGEMA_signal_3776) ) ;
    buf_clk new_AGEMA_reg_buffer_1002 ( .C (clk), .D (new_AGEMA_signal_3777), .Q (new_AGEMA_signal_3778) ) ;
    buf_clk new_AGEMA_reg_buffer_1004 ( .C (clk), .D (new_AGEMA_signal_3779), .Q (new_AGEMA_signal_3780) ) ;
    buf_clk new_AGEMA_reg_buffer_1006 ( .C (clk), .D (new_AGEMA_signal_3781), .Q (new_AGEMA_signal_3782) ) ;
    buf_clk new_AGEMA_reg_buffer_1008 ( .C (clk), .D (new_AGEMA_signal_3783), .Q (new_AGEMA_signal_3784) ) ;
    buf_clk new_AGEMA_reg_buffer_1010 ( .C (clk), .D (new_AGEMA_signal_3785), .Q (new_AGEMA_signal_3786) ) ;
    buf_clk new_AGEMA_reg_buffer_1012 ( .C (clk), .D (new_AGEMA_signal_3787), .Q (new_AGEMA_signal_3788) ) ;
    buf_clk new_AGEMA_reg_buffer_1014 ( .C (clk), .D (new_AGEMA_signal_3789), .Q (new_AGEMA_signal_3790) ) ;
    buf_clk new_AGEMA_reg_buffer_1016 ( .C (clk), .D (new_AGEMA_signal_3791), .Q (new_AGEMA_signal_3792) ) ;
    buf_clk new_AGEMA_reg_buffer_1018 ( .C (clk), .D (new_AGEMA_signal_3793), .Q (new_AGEMA_signal_3794) ) ;
    buf_clk new_AGEMA_reg_buffer_1020 ( .C (clk), .D (new_AGEMA_signal_3795), .Q (new_AGEMA_signal_3796) ) ;
    buf_clk new_AGEMA_reg_buffer_1022 ( .C (clk), .D (new_AGEMA_signal_3797), .Q (new_AGEMA_signal_3798) ) ;
    buf_clk new_AGEMA_reg_buffer_1024 ( .C (clk), .D (new_AGEMA_signal_3799), .Q (new_AGEMA_signal_3800) ) ;
    buf_clk new_AGEMA_reg_buffer_1026 ( .C (clk), .D (new_AGEMA_signal_3801), .Q (new_AGEMA_signal_3802) ) ;
    buf_clk new_AGEMA_reg_buffer_1028 ( .C (clk), .D (new_AGEMA_signal_3803), .Q (new_AGEMA_signal_3804) ) ;
    buf_clk new_AGEMA_reg_buffer_1030 ( .C (clk), .D (new_AGEMA_signal_3805), .Q (new_AGEMA_signal_3806) ) ;
    buf_clk new_AGEMA_reg_buffer_1032 ( .C (clk), .D (new_AGEMA_signal_3807), .Q (new_AGEMA_signal_3808) ) ;
    buf_clk new_AGEMA_reg_buffer_1034 ( .C (clk), .D (new_AGEMA_signal_3809), .Q (new_AGEMA_signal_3810) ) ;
    buf_clk new_AGEMA_reg_buffer_1036 ( .C (clk), .D (new_AGEMA_signal_3811), .Q (new_AGEMA_signal_3812) ) ;
    buf_clk new_AGEMA_reg_buffer_1038 ( .C (clk), .D (new_AGEMA_signal_3813), .Q (new_AGEMA_signal_3814) ) ;
    buf_clk new_AGEMA_reg_buffer_1040 ( .C (clk), .D (new_AGEMA_signal_3815), .Q (new_AGEMA_signal_3816) ) ;
    buf_clk new_AGEMA_reg_buffer_1042 ( .C (clk), .D (new_AGEMA_signal_3817), .Q (new_AGEMA_signal_3818) ) ;
    buf_clk new_AGEMA_reg_buffer_1044 ( .C (clk), .D (new_AGEMA_signal_3819), .Q (new_AGEMA_signal_3820) ) ;
    buf_clk new_AGEMA_reg_buffer_1046 ( .C (clk), .D (new_AGEMA_signal_3821), .Q (new_AGEMA_signal_3822) ) ;
    buf_clk new_AGEMA_reg_buffer_1048 ( .C (clk), .D (new_AGEMA_signal_3823), .Q (new_AGEMA_signal_3824) ) ;
    buf_clk new_AGEMA_reg_buffer_1050 ( .C (clk), .D (new_AGEMA_signal_3825), .Q (new_AGEMA_signal_3826) ) ;
    buf_clk new_AGEMA_reg_buffer_1052 ( .C (clk), .D (new_AGEMA_signal_3827), .Q (new_AGEMA_signal_3828) ) ;
    buf_clk new_AGEMA_reg_buffer_1054 ( .C (clk), .D (new_AGEMA_signal_3829), .Q (new_AGEMA_signal_3830) ) ;
    buf_clk new_AGEMA_reg_buffer_1056 ( .C (clk), .D (new_AGEMA_signal_3831), .Q (new_AGEMA_signal_3832) ) ;
    buf_clk new_AGEMA_reg_buffer_1058 ( .C (clk), .D (new_AGEMA_signal_3833), .Q (new_AGEMA_signal_3834) ) ;
    buf_clk new_AGEMA_reg_buffer_1060 ( .C (clk), .D (new_AGEMA_signal_3835), .Q (new_AGEMA_signal_3836) ) ;
    buf_clk new_AGEMA_reg_buffer_1062 ( .C (clk), .D (new_AGEMA_signal_3837), .Q (new_AGEMA_signal_3838) ) ;
    buf_clk new_AGEMA_reg_buffer_1064 ( .C (clk), .D (new_AGEMA_signal_3839), .Q (new_AGEMA_signal_3840) ) ;
    buf_clk new_AGEMA_reg_buffer_1066 ( .C (clk), .D (new_AGEMA_signal_3841), .Q (new_AGEMA_signal_3842) ) ;
    buf_clk new_AGEMA_reg_buffer_1068 ( .C (clk), .D (new_AGEMA_signal_3843), .Q (new_AGEMA_signal_3844) ) ;
    buf_clk new_AGEMA_reg_buffer_1070 ( .C (clk), .D (new_AGEMA_signal_3845), .Q (new_AGEMA_signal_3846) ) ;
    buf_clk new_AGEMA_reg_buffer_1072 ( .C (clk), .D (new_AGEMA_signal_3847), .Q (new_AGEMA_signal_3848) ) ;
    buf_clk new_AGEMA_reg_buffer_1074 ( .C (clk), .D (new_AGEMA_signal_3849), .Q (new_AGEMA_signal_3850) ) ;
    buf_clk new_AGEMA_reg_buffer_1076 ( .C (clk), .D (new_AGEMA_signal_3851), .Q (new_AGEMA_signal_3852) ) ;
    buf_clk new_AGEMA_reg_buffer_1078 ( .C (clk), .D (new_AGEMA_signal_3853), .Q (new_AGEMA_signal_3854) ) ;
    buf_clk new_AGEMA_reg_buffer_1080 ( .C (clk), .D (new_AGEMA_signal_3855), .Q (new_AGEMA_signal_3856) ) ;
    buf_clk new_AGEMA_reg_buffer_1082 ( .C (clk), .D (new_AGEMA_signal_3857), .Q (new_AGEMA_signal_3858) ) ;
    buf_clk new_AGEMA_reg_buffer_1084 ( .C (clk), .D (new_AGEMA_signal_3859), .Q (new_AGEMA_signal_3860) ) ;
    buf_clk new_AGEMA_reg_buffer_1086 ( .C (clk), .D (new_AGEMA_signal_3861), .Q (new_AGEMA_signal_3862) ) ;
    buf_clk new_AGEMA_reg_buffer_1088 ( .C (clk), .D (new_AGEMA_signal_3863), .Q (new_AGEMA_signal_3864) ) ;
    buf_clk new_AGEMA_reg_buffer_1090 ( .C (clk), .D (new_AGEMA_signal_3865), .Q (new_AGEMA_signal_3866) ) ;
    buf_clk new_AGEMA_reg_buffer_1092 ( .C (clk), .D (new_AGEMA_signal_3867), .Q (new_AGEMA_signal_3868) ) ;
    buf_clk new_AGEMA_reg_buffer_1094 ( .C (clk), .D (new_AGEMA_signal_3869), .Q (new_AGEMA_signal_3870) ) ;
    buf_clk new_AGEMA_reg_buffer_1096 ( .C (clk), .D (new_AGEMA_signal_3871), .Q (new_AGEMA_signal_3872) ) ;
    buf_clk new_AGEMA_reg_buffer_1098 ( .C (clk), .D (new_AGEMA_signal_3873), .Q (new_AGEMA_signal_3874) ) ;
    buf_clk new_AGEMA_reg_buffer_1100 ( .C (clk), .D (new_AGEMA_signal_3875), .Q (new_AGEMA_signal_3876) ) ;
    buf_clk new_AGEMA_reg_buffer_1102 ( .C (clk), .D (new_AGEMA_signal_3877), .Q (new_AGEMA_signal_3878) ) ;
    buf_clk new_AGEMA_reg_buffer_1104 ( .C (clk), .D (new_AGEMA_signal_3879), .Q (new_AGEMA_signal_3880) ) ;
    buf_clk new_AGEMA_reg_buffer_1106 ( .C (clk), .D (new_AGEMA_signal_3881), .Q (new_AGEMA_signal_3882) ) ;
    buf_clk new_AGEMA_reg_buffer_1108 ( .C (clk), .D (new_AGEMA_signal_3883), .Q (new_AGEMA_signal_3884) ) ;
    buf_clk new_AGEMA_reg_buffer_1110 ( .C (clk), .D (new_AGEMA_signal_3885), .Q (new_AGEMA_signal_3886) ) ;
    buf_clk new_AGEMA_reg_buffer_1112 ( .C (clk), .D (new_AGEMA_signal_3887), .Q (new_AGEMA_signal_3888) ) ;
    buf_clk new_AGEMA_reg_buffer_1114 ( .C (clk), .D (new_AGEMA_signal_3889), .Q (new_AGEMA_signal_3890) ) ;
    buf_clk new_AGEMA_reg_buffer_1116 ( .C (clk), .D (new_AGEMA_signal_3891), .Q (new_AGEMA_signal_3892) ) ;
    buf_clk new_AGEMA_reg_buffer_1118 ( .C (clk), .D (new_AGEMA_signal_3893), .Q (new_AGEMA_signal_3894) ) ;
    buf_clk new_AGEMA_reg_buffer_1120 ( .C (clk), .D (new_AGEMA_signal_3895), .Q (new_AGEMA_signal_3896) ) ;
    buf_clk new_AGEMA_reg_buffer_1122 ( .C (clk), .D (new_AGEMA_signal_3897), .Q (new_AGEMA_signal_3898) ) ;
    buf_clk new_AGEMA_reg_buffer_1124 ( .C (clk), .D (new_AGEMA_signal_3899), .Q (new_AGEMA_signal_3900) ) ;
    buf_clk new_AGEMA_reg_buffer_1126 ( .C (clk), .D (new_AGEMA_signal_3901), .Q (new_AGEMA_signal_3902) ) ;
    buf_clk new_AGEMA_reg_buffer_1128 ( .C (clk), .D (new_AGEMA_signal_3903), .Q (new_AGEMA_signal_3904) ) ;
    buf_clk new_AGEMA_reg_buffer_1130 ( .C (clk), .D (new_AGEMA_signal_3905), .Q (new_AGEMA_signal_3906) ) ;
    buf_clk new_AGEMA_reg_buffer_1132 ( .C (clk), .D (new_AGEMA_signal_3907), .Q (new_AGEMA_signal_3908) ) ;
    buf_clk new_AGEMA_reg_buffer_1134 ( .C (clk), .D (new_AGEMA_signal_3909), .Q (new_AGEMA_signal_3910) ) ;
    buf_clk new_AGEMA_reg_buffer_1136 ( .C (clk), .D (new_AGEMA_signal_3911), .Q (new_AGEMA_signal_3912) ) ;
    buf_clk new_AGEMA_reg_buffer_1138 ( .C (clk), .D (new_AGEMA_signal_3913), .Q (new_AGEMA_signal_3914) ) ;
    buf_clk new_AGEMA_reg_buffer_1140 ( .C (clk), .D (new_AGEMA_signal_3915), .Q (new_AGEMA_signal_3916) ) ;
    buf_clk new_AGEMA_reg_buffer_1142 ( .C (clk), .D (new_AGEMA_signal_3917), .Q (new_AGEMA_signal_3918) ) ;
    buf_clk new_AGEMA_reg_buffer_1144 ( .C (clk), .D (new_AGEMA_signal_3919), .Q (new_AGEMA_signal_3920) ) ;
    buf_clk new_AGEMA_reg_buffer_1146 ( .C (clk), .D (new_AGEMA_signal_3921), .Q (new_AGEMA_signal_3922) ) ;
    buf_clk new_AGEMA_reg_buffer_1148 ( .C (clk), .D (new_AGEMA_signal_3923), .Q (new_AGEMA_signal_3924) ) ;
    buf_clk new_AGEMA_reg_buffer_1150 ( .C (clk), .D (new_AGEMA_signal_3925), .Q (new_AGEMA_signal_3926) ) ;
    buf_clk new_AGEMA_reg_buffer_1152 ( .C (clk), .D (new_AGEMA_signal_3927), .Q (new_AGEMA_signal_3928) ) ;
    buf_clk new_AGEMA_reg_buffer_1154 ( .C (clk), .D (new_AGEMA_signal_3929), .Q (new_AGEMA_signal_3930) ) ;
    buf_clk new_AGEMA_reg_buffer_1156 ( .C (clk), .D (new_AGEMA_signal_3931), .Q (new_AGEMA_signal_3932) ) ;
    buf_clk new_AGEMA_reg_buffer_1158 ( .C (clk), .D (new_AGEMA_signal_3933), .Q (new_AGEMA_signal_3934) ) ;
    buf_clk new_AGEMA_reg_buffer_1160 ( .C (clk), .D (new_AGEMA_signal_3935), .Q (new_AGEMA_signal_3936) ) ;
    buf_clk new_AGEMA_reg_buffer_1162 ( .C (clk), .D (new_AGEMA_signal_3937), .Q (new_AGEMA_signal_3938) ) ;
    buf_clk new_AGEMA_reg_buffer_1164 ( .C (clk), .D (new_AGEMA_signal_3939), .Q (new_AGEMA_signal_3940) ) ;
    buf_clk new_AGEMA_reg_buffer_1166 ( .C (clk), .D (new_AGEMA_signal_3941), .Q (new_AGEMA_signal_3942) ) ;
    buf_clk new_AGEMA_reg_buffer_1168 ( .C (clk), .D (new_AGEMA_signal_3943), .Q (new_AGEMA_signal_3944) ) ;
    buf_clk new_AGEMA_reg_buffer_1170 ( .C (clk), .D (new_AGEMA_signal_3945), .Q (new_AGEMA_signal_3946) ) ;
    buf_clk new_AGEMA_reg_buffer_1172 ( .C (clk), .D (new_AGEMA_signal_3947), .Q (new_AGEMA_signal_3948) ) ;
    buf_clk new_AGEMA_reg_buffer_1174 ( .C (clk), .D (new_AGEMA_signal_3949), .Q (new_AGEMA_signal_3950) ) ;
    buf_clk new_AGEMA_reg_buffer_1176 ( .C (clk), .D (new_AGEMA_signal_3951), .Q (new_AGEMA_signal_3952) ) ;
    buf_clk new_AGEMA_reg_buffer_1178 ( .C (clk), .D (new_AGEMA_signal_3953), .Q (new_AGEMA_signal_3954) ) ;
    buf_clk new_AGEMA_reg_buffer_1180 ( .C (clk), .D (new_AGEMA_signal_3955), .Q (new_AGEMA_signal_3956) ) ;
    buf_clk new_AGEMA_reg_buffer_1182 ( .C (clk), .D (new_AGEMA_signal_3957), .Q (new_AGEMA_signal_3958) ) ;
    buf_clk new_AGEMA_reg_buffer_1184 ( .C (clk), .D (new_AGEMA_signal_3959), .Q (new_AGEMA_signal_3960) ) ;
    buf_clk new_AGEMA_reg_buffer_1186 ( .C (clk), .D (new_AGEMA_signal_3961), .Q (new_AGEMA_signal_3962) ) ;
    buf_clk new_AGEMA_reg_buffer_1188 ( .C (clk), .D (new_AGEMA_signal_3963), .Q (new_AGEMA_signal_3964) ) ;
    buf_clk new_AGEMA_reg_buffer_1190 ( .C (clk), .D (new_AGEMA_signal_3965), .Q (new_AGEMA_signal_3966) ) ;
    buf_clk new_AGEMA_reg_buffer_1192 ( .C (clk), .D (new_AGEMA_signal_3967), .Q (new_AGEMA_signal_3968) ) ;
    buf_clk new_AGEMA_reg_buffer_1194 ( .C (clk), .D (new_AGEMA_signal_3969), .Q (new_AGEMA_signal_3970) ) ;
    buf_clk new_AGEMA_reg_buffer_1196 ( .C (clk), .D (new_AGEMA_signal_3971), .Q (new_AGEMA_signal_3972) ) ;
    buf_clk new_AGEMA_reg_buffer_1198 ( .C (clk), .D (new_AGEMA_signal_3973), .Q (new_AGEMA_signal_3974) ) ;
    buf_clk new_AGEMA_reg_buffer_1200 ( .C (clk), .D (new_AGEMA_signal_3975), .Q (new_AGEMA_signal_3976) ) ;
    buf_clk new_AGEMA_reg_buffer_1202 ( .C (clk), .D (new_AGEMA_signal_3977), .Q (new_AGEMA_signal_3978) ) ;
    buf_clk new_AGEMA_reg_buffer_1204 ( .C (clk), .D (new_AGEMA_signal_3979), .Q (new_AGEMA_signal_3980) ) ;
    buf_clk new_AGEMA_reg_buffer_1210 ( .C (clk), .D (new_AGEMA_signal_3985), .Q (new_AGEMA_signal_3986) ) ;
    buf_clk new_AGEMA_reg_buffer_1216 ( .C (clk), .D (new_AGEMA_signal_3991), .Q (new_AGEMA_signal_3992) ) ;
    buf_clk new_AGEMA_reg_buffer_1222 ( .C (clk), .D (new_AGEMA_signal_3997), .Q (new_AGEMA_signal_3998) ) ;
    buf_clk new_AGEMA_reg_buffer_1228 ( .C (clk), .D (new_AGEMA_signal_4003), .Q (new_AGEMA_signal_4004) ) ;
    buf_clk new_AGEMA_reg_buffer_1234 ( .C (clk), .D (new_AGEMA_signal_4009), .Q (new_AGEMA_signal_4010) ) ;
    buf_clk new_AGEMA_reg_buffer_1240 ( .C (clk), .D (new_AGEMA_signal_4015), .Q (new_AGEMA_signal_4016) ) ;
    buf_clk new_AGEMA_reg_buffer_1246 ( .C (clk), .D (new_AGEMA_signal_4021), .Q (new_AGEMA_signal_4022) ) ;
    buf_clk new_AGEMA_reg_buffer_1252 ( .C (clk), .D (new_AGEMA_signal_4027), .Q (new_AGEMA_signal_4028) ) ;
    buf_clk new_AGEMA_reg_buffer_1258 ( .C (clk), .D (new_AGEMA_signal_4033), .Q (new_AGEMA_signal_4034) ) ;
    buf_clk new_AGEMA_reg_buffer_1264 ( .C (clk), .D (new_AGEMA_signal_4039), .Q (new_AGEMA_signal_4040) ) ;
    buf_clk new_AGEMA_reg_buffer_1270 ( .C (clk), .D (new_AGEMA_signal_4045), .Q (new_AGEMA_signal_4046) ) ;
    buf_clk new_AGEMA_reg_buffer_1276 ( .C (clk), .D (new_AGEMA_signal_4051), .Q (new_AGEMA_signal_4052) ) ;
    buf_clk new_AGEMA_reg_buffer_1282 ( .C (clk), .D (new_AGEMA_signal_4057), .Q (new_AGEMA_signal_4058) ) ;
    buf_clk new_AGEMA_reg_buffer_1288 ( .C (clk), .D (new_AGEMA_signal_4063), .Q (new_AGEMA_signal_4064) ) ;
    buf_clk new_AGEMA_reg_buffer_1294 ( .C (clk), .D (new_AGEMA_signal_4069), .Q (new_AGEMA_signal_4070) ) ;
    buf_clk new_AGEMA_reg_buffer_1300 ( .C (clk), .D (new_AGEMA_signal_4075), .Q (new_AGEMA_signal_4076) ) ;
    buf_clk new_AGEMA_reg_buffer_1306 ( .C (clk), .D (new_AGEMA_signal_4081), .Q (new_AGEMA_signal_4082) ) ;
    buf_clk new_AGEMA_reg_buffer_1312 ( .C (clk), .D (new_AGEMA_signal_4087), .Q (new_AGEMA_signal_4088) ) ;
    buf_clk new_AGEMA_reg_buffer_1318 ( .C (clk), .D (new_AGEMA_signal_4093), .Q (new_AGEMA_signal_4094) ) ;
    buf_clk new_AGEMA_reg_buffer_1324 ( .C (clk), .D (new_AGEMA_signal_4099), .Q (new_AGEMA_signal_4100) ) ;
    buf_clk new_AGEMA_reg_buffer_1330 ( .C (clk), .D (new_AGEMA_signal_4105), .Q (new_AGEMA_signal_4106) ) ;
    buf_clk new_AGEMA_reg_buffer_1336 ( .C (clk), .D (new_AGEMA_signal_4111), .Q (new_AGEMA_signal_4112) ) ;
    buf_clk new_AGEMA_reg_buffer_1342 ( .C (clk), .D (new_AGEMA_signal_4117), .Q (new_AGEMA_signal_4118) ) ;
    buf_clk new_AGEMA_reg_buffer_1348 ( .C (clk), .D (new_AGEMA_signal_4123), .Q (new_AGEMA_signal_4124) ) ;
    buf_clk new_AGEMA_reg_buffer_1354 ( .C (clk), .D (new_AGEMA_signal_4129), .Q (new_AGEMA_signal_4130) ) ;
    buf_clk new_AGEMA_reg_buffer_1360 ( .C (clk), .D (new_AGEMA_signal_4135), .Q (new_AGEMA_signal_4136) ) ;
    buf_clk new_AGEMA_reg_buffer_1366 ( .C (clk), .D (new_AGEMA_signal_4141), .Q (new_AGEMA_signal_4142) ) ;
    buf_clk new_AGEMA_reg_buffer_1372 ( .C (clk), .D (new_AGEMA_signal_4147), .Q (new_AGEMA_signal_4148) ) ;
    buf_clk new_AGEMA_reg_buffer_1378 ( .C (clk), .D (new_AGEMA_signal_4153), .Q (new_AGEMA_signal_4154) ) ;
    buf_clk new_AGEMA_reg_buffer_1384 ( .C (clk), .D (new_AGEMA_signal_4159), .Q (new_AGEMA_signal_4160) ) ;
    buf_clk new_AGEMA_reg_buffer_1390 ( .C (clk), .D (new_AGEMA_signal_4165), .Q (new_AGEMA_signal_4166) ) ;
    buf_clk new_AGEMA_reg_buffer_1396 ( .C (clk), .D (new_AGEMA_signal_4171), .Q (new_AGEMA_signal_4172) ) ;
    buf_clk new_AGEMA_reg_buffer_1402 ( .C (clk), .D (new_AGEMA_signal_4177), .Q (new_AGEMA_signal_4178) ) ;
    buf_clk new_AGEMA_reg_buffer_1408 ( .C (clk), .D (new_AGEMA_signal_4183), .Q (new_AGEMA_signal_4184) ) ;
    buf_clk new_AGEMA_reg_buffer_1414 ( .C (clk), .D (new_AGEMA_signal_4189), .Q (new_AGEMA_signal_4190) ) ;
    buf_clk new_AGEMA_reg_buffer_1420 ( .C (clk), .D (new_AGEMA_signal_4195), .Q (new_AGEMA_signal_4196) ) ;
    buf_clk new_AGEMA_reg_buffer_1426 ( .C (clk), .D (new_AGEMA_signal_4201), .Q (new_AGEMA_signal_4202) ) ;
    buf_clk new_AGEMA_reg_buffer_1432 ( .C (clk), .D (new_AGEMA_signal_4207), .Q (new_AGEMA_signal_4208) ) ;
    buf_clk new_AGEMA_reg_buffer_1438 ( .C (clk), .D (new_AGEMA_signal_4213), .Q (new_AGEMA_signal_4214) ) ;
    buf_clk new_AGEMA_reg_buffer_1444 ( .C (clk), .D (new_AGEMA_signal_4219), .Q (new_AGEMA_signal_4220) ) ;
    buf_clk new_AGEMA_reg_buffer_1450 ( .C (clk), .D (new_AGEMA_signal_4225), .Q (new_AGEMA_signal_4226) ) ;
    buf_clk new_AGEMA_reg_buffer_1456 ( .C (clk), .D (new_AGEMA_signal_4231), .Q (new_AGEMA_signal_4232) ) ;
    buf_clk new_AGEMA_reg_buffer_1462 ( .C (clk), .D (new_AGEMA_signal_4237), .Q (new_AGEMA_signal_4238) ) ;
    buf_clk new_AGEMA_reg_buffer_1468 ( .C (clk), .D (new_AGEMA_signal_4243), .Q (new_AGEMA_signal_4244) ) ;
    buf_clk new_AGEMA_reg_buffer_1474 ( .C (clk), .D (new_AGEMA_signal_4249), .Q (new_AGEMA_signal_4250) ) ;
    buf_clk new_AGEMA_reg_buffer_1480 ( .C (clk), .D (new_AGEMA_signal_4255), .Q (new_AGEMA_signal_4256) ) ;
    buf_clk new_AGEMA_reg_buffer_1486 ( .C (clk), .D (new_AGEMA_signal_4261), .Q (new_AGEMA_signal_4262) ) ;
    buf_clk new_AGEMA_reg_buffer_1492 ( .C (clk), .D (new_AGEMA_signal_4267), .Q (new_AGEMA_signal_4268) ) ;
    buf_clk new_AGEMA_reg_buffer_1498 ( .C (clk), .D (new_AGEMA_signal_4273), .Q (new_AGEMA_signal_4274) ) ;
    buf_clk new_AGEMA_reg_buffer_1504 ( .C (clk), .D (new_AGEMA_signal_4279), .Q (new_AGEMA_signal_4280) ) ;
    buf_clk new_AGEMA_reg_buffer_1510 ( .C (clk), .D (new_AGEMA_signal_4285), .Q (new_AGEMA_signal_4286) ) ;
    buf_clk new_AGEMA_reg_buffer_1516 ( .C (clk), .D (new_AGEMA_signal_4291), .Q (new_AGEMA_signal_4292) ) ;
    buf_clk new_AGEMA_reg_buffer_1522 ( .C (clk), .D (new_AGEMA_signal_4297), .Q (new_AGEMA_signal_4298) ) ;
    buf_clk new_AGEMA_reg_buffer_1528 ( .C (clk), .D (new_AGEMA_signal_4303), .Q (new_AGEMA_signal_4304) ) ;
    buf_clk new_AGEMA_reg_buffer_1534 ( .C (clk), .D (new_AGEMA_signal_4309), .Q (new_AGEMA_signal_4310) ) ;
    buf_clk new_AGEMA_reg_buffer_1540 ( .C (clk), .D (new_AGEMA_signal_4315), .Q (new_AGEMA_signal_4316) ) ;
    buf_clk new_AGEMA_reg_buffer_1546 ( .C (clk), .D (new_AGEMA_signal_4321), .Q (new_AGEMA_signal_4322) ) ;
    buf_clk new_AGEMA_reg_buffer_1552 ( .C (clk), .D (new_AGEMA_signal_4327), .Q (new_AGEMA_signal_4328) ) ;
    buf_clk new_AGEMA_reg_buffer_1558 ( .C (clk), .D (new_AGEMA_signal_4333), .Q (new_AGEMA_signal_4334) ) ;
    buf_clk new_AGEMA_reg_buffer_1564 ( .C (clk), .D (new_AGEMA_signal_4339), .Q (new_AGEMA_signal_4340) ) ;
    buf_clk new_AGEMA_reg_buffer_1570 ( .C (clk), .D (new_AGEMA_signal_4345), .Q (new_AGEMA_signal_4346) ) ;
    buf_clk new_AGEMA_reg_buffer_1576 ( .C (clk), .D (new_AGEMA_signal_4351), .Q (new_AGEMA_signal_4352) ) ;
    buf_clk new_AGEMA_reg_buffer_1582 ( .C (clk), .D (new_AGEMA_signal_4357), .Q (new_AGEMA_signal_4358) ) ;
    buf_clk new_AGEMA_reg_buffer_1588 ( .C (clk), .D (new_AGEMA_signal_4363), .Q (new_AGEMA_signal_4364) ) ;
    buf_clk new_AGEMA_reg_buffer_1594 ( .C (clk), .D (new_AGEMA_signal_4369), .Q (new_AGEMA_signal_4370) ) ;
    buf_clk new_AGEMA_reg_buffer_1600 ( .C (clk), .D (new_AGEMA_signal_4375), .Q (new_AGEMA_signal_4376) ) ;
    buf_clk new_AGEMA_reg_buffer_1606 ( .C (clk), .D (new_AGEMA_signal_4381), .Q (new_AGEMA_signal_4382) ) ;
    buf_clk new_AGEMA_reg_buffer_1612 ( .C (clk), .D (new_AGEMA_signal_4387), .Q (new_AGEMA_signal_4388) ) ;
    buf_clk new_AGEMA_reg_buffer_1618 ( .C (clk), .D (new_AGEMA_signal_4393), .Q (new_AGEMA_signal_4394) ) ;
    buf_clk new_AGEMA_reg_buffer_1624 ( .C (clk), .D (new_AGEMA_signal_4399), .Q (new_AGEMA_signal_4400) ) ;
    buf_clk new_AGEMA_reg_buffer_1630 ( .C (clk), .D (new_AGEMA_signal_4405), .Q (new_AGEMA_signal_4406) ) ;
    buf_clk new_AGEMA_reg_buffer_1636 ( .C (clk), .D (new_AGEMA_signal_4411), .Q (new_AGEMA_signal_4412) ) ;
    buf_clk new_AGEMA_reg_buffer_1642 ( .C (clk), .D (new_AGEMA_signal_4417), .Q (new_AGEMA_signal_4418) ) ;
    buf_clk new_AGEMA_reg_buffer_1648 ( .C (clk), .D (new_AGEMA_signal_4423), .Q (new_AGEMA_signal_4424) ) ;
    buf_clk new_AGEMA_reg_buffer_1654 ( .C (clk), .D (new_AGEMA_signal_4429), .Q (new_AGEMA_signal_4430) ) ;
    buf_clk new_AGEMA_reg_buffer_1660 ( .C (clk), .D (new_AGEMA_signal_4435), .Q (new_AGEMA_signal_4436) ) ;
    buf_clk new_AGEMA_reg_buffer_1666 ( .C (clk), .D (new_AGEMA_signal_4441), .Q (new_AGEMA_signal_4442) ) ;
    buf_clk new_AGEMA_reg_buffer_1672 ( .C (clk), .D (new_AGEMA_signal_4447), .Q (new_AGEMA_signal_4448) ) ;
    buf_clk new_AGEMA_reg_buffer_1678 ( .C (clk), .D (new_AGEMA_signal_4453), .Q (new_AGEMA_signal_4454) ) ;
    buf_clk new_AGEMA_reg_buffer_1684 ( .C (clk), .D (new_AGEMA_signal_4459), .Q (new_AGEMA_signal_4460) ) ;
    buf_clk new_AGEMA_reg_buffer_1690 ( .C (clk), .D (new_AGEMA_signal_4465), .Q (new_AGEMA_signal_4466) ) ;
    buf_clk new_AGEMA_reg_buffer_1696 ( .C (clk), .D (new_AGEMA_signal_4471), .Q (new_AGEMA_signal_4472) ) ;
    buf_clk new_AGEMA_reg_buffer_1702 ( .C (clk), .D (new_AGEMA_signal_4477), .Q (new_AGEMA_signal_4478) ) ;
    buf_clk new_AGEMA_reg_buffer_1708 ( .C (clk), .D (new_AGEMA_signal_4483), .Q (new_AGEMA_signal_4484) ) ;
    buf_clk new_AGEMA_reg_buffer_1714 ( .C (clk), .D (new_AGEMA_signal_4489), .Q (new_AGEMA_signal_4490) ) ;
    buf_clk new_AGEMA_reg_buffer_1720 ( .C (clk), .D (new_AGEMA_signal_4495), .Q (new_AGEMA_signal_4496) ) ;
    buf_clk new_AGEMA_reg_buffer_1726 ( .C (clk), .D (new_AGEMA_signal_4501), .Q (new_AGEMA_signal_4502) ) ;
    buf_clk new_AGEMA_reg_buffer_1732 ( .C (clk), .D (new_AGEMA_signal_4507), .Q (new_AGEMA_signal_4508) ) ;
    buf_clk new_AGEMA_reg_buffer_1738 ( .C (clk), .D (new_AGEMA_signal_4513), .Q (new_AGEMA_signal_4514) ) ;
    buf_clk new_AGEMA_reg_buffer_1744 ( .C (clk), .D (new_AGEMA_signal_4519), .Q (new_AGEMA_signal_4520) ) ;
    buf_clk new_AGEMA_reg_buffer_1750 ( .C (clk), .D (new_AGEMA_signal_4525), .Q (new_AGEMA_signal_4526) ) ;
    buf_clk new_AGEMA_reg_buffer_1756 ( .C (clk), .D (new_AGEMA_signal_4531), .Q (new_AGEMA_signal_4532) ) ;
    buf_clk new_AGEMA_reg_buffer_1762 ( .C (clk), .D (new_AGEMA_signal_4537), .Q (new_AGEMA_signal_4538) ) ;
    buf_clk new_AGEMA_reg_buffer_1768 ( .C (clk), .D (new_AGEMA_signal_4543), .Q (new_AGEMA_signal_4544) ) ;
    buf_clk new_AGEMA_reg_buffer_1774 ( .C (clk), .D (new_AGEMA_signal_4549), .Q (new_AGEMA_signal_4550) ) ;
    buf_clk new_AGEMA_reg_buffer_1780 ( .C (clk), .D (new_AGEMA_signal_4555), .Q (new_AGEMA_signal_4556) ) ;
    buf_clk new_AGEMA_reg_buffer_1786 ( .C (clk), .D (new_AGEMA_signal_4561), .Q (new_AGEMA_signal_4562) ) ;
    buf_clk new_AGEMA_reg_buffer_1792 ( .C (clk), .D (new_AGEMA_signal_4567), .Q (new_AGEMA_signal_4568) ) ;
    buf_clk new_AGEMA_reg_buffer_1798 ( .C (clk), .D (new_AGEMA_signal_4573), .Q (new_AGEMA_signal_4574) ) ;
    buf_clk new_AGEMA_reg_buffer_1804 ( .C (clk), .D (new_AGEMA_signal_4579), .Q (new_AGEMA_signal_4580) ) ;
    buf_clk new_AGEMA_reg_buffer_1810 ( .C (clk), .D (new_AGEMA_signal_4585), .Q (new_AGEMA_signal_4586) ) ;
    buf_clk new_AGEMA_reg_buffer_1816 ( .C (clk), .D (new_AGEMA_signal_4591), .Q (new_AGEMA_signal_4592) ) ;
    buf_clk new_AGEMA_reg_buffer_1822 ( .C (clk), .D (new_AGEMA_signal_4597), .Q (new_AGEMA_signal_4598) ) ;
    buf_clk new_AGEMA_reg_buffer_1828 ( .C (clk), .D (new_AGEMA_signal_4603), .Q (new_AGEMA_signal_4604) ) ;
    buf_clk new_AGEMA_reg_buffer_1834 ( .C (clk), .D (new_AGEMA_signal_4609), .Q (new_AGEMA_signal_4610) ) ;
    buf_clk new_AGEMA_reg_buffer_1840 ( .C (clk), .D (new_AGEMA_signal_4615), .Q (new_AGEMA_signal_4616) ) ;
    buf_clk new_AGEMA_reg_buffer_1846 ( .C (clk), .D (new_AGEMA_signal_4621), .Q (new_AGEMA_signal_4622) ) ;
    buf_clk new_AGEMA_reg_buffer_1852 ( .C (clk), .D (new_AGEMA_signal_4627), .Q (new_AGEMA_signal_4628) ) ;
    buf_clk new_AGEMA_reg_buffer_1858 ( .C (clk), .D (new_AGEMA_signal_4633), .Q (new_AGEMA_signal_4634) ) ;
    buf_clk new_AGEMA_reg_buffer_1864 ( .C (clk), .D (new_AGEMA_signal_4639), .Q (new_AGEMA_signal_4640) ) ;
    buf_clk new_AGEMA_reg_buffer_1870 ( .C (clk), .D (new_AGEMA_signal_4645), .Q (new_AGEMA_signal_4646) ) ;
    buf_clk new_AGEMA_reg_buffer_1876 ( .C (clk), .D (new_AGEMA_signal_4651), .Q (new_AGEMA_signal_4652) ) ;
    buf_clk new_AGEMA_reg_buffer_1882 ( .C (clk), .D (new_AGEMA_signal_4657), .Q (new_AGEMA_signal_4658) ) ;
    buf_clk new_AGEMA_reg_buffer_1888 ( .C (clk), .D (new_AGEMA_signal_4663), .Q (new_AGEMA_signal_4664) ) ;
    buf_clk new_AGEMA_reg_buffer_1894 ( .C (clk), .D (new_AGEMA_signal_4669), .Q (new_AGEMA_signal_4670) ) ;
    buf_clk new_AGEMA_reg_buffer_1900 ( .C (clk), .D (new_AGEMA_signal_4675), .Q (new_AGEMA_signal_4676) ) ;
    buf_clk new_AGEMA_reg_buffer_1906 ( .C (clk), .D (new_AGEMA_signal_4681), .Q (new_AGEMA_signal_4682) ) ;
    buf_clk new_AGEMA_reg_buffer_1912 ( .C (clk), .D (new_AGEMA_signal_4687), .Q (new_AGEMA_signal_4688) ) ;
    buf_clk new_AGEMA_reg_buffer_1918 ( .C (clk), .D (new_AGEMA_signal_4693), .Q (new_AGEMA_signal_4694) ) ;
    buf_clk new_AGEMA_reg_buffer_1924 ( .C (clk), .D (new_AGEMA_signal_4699), .Q (new_AGEMA_signal_4700) ) ;
    buf_clk new_AGEMA_reg_buffer_1930 ( .C (clk), .D (new_AGEMA_signal_4705), .Q (new_AGEMA_signal_4706) ) ;
    buf_clk new_AGEMA_reg_buffer_1936 ( .C (clk), .D (new_AGEMA_signal_4711), .Q (new_AGEMA_signal_4712) ) ;
    buf_clk new_AGEMA_reg_buffer_1942 ( .C (clk), .D (new_AGEMA_signal_4717), .Q (new_AGEMA_signal_4718) ) ;
    buf_clk new_AGEMA_reg_buffer_1948 ( .C (clk), .D (new_AGEMA_signal_4723), .Q (new_AGEMA_signal_4724) ) ;
    buf_clk new_AGEMA_reg_buffer_1954 ( .C (clk), .D (new_AGEMA_signal_4729), .Q (new_AGEMA_signal_4730) ) ;
    buf_clk new_AGEMA_reg_buffer_1960 ( .C (clk), .D (new_AGEMA_signal_4735), .Q (new_AGEMA_signal_4736) ) ;
    buf_clk new_AGEMA_reg_buffer_1966 ( .C (clk), .D (new_AGEMA_signal_4741), .Q (new_AGEMA_signal_4742) ) ;
    buf_clk new_AGEMA_reg_buffer_1972 ( .C (clk), .D (new_AGEMA_signal_4747), .Q (new_AGEMA_signal_4748) ) ;
    buf_clk new_AGEMA_reg_buffer_1978 ( .C (clk), .D (new_AGEMA_signal_4753), .Q (new_AGEMA_signal_4754) ) ;
    buf_clk new_AGEMA_reg_buffer_1984 ( .C (clk), .D (new_AGEMA_signal_4759), .Q (new_AGEMA_signal_4760) ) ;
    buf_clk new_AGEMA_reg_buffer_1990 ( .C (clk), .D (new_AGEMA_signal_4765), .Q (new_AGEMA_signal_4766) ) ;
    buf_clk new_AGEMA_reg_buffer_1996 ( .C (clk), .D (new_AGEMA_signal_4771), .Q (new_AGEMA_signal_4772) ) ;
    buf_clk new_AGEMA_reg_buffer_2002 ( .C (clk), .D (new_AGEMA_signal_4777), .Q (new_AGEMA_signal_4778) ) ;
    buf_clk new_AGEMA_reg_buffer_2008 ( .C (clk), .D (new_AGEMA_signal_4783), .Q (new_AGEMA_signal_4784) ) ;
    buf_clk new_AGEMA_reg_buffer_2014 ( .C (clk), .D (new_AGEMA_signal_4789), .Q (new_AGEMA_signal_4790) ) ;
    buf_clk new_AGEMA_reg_buffer_2020 ( .C (clk), .D (new_AGEMA_signal_4795), .Q (new_AGEMA_signal_4796) ) ;
    buf_clk new_AGEMA_reg_buffer_2026 ( .C (clk), .D (new_AGEMA_signal_4801), .Q (new_AGEMA_signal_4802) ) ;
    buf_clk new_AGEMA_reg_buffer_2032 ( .C (clk), .D (new_AGEMA_signal_4807), .Q (new_AGEMA_signal_4808) ) ;
    buf_clk new_AGEMA_reg_buffer_2038 ( .C (clk), .D (new_AGEMA_signal_4813), .Q (new_AGEMA_signal_4814) ) ;
    buf_clk new_AGEMA_reg_buffer_2044 ( .C (clk), .D (new_AGEMA_signal_4819), .Q (new_AGEMA_signal_4820) ) ;
    buf_clk new_AGEMA_reg_buffer_2050 ( .C (clk), .D (new_AGEMA_signal_4825), .Q (new_AGEMA_signal_4826) ) ;
    buf_clk new_AGEMA_reg_buffer_2056 ( .C (clk), .D (new_AGEMA_signal_4831), .Q (new_AGEMA_signal_4832) ) ;
    buf_clk new_AGEMA_reg_buffer_2062 ( .C (clk), .D (new_AGEMA_signal_4837), .Q (new_AGEMA_signal_4838) ) ;
    buf_clk new_AGEMA_reg_buffer_2068 ( .C (clk), .D (new_AGEMA_signal_4843), .Q (new_AGEMA_signal_4844) ) ;
    buf_clk new_AGEMA_reg_buffer_2074 ( .C (clk), .D (new_AGEMA_signal_4849), .Q (new_AGEMA_signal_4850) ) ;
    buf_clk new_AGEMA_reg_buffer_2080 ( .C (clk), .D (new_AGEMA_signal_4855), .Q (new_AGEMA_signal_4856) ) ;
    buf_clk new_AGEMA_reg_buffer_2086 ( .C (clk), .D (new_AGEMA_signal_4861), .Q (new_AGEMA_signal_4862) ) ;
    buf_clk new_AGEMA_reg_buffer_2092 ( .C (clk), .D (new_AGEMA_signal_4867), .Q (new_AGEMA_signal_4868) ) ;
    buf_clk new_AGEMA_reg_buffer_2098 ( .C (clk), .D (new_AGEMA_signal_4873), .Q (new_AGEMA_signal_4874) ) ;
    buf_clk new_AGEMA_reg_buffer_2104 ( .C (clk), .D (new_AGEMA_signal_4879), .Q (new_AGEMA_signal_4880) ) ;
    buf_clk new_AGEMA_reg_buffer_2110 ( .C (clk), .D (new_AGEMA_signal_4885), .Q (new_AGEMA_signal_4886) ) ;
    buf_clk new_AGEMA_reg_buffer_2116 ( .C (clk), .D (new_AGEMA_signal_4891), .Q (new_AGEMA_signal_4892) ) ;
    buf_clk new_AGEMA_reg_buffer_2122 ( .C (clk), .D (new_AGEMA_signal_4897), .Q (new_AGEMA_signal_4898) ) ;
    buf_clk new_AGEMA_reg_buffer_2128 ( .C (clk), .D (new_AGEMA_signal_4903), .Q (new_AGEMA_signal_4904) ) ;
    buf_clk new_AGEMA_reg_buffer_2134 ( .C (clk), .D (new_AGEMA_signal_4909), .Q (new_AGEMA_signal_4910) ) ;
    buf_clk new_AGEMA_reg_buffer_2140 ( .C (clk), .D (new_AGEMA_signal_4915), .Q (new_AGEMA_signal_4916) ) ;
    buf_clk new_AGEMA_reg_buffer_2146 ( .C (clk), .D (new_AGEMA_signal_4921), .Q (new_AGEMA_signal_4922) ) ;
    buf_clk new_AGEMA_reg_buffer_2152 ( .C (clk), .D (new_AGEMA_signal_4927), .Q (new_AGEMA_signal_4928) ) ;
    buf_clk new_AGEMA_reg_buffer_2158 ( .C (clk), .D (new_AGEMA_signal_4933), .Q (new_AGEMA_signal_4934) ) ;
    buf_clk new_AGEMA_reg_buffer_2164 ( .C (clk), .D (new_AGEMA_signal_4939), .Q (new_AGEMA_signal_4940) ) ;
    buf_clk new_AGEMA_reg_buffer_2170 ( .C (clk), .D (new_AGEMA_signal_4945), .Q (new_AGEMA_signal_4946) ) ;
    buf_clk new_AGEMA_reg_buffer_2176 ( .C (clk), .D (new_AGEMA_signal_4951), .Q (new_AGEMA_signal_4952) ) ;
    buf_clk new_AGEMA_reg_buffer_2182 ( .C (clk), .D (new_AGEMA_signal_4957), .Q (new_AGEMA_signal_4958) ) ;
    buf_clk new_AGEMA_reg_buffer_2188 ( .C (clk), .D (new_AGEMA_signal_4963), .Q (new_AGEMA_signal_4964) ) ;
    buf_clk new_AGEMA_reg_buffer_2194 ( .C (clk), .D (new_AGEMA_signal_4969), .Q (new_AGEMA_signal_4970) ) ;
    buf_clk new_AGEMA_reg_buffer_2200 ( .C (clk), .D (new_AGEMA_signal_4975), .Q (new_AGEMA_signal_4976) ) ;
    buf_clk new_AGEMA_reg_buffer_2206 ( .C (clk), .D (new_AGEMA_signal_4981), .Q (new_AGEMA_signal_4982) ) ;
    buf_clk new_AGEMA_reg_buffer_2212 ( .C (clk), .D (new_AGEMA_signal_4987), .Q (new_AGEMA_signal_4988) ) ;
    buf_clk new_AGEMA_reg_buffer_2218 ( .C (clk), .D (new_AGEMA_signal_4993), .Q (new_AGEMA_signal_4994) ) ;
    buf_clk new_AGEMA_reg_buffer_2224 ( .C (clk), .D (new_AGEMA_signal_4999), .Q (new_AGEMA_signal_5000) ) ;
    buf_clk new_AGEMA_reg_buffer_2230 ( .C (clk), .D (new_AGEMA_signal_5005), .Q (new_AGEMA_signal_5006) ) ;
    buf_clk new_AGEMA_reg_buffer_2236 ( .C (clk), .D (new_AGEMA_signal_5011), .Q (new_AGEMA_signal_5012) ) ;
    buf_clk new_AGEMA_reg_buffer_2242 ( .C (clk), .D (new_AGEMA_signal_5017), .Q (new_AGEMA_signal_5018) ) ;
    buf_clk new_AGEMA_reg_buffer_2248 ( .C (clk), .D (new_AGEMA_signal_5023), .Q (new_AGEMA_signal_5024) ) ;
    buf_clk new_AGEMA_reg_buffer_2254 ( .C (clk), .D (new_AGEMA_signal_5029), .Q (new_AGEMA_signal_5030) ) ;
    buf_clk new_AGEMA_reg_buffer_2260 ( .C (clk), .D (new_AGEMA_signal_5035), .Q (new_AGEMA_signal_5036) ) ;
    buf_clk new_AGEMA_reg_buffer_2266 ( .C (clk), .D (new_AGEMA_signal_5041), .Q (new_AGEMA_signal_5042) ) ;
    buf_clk new_AGEMA_reg_buffer_2272 ( .C (clk), .D (new_AGEMA_signal_5047), .Q (new_AGEMA_signal_5048) ) ;
    buf_clk new_AGEMA_reg_buffer_2278 ( .C (clk), .D (new_AGEMA_signal_5053), .Q (new_AGEMA_signal_5054) ) ;
    buf_clk new_AGEMA_reg_buffer_2284 ( .C (clk), .D (new_AGEMA_signal_5059), .Q (new_AGEMA_signal_5060) ) ;
    buf_clk new_AGEMA_reg_buffer_2290 ( .C (clk), .D (new_AGEMA_signal_5065), .Q (new_AGEMA_signal_5066) ) ;
    buf_clk new_AGEMA_reg_buffer_2296 ( .C (clk), .D (new_AGEMA_signal_5071), .Q (new_AGEMA_signal_5072) ) ;
    buf_clk new_AGEMA_reg_buffer_2302 ( .C (clk), .D (new_AGEMA_signal_5077), .Q (new_AGEMA_signal_5078) ) ;
    buf_clk new_AGEMA_reg_buffer_2308 ( .C (clk), .D (new_AGEMA_signal_5083), .Q (new_AGEMA_signal_5084) ) ;
    buf_clk new_AGEMA_reg_buffer_2314 ( .C (clk), .D (new_AGEMA_signal_5089), .Q (new_AGEMA_signal_5090) ) ;
    buf_clk new_AGEMA_reg_buffer_2320 ( .C (clk), .D (new_AGEMA_signal_5095), .Q (new_AGEMA_signal_5096) ) ;
    buf_clk new_AGEMA_reg_buffer_2326 ( .C (clk), .D (new_AGEMA_signal_5101), .Q (new_AGEMA_signal_5102) ) ;
    buf_clk new_AGEMA_reg_buffer_2332 ( .C (clk), .D (new_AGEMA_signal_5107), .Q (new_AGEMA_signal_5108) ) ;
    buf_clk new_AGEMA_reg_buffer_2338 ( .C (clk), .D (new_AGEMA_signal_5113), .Q (new_AGEMA_signal_5114) ) ;
    buf_clk new_AGEMA_reg_buffer_2344 ( .C (clk), .D (new_AGEMA_signal_5119), .Q (new_AGEMA_signal_5120) ) ;
    buf_clk new_AGEMA_reg_buffer_2350 ( .C (clk), .D (new_AGEMA_signal_5125), .Q (new_AGEMA_signal_5126) ) ;
    buf_clk new_AGEMA_reg_buffer_2356 ( .C (clk), .D (new_AGEMA_signal_5131), .Q (new_AGEMA_signal_5132) ) ;
    buf_clk new_AGEMA_reg_buffer_2652 ( .C (clk), .D (new_AGEMA_signal_5427), .Q (new_AGEMA_signal_5428) ) ;
    buf_clk new_AGEMA_reg_buffer_2660 ( .C (clk), .D (new_AGEMA_signal_5435), .Q (new_AGEMA_signal_5436) ) ;
    buf_clk new_AGEMA_reg_buffer_2668 ( .C (clk), .D (new_AGEMA_signal_5443), .Q (new_AGEMA_signal_5444) ) ;
    buf_clk new_AGEMA_reg_buffer_2676 ( .C (clk), .D (new_AGEMA_signal_5451), .Q (new_AGEMA_signal_5452) ) ;
    buf_clk new_AGEMA_reg_buffer_2684 ( .C (clk), .D (new_AGEMA_signal_5459), .Q (new_AGEMA_signal_5460) ) ;
    buf_clk new_AGEMA_reg_buffer_2692 ( .C (clk), .D (new_AGEMA_signal_5467), .Q (new_AGEMA_signal_5468) ) ;
    buf_clk new_AGEMA_reg_buffer_2700 ( .C (clk), .D (new_AGEMA_signal_5475), .Q (new_AGEMA_signal_5476) ) ;
    buf_clk new_AGEMA_reg_buffer_2708 ( .C (clk), .D (new_AGEMA_signal_5483), .Q (new_AGEMA_signal_5484) ) ;
    buf_clk new_AGEMA_reg_buffer_2716 ( .C (clk), .D (new_AGEMA_signal_5491), .Q (new_AGEMA_signal_5492) ) ;
    buf_clk new_AGEMA_reg_buffer_2724 ( .C (clk), .D (new_AGEMA_signal_5499), .Q (new_AGEMA_signal_5500) ) ;
    buf_clk new_AGEMA_reg_buffer_2732 ( .C (clk), .D (new_AGEMA_signal_5507), .Q (new_AGEMA_signal_5508) ) ;
    buf_clk new_AGEMA_reg_buffer_2740 ( .C (clk), .D (new_AGEMA_signal_5515), .Q (new_AGEMA_signal_5516) ) ;
    buf_clk new_AGEMA_reg_buffer_2748 ( .C (clk), .D (new_AGEMA_signal_5523), .Q (new_AGEMA_signal_5524) ) ;
    buf_clk new_AGEMA_reg_buffer_2756 ( .C (clk), .D (new_AGEMA_signal_5531), .Q (new_AGEMA_signal_5532) ) ;
    buf_clk new_AGEMA_reg_buffer_2764 ( .C (clk), .D (new_AGEMA_signal_5539), .Q (new_AGEMA_signal_5540) ) ;
    buf_clk new_AGEMA_reg_buffer_2772 ( .C (clk), .D (new_AGEMA_signal_5547), .Q (new_AGEMA_signal_5548) ) ;
    buf_clk new_AGEMA_reg_buffer_2780 ( .C (clk), .D (new_AGEMA_signal_5555), .Q (new_AGEMA_signal_5556) ) ;
    buf_clk new_AGEMA_reg_buffer_2788 ( .C (clk), .D (new_AGEMA_signal_5563), .Q (new_AGEMA_signal_5564) ) ;
    buf_clk new_AGEMA_reg_buffer_2796 ( .C (clk), .D (new_AGEMA_signal_5571), .Q (new_AGEMA_signal_5572) ) ;
    buf_clk new_AGEMA_reg_buffer_2804 ( .C (clk), .D (new_AGEMA_signal_5579), .Q (new_AGEMA_signal_5580) ) ;
    buf_clk new_AGEMA_reg_buffer_2812 ( .C (clk), .D (new_AGEMA_signal_5587), .Q (new_AGEMA_signal_5588) ) ;
    buf_clk new_AGEMA_reg_buffer_2820 ( .C (clk), .D (new_AGEMA_signal_5595), .Q (new_AGEMA_signal_5596) ) ;
    buf_clk new_AGEMA_reg_buffer_2828 ( .C (clk), .D (new_AGEMA_signal_5603), .Q (new_AGEMA_signal_5604) ) ;
    buf_clk new_AGEMA_reg_buffer_2836 ( .C (clk), .D (new_AGEMA_signal_5611), .Q (new_AGEMA_signal_5612) ) ;
    buf_clk new_AGEMA_reg_buffer_2844 ( .C (clk), .D (new_AGEMA_signal_5619), .Q (new_AGEMA_signal_5620) ) ;
    buf_clk new_AGEMA_reg_buffer_2852 ( .C (clk), .D (new_AGEMA_signal_5627), .Q (new_AGEMA_signal_5628) ) ;
    buf_clk new_AGEMA_reg_buffer_2860 ( .C (clk), .D (new_AGEMA_signal_5635), .Q (new_AGEMA_signal_5636) ) ;
    buf_clk new_AGEMA_reg_buffer_2868 ( .C (clk), .D (new_AGEMA_signal_5643), .Q (new_AGEMA_signal_5644) ) ;
    buf_clk new_AGEMA_reg_buffer_2876 ( .C (clk), .D (new_AGEMA_signal_5651), .Q (new_AGEMA_signal_5652) ) ;
    buf_clk new_AGEMA_reg_buffer_2884 ( .C (clk), .D (new_AGEMA_signal_5659), .Q (new_AGEMA_signal_5660) ) ;
    buf_clk new_AGEMA_reg_buffer_2892 ( .C (clk), .D (new_AGEMA_signal_5667), .Q (new_AGEMA_signal_5668) ) ;
    buf_clk new_AGEMA_reg_buffer_2900 ( .C (clk), .D (new_AGEMA_signal_5675), .Q (new_AGEMA_signal_5676) ) ;
    buf_clk new_AGEMA_reg_buffer_2908 ( .C (clk), .D (new_AGEMA_signal_5683), .Q (new_AGEMA_signal_5684) ) ;
    buf_clk new_AGEMA_reg_buffer_2916 ( .C (clk), .D (new_AGEMA_signal_5691), .Q (new_AGEMA_signal_5692) ) ;
    buf_clk new_AGEMA_reg_buffer_2924 ( .C (clk), .D (new_AGEMA_signal_5699), .Q (new_AGEMA_signal_5700) ) ;
    buf_clk new_AGEMA_reg_buffer_2932 ( .C (clk), .D (new_AGEMA_signal_5707), .Q (new_AGEMA_signal_5708) ) ;
    buf_clk new_AGEMA_reg_buffer_2940 ( .C (clk), .D (new_AGEMA_signal_5715), .Q (new_AGEMA_signal_5716) ) ;
    buf_clk new_AGEMA_reg_buffer_2948 ( .C (clk), .D (new_AGEMA_signal_5723), .Q (new_AGEMA_signal_5724) ) ;
    buf_clk new_AGEMA_reg_buffer_2956 ( .C (clk), .D (new_AGEMA_signal_5731), .Q (new_AGEMA_signal_5732) ) ;
    buf_clk new_AGEMA_reg_buffer_2964 ( .C (clk), .D (new_AGEMA_signal_5739), .Q (new_AGEMA_signal_5740) ) ;
    buf_clk new_AGEMA_reg_buffer_2972 ( .C (clk), .D (new_AGEMA_signal_5747), .Q (new_AGEMA_signal_5748) ) ;
    buf_clk new_AGEMA_reg_buffer_2980 ( .C (clk), .D (new_AGEMA_signal_5755), .Q (new_AGEMA_signal_5756) ) ;
    buf_clk new_AGEMA_reg_buffer_2988 ( .C (clk), .D (new_AGEMA_signal_5763), .Q (new_AGEMA_signal_5764) ) ;
    buf_clk new_AGEMA_reg_buffer_2996 ( .C (clk), .D (new_AGEMA_signal_5771), .Q (new_AGEMA_signal_5772) ) ;
    buf_clk new_AGEMA_reg_buffer_3004 ( .C (clk), .D (new_AGEMA_signal_5779), .Q (new_AGEMA_signal_5780) ) ;
    buf_clk new_AGEMA_reg_buffer_3012 ( .C (clk), .D (new_AGEMA_signal_5787), .Q (new_AGEMA_signal_5788) ) ;
    buf_clk new_AGEMA_reg_buffer_3020 ( .C (clk), .D (new_AGEMA_signal_5795), .Q (new_AGEMA_signal_5796) ) ;
    buf_clk new_AGEMA_reg_buffer_3028 ( .C (clk), .D (new_AGEMA_signal_5803), .Q (new_AGEMA_signal_5804) ) ;
    buf_clk new_AGEMA_reg_buffer_3036 ( .C (clk), .D (new_AGEMA_signal_5811), .Q (new_AGEMA_signal_5812) ) ;
    buf_clk new_AGEMA_reg_buffer_3044 ( .C (clk), .D (new_AGEMA_signal_5819), .Q (new_AGEMA_signal_5820) ) ;
    buf_clk new_AGEMA_reg_buffer_3052 ( .C (clk), .D (new_AGEMA_signal_5827), .Q (new_AGEMA_signal_5828) ) ;
    buf_clk new_AGEMA_reg_buffer_3060 ( .C (clk), .D (new_AGEMA_signal_5835), .Q (new_AGEMA_signal_5836) ) ;
    buf_clk new_AGEMA_reg_buffer_3068 ( .C (clk), .D (new_AGEMA_signal_5843), .Q (new_AGEMA_signal_5844) ) ;
    buf_clk new_AGEMA_reg_buffer_3076 ( .C (clk), .D (new_AGEMA_signal_5851), .Q (new_AGEMA_signal_5852) ) ;
    buf_clk new_AGEMA_reg_buffer_3084 ( .C (clk), .D (new_AGEMA_signal_5859), .Q (new_AGEMA_signal_5860) ) ;
    buf_clk new_AGEMA_reg_buffer_3092 ( .C (clk), .D (new_AGEMA_signal_5867), .Q (new_AGEMA_signal_5868) ) ;
    buf_clk new_AGEMA_reg_buffer_3100 ( .C (clk), .D (new_AGEMA_signal_5875), .Q (new_AGEMA_signal_5876) ) ;
    buf_clk new_AGEMA_reg_buffer_3108 ( .C (clk), .D (new_AGEMA_signal_5883), .Q (new_AGEMA_signal_5884) ) ;
    buf_clk new_AGEMA_reg_buffer_3116 ( .C (clk), .D (new_AGEMA_signal_5891), .Q (new_AGEMA_signal_5892) ) ;
    buf_clk new_AGEMA_reg_buffer_3124 ( .C (clk), .D (new_AGEMA_signal_5899), .Q (new_AGEMA_signal_5900) ) ;
    buf_clk new_AGEMA_reg_buffer_3132 ( .C (clk), .D (new_AGEMA_signal_5907), .Q (new_AGEMA_signal_5908) ) ;
    buf_clk new_AGEMA_reg_buffer_3140 ( .C (clk), .D (new_AGEMA_signal_5915), .Q (new_AGEMA_signal_5916) ) ;
    buf_clk new_AGEMA_reg_buffer_3148 ( .C (clk), .D (new_AGEMA_signal_5923), .Q (new_AGEMA_signal_5924) ) ;
    buf_clk new_AGEMA_reg_buffer_3156 ( .C (clk), .D (new_AGEMA_signal_5931), .Q (new_AGEMA_signal_5932) ) ;
    buf_clk new_AGEMA_reg_buffer_3164 ( .C (clk), .D (new_AGEMA_signal_5939), .Q (new_AGEMA_signal_5940) ) ;
    buf_clk new_AGEMA_reg_buffer_3172 ( .C (clk), .D (new_AGEMA_signal_5947), .Q (new_AGEMA_signal_5948) ) ;
    buf_clk new_AGEMA_reg_buffer_3180 ( .C (clk), .D (new_AGEMA_signal_5955), .Q (new_AGEMA_signal_5956) ) ;
    buf_clk new_AGEMA_reg_buffer_3188 ( .C (clk), .D (new_AGEMA_signal_5963), .Q (new_AGEMA_signal_5964) ) ;
    buf_clk new_AGEMA_reg_buffer_3196 ( .C (clk), .D (new_AGEMA_signal_5971), .Q (new_AGEMA_signal_5972) ) ;
    buf_clk new_AGEMA_reg_buffer_3204 ( .C (clk), .D (new_AGEMA_signal_5979), .Q (new_AGEMA_signal_5980) ) ;
    buf_clk new_AGEMA_reg_buffer_3212 ( .C (clk), .D (new_AGEMA_signal_5987), .Q (new_AGEMA_signal_5988) ) ;
    buf_clk new_AGEMA_reg_buffer_3220 ( .C (clk), .D (new_AGEMA_signal_5995), .Q (new_AGEMA_signal_5996) ) ;
    buf_clk new_AGEMA_reg_buffer_3228 ( .C (clk), .D (new_AGEMA_signal_6003), .Q (new_AGEMA_signal_6004) ) ;
    buf_clk new_AGEMA_reg_buffer_3236 ( .C (clk), .D (new_AGEMA_signal_6011), .Q (new_AGEMA_signal_6012) ) ;
    buf_clk new_AGEMA_reg_buffer_3244 ( .C (clk), .D (new_AGEMA_signal_6019), .Q (new_AGEMA_signal_6020) ) ;
    buf_clk new_AGEMA_reg_buffer_3252 ( .C (clk), .D (new_AGEMA_signal_6027), .Q (new_AGEMA_signal_6028) ) ;
    buf_clk new_AGEMA_reg_buffer_3260 ( .C (clk), .D (new_AGEMA_signal_6035), .Q (new_AGEMA_signal_6036) ) ;
    buf_clk new_AGEMA_reg_buffer_3268 ( .C (clk), .D (new_AGEMA_signal_6043), .Q (new_AGEMA_signal_6044) ) ;
    buf_clk new_AGEMA_reg_buffer_3276 ( .C (clk), .D (new_AGEMA_signal_6051), .Q (new_AGEMA_signal_6052) ) ;
    buf_clk new_AGEMA_reg_buffer_3284 ( .C (clk), .D (new_AGEMA_signal_6059), .Q (new_AGEMA_signal_6060) ) ;
    buf_clk new_AGEMA_reg_buffer_3292 ( .C (clk), .D (new_AGEMA_signal_6067), .Q (new_AGEMA_signal_6068) ) ;
    buf_clk new_AGEMA_reg_buffer_3300 ( .C (clk), .D (new_AGEMA_signal_6075), .Q (new_AGEMA_signal_6076) ) ;
    buf_clk new_AGEMA_reg_buffer_3308 ( .C (clk), .D (new_AGEMA_signal_6083), .Q (new_AGEMA_signal_6084) ) ;
    buf_clk new_AGEMA_reg_buffer_3316 ( .C (clk), .D (new_AGEMA_signal_6091), .Q (new_AGEMA_signal_6092) ) ;
    buf_clk new_AGEMA_reg_buffer_3324 ( .C (clk), .D (new_AGEMA_signal_6099), .Q (new_AGEMA_signal_6100) ) ;
    buf_clk new_AGEMA_reg_buffer_3332 ( .C (clk), .D (new_AGEMA_signal_6107), .Q (new_AGEMA_signal_6108) ) ;
    buf_clk new_AGEMA_reg_buffer_3340 ( .C (clk), .D (new_AGEMA_signal_6115), .Q (new_AGEMA_signal_6116) ) ;
    buf_clk new_AGEMA_reg_buffer_3348 ( .C (clk), .D (new_AGEMA_signal_6123), .Q (new_AGEMA_signal_6124) ) ;
    buf_clk new_AGEMA_reg_buffer_3356 ( .C (clk), .D (new_AGEMA_signal_6131), .Q (new_AGEMA_signal_6132) ) ;
    buf_clk new_AGEMA_reg_buffer_3364 ( .C (clk), .D (new_AGEMA_signal_6139), .Q (new_AGEMA_signal_6140) ) ;
    buf_clk new_AGEMA_reg_buffer_3372 ( .C (clk), .D (new_AGEMA_signal_6147), .Q (new_AGEMA_signal_6148) ) ;
    buf_clk new_AGEMA_reg_buffer_3380 ( .C (clk), .D (new_AGEMA_signal_6155), .Q (new_AGEMA_signal_6156) ) ;
    buf_clk new_AGEMA_reg_buffer_3388 ( .C (clk), .D (new_AGEMA_signal_6163), .Q (new_AGEMA_signal_6164) ) ;
    buf_clk new_AGEMA_reg_buffer_3396 ( .C (clk), .D (new_AGEMA_signal_6171), .Q (new_AGEMA_signal_6172) ) ;
    buf_clk new_AGEMA_reg_buffer_3404 ( .C (clk), .D (new_AGEMA_signal_6179), .Q (new_AGEMA_signal_6180) ) ;
    buf_clk new_AGEMA_reg_buffer_3412 ( .C (clk), .D (new_AGEMA_signal_6187), .Q (new_AGEMA_signal_6188) ) ;
    buf_clk new_AGEMA_reg_buffer_3420 ( .C (clk), .D (new_AGEMA_signal_6195), .Q (new_AGEMA_signal_6196) ) ;
    buf_clk new_AGEMA_reg_buffer_3428 ( .C (clk), .D (new_AGEMA_signal_6203), .Q (new_AGEMA_signal_6204) ) ;
    buf_clk new_AGEMA_reg_buffer_3436 ( .C (clk), .D (new_AGEMA_signal_6211), .Q (new_AGEMA_signal_6212) ) ;
    buf_clk new_AGEMA_reg_buffer_3444 ( .C (clk), .D (new_AGEMA_signal_6219), .Q (new_AGEMA_signal_6220) ) ;
    buf_clk new_AGEMA_reg_buffer_3452 ( .C (clk), .D (new_AGEMA_signal_6227), .Q (new_AGEMA_signal_6228) ) ;
    buf_clk new_AGEMA_reg_buffer_3460 ( .C (clk), .D (new_AGEMA_signal_6235), .Q (new_AGEMA_signal_6236) ) ;
    buf_clk new_AGEMA_reg_buffer_3468 ( .C (clk), .D (new_AGEMA_signal_6243), .Q (new_AGEMA_signal_6244) ) ;
    buf_clk new_AGEMA_reg_buffer_3476 ( .C (clk), .D (new_AGEMA_signal_6251), .Q (new_AGEMA_signal_6252) ) ;
    buf_clk new_AGEMA_reg_buffer_3484 ( .C (clk), .D (new_AGEMA_signal_6259), .Q (new_AGEMA_signal_6260) ) ;
    buf_clk new_AGEMA_reg_buffer_3492 ( .C (clk), .D (new_AGEMA_signal_6267), .Q (new_AGEMA_signal_6268) ) ;
    buf_clk new_AGEMA_reg_buffer_3500 ( .C (clk), .D (new_AGEMA_signal_6275), .Q (new_AGEMA_signal_6276) ) ;
    buf_clk new_AGEMA_reg_buffer_3508 ( .C (clk), .D (new_AGEMA_signal_6283), .Q (new_AGEMA_signal_6284) ) ;
    buf_clk new_AGEMA_reg_buffer_3516 ( .C (clk), .D (new_AGEMA_signal_6291), .Q (new_AGEMA_signal_6292) ) ;
    buf_clk new_AGEMA_reg_buffer_3524 ( .C (clk), .D (new_AGEMA_signal_6299), .Q (new_AGEMA_signal_6300) ) ;
    buf_clk new_AGEMA_reg_buffer_3532 ( .C (clk), .D (new_AGEMA_signal_6307), .Q (new_AGEMA_signal_6308) ) ;
    buf_clk new_AGEMA_reg_buffer_3540 ( .C (clk), .D (new_AGEMA_signal_6315), .Q (new_AGEMA_signal_6316) ) ;
    buf_clk new_AGEMA_reg_buffer_3548 ( .C (clk), .D (new_AGEMA_signal_6323), .Q (new_AGEMA_signal_6324) ) ;
    buf_clk new_AGEMA_reg_buffer_3556 ( .C (clk), .D (new_AGEMA_signal_6331), .Q (new_AGEMA_signal_6332) ) ;
    buf_clk new_AGEMA_reg_buffer_3564 ( .C (clk), .D (new_AGEMA_signal_6339), .Q (new_AGEMA_signal_6340) ) ;
    buf_clk new_AGEMA_reg_buffer_3572 ( .C (clk), .D (new_AGEMA_signal_6347), .Q (new_AGEMA_signal_6348) ) ;
    buf_clk new_AGEMA_reg_buffer_3580 ( .C (clk), .D (new_AGEMA_signal_6355), .Q (new_AGEMA_signal_6356) ) ;
    buf_clk new_AGEMA_reg_buffer_3588 ( .C (clk), .D (new_AGEMA_signal_6363), .Q (new_AGEMA_signal_6364) ) ;
    buf_clk new_AGEMA_reg_buffer_3596 ( .C (clk), .D (new_AGEMA_signal_6371), .Q (new_AGEMA_signal_6372) ) ;
    buf_clk new_AGEMA_reg_buffer_3604 ( .C (clk), .D (new_AGEMA_signal_6379), .Q (new_AGEMA_signal_6380) ) ;
    buf_clk new_AGEMA_reg_buffer_3612 ( .C (clk), .D (new_AGEMA_signal_6387), .Q (new_AGEMA_signal_6388) ) ;
    buf_clk new_AGEMA_reg_buffer_3620 ( .C (clk), .D (new_AGEMA_signal_6395), .Q (new_AGEMA_signal_6396) ) ;
    buf_clk new_AGEMA_reg_buffer_3628 ( .C (clk), .D (new_AGEMA_signal_6403), .Q (new_AGEMA_signal_6404) ) ;
    buf_clk new_AGEMA_reg_buffer_3636 ( .C (clk), .D (new_AGEMA_signal_6411), .Q (new_AGEMA_signal_6412) ) ;
    buf_clk new_AGEMA_reg_buffer_3644 ( .C (clk), .D (new_AGEMA_signal_6419), .Q (new_AGEMA_signal_6420) ) ;
    buf_clk new_AGEMA_reg_buffer_3652 ( .C (clk), .D (new_AGEMA_signal_6427), .Q (new_AGEMA_signal_6428) ) ;
    buf_clk new_AGEMA_reg_buffer_3660 ( .C (clk), .D (new_AGEMA_signal_6435), .Q (new_AGEMA_signal_6436) ) ;
    buf_clk new_AGEMA_reg_buffer_3668 ( .C (clk), .D (new_AGEMA_signal_6443), .Q (new_AGEMA_signal_6444) ) ;
    buf_clk new_AGEMA_reg_buffer_3676 ( .C (clk), .D (new_AGEMA_signal_6451), .Q (new_AGEMA_signal_6452) ) ;
    buf_clk new_AGEMA_reg_buffer_3684 ( .C (clk), .D (new_AGEMA_signal_6459), .Q (new_AGEMA_signal_6460) ) ;
    buf_clk new_AGEMA_reg_buffer_3692 ( .C (clk), .D (new_AGEMA_signal_6467), .Q (new_AGEMA_signal_6468) ) ;
    buf_clk new_AGEMA_reg_buffer_3700 ( .C (clk), .D (new_AGEMA_signal_6475), .Q (new_AGEMA_signal_6476) ) ;
    buf_clk new_AGEMA_reg_buffer_3708 ( .C (clk), .D (new_AGEMA_signal_6483), .Q (new_AGEMA_signal_6484) ) ;
    buf_clk new_AGEMA_reg_buffer_3716 ( .C (clk), .D (new_AGEMA_signal_6491), .Q (new_AGEMA_signal_6492) ) ;
    buf_clk new_AGEMA_reg_buffer_3724 ( .C (clk), .D (new_AGEMA_signal_6499), .Q (new_AGEMA_signal_6500) ) ;
    buf_clk new_AGEMA_reg_buffer_3732 ( .C (clk), .D (new_AGEMA_signal_6507), .Q (new_AGEMA_signal_6508) ) ;
    buf_clk new_AGEMA_reg_buffer_3740 ( .C (clk), .D (new_AGEMA_signal_6515), .Q (new_AGEMA_signal_6516) ) ;
    buf_clk new_AGEMA_reg_buffer_3748 ( .C (clk), .D (new_AGEMA_signal_6523), .Q (new_AGEMA_signal_6524) ) ;
    buf_clk new_AGEMA_reg_buffer_3756 ( .C (clk), .D (new_AGEMA_signal_6531), .Q (new_AGEMA_signal_6532) ) ;
    buf_clk new_AGEMA_reg_buffer_3764 ( .C (clk), .D (new_AGEMA_signal_6539), .Q (new_AGEMA_signal_6540) ) ;
    buf_clk new_AGEMA_reg_buffer_3772 ( .C (clk), .D (new_AGEMA_signal_6547), .Q (new_AGEMA_signal_6548) ) ;
    buf_clk new_AGEMA_reg_buffer_3780 ( .C (clk), .D (new_AGEMA_signal_6555), .Q (new_AGEMA_signal_6556) ) ;
    buf_clk new_AGEMA_reg_buffer_3788 ( .C (clk), .D (new_AGEMA_signal_6563), .Q (new_AGEMA_signal_6564) ) ;
    buf_clk new_AGEMA_reg_buffer_3796 ( .C (clk), .D (new_AGEMA_signal_6571), .Q (new_AGEMA_signal_6572) ) ;
    buf_clk new_AGEMA_reg_buffer_3804 ( .C (clk), .D (new_AGEMA_signal_6579), .Q (new_AGEMA_signal_6580) ) ;
    buf_clk new_AGEMA_reg_buffer_3812 ( .C (clk), .D (new_AGEMA_signal_6587), .Q (new_AGEMA_signal_6588) ) ;
    buf_clk new_AGEMA_reg_buffer_3820 ( .C (clk), .D (new_AGEMA_signal_6595), .Q (new_AGEMA_signal_6596) ) ;
    buf_clk new_AGEMA_reg_buffer_3828 ( .C (clk), .D (new_AGEMA_signal_6603), .Q (new_AGEMA_signal_6604) ) ;
    buf_clk new_AGEMA_reg_buffer_3836 ( .C (clk), .D (new_AGEMA_signal_6611), .Q (new_AGEMA_signal_6612) ) ;
    buf_clk new_AGEMA_reg_buffer_3844 ( .C (clk), .D (new_AGEMA_signal_6619), .Q (new_AGEMA_signal_6620) ) ;
    buf_clk new_AGEMA_reg_buffer_3852 ( .C (clk), .D (new_AGEMA_signal_6627), .Q (new_AGEMA_signal_6628) ) ;
    buf_clk new_AGEMA_reg_buffer_3860 ( .C (clk), .D (new_AGEMA_signal_6635), .Q (new_AGEMA_signal_6636) ) ;
    buf_clk new_AGEMA_reg_buffer_3868 ( .C (clk), .D (new_AGEMA_signal_6643), .Q (new_AGEMA_signal_6644) ) ;
    buf_clk new_AGEMA_reg_buffer_3876 ( .C (clk), .D (new_AGEMA_signal_6651), .Q (new_AGEMA_signal_6652) ) ;
    buf_clk new_AGEMA_reg_buffer_3884 ( .C (clk), .D (new_AGEMA_signal_6659), .Q (new_AGEMA_signal_6660) ) ;
    buf_clk new_AGEMA_reg_buffer_3892 ( .C (clk), .D (new_AGEMA_signal_6667), .Q (new_AGEMA_signal_6668) ) ;
    buf_clk new_AGEMA_reg_buffer_3900 ( .C (clk), .D (new_AGEMA_signal_6675), .Q (new_AGEMA_signal_6676) ) ;
    buf_clk new_AGEMA_reg_buffer_3908 ( .C (clk), .D (new_AGEMA_signal_6683), .Q (new_AGEMA_signal_6684) ) ;
    buf_clk new_AGEMA_reg_buffer_3916 ( .C (clk), .D (new_AGEMA_signal_6691), .Q (new_AGEMA_signal_6692) ) ;
    buf_clk new_AGEMA_reg_buffer_3924 ( .C (clk), .D (new_AGEMA_signal_6699), .Q (new_AGEMA_signal_6700) ) ;
    buf_clk new_AGEMA_reg_buffer_3932 ( .C (clk), .D (new_AGEMA_signal_6707), .Q (new_AGEMA_signal_6708) ) ;
    buf_clk new_AGEMA_reg_buffer_3940 ( .C (clk), .D (new_AGEMA_signal_6715), .Q (new_AGEMA_signal_6716) ) ;
    buf_clk new_AGEMA_reg_buffer_3948 ( .C (clk), .D (new_AGEMA_signal_6723), .Q (new_AGEMA_signal_6724) ) ;
    buf_clk new_AGEMA_reg_buffer_3956 ( .C (clk), .D (new_AGEMA_signal_6731), .Q (new_AGEMA_signal_6732) ) ;
    buf_clk new_AGEMA_reg_buffer_3964 ( .C (clk), .D (new_AGEMA_signal_6739), .Q (new_AGEMA_signal_6740) ) ;
    buf_clk new_AGEMA_reg_buffer_3972 ( .C (clk), .D (new_AGEMA_signal_6747), .Q (new_AGEMA_signal_6748) ) ;
    buf_clk new_AGEMA_reg_buffer_3980 ( .C (clk), .D (new_AGEMA_signal_6755), .Q (new_AGEMA_signal_6756) ) ;
    buf_clk new_AGEMA_reg_buffer_3988 ( .C (clk), .D (new_AGEMA_signal_6763), .Q (new_AGEMA_signal_6764) ) ;
    buf_clk new_AGEMA_reg_buffer_3996 ( .C (clk), .D (new_AGEMA_signal_6771), .Q (new_AGEMA_signal_6772) ) ;
    buf_clk new_AGEMA_reg_buffer_4004 ( .C (clk), .D (new_AGEMA_signal_6779), .Q (new_AGEMA_signal_6780) ) ;
    buf_clk new_AGEMA_reg_buffer_4012 ( .C (clk), .D (new_AGEMA_signal_6787), .Q (new_AGEMA_signal_6788) ) ;
    buf_clk new_AGEMA_reg_buffer_4020 ( .C (clk), .D (new_AGEMA_signal_6795), .Q (new_AGEMA_signal_6796) ) ;
    buf_clk new_AGEMA_reg_buffer_4028 ( .C (clk), .D (new_AGEMA_signal_6803), .Q (new_AGEMA_signal_6804) ) ;
    buf_clk new_AGEMA_reg_buffer_4036 ( .C (clk), .D (new_AGEMA_signal_6811), .Q (new_AGEMA_signal_6812) ) ;
    buf_clk new_AGEMA_reg_buffer_4044 ( .C (clk), .D (new_AGEMA_signal_6819), .Q (new_AGEMA_signal_6820) ) ;
    buf_clk new_AGEMA_reg_buffer_4052 ( .C (clk), .D (new_AGEMA_signal_6827), .Q (new_AGEMA_signal_6828) ) ;
    buf_clk new_AGEMA_reg_buffer_4060 ( .C (clk), .D (new_AGEMA_signal_6835), .Q (new_AGEMA_signal_6836) ) ;
    buf_clk new_AGEMA_reg_buffer_4068 ( .C (clk), .D (new_AGEMA_signal_6843), .Q (new_AGEMA_signal_6844) ) ;
    buf_clk new_AGEMA_reg_buffer_4076 ( .C (clk), .D (new_AGEMA_signal_6851), .Q (new_AGEMA_signal_6852) ) ;
    buf_clk new_AGEMA_reg_buffer_4084 ( .C (clk), .D (new_AGEMA_signal_6859), .Q (new_AGEMA_signal_6860) ) ;
    buf_clk new_AGEMA_reg_buffer_4092 ( .C (clk), .D (new_AGEMA_signal_6867), .Q (new_AGEMA_signal_6868) ) ;
    buf_clk new_AGEMA_reg_buffer_4100 ( .C (clk), .D (new_AGEMA_signal_6875), .Q (new_AGEMA_signal_6876) ) ;
    buf_clk new_AGEMA_reg_buffer_4108 ( .C (clk), .D (new_AGEMA_signal_6883), .Q (new_AGEMA_signal_6884) ) ;
    buf_clk new_AGEMA_reg_buffer_4116 ( .C (clk), .D (new_AGEMA_signal_6891), .Q (new_AGEMA_signal_6892) ) ;
    buf_clk new_AGEMA_reg_buffer_4124 ( .C (clk), .D (new_AGEMA_signal_6899), .Q (new_AGEMA_signal_6900) ) ;
    buf_clk new_AGEMA_reg_buffer_4132 ( .C (clk), .D (new_AGEMA_signal_6907), .Q (new_AGEMA_signal_6908) ) ;
    buf_clk new_AGEMA_reg_buffer_4140 ( .C (clk), .D (new_AGEMA_signal_6915), .Q (new_AGEMA_signal_6916) ) ;
    buf_clk new_AGEMA_reg_buffer_4148 ( .C (clk), .D (new_AGEMA_signal_6923), .Q (new_AGEMA_signal_6924) ) ;
    buf_clk new_AGEMA_reg_buffer_4156 ( .C (clk), .D (new_AGEMA_signal_6931), .Q (new_AGEMA_signal_6932) ) ;
    buf_clk new_AGEMA_reg_buffer_4164 ( .C (clk), .D (new_AGEMA_signal_6939), .Q (new_AGEMA_signal_6940) ) ;
    buf_clk new_AGEMA_reg_buffer_4172 ( .C (clk), .D (new_AGEMA_signal_6947), .Q (new_AGEMA_signal_6948) ) ;
    buf_clk new_AGEMA_reg_buffer_4180 ( .C (clk), .D (new_AGEMA_signal_6955), .Q (new_AGEMA_signal_6956) ) ;
    buf_clk new_AGEMA_reg_buffer_4668 ( .C (clk), .D (new_AGEMA_signal_7443), .Q (new_AGEMA_signal_7444) ) ;
    buf_clk new_AGEMA_reg_buffer_4676 ( .C (clk), .D (new_AGEMA_signal_7451), .Q (new_AGEMA_signal_7452) ) ;
    buf_clk new_AGEMA_reg_buffer_4684 ( .C (clk), .D (new_AGEMA_signal_7459), .Q (new_AGEMA_signal_7460) ) ;
    buf_clk new_AGEMA_reg_buffer_4692 ( .C (clk), .D (new_AGEMA_signal_7467), .Q (new_AGEMA_signal_7468) ) ;
    buf_clk new_AGEMA_reg_buffer_4700 ( .C (clk), .D (new_AGEMA_signal_7475), .Q (new_AGEMA_signal_7476) ) ;
    buf_clk new_AGEMA_reg_buffer_4708 ( .C (clk), .D (new_AGEMA_signal_7483), .Q (new_AGEMA_signal_7484) ) ;
    buf_clk new_AGEMA_reg_buffer_4716 ( .C (clk), .D (new_AGEMA_signal_7491), .Q (new_AGEMA_signal_7492) ) ;
    buf_clk new_AGEMA_reg_buffer_4724 ( .C (clk), .D (new_AGEMA_signal_7499), .Q (new_AGEMA_signal_7500) ) ;
    buf_clk new_AGEMA_reg_buffer_4732 ( .C (clk), .D (new_AGEMA_signal_7507), .Q (new_AGEMA_signal_7508) ) ;
    buf_clk new_AGEMA_reg_buffer_4740 ( .C (clk), .D (new_AGEMA_signal_7515), .Q (new_AGEMA_signal_7516) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_1205 ( .C (clk), .D (new_AGEMA_signal_3980), .Q (new_AGEMA_signal_3981) ) ;
    buf_clk new_AGEMA_reg_buffer_1211 ( .C (clk), .D (new_AGEMA_signal_3986), .Q (new_AGEMA_signal_3987) ) ;
    buf_clk new_AGEMA_reg_buffer_1217 ( .C (clk), .D (new_AGEMA_signal_3992), .Q (new_AGEMA_signal_3993) ) ;
    buf_clk new_AGEMA_reg_buffer_1223 ( .C (clk), .D (new_AGEMA_signal_3998), .Q (new_AGEMA_signal_3999) ) ;
    buf_clk new_AGEMA_reg_buffer_1229 ( .C (clk), .D (new_AGEMA_signal_4004), .Q (new_AGEMA_signal_4005) ) ;
    buf_clk new_AGEMA_reg_buffer_1235 ( .C (clk), .D (new_AGEMA_signal_4010), .Q (new_AGEMA_signal_4011) ) ;
    buf_clk new_AGEMA_reg_buffer_1241 ( .C (clk), .D (new_AGEMA_signal_4016), .Q (new_AGEMA_signal_4017) ) ;
    buf_clk new_AGEMA_reg_buffer_1247 ( .C (clk), .D (new_AGEMA_signal_4022), .Q (new_AGEMA_signal_4023) ) ;
    buf_clk new_AGEMA_reg_buffer_1253 ( .C (clk), .D (new_AGEMA_signal_4028), .Q (new_AGEMA_signal_4029) ) ;
    buf_clk new_AGEMA_reg_buffer_1259 ( .C (clk), .D (new_AGEMA_signal_4034), .Q (new_AGEMA_signal_4035) ) ;
    buf_clk new_AGEMA_reg_buffer_1265 ( .C (clk), .D (new_AGEMA_signal_4040), .Q (new_AGEMA_signal_4041) ) ;
    buf_clk new_AGEMA_reg_buffer_1271 ( .C (clk), .D (new_AGEMA_signal_4046), .Q (new_AGEMA_signal_4047) ) ;
    buf_clk new_AGEMA_reg_buffer_1277 ( .C (clk), .D (new_AGEMA_signal_4052), .Q (new_AGEMA_signal_4053) ) ;
    buf_clk new_AGEMA_reg_buffer_1283 ( .C (clk), .D (new_AGEMA_signal_4058), .Q (new_AGEMA_signal_4059) ) ;
    buf_clk new_AGEMA_reg_buffer_1289 ( .C (clk), .D (new_AGEMA_signal_4064), .Q (new_AGEMA_signal_4065) ) ;
    buf_clk new_AGEMA_reg_buffer_1295 ( .C (clk), .D (new_AGEMA_signal_4070), .Q (new_AGEMA_signal_4071) ) ;
    buf_clk new_AGEMA_reg_buffer_1301 ( .C (clk), .D (new_AGEMA_signal_4076), .Q (new_AGEMA_signal_4077) ) ;
    buf_clk new_AGEMA_reg_buffer_1307 ( .C (clk), .D (new_AGEMA_signal_4082), .Q (new_AGEMA_signal_4083) ) ;
    buf_clk new_AGEMA_reg_buffer_1313 ( .C (clk), .D (new_AGEMA_signal_4088), .Q (new_AGEMA_signal_4089) ) ;
    buf_clk new_AGEMA_reg_buffer_1319 ( .C (clk), .D (new_AGEMA_signal_4094), .Q (new_AGEMA_signal_4095) ) ;
    buf_clk new_AGEMA_reg_buffer_1325 ( .C (clk), .D (new_AGEMA_signal_4100), .Q (new_AGEMA_signal_4101) ) ;
    buf_clk new_AGEMA_reg_buffer_1331 ( .C (clk), .D (new_AGEMA_signal_4106), .Q (new_AGEMA_signal_4107) ) ;
    buf_clk new_AGEMA_reg_buffer_1337 ( .C (clk), .D (new_AGEMA_signal_4112), .Q (new_AGEMA_signal_4113) ) ;
    buf_clk new_AGEMA_reg_buffer_1343 ( .C (clk), .D (new_AGEMA_signal_4118), .Q (new_AGEMA_signal_4119) ) ;
    buf_clk new_AGEMA_reg_buffer_1349 ( .C (clk), .D (new_AGEMA_signal_4124), .Q (new_AGEMA_signal_4125) ) ;
    buf_clk new_AGEMA_reg_buffer_1355 ( .C (clk), .D (new_AGEMA_signal_4130), .Q (new_AGEMA_signal_4131) ) ;
    buf_clk new_AGEMA_reg_buffer_1361 ( .C (clk), .D (new_AGEMA_signal_4136), .Q (new_AGEMA_signal_4137) ) ;
    buf_clk new_AGEMA_reg_buffer_1367 ( .C (clk), .D (new_AGEMA_signal_4142), .Q (new_AGEMA_signal_4143) ) ;
    buf_clk new_AGEMA_reg_buffer_1373 ( .C (clk), .D (new_AGEMA_signal_4148), .Q (new_AGEMA_signal_4149) ) ;
    buf_clk new_AGEMA_reg_buffer_1379 ( .C (clk), .D (new_AGEMA_signal_4154), .Q (new_AGEMA_signal_4155) ) ;
    buf_clk new_AGEMA_reg_buffer_1385 ( .C (clk), .D (new_AGEMA_signal_4160), .Q (new_AGEMA_signal_4161) ) ;
    buf_clk new_AGEMA_reg_buffer_1391 ( .C (clk), .D (new_AGEMA_signal_4166), .Q (new_AGEMA_signal_4167) ) ;
    buf_clk new_AGEMA_reg_buffer_1397 ( .C (clk), .D (new_AGEMA_signal_4172), .Q (new_AGEMA_signal_4173) ) ;
    buf_clk new_AGEMA_reg_buffer_1403 ( .C (clk), .D (new_AGEMA_signal_4178), .Q (new_AGEMA_signal_4179) ) ;
    buf_clk new_AGEMA_reg_buffer_1409 ( .C (clk), .D (new_AGEMA_signal_4184), .Q (new_AGEMA_signal_4185) ) ;
    buf_clk new_AGEMA_reg_buffer_1415 ( .C (clk), .D (new_AGEMA_signal_4190), .Q (new_AGEMA_signal_4191) ) ;
    buf_clk new_AGEMA_reg_buffer_1421 ( .C (clk), .D (new_AGEMA_signal_4196), .Q (new_AGEMA_signal_4197) ) ;
    buf_clk new_AGEMA_reg_buffer_1427 ( .C (clk), .D (new_AGEMA_signal_4202), .Q (new_AGEMA_signal_4203) ) ;
    buf_clk new_AGEMA_reg_buffer_1433 ( .C (clk), .D (new_AGEMA_signal_4208), .Q (new_AGEMA_signal_4209) ) ;
    buf_clk new_AGEMA_reg_buffer_1439 ( .C (clk), .D (new_AGEMA_signal_4214), .Q (new_AGEMA_signal_4215) ) ;
    buf_clk new_AGEMA_reg_buffer_1445 ( .C (clk), .D (new_AGEMA_signal_4220), .Q (new_AGEMA_signal_4221) ) ;
    buf_clk new_AGEMA_reg_buffer_1451 ( .C (clk), .D (new_AGEMA_signal_4226), .Q (new_AGEMA_signal_4227) ) ;
    buf_clk new_AGEMA_reg_buffer_1457 ( .C (clk), .D (new_AGEMA_signal_4232), .Q (new_AGEMA_signal_4233) ) ;
    buf_clk new_AGEMA_reg_buffer_1463 ( .C (clk), .D (new_AGEMA_signal_4238), .Q (new_AGEMA_signal_4239) ) ;
    buf_clk new_AGEMA_reg_buffer_1469 ( .C (clk), .D (new_AGEMA_signal_4244), .Q (new_AGEMA_signal_4245) ) ;
    buf_clk new_AGEMA_reg_buffer_1475 ( .C (clk), .D (new_AGEMA_signal_4250), .Q (new_AGEMA_signal_4251) ) ;
    buf_clk new_AGEMA_reg_buffer_1481 ( .C (clk), .D (new_AGEMA_signal_4256), .Q (new_AGEMA_signal_4257) ) ;
    buf_clk new_AGEMA_reg_buffer_1487 ( .C (clk), .D (new_AGEMA_signal_4262), .Q (new_AGEMA_signal_4263) ) ;
    buf_clk new_AGEMA_reg_buffer_1493 ( .C (clk), .D (new_AGEMA_signal_4268), .Q (new_AGEMA_signal_4269) ) ;
    buf_clk new_AGEMA_reg_buffer_1499 ( .C (clk), .D (new_AGEMA_signal_4274), .Q (new_AGEMA_signal_4275) ) ;
    buf_clk new_AGEMA_reg_buffer_1505 ( .C (clk), .D (new_AGEMA_signal_4280), .Q (new_AGEMA_signal_4281) ) ;
    buf_clk new_AGEMA_reg_buffer_1511 ( .C (clk), .D (new_AGEMA_signal_4286), .Q (new_AGEMA_signal_4287) ) ;
    buf_clk new_AGEMA_reg_buffer_1517 ( .C (clk), .D (new_AGEMA_signal_4292), .Q (new_AGEMA_signal_4293) ) ;
    buf_clk new_AGEMA_reg_buffer_1523 ( .C (clk), .D (new_AGEMA_signal_4298), .Q (new_AGEMA_signal_4299) ) ;
    buf_clk new_AGEMA_reg_buffer_1529 ( .C (clk), .D (new_AGEMA_signal_4304), .Q (new_AGEMA_signal_4305) ) ;
    buf_clk new_AGEMA_reg_buffer_1535 ( .C (clk), .D (new_AGEMA_signal_4310), .Q (new_AGEMA_signal_4311) ) ;
    buf_clk new_AGEMA_reg_buffer_1541 ( .C (clk), .D (new_AGEMA_signal_4316), .Q (new_AGEMA_signal_4317) ) ;
    buf_clk new_AGEMA_reg_buffer_1547 ( .C (clk), .D (new_AGEMA_signal_4322), .Q (new_AGEMA_signal_4323) ) ;
    buf_clk new_AGEMA_reg_buffer_1553 ( .C (clk), .D (new_AGEMA_signal_4328), .Q (new_AGEMA_signal_4329) ) ;
    buf_clk new_AGEMA_reg_buffer_1559 ( .C (clk), .D (new_AGEMA_signal_4334), .Q (new_AGEMA_signal_4335) ) ;
    buf_clk new_AGEMA_reg_buffer_1565 ( .C (clk), .D (new_AGEMA_signal_4340), .Q (new_AGEMA_signal_4341) ) ;
    buf_clk new_AGEMA_reg_buffer_1571 ( .C (clk), .D (new_AGEMA_signal_4346), .Q (new_AGEMA_signal_4347) ) ;
    buf_clk new_AGEMA_reg_buffer_1577 ( .C (clk), .D (new_AGEMA_signal_4352), .Q (new_AGEMA_signal_4353) ) ;
    buf_clk new_AGEMA_reg_buffer_1583 ( .C (clk), .D (new_AGEMA_signal_4358), .Q (new_AGEMA_signal_4359) ) ;
    buf_clk new_AGEMA_reg_buffer_1589 ( .C (clk), .D (new_AGEMA_signal_4364), .Q (new_AGEMA_signal_4365) ) ;
    buf_clk new_AGEMA_reg_buffer_1595 ( .C (clk), .D (new_AGEMA_signal_4370), .Q (new_AGEMA_signal_4371) ) ;
    buf_clk new_AGEMA_reg_buffer_1601 ( .C (clk), .D (new_AGEMA_signal_4376), .Q (new_AGEMA_signal_4377) ) ;
    buf_clk new_AGEMA_reg_buffer_1607 ( .C (clk), .D (new_AGEMA_signal_4382), .Q (new_AGEMA_signal_4383) ) ;
    buf_clk new_AGEMA_reg_buffer_1613 ( .C (clk), .D (new_AGEMA_signal_4388), .Q (new_AGEMA_signal_4389) ) ;
    buf_clk new_AGEMA_reg_buffer_1619 ( .C (clk), .D (new_AGEMA_signal_4394), .Q (new_AGEMA_signal_4395) ) ;
    buf_clk new_AGEMA_reg_buffer_1625 ( .C (clk), .D (new_AGEMA_signal_4400), .Q (new_AGEMA_signal_4401) ) ;
    buf_clk new_AGEMA_reg_buffer_1631 ( .C (clk), .D (new_AGEMA_signal_4406), .Q (new_AGEMA_signal_4407) ) ;
    buf_clk new_AGEMA_reg_buffer_1637 ( .C (clk), .D (new_AGEMA_signal_4412), .Q (new_AGEMA_signal_4413) ) ;
    buf_clk new_AGEMA_reg_buffer_1643 ( .C (clk), .D (new_AGEMA_signal_4418), .Q (new_AGEMA_signal_4419) ) ;
    buf_clk new_AGEMA_reg_buffer_1649 ( .C (clk), .D (new_AGEMA_signal_4424), .Q (new_AGEMA_signal_4425) ) ;
    buf_clk new_AGEMA_reg_buffer_1655 ( .C (clk), .D (new_AGEMA_signal_4430), .Q (new_AGEMA_signal_4431) ) ;
    buf_clk new_AGEMA_reg_buffer_1661 ( .C (clk), .D (new_AGEMA_signal_4436), .Q (new_AGEMA_signal_4437) ) ;
    buf_clk new_AGEMA_reg_buffer_1667 ( .C (clk), .D (new_AGEMA_signal_4442), .Q (new_AGEMA_signal_4443) ) ;
    buf_clk new_AGEMA_reg_buffer_1673 ( .C (clk), .D (new_AGEMA_signal_4448), .Q (new_AGEMA_signal_4449) ) ;
    buf_clk new_AGEMA_reg_buffer_1679 ( .C (clk), .D (new_AGEMA_signal_4454), .Q (new_AGEMA_signal_4455) ) ;
    buf_clk new_AGEMA_reg_buffer_1685 ( .C (clk), .D (new_AGEMA_signal_4460), .Q (new_AGEMA_signal_4461) ) ;
    buf_clk new_AGEMA_reg_buffer_1691 ( .C (clk), .D (new_AGEMA_signal_4466), .Q (new_AGEMA_signal_4467) ) ;
    buf_clk new_AGEMA_reg_buffer_1697 ( .C (clk), .D (new_AGEMA_signal_4472), .Q (new_AGEMA_signal_4473) ) ;
    buf_clk new_AGEMA_reg_buffer_1703 ( .C (clk), .D (new_AGEMA_signal_4478), .Q (new_AGEMA_signal_4479) ) ;
    buf_clk new_AGEMA_reg_buffer_1709 ( .C (clk), .D (new_AGEMA_signal_4484), .Q (new_AGEMA_signal_4485) ) ;
    buf_clk new_AGEMA_reg_buffer_1715 ( .C (clk), .D (new_AGEMA_signal_4490), .Q (new_AGEMA_signal_4491) ) ;
    buf_clk new_AGEMA_reg_buffer_1721 ( .C (clk), .D (new_AGEMA_signal_4496), .Q (new_AGEMA_signal_4497) ) ;
    buf_clk new_AGEMA_reg_buffer_1727 ( .C (clk), .D (new_AGEMA_signal_4502), .Q (new_AGEMA_signal_4503) ) ;
    buf_clk new_AGEMA_reg_buffer_1733 ( .C (clk), .D (new_AGEMA_signal_4508), .Q (new_AGEMA_signal_4509) ) ;
    buf_clk new_AGEMA_reg_buffer_1739 ( .C (clk), .D (new_AGEMA_signal_4514), .Q (new_AGEMA_signal_4515) ) ;
    buf_clk new_AGEMA_reg_buffer_1745 ( .C (clk), .D (new_AGEMA_signal_4520), .Q (new_AGEMA_signal_4521) ) ;
    buf_clk new_AGEMA_reg_buffer_1751 ( .C (clk), .D (new_AGEMA_signal_4526), .Q (new_AGEMA_signal_4527) ) ;
    buf_clk new_AGEMA_reg_buffer_1757 ( .C (clk), .D (new_AGEMA_signal_4532), .Q (new_AGEMA_signal_4533) ) ;
    buf_clk new_AGEMA_reg_buffer_1763 ( .C (clk), .D (new_AGEMA_signal_4538), .Q (new_AGEMA_signal_4539) ) ;
    buf_clk new_AGEMA_reg_buffer_1769 ( .C (clk), .D (new_AGEMA_signal_4544), .Q (new_AGEMA_signal_4545) ) ;
    buf_clk new_AGEMA_reg_buffer_1775 ( .C (clk), .D (new_AGEMA_signal_4550), .Q (new_AGEMA_signal_4551) ) ;
    buf_clk new_AGEMA_reg_buffer_1781 ( .C (clk), .D (new_AGEMA_signal_4556), .Q (new_AGEMA_signal_4557) ) ;
    buf_clk new_AGEMA_reg_buffer_1787 ( .C (clk), .D (new_AGEMA_signal_4562), .Q (new_AGEMA_signal_4563) ) ;
    buf_clk new_AGEMA_reg_buffer_1793 ( .C (clk), .D (new_AGEMA_signal_4568), .Q (new_AGEMA_signal_4569) ) ;
    buf_clk new_AGEMA_reg_buffer_1799 ( .C (clk), .D (new_AGEMA_signal_4574), .Q (new_AGEMA_signal_4575) ) ;
    buf_clk new_AGEMA_reg_buffer_1805 ( .C (clk), .D (new_AGEMA_signal_4580), .Q (new_AGEMA_signal_4581) ) ;
    buf_clk new_AGEMA_reg_buffer_1811 ( .C (clk), .D (new_AGEMA_signal_4586), .Q (new_AGEMA_signal_4587) ) ;
    buf_clk new_AGEMA_reg_buffer_1817 ( .C (clk), .D (new_AGEMA_signal_4592), .Q (new_AGEMA_signal_4593) ) ;
    buf_clk new_AGEMA_reg_buffer_1823 ( .C (clk), .D (new_AGEMA_signal_4598), .Q (new_AGEMA_signal_4599) ) ;
    buf_clk new_AGEMA_reg_buffer_1829 ( .C (clk), .D (new_AGEMA_signal_4604), .Q (new_AGEMA_signal_4605) ) ;
    buf_clk new_AGEMA_reg_buffer_1835 ( .C (clk), .D (new_AGEMA_signal_4610), .Q (new_AGEMA_signal_4611) ) ;
    buf_clk new_AGEMA_reg_buffer_1841 ( .C (clk), .D (new_AGEMA_signal_4616), .Q (new_AGEMA_signal_4617) ) ;
    buf_clk new_AGEMA_reg_buffer_1847 ( .C (clk), .D (new_AGEMA_signal_4622), .Q (new_AGEMA_signal_4623) ) ;
    buf_clk new_AGEMA_reg_buffer_1853 ( .C (clk), .D (new_AGEMA_signal_4628), .Q (new_AGEMA_signal_4629) ) ;
    buf_clk new_AGEMA_reg_buffer_1859 ( .C (clk), .D (new_AGEMA_signal_4634), .Q (new_AGEMA_signal_4635) ) ;
    buf_clk new_AGEMA_reg_buffer_1865 ( .C (clk), .D (new_AGEMA_signal_4640), .Q (new_AGEMA_signal_4641) ) ;
    buf_clk new_AGEMA_reg_buffer_1871 ( .C (clk), .D (new_AGEMA_signal_4646), .Q (new_AGEMA_signal_4647) ) ;
    buf_clk new_AGEMA_reg_buffer_1877 ( .C (clk), .D (new_AGEMA_signal_4652), .Q (new_AGEMA_signal_4653) ) ;
    buf_clk new_AGEMA_reg_buffer_1883 ( .C (clk), .D (new_AGEMA_signal_4658), .Q (new_AGEMA_signal_4659) ) ;
    buf_clk new_AGEMA_reg_buffer_1889 ( .C (clk), .D (new_AGEMA_signal_4664), .Q (new_AGEMA_signal_4665) ) ;
    buf_clk new_AGEMA_reg_buffer_1895 ( .C (clk), .D (new_AGEMA_signal_4670), .Q (new_AGEMA_signal_4671) ) ;
    buf_clk new_AGEMA_reg_buffer_1901 ( .C (clk), .D (new_AGEMA_signal_4676), .Q (new_AGEMA_signal_4677) ) ;
    buf_clk new_AGEMA_reg_buffer_1907 ( .C (clk), .D (new_AGEMA_signal_4682), .Q (new_AGEMA_signal_4683) ) ;
    buf_clk new_AGEMA_reg_buffer_1913 ( .C (clk), .D (new_AGEMA_signal_4688), .Q (new_AGEMA_signal_4689) ) ;
    buf_clk new_AGEMA_reg_buffer_1919 ( .C (clk), .D (new_AGEMA_signal_4694), .Q (new_AGEMA_signal_4695) ) ;
    buf_clk new_AGEMA_reg_buffer_1925 ( .C (clk), .D (new_AGEMA_signal_4700), .Q (new_AGEMA_signal_4701) ) ;
    buf_clk new_AGEMA_reg_buffer_1931 ( .C (clk), .D (new_AGEMA_signal_4706), .Q (new_AGEMA_signal_4707) ) ;
    buf_clk new_AGEMA_reg_buffer_1937 ( .C (clk), .D (new_AGEMA_signal_4712), .Q (new_AGEMA_signal_4713) ) ;
    buf_clk new_AGEMA_reg_buffer_1943 ( .C (clk), .D (new_AGEMA_signal_4718), .Q (new_AGEMA_signal_4719) ) ;
    buf_clk new_AGEMA_reg_buffer_1949 ( .C (clk), .D (new_AGEMA_signal_4724), .Q (new_AGEMA_signal_4725) ) ;
    buf_clk new_AGEMA_reg_buffer_1955 ( .C (clk), .D (new_AGEMA_signal_4730), .Q (new_AGEMA_signal_4731) ) ;
    buf_clk new_AGEMA_reg_buffer_1961 ( .C (clk), .D (new_AGEMA_signal_4736), .Q (new_AGEMA_signal_4737) ) ;
    buf_clk new_AGEMA_reg_buffer_1967 ( .C (clk), .D (new_AGEMA_signal_4742), .Q (new_AGEMA_signal_4743) ) ;
    buf_clk new_AGEMA_reg_buffer_1973 ( .C (clk), .D (new_AGEMA_signal_4748), .Q (new_AGEMA_signal_4749) ) ;
    buf_clk new_AGEMA_reg_buffer_1979 ( .C (clk), .D (new_AGEMA_signal_4754), .Q (new_AGEMA_signal_4755) ) ;
    buf_clk new_AGEMA_reg_buffer_1985 ( .C (clk), .D (new_AGEMA_signal_4760), .Q (new_AGEMA_signal_4761) ) ;
    buf_clk new_AGEMA_reg_buffer_1991 ( .C (clk), .D (new_AGEMA_signal_4766), .Q (new_AGEMA_signal_4767) ) ;
    buf_clk new_AGEMA_reg_buffer_1997 ( .C (clk), .D (new_AGEMA_signal_4772), .Q (new_AGEMA_signal_4773) ) ;
    buf_clk new_AGEMA_reg_buffer_2003 ( .C (clk), .D (new_AGEMA_signal_4778), .Q (new_AGEMA_signal_4779) ) ;
    buf_clk new_AGEMA_reg_buffer_2009 ( .C (clk), .D (new_AGEMA_signal_4784), .Q (new_AGEMA_signal_4785) ) ;
    buf_clk new_AGEMA_reg_buffer_2015 ( .C (clk), .D (new_AGEMA_signal_4790), .Q (new_AGEMA_signal_4791) ) ;
    buf_clk new_AGEMA_reg_buffer_2021 ( .C (clk), .D (new_AGEMA_signal_4796), .Q (new_AGEMA_signal_4797) ) ;
    buf_clk new_AGEMA_reg_buffer_2027 ( .C (clk), .D (new_AGEMA_signal_4802), .Q (new_AGEMA_signal_4803) ) ;
    buf_clk new_AGEMA_reg_buffer_2033 ( .C (clk), .D (new_AGEMA_signal_4808), .Q (new_AGEMA_signal_4809) ) ;
    buf_clk new_AGEMA_reg_buffer_2039 ( .C (clk), .D (new_AGEMA_signal_4814), .Q (new_AGEMA_signal_4815) ) ;
    buf_clk new_AGEMA_reg_buffer_2045 ( .C (clk), .D (new_AGEMA_signal_4820), .Q (new_AGEMA_signal_4821) ) ;
    buf_clk new_AGEMA_reg_buffer_2051 ( .C (clk), .D (new_AGEMA_signal_4826), .Q (new_AGEMA_signal_4827) ) ;
    buf_clk new_AGEMA_reg_buffer_2057 ( .C (clk), .D (new_AGEMA_signal_4832), .Q (new_AGEMA_signal_4833) ) ;
    buf_clk new_AGEMA_reg_buffer_2063 ( .C (clk), .D (new_AGEMA_signal_4838), .Q (new_AGEMA_signal_4839) ) ;
    buf_clk new_AGEMA_reg_buffer_2069 ( .C (clk), .D (new_AGEMA_signal_4844), .Q (new_AGEMA_signal_4845) ) ;
    buf_clk new_AGEMA_reg_buffer_2075 ( .C (clk), .D (new_AGEMA_signal_4850), .Q (new_AGEMA_signal_4851) ) ;
    buf_clk new_AGEMA_reg_buffer_2081 ( .C (clk), .D (new_AGEMA_signal_4856), .Q (new_AGEMA_signal_4857) ) ;
    buf_clk new_AGEMA_reg_buffer_2087 ( .C (clk), .D (new_AGEMA_signal_4862), .Q (new_AGEMA_signal_4863) ) ;
    buf_clk new_AGEMA_reg_buffer_2093 ( .C (clk), .D (new_AGEMA_signal_4868), .Q (new_AGEMA_signal_4869) ) ;
    buf_clk new_AGEMA_reg_buffer_2099 ( .C (clk), .D (new_AGEMA_signal_4874), .Q (new_AGEMA_signal_4875) ) ;
    buf_clk new_AGEMA_reg_buffer_2105 ( .C (clk), .D (new_AGEMA_signal_4880), .Q (new_AGEMA_signal_4881) ) ;
    buf_clk new_AGEMA_reg_buffer_2111 ( .C (clk), .D (new_AGEMA_signal_4886), .Q (new_AGEMA_signal_4887) ) ;
    buf_clk new_AGEMA_reg_buffer_2117 ( .C (clk), .D (new_AGEMA_signal_4892), .Q (new_AGEMA_signal_4893) ) ;
    buf_clk new_AGEMA_reg_buffer_2123 ( .C (clk), .D (new_AGEMA_signal_4898), .Q (new_AGEMA_signal_4899) ) ;
    buf_clk new_AGEMA_reg_buffer_2129 ( .C (clk), .D (new_AGEMA_signal_4904), .Q (new_AGEMA_signal_4905) ) ;
    buf_clk new_AGEMA_reg_buffer_2135 ( .C (clk), .D (new_AGEMA_signal_4910), .Q (new_AGEMA_signal_4911) ) ;
    buf_clk new_AGEMA_reg_buffer_2141 ( .C (clk), .D (new_AGEMA_signal_4916), .Q (new_AGEMA_signal_4917) ) ;
    buf_clk new_AGEMA_reg_buffer_2147 ( .C (clk), .D (new_AGEMA_signal_4922), .Q (new_AGEMA_signal_4923) ) ;
    buf_clk new_AGEMA_reg_buffer_2153 ( .C (clk), .D (new_AGEMA_signal_4928), .Q (new_AGEMA_signal_4929) ) ;
    buf_clk new_AGEMA_reg_buffer_2159 ( .C (clk), .D (new_AGEMA_signal_4934), .Q (new_AGEMA_signal_4935) ) ;
    buf_clk new_AGEMA_reg_buffer_2165 ( .C (clk), .D (new_AGEMA_signal_4940), .Q (new_AGEMA_signal_4941) ) ;
    buf_clk new_AGEMA_reg_buffer_2171 ( .C (clk), .D (new_AGEMA_signal_4946), .Q (new_AGEMA_signal_4947) ) ;
    buf_clk new_AGEMA_reg_buffer_2177 ( .C (clk), .D (new_AGEMA_signal_4952), .Q (new_AGEMA_signal_4953) ) ;
    buf_clk new_AGEMA_reg_buffer_2183 ( .C (clk), .D (new_AGEMA_signal_4958), .Q (new_AGEMA_signal_4959) ) ;
    buf_clk new_AGEMA_reg_buffer_2189 ( .C (clk), .D (new_AGEMA_signal_4964), .Q (new_AGEMA_signal_4965) ) ;
    buf_clk new_AGEMA_reg_buffer_2195 ( .C (clk), .D (new_AGEMA_signal_4970), .Q (new_AGEMA_signal_4971) ) ;
    buf_clk new_AGEMA_reg_buffer_2201 ( .C (clk), .D (new_AGEMA_signal_4976), .Q (new_AGEMA_signal_4977) ) ;
    buf_clk new_AGEMA_reg_buffer_2207 ( .C (clk), .D (new_AGEMA_signal_4982), .Q (new_AGEMA_signal_4983) ) ;
    buf_clk new_AGEMA_reg_buffer_2213 ( .C (clk), .D (new_AGEMA_signal_4988), .Q (new_AGEMA_signal_4989) ) ;
    buf_clk new_AGEMA_reg_buffer_2219 ( .C (clk), .D (new_AGEMA_signal_4994), .Q (new_AGEMA_signal_4995) ) ;
    buf_clk new_AGEMA_reg_buffer_2225 ( .C (clk), .D (new_AGEMA_signal_5000), .Q (new_AGEMA_signal_5001) ) ;
    buf_clk new_AGEMA_reg_buffer_2231 ( .C (clk), .D (new_AGEMA_signal_5006), .Q (new_AGEMA_signal_5007) ) ;
    buf_clk new_AGEMA_reg_buffer_2237 ( .C (clk), .D (new_AGEMA_signal_5012), .Q (new_AGEMA_signal_5013) ) ;
    buf_clk new_AGEMA_reg_buffer_2243 ( .C (clk), .D (new_AGEMA_signal_5018), .Q (new_AGEMA_signal_5019) ) ;
    buf_clk new_AGEMA_reg_buffer_2249 ( .C (clk), .D (new_AGEMA_signal_5024), .Q (new_AGEMA_signal_5025) ) ;
    buf_clk new_AGEMA_reg_buffer_2255 ( .C (clk), .D (new_AGEMA_signal_5030), .Q (new_AGEMA_signal_5031) ) ;
    buf_clk new_AGEMA_reg_buffer_2261 ( .C (clk), .D (new_AGEMA_signal_5036), .Q (new_AGEMA_signal_5037) ) ;
    buf_clk new_AGEMA_reg_buffer_2267 ( .C (clk), .D (new_AGEMA_signal_5042), .Q (new_AGEMA_signal_5043) ) ;
    buf_clk new_AGEMA_reg_buffer_2273 ( .C (clk), .D (new_AGEMA_signal_5048), .Q (new_AGEMA_signal_5049) ) ;
    buf_clk new_AGEMA_reg_buffer_2279 ( .C (clk), .D (new_AGEMA_signal_5054), .Q (new_AGEMA_signal_5055) ) ;
    buf_clk new_AGEMA_reg_buffer_2285 ( .C (clk), .D (new_AGEMA_signal_5060), .Q (new_AGEMA_signal_5061) ) ;
    buf_clk new_AGEMA_reg_buffer_2291 ( .C (clk), .D (new_AGEMA_signal_5066), .Q (new_AGEMA_signal_5067) ) ;
    buf_clk new_AGEMA_reg_buffer_2297 ( .C (clk), .D (new_AGEMA_signal_5072), .Q (new_AGEMA_signal_5073) ) ;
    buf_clk new_AGEMA_reg_buffer_2303 ( .C (clk), .D (new_AGEMA_signal_5078), .Q (new_AGEMA_signal_5079) ) ;
    buf_clk new_AGEMA_reg_buffer_2309 ( .C (clk), .D (new_AGEMA_signal_5084), .Q (new_AGEMA_signal_5085) ) ;
    buf_clk new_AGEMA_reg_buffer_2315 ( .C (clk), .D (new_AGEMA_signal_5090), .Q (new_AGEMA_signal_5091) ) ;
    buf_clk new_AGEMA_reg_buffer_2321 ( .C (clk), .D (new_AGEMA_signal_5096), .Q (new_AGEMA_signal_5097) ) ;
    buf_clk new_AGEMA_reg_buffer_2327 ( .C (clk), .D (new_AGEMA_signal_5102), .Q (new_AGEMA_signal_5103) ) ;
    buf_clk new_AGEMA_reg_buffer_2333 ( .C (clk), .D (new_AGEMA_signal_5108), .Q (new_AGEMA_signal_5109) ) ;
    buf_clk new_AGEMA_reg_buffer_2339 ( .C (clk), .D (new_AGEMA_signal_5114), .Q (new_AGEMA_signal_5115) ) ;
    buf_clk new_AGEMA_reg_buffer_2345 ( .C (clk), .D (new_AGEMA_signal_5120), .Q (new_AGEMA_signal_5121) ) ;
    buf_clk new_AGEMA_reg_buffer_2351 ( .C (clk), .D (new_AGEMA_signal_5126), .Q (new_AGEMA_signal_5127) ) ;
    buf_clk new_AGEMA_reg_buffer_2357 ( .C (clk), .D (new_AGEMA_signal_5132), .Q (new_AGEMA_signal_5133) ) ;
    buf_clk new_AGEMA_reg_buffer_2361 ( .C (clk), .D (SubCellInst_SboxInst_0_n15), .Q (new_AGEMA_signal_5137) ) ;
    buf_clk new_AGEMA_reg_buffer_2363 ( .C (clk), .D (new_AGEMA_signal_1277), .Q (new_AGEMA_signal_5139) ) ;
    buf_clk new_AGEMA_reg_buffer_2365 ( .C (clk), .D (new_AGEMA_signal_1278), .Q (new_AGEMA_signal_5141) ) ;
    buf_clk new_AGEMA_reg_buffer_2367 ( .C (clk), .D (new_AGEMA_signal_3596), .Q (new_AGEMA_signal_5143) ) ;
    buf_clk new_AGEMA_reg_buffer_2369 ( .C (clk), .D (new_AGEMA_signal_3598), .Q (new_AGEMA_signal_5145) ) ;
    buf_clk new_AGEMA_reg_buffer_2371 ( .C (clk), .D (new_AGEMA_signal_3600), .Q (new_AGEMA_signal_5147) ) ;
    buf_clk new_AGEMA_reg_buffer_2373 ( .C (clk), .D (SubCellInst_SboxInst_0_n6), .Q (new_AGEMA_signal_5149) ) ;
    buf_clk new_AGEMA_reg_buffer_2375 ( .C (clk), .D (new_AGEMA_signal_1281), .Q (new_AGEMA_signal_5151) ) ;
    buf_clk new_AGEMA_reg_buffer_2377 ( .C (clk), .D (new_AGEMA_signal_1282), .Q (new_AGEMA_signal_5153) ) ;
    buf_clk new_AGEMA_reg_buffer_2379 ( .C (clk), .D (SubCellInst_SboxInst_1_n15), .Q (new_AGEMA_signal_5155) ) ;
    buf_clk new_AGEMA_reg_buffer_2381 ( .C (clk), .D (new_AGEMA_signal_1289), .Q (new_AGEMA_signal_5157) ) ;
    buf_clk new_AGEMA_reg_buffer_2383 ( .C (clk), .D (new_AGEMA_signal_1290), .Q (new_AGEMA_signal_5159) ) ;
    buf_clk new_AGEMA_reg_buffer_2385 ( .C (clk), .D (new_AGEMA_signal_3620), .Q (new_AGEMA_signal_5161) ) ;
    buf_clk new_AGEMA_reg_buffer_2387 ( .C (clk), .D (new_AGEMA_signal_3622), .Q (new_AGEMA_signal_5163) ) ;
    buf_clk new_AGEMA_reg_buffer_2389 ( .C (clk), .D (new_AGEMA_signal_3624), .Q (new_AGEMA_signal_5165) ) ;
    buf_clk new_AGEMA_reg_buffer_2391 ( .C (clk), .D (SubCellInst_SboxInst_1_n6), .Q (new_AGEMA_signal_5167) ) ;
    buf_clk new_AGEMA_reg_buffer_2393 ( .C (clk), .D (new_AGEMA_signal_1293), .Q (new_AGEMA_signal_5169) ) ;
    buf_clk new_AGEMA_reg_buffer_2395 ( .C (clk), .D (new_AGEMA_signal_1294), .Q (new_AGEMA_signal_5171) ) ;
    buf_clk new_AGEMA_reg_buffer_2397 ( .C (clk), .D (SubCellInst_SboxInst_2_n15), .Q (new_AGEMA_signal_5173) ) ;
    buf_clk new_AGEMA_reg_buffer_2399 ( .C (clk), .D (new_AGEMA_signal_1301), .Q (new_AGEMA_signal_5175) ) ;
    buf_clk new_AGEMA_reg_buffer_2401 ( .C (clk), .D (new_AGEMA_signal_1302), .Q (new_AGEMA_signal_5177) ) ;
    buf_clk new_AGEMA_reg_buffer_2403 ( .C (clk), .D (new_AGEMA_signal_3644), .Q (new_AGEMA_signal_5179) ) ;
    buf_clk new_AGEMA_reg_buffer_2405 ( .C (clk), .D (new_AGEMA_signal_3646), .Q (new_AGEMA_signal_5181) ) ;
    buf_clk new_AGEMA_reg_buffer_2407 ( .C (clk), .D (new_AGEMA_signal_3648), .Q (new_AGEMA_signal_5183) ) ;
    buf_clk new_AGEMA_reg_buffer_2409 ( .C (clk), .D (SubCellInst_SboxInst_2_n6), .Q (new_AGEMA_signal_5185) ) ;
    buf_clk new_AGEMA_reg_buffer_2411 ( .C (clk), .D (new_AGEMA_signal_1305), .Q (new_AGEMA_signal_5187) ) ;
    buf_clk new_AGEMA_reg_buffer_2413 ( .C (clk), .D (new_AGEMA_signal_1306), .Q (new_AGEMA_signal_5189) ) ;
    buf_clk new_AGEMA_reg_buffer_2415 ( .C (clk), .D (SubCellInst_SboxInst_3_n15), .Q (new_AGEMA_signal_5191) ) ;
    buf_clk new_AGEMA_reg_buffer_2417 ( .C (clk), .D (new_AGEMA_signal_1313), .Q (new_AGEMA_signal_5193) ) ;
    buf_clk new_AGEMA_reg_buffer_2419 ( .C (clk), .D (new_AGEMA_signal_1314), .Q (new_AGEMA_signal_5195) ) ;
    buf_clk new_AGEMA_reg_buffer_2421 ( .C (clk), .D (new_AGEMA_signal_3668), .Q (new_AGEMA_signal_5197) ) ;
    buf_clk new_AGEMA_reg_buffer_2423 ( .C (clk), .D (new_AGEMA_signal_3670), .Q (new_AGEMA_signal_5199) ) ;
    buf_clk new_AGEMA_reg_buffer_2425 ( .C (clk), .D (new_AGEMA_signal_3672), .Q (new_AGEMA_signal_5201) ) ;
    buf_clk new_AGEMA_reg_buffer_2427 ( .C (clk), .D (SubCellInst_SboxInst_3_n6), .Q (new_AGEMA_signal_5203) ) ;
    buf_clk new_AGEMA_reg_buffer_2429 ( .C (clk), .D (new_AGEMA_signal_1317), .Q (new_AGEMA_signal_5205) ) ;
    buf_clk new_AGEMA_reg_buffer_2431 ( .C (clk), .D (new_AGEMA_signal_1318), .Q (new_AGEMA_signal_5207) ) ;
    buf_clk new_AGEMA_reg_buffer_2433 ( .C (clk), .D (SubCellInst_SboxInst_4_n15), .Q (new_AGEMA_signal_5209) ) ;
    buf_clk new_AGEMA_reg_buffer_2435 ( .C (clk), .D (new_AGEMA_signal_1325), .Q (new_AGEMA_signal_5211) ) ;
    buf_clk new_AGEMA_reg_buffer_2437 ( .C (clk), .D (new_AGEMA_signal_1326), .Q (new_AGEMA_signal_5213) ) ;
    buf_clk new_AGEMA_reg_buffer_2439 ( .C (clk), .D (new_AGEMA_signal_3692), .Q (new_AGEMA_signal_5215) ) ;
    buf_clk new_AGEMA_reg_buffer_2441 ( .C (clk), .D (new_AGEMA_signal_3694), .Q (new_AGEMA_signal_5217) ) ;
    buf_clk new_AGEMA_reg_buffer_2443 ( .C (clk), .D (new_AGEMA_signal_3696), .Q (new_AGEMA_signal_5219) ) ;
    buf_clk new_AGEMA_reg_buffer_2445 ( .C (clk), .D (SubCellInst_SboxInst_4_n6), .Q (new_AGEMA_signal_5221) ) ;
    buf_clk new_AGEMA_reg_buffer_2447 ( .C (clk), .D (new_AGEMA_signal_1329), .Q (new_AGEMA_signal_5223) ) ;
    buf_clk new_AGEMA_reg_buffer_2449 ( .C (clk), .D (new_AGEMA_signal_1330), .Q (new_AGEMA_signal_5225) ) ;
    buf_clk new_AGEMA_reg_buffer_2451 ( .C (clk), .D (SubCellInst_SboxInst_5_n15), .Q (new_AGEMA_signal_5227) ) ;
    buf_clk new_AGEMA_reg_buffer_2453 ( .C (clk), .D (new_AGEMA_signal_1337), .Q (new_AGEMA_signal_5229) ) ;
    buf_clk new_AGEMA_reg_buffer_2455 ( .C (clk), .D (new_AGEMA_signal_1338), .Q (new_AGEMA_signal_5231) ) ;
    buf_clk new_AGEMA_reg_buffer_2457 ( .C (clk), .D (new_AGEMA_signal_3716), .Q (new_AGEMA_signal_5233) ) ;
    buf_clk new_AGEMA_reg_buffer_2459 ( .C (clk), .D (new_AGEMA_signal_3718), .Q (new_AGEMA_signal_5235) ) ;
    buf_clk new_AGEMA_reg_buffer_2461 ( .C (clk), .D (new_AGEMA_signal_3720), .Q (new_AGEMA_signal_5237) ) ;
    buf_clk new_AGEMA_reg_buffer_2463 ( .C (clk), .D (SubCellInst_SboxInst_5_n6), .Q (new_AGEMA_signal_5239) ) ;
    buf_clk new_AGEMA_reg_buffer_2465 ( .C (clk), .D (new_AGEMA_signal_1341), .Q (new_AGEMA_signal_5241) ) ;
    buf_clk new_AGEMA_reg_buffer_2467 ( .C (clk), .D (new_AGEMA_signal_1342), .Q (new_AGEMA_signal_5243) ) ;
    buf_clk new_AGEMA_reg_buffer_2469 ( .C (clk), .D (SubCellInst_SboxInst_6_n15), .Q (new_AGEMA_signal_5245) ) ;
    buf_clk new_AGEMA_reg_buffer_2471 ( .C (clk), .D (new_AGEMA_signal_1349), .Q (new_AGEMA_signal_5247) ) ;
    buf_clk new_AGEMA_reg_buffer_2473 ( .C (clk), .D (new_AGEMA_signal_1350), .Q (new_AGEMA_signal_5249) ) ;
    buf_clk new_AGEMA_reg_buffer_2475 ( .C (clk), .D (new_AGEMA_signal_3740), .Q (new_AGEMA_signal_5251) ) ;
    buf_clk new_AGEMA_reg_buffer_2477 ( .C (clk), .D (new_AGEMA_signal_3742), .Q (new_AGEMA_signal_5253) ) ;
    buf_clk new_AGEMA_reg_buffer_2479 ( .C (clk), .D (new_AGEMA_signal_3744), .Q (new_AGEMA_signal_5255) ) ;
    buf_clk new_AGEMA_reg_buffer_2481 ( .C (clk), .D (SubCellInst_SboxInst_6_n6), .Q (new_AGEMA_signal_5257) ) ;
    buf_clk new_AGEMA_reg_buffer_2483 ( .C (clk), .D (new_AGEMA_signal_1353), .Q (new_AGEMA_signal_5259) ) ;
    buf_clk new_AGEMA_reg_buffer_2485 ( .C (clk), .D (new_AGEMA_signal_1354), .Q (new_AGEMA_signal_5261) ) ;
    buf_clk new_AGEMA_reg_buffer_2487 ( .C (clk), .D (SubCellInst_SboxInst_7_n15), .Q (new_AGEMA_signal_5263) ) ;
    buf_clk new_AGEMA_reg_buffer_2489 ( .C (clk), .D (new_AGEMA_signal_1361), .Q (new_AGEMA_signal_5265) ) ;
    buf_clk new_AGEMA_reg_buffer_2491 ( .C (clk), .D (new_AGEMA_signal_1362), .Q (new_AGEMA_signal_5267) ) ;
    buf_clk new_AGEMA_reg_buffer_2493 ( .C (clk), .D (new_AGEMA_signal_3764), .Q (new_AGEMA_signal_5269) ) ;
    buf_clk new_AGEMA_reg_buffer_2495 ( .C (clk), .D (new_AGEMA_signal_3766), .Q (new_AGEMA_signal_5271) ) ;
    buf_clk new_AGEMA_reg_buffer_2497 ( .C (clk), .D (new_AGEMA_signal_3768), .Q (new_AGEMA_signal_5273) ) ;
    buf_clk new_AGEMA_reg_buffer_2499 ( .C (clk), .D (SubCellInst_SboxInst_7_n6), .Q (new_AGEMA_signal_5275) ) ;
    buf_clk new_AGEMA_reg_buffer_2501 ( .C (clk), .D (new_AGEMA_signal_1365), .Q (new_AGEMA_signal_5277) ) ;
    buf_clk new_AGEMA_reg_buffer_2503 ( .C (clk), .D (new_AGEMA_signal_1366), .Q (new_AGEMA_signal_5279) ) ;
    buf_clk new_AGEMA_reg_buffer_2505 ( .C (clk), .D (SubCellInst_SboxInst_8_n15), .Q (new_AGEMA_signal_5281) ) ;
    buf_clk new_AGEMA_reg_buffer_2507 ( .C (clk), .D (new_AGEMA_signal_1373), .Q (new_AGEMA_signal_5283) ) ;
    buf_clk new_AGEMA_reg_buffer_2509 ( .C (clk), .D (new_AGEMA_signal_1374), .Q (new_AGEMA_signal_5285) ) ;
    buf_clk new_AGEMA_reg_buffer_2511 ( .C (clk), .D (new_AGEMA_signal_3788), .Q (new_AGEMA_signal_5287) ) ;
    buf_clk new_AGEMA_reg_buffer_2513 ( .C (clk), .D (new_AGEMA_signal_3790), .Q (new_AGEMA_signal_5289) ) ;
    buf_clk new_AGEMA_reg_buffer_2515 ( .C (clk), .D (new_AGEMA_signal_3792), .Q (new_AGEMA_signal_5291) ) ;
    buf_clk new_AGEMA_reg_buffer_2517 ( .C (clk), .D (SubCellInst_SboxInst_8_n6), .Q (new_AGEMA_signal_5293) ) ;
    buf_clk new_AGEMA_reg_buffer_2519 ( .C (clk), .D (new_AGEMA_signal_1377), .Q (new_AGEMA_signal_5295) ) ;
    buf_clk new_AGEMA_reg_buffer_2521 ( .C (clk), .D (new_AGEMA_signal_1378), .Q (new_AGEMA_signal_5297) ) ;
    buf_clk new_AGEMA_reg_buffer_2523 ( .C (clk), .D (SubCellInst_SboxInst_9_n15), .Q (new_AGEMA_signal_5299) ) ;
    buf_clk new_AGEMA_reg_buffer_2525 ( .C (clk), .D (new_AGEMA_signal_1385), .Q (new_AGEMA_signal_5301) ) ;
    buf_clk new_AGEMA_reg_buffer_2527 ( .C (clk), .D (new_AGEMA_signal_1386), .Q (new_AGEMA_signal_5303) ) ;
    buf_clk new_AGEMA_reg_buffer_2529 ( .C (clk), .D (new_AGEMA_signal_3812), .Q (new_AGEMA_signal_5305) ) ;
    buf_clk new_AGEMA_reg_buffer_2531 ( .C (clk), .D (new_AGEMA_signal_3814), .Q (new_AGEMA_signal_5307) ) ;
    buf_clk new_AGEMA_reg_buffer_2533 ( .C (clk), .D (new_AGEMA_signal_3816), .Q (new_AGEMA_signal_5309) ) ;
    buf_clk new_AGEMA_reg_buffer_2535 ( .C (clk), .D (SubCellInst_SboxInst_9_n6), .Q (new_AGEMA_signal_5311) ) ;
    buf_clk new_AGEMA_reg_buffer_2537 ( .C (clk), .D (new_AGEMA_signal_1389), .Q (new_AGEMA_signal_5313) ) ;
    buf_clk new_AGEMA_reg_buffer_2539 ( .C (clk), .D (new_AGEMA_signal_1390), .Q (new_AGEMA_signal_5315) ) ;
    buf_clk new_AGEMA_reg_buffer_2541 ( .C (clk), .D (SubCellInst_SboxInst_10_n15), .Q (new_AGEMA_signal_5317) ) ;
    buf_clk new_AGEMA_reg_buffer_2543 ( .C (clk), .D (new_AGEMA_signal_1397), .Q (new_AGEMA_signal_5319) ) ;
    buf_clk new_AGEMA_reg_buffer_2545 ( .C (clk), .D (new_AGEMA_signal_1398), .Q (new_AGEMA_signal_5321) ) ;
    buf_clk new_AGEMA_reg_buffer_2547 ( .C (clk), .D (new_AGEMA_signal_3836), .Q (new_AGEMA_signal_5323) ) ;
    buf_clk new_AGEMA_reg_buffer_2549 ( .C (clk), .D (new_AGEMA_signal_3838), .Q (new_AGEMA_signal_5325) ) ;
    buf_clk new_AGEMA_reg_buffer_2551 ( .C (clk), .D (new_AGEMA_signal_3840), .Q (new_AGEMA_signal_5327) ) ;
    buf_clk new_AGEMA_reg_buffer_2553 ( .C (clk), .D (SubCellInst_SboxInst_10_n6), .Q (new_AGEMA_signal_5329) ) ;
    buf_clk new_AGEMA_reg_buffer_2555 ( .C (clk), .D (new_AGEMA_signal_1401), .Q (new_AGEMA_signal_5331) ) ;
    buf_clk new_AGEMA_reg_buffer_2557 ( .C (clk), .D (new_AGEMA_signal_1402), .Q (new_AGEMA_signal_5333) ) ;
    buf_clk new_AGEMA_reg_buffer_2559 ( .C (clk), .D (SubCellInst_SboxInst_11_n15), .Q (new_AGEMA_signal_5335) ) ;
    buf_clk new_AGEMA_reg_buffer_2561 ( .C (clk), .D (new_AGEMA_signal_1409), .Q (new_AGEMA_signal_5337) ) ;
    buf_clk new_AGEMA_reg_buffer_2563 ( .C (clk), .D (new_AGEMA_signal_1410), .Q (new_AGEMA_signal_5339) ) ;
    buf_clk new_AGEMA_reg_buffer_2565 ( .C (clk), .D (new_AGEMA_signal_3860), .Q (new_AGEMA_signal_5341) ) ;
    buf_clk new_AGEMA_reg_buffer_2567 ( .C (clk), .D (new_AGEMA_signal_3862), .Q (new_AGEMA_signal_5343) ) ;
    buf_clk new_AGEMA_reg_buffer_2569 ( .C (clk), .D (new_AGEMA_signal_3864), .Q (new_AGEMA_signal_5345) ) ;
    buf_clk new_AGEMA_reg_buffer_2571 ( .C (clk), .D (SubCellInst_SboxInst_11_n6), .Q (new_AGEMA_signal_5347) ) ;
    buf_clk new_AGEMA_reg_buffer_2573 ( .C (clk), .D (new_AGEMA_signal_1413), .Q (new_AGEMA_signal_5349) ) ;
    buf_clk new_AGEMA_reg_buffer_2575 ( .C (clk), .D (new_AGEMA_signal_1414), .Q (new_AGEMA_signal_5351) ) ;
    buf_clk new_AGEMA_reg_buffer_2577 ( .C (clk), .D (SubCellInst_SboxInst_12_n15), .Q (new_AGEMA_signal_5353) ) ;
    buf_clk new_AGEMA_reg_buffer_2579 ( .C (clk), .D (new_AGEMA_signal_1421), .Q (new_AGEMA_signal_5355) ) ;
    buf_clk new_AGEMA_reg_buffer_2581 ( .C (clk), .D (new_AGEMA_signal_1422), .Q (new_AGEMA_signal_5357) ) ;
    buf_clk new_AGEMA_reg_buffer_2583 ( .C (clk), .D (new_AGEMA_signal_3884), .Q (new_AGEMA_signal_5359) ) ;
    buf_clk new_AGEMA_reg_buffer_2585 ( .C (clk), .D (new_AGEMA_signal_3886), .Q (new_AGEMA_signal_5361) ) ;
    buf_clk new_AGEMA_reg_buffer_2587 ( .C (clk), .D (new_AGEMA_signal_3888), .Q (new_AGEMA_signal_5363) ) ;
    buf_clk new_AGEMA_reg_buffer_2589 ( .C (clk), .D (SubCellInst_SboxInst_12_n6), .Q (new_AGEMA_signal_5365) ) ;
    buf_clk new_AGEMA_reg_buffer_2591 ( .C (clk), .D (new_AGEMA_signal_1425), .Q (new_AGEMA_signal_5367) ) ;
    buf_clk new_AGEMA_reg_buffer_2593 ( .C (clk), .D (new_AGEMA_signal_1426), .Q (new_AGEMA_signal_5369) ) ;
    buf_clk new_AGEMA_reg_buffer_2595 ( .C (clk), .D (SubCellInst_SboxInst_13_n15), .Q (new_AGEMA_signal_5371) ) ;
    buf_clk new_AGEMA_reg_buffer_2597 ( .C (clk), .D (new_AGEMA_signal_1433), .Q (new_AGEMA_signal_5373) ) ;
    buf_clk new_AGEMA_reg_buffer_2599 ( .C (clk), .D (new_AGEMA_signal_1434), .Q (new_AGEMA_signal_5375) ) ;
    buf_clk new_AGEMA_reg_buffer_2601 ( .C (clk), .D (new_AGEMA_signal_3908), .Q (new_AGEMA_signal_5377) ) ;
    buf_clk new_AGEMA_reg_buffer_2603 ( .C (clk), .D (new_AGEMA_signal_3910), .Q (new_AGEMA_signal_5379) ) ;
    buf_clk new_AGEMA_reg_buffer_2605 ( .C (clk), .D (new_AGEMA_signal_3912), .Q (new_AGEMA_signal_5381) ) ;
    buf_clk new_AGEMA_reg_buffer_2607 ( .C (clk), .D (SubCellInst_SboxInst_13_n6), .Q (new_AGEMA_signal_5383) ) ;
    buf_clk new_AGEMA_reg_buffer_2609 ( .C (clk), .D (new_AGEMA_signal_1437), .Q (new_AGEMA_signal_5385) ) ;
    buf_clk new_AGEMA_reg_buffer_2611 ( .C (clk), .D (new_AGEMA_signal_1438), .Q (new_AGEMA_signal_5387) ) ;
    buf_clk new_AGEMA_reg_buffer_2613 ( .C (clk), .D (SubCellInst_SboxInst_14_n15), .Q (new_AGEMA_signal_5389) ) ;
    buf_clk new_AGEMA_reg_buffer_2615 ( .C (clk), .D (new_AGEMA_signal_1445), .Q (new_AGEMA_signal_5391) ) ;
    buf_clk new_AGEMA_reg_buffer_2617 ( .C (clk), .D (new_AGEMA_signal_1446), .Q (new_AGEMA_signal_5393) ) ;
    buf_clk new_AGEMA_reg_buffer_2619 ( .C (clk), .D (new_AGEMA_signal_3932), .Q (new_AGEMA_signal_5395) ) ;
    buf_clk new_AGEMA_reg_buffer_2621 ( .C (clk), .D (new_AGEMA_signal_3934), .Q (new_AGEMA_signal_5397) ) ;
    buf_clk new_AGEMA_reg_buffer_2623 ( .C (clk), .D (new_AGEMA_signal_3936), .Q (new_AGEMA_signal_5399) ) ;
    buf_clk new_AGEMA_reg_buffer_2625 ( .C (clk), .D (SubCellInst_SboxInst_14_n6), .Q (new_AGEMA_signal_5401) ) ;
    buf_clk new_AGEMA_reg_buffer_2627 ( .C (clk), .D (new_AGEMA_signal_1449), .Q (new_AGEMA_signal_5403) ) ;
    buf_clk new_AGEMA_reg_buffer_2629 ( .C (clk), .D (new_AGEMA_signal_1450), .Q (new_AGEMA_signal_5405) ) ;
    buf_clk new_AGEMA_reg_buffer_2631 ( .C (clk), .D (SubCellInst_SboxInst_15_n15), .Q (new_AGEMA_signal_5407) ) ;
    buf_clk new_AGEMA_reg_buffer_2633 ( .C (clk), .D (new_AGEMA_signal_1457), .Q (new_AGEMA_signal_5409) ) ;
    buf_clk new_AGEMA_reg_buffer_2635 ( .C (clk), .D (new_AGEMA_signal_1458), .Q (new_AGEMA_signal_5411) ) ;
    buf_clk new_AGEMA_reg_buffer_2637 ( .C (clk), .D (new_AGEMA_signal_3956), .Q (new_AGEMA_signal_5413) ) ;
    buf_clk new_AGEMA_reg_buffer_2639 ( .C (clk), .D (new_AGEMA_signal_3958), .Q (new_AGEMA_signal_5415) ) ;
    buf_clk new_AGEMA_reg_buffer_2641 ( .C (clk), .D (new_AGEMA_signal_3960), .Q (new_AGEMA_signal_5417) ) ;
    buf_clk new_AGEMA_reg_buffer_2643 ( .C (clk), .D (SubCellInst_SboxInst_15_n6), .Q (new_AGEMA_signal_5419) ) ;
    buf_clk new_AGEMA_reg_buffer_2645 ( .C (clk), .D (new_AGEMA_signal_1461), .Q (new_AGEMA_signal_5421) ) ;
    buf_clk new_AGEMA_reg_buffer_2647 ( .C (clk), .D (new_AGEMA_signal_1462), .Q (new_AGEMA_signal_5423) ) ;
    buf_clk new_AGEMA_reg_buffer_2653 ( .C (clk), .D (new_AGEMA_signal_5428), .Q (new_AGEMA_signal_5429) ) ;
    buf_clk new_AGEMA_reg_buffer_2661 ( .C (clk), .D (new_AGEMA_signal_5436), .Q (new_AGEMA_signal_5437) ) ;
    buf_clk new_AGEMA_reg_buffer_2669 ( .C (clk), .D (new_AGEMA_signal_5444), .Q (new_AGEMA_signal_5445) ) ;
    buf_clk new_AGEMA_reg_buffer_2677 ( .C (clk), .D (new_AGEMA_signal_5452), .Q (new_AGEMA_signal_5453) ) ;
    buf_clk new_AGEMA_reg_buffer_2685 ( .C (clk), .D (new_AGEMA_signal_5460), .Q (new_AGEMA_signal_5461) ) ;
    buf_clk new_AGEMA_reg_buffer_2693 ( .C (clk), .D (new_AGEMA_signal_5468), .Q (new_AGEMA_signal_5469) ) ;
    buf_clk new_AGEMA_reg_buffer_2701 ( .C (clk), .D (new_AGEMA_signal_5476), .Q (new_AGEMA_signal_5477) ) ;
    buf_clk new_AGEMA_reg_buffer_2709 ( .C (clk), .D (new_AGEMA_signal_5484), .Q (new_AGEMA_signal_5485) ) ;
    buf_clk new_AGEMA_reg_buffer_2717 ( .C (clk), .D (new_AGEMA_signal_5492), .Q (new_AGEMA_signal_5493) ) ;
    buf_clk new_AGEMA_reg_buffer_2725 ( .C (clk), .D (new_AGEMA_signal_5500), .Q (new_AGEMA_signal_5501) ) ;
    buf_clk new_AGEMA_reg_buffer_2733 ( .C (clk), .D (new_AGEMA_signal_5508), .Q (new_AGEMA_signal_5509) ) ;
    buf_clk new_AGEMA_reg_buffer_2741 ( .C (clk), .D (new_AGEMA_signal_5516), .Q (new_AGEMA_signal_5517) ) ;
    buf_clk new_AGEMA_reg_buffer_2749 ( .C (clk), .D (new_AGEMA_signal_5524), .Q (new_AGEMA_signal_5525) ) ;
    buf_clk new_AGEMA_reg_buffer_2757 ( .C (clk), .D (new_AGEMA_signal_5532), .Q (new_AGEMA_signal_5533) ) ;
    buf_clk new_AGEMA_reg_buffer_2765 ( .C (clk), .D (new_AGEMA_signal_5540), .Q (new_AGEMA_signal_5541) ) ;
    buf_clk new_AGEMA_reg_buffer_2773 ( .C (clk), .D (new_AGEMA_signal_5548), .Q (new_AGEMA_signal_5549) ) ;
    buf_clk new_AGEMA_reg_buffer_2781 ( .C (clk), .D (new_AGEMA_signal_5556), .Q (new_AGEMA_signal_5557) ) ;
    buf_clk new_AGEMA_reg_buffer_2789 ( .C (clk), .D (new_AGEMA_signal_5564), .Q (new_AGEMA_signal_5565) ) ;
    buf_clk new_AGEMA_reg_buffer_2797 ( .C (clk), .D (new_AGEMA_signal_5572), .Q (new_AGEMA_signal_5573) ) ;
    buf_clk new_AGEMA_reg_buffer_2805 ( .C (clk), .D (new_AGEMA_signal_5580), .Q (new_AGEMA_signal_5581) ) ;
    buf_clk new_AGEMA_reg_buffer_2813 ( .C (clk), .D (new_AGEMA_signal_5588), .Q (new_AGEMA_signal_5589) ) ;
    buf_clk new_AGEMA_reg_buffer_2821 ( .C (clk), .D (new_AGEMA_signal_5596), .Q (new_AGEMA_signal_5597) ) ;
    buf_clk new_AGEMA_reg_buffer_2829 ( .C (clk), .D (new_AGEMA_signal_5604), .Q (new_AGEMA_signal_5605) ) ;
    buf_clk new_AGEMA_reg_buffer_2837 ( .C (clk), .D (new_AGEMA_signal_5612), .Q (new_AGEMA_signal_5613) ) ;
    buf_clk new_AGEMA_reg_buffer_2845 ( .C (clk), .D (new_AGEMA_signal_5620), .Q (new_AGEMA_signal_5621) ) ;
    buf_clk new_AGEMA_reg_buffer_2853 ( .C (clk), .D (new_AGEMA_signal_5628), .Q (new_AGEMA_signal_5629) ) ;
    buf_clk new_AGEMA_reg_buffer_2861 ( .C (clk), .D (new_AGEMA_signal_5636), .Q (new_AGEMA_signal_5637) ) ;
    buf_clk new_AGEMA_reg_buffer_2869 ( .C (clk), .D (new_AGEMA_signal_5644), .Q (new_AGEMA_signal_5645) ) ;
    buf_clk new_AGEMA_reg_buffer_2877 ( .C (clk), .D (new_AGEMA_signal_5652), .Q (new_AGEMA_signal_5653) ) ;
    buf_clk new_AGEMA_reg_buffer_2885 ( .C (clk), .D (new_AGEMA_signal_5660), .Q (new_AGEMA_signal_5661) ) ;
    buf_clk new_AGEMA_reg_buffer_2893 ( .C (clk), .D (new_AGEMA_signal_5668), .Q (new_AGEMA_signal_5669) ) ;
    buf_clk new_AGEMA_reg_buffer_2901 ( .C (clk), .D (new_AGEMA_signal_5676), .Q (new_AGEMA_signal_5677) ) ;
    buf_clk new_AGEMA_reg_buffer_2909 ( .C (clk), .D (new_AGEMA_signal_5684), .Q (new_AGEMA_signal_5685) ) ;
    buf_clk new_AGEMA_reg_buffer_2917 ( .C (clk), .D (new_AGEMA_signal_5692), .Q (new_AGEMA_signal_5693) ) ;
    buf_clk new_AGEMA_reg_buffer_2925 ( .C (clk), .D (new_AGEMA_signal_5700), .Q (new_AGEMA_signal_5701) ) ;
    buf_clk new_AGEMA_reg_buffer_2933 ( .C (clk), .D (new_AGEMA_signal_5708), .Q (new_AGEMA_signal_5709) ) ;
    buf_clk new_AGEMA_reg_buffer_2941 ( .C (clk), .D (new_AGEMA_signal_5716), .Q (new_AGEMA_signal_5717) ) ;
    buf_clk new_AGEMA_reg_buffer_2949 ( .C (clk), .D (new_AGEMA_signal_5724), .Q (new_AGEMA_signal_5725) ) ;
    buf_clk new_AGEMA_reg_buffer_2957 ( .C (clk), .D (new_AGEMA_signal_5732), .Q (new_AGEMA_signal_5733) ) ;
    buf_clk new_AGEMA_reg_buffer_2965 ( .C (clk), .D (new_AGEMA_signal_5740), .Q (new_AGEMA_signal_5741) ) ;
    buf_clk new_AGEMA_reg_buffer_2973 ( .C (clk), .D (new_AGEMA_signal_5748), .Q (new_AGEMA_signal_5749) ) ;
    buf_clk new_AGEMA_reg_buffer_2981 ( .C (clk), .D (new_AGEMA_signal_5756), .Q (new_AGEMA_signal_5757) ) ;
    buf_clk new_AGEMA_reg_buffer_2989 ( .C (clk), .D (new_AGEMA_signal_5764), .Q (new_AGEMA_signal_5765) ) ;
    buf_clk new_AGEMA_reg_buffer_2997 ( .C (clk), .D (new_AGEMA_signal_5772), .Q (new_AGEMA_signal_5773) ) ;
    buf_clk new_AGEMA_reg_buffer_3005 ( .C (clk), .D (new_AGEMA_signal_5780), .Q (new_AGEMA_signal_5781) ) ;
    buf_clk new_AGEMA_reg_buffer_3013 ( .C (clk), .D (new_AGEMA_signal_5788), .Q (new_AGEMA_signal_5789) ) ;
    buf_clk new_AGEMA_reg_buffer_3021 ( .C (clk), .D (new_AGEMA_signal_5796), .Q (new_AGEMA_signal_5797) ) ;
    buf_clk new_AGEMA_reg_buffer_3029 ( .C (clk), .D (new_AGEMA_signal_5804), .Q (new_AGEMA_signal_5805) ) ;
    buf_clk new_AGEMA_reg_buffer_3037 ( .C (clk), .D (new_AGEMA_signal_5812), .Q (new_AGEMA_signal_5813) ) ;
    buf_clk new_AGEMA_reg_buffer_3045 ( .C (clk), .D (new_AGEMA_signal_5820), .Q (new_AGEMA_signal_5821) ) ;
    buf_clk new_AGEMA_reg_buffer_3053 ( .C (clk), .D (new_AGEMA_signal_5828), .Q (new_AGEMA_signal_5829) ) ;
    buf_clk new_AGEMA_reg_buffer_3061 ( .C (clk), .D (new_AGEMA_signal_5836), .Q (new_AGEMA_signal_5837) ) ;
    buf_clk new_AGEMA_reg_buffer_3069 ( .C (clk), .D (new_AGEMA_signal_5844), .Q (new_AGEMA_signal_5845) ) ;
    buf_clk new_AGEMA_reg_buffer_3077 ( .C (clk), .D (new_AGEMA_signal_5852), .Q (new_AGEMA_signal_5853) ) ;
    buf_clk new_AGEMA_reg_buffer_3085 ( .C (clk), .D (new_AGEMA_signal_5860), .Q (new_AGEMA_signal_5861) ) ;
    buf_clk new_AGEMA_reg_buffer_3093 ( .C (clk), .D (new_AGEMA_signal_5868), .Q (new_AGEMA_signal_5869) ) ;
    buf_clk new_AGEMA_reg_buffer_3101 ( .C (clk), .D (new_AGEMA_signal_5876), .Q (new_AGEMA_signal_5877) ) ;
    buf_clk new_AGEMA_reg_buffer_3109 ( .C (clk), .D (new_AGEMA_signal_5884), .Q (new_AGEMA_signal_5885) ) ;
    buf_clk new_AGEMA_reg_buffer_3117 ( .C (clk), .D (new_AGEMA_signal_5892), .Q (new_AGEMA_signal_5893) ) ;
    buf_clk new_AGEMA_reg_buffer_3125 ( .C (clk), .D (new_AGEMA_signal_5900), .Q (new_AGEMA_signal_5901) ) ;
    buf_clk new_AGEMA_reg_buffer_3133 ( .C (clk), .D (new_AGEMA_signal_5908), .Q (new_AGEMA_signal_5909) ) ;
    buf_clk new_AGEMA_reg_buffer_3141 ( .C (clk), .D (new_AGEMA_signal_5916), .Q (new_AGEMA_signal_5917) ) ;
    buf_clk new_AGEMA_reg_buffer_3149 ( .C (clk), .D (new_AGEMA_signal_5924), .Q (new_AGEMA_signal_5925) ) ;
    buf_clk new_AGEMA_reg_buffer_3157 ( .C (clk), .D (new_AGEMA_signal_5932), .Q (new_AGEMA_signal_5933) ) ;
    buf_clk new_AGEMA_reg_buffer_3165 ( .C (clk), .D (new_AGEMA_signal_5940), .Q (new_AGEMA_signal_5941) ) ;
    buf_clk new_AGEMA_reg_buffer_3173 ( .C (clk), .D (new_AGEMA_signal_5948), .Q (new_AGEMA_signal_5949) ) ;
    buf_clk new_AGEMA_reg_buffer_3181 ( .C (clk), .D (new_AGEMA_signal_5956), .Q (new_AGEMA_signal_5957) ) ;
    buf_clk new_AGEMA_reg_buffer_3189 ( .C (clk), .D (new_AGEMA_signal_5964), .Q (new_AGEMA_signal_5965) ) ;
    buf_clk new_AGEMA_reg_buffer_3197 ( .C (clk), .D (new_AGEMA_signal_5972), .Q (new_AGEMA_signal_5973) ) ;
    buf_clk new_AGEMA_reg_buffer_3205 ( .C (clk), .D (new_AGEMA_signal_5980), .Q (new_AGEMA_signal_5981) ) ;
    buf_clk new_AGEMA_reg_buffer_3213 ( .C (clk), .D (new_AGEMA_signal_5988), .Q (new_AGEMA_signal_5989) ) ;
    buf_clk new_AGEMA_reg_buffer_3221 ( .C (clk), .D (new_AGEMA_signal_5996), .Q (new_AGEMA_signal_5997) ) ;
    buf_clk new_AGEMA_reg_buffer_3229 ( .C (clk), .D (new_AGEMA_signal_6004), .Q (new_AGEMA_signal_6005) ) ;
    buf_clk new_AGEMA_reg_buffer_3237 ( .C (clk), .D (new_AGEMA_signal_6012), .Q (new_AGEMA_signal_6013) ) ;
    buf_clk new_AGEMA_reg_buffer_3245 ( .C (clk), .D (new_AGEMA_signal_6020), .Q (new_AGEMA_signal_6021) ) ;
    buf_clk new_AGEMA_reg_buffer_3253 ( .C (clk), .D (new_AGEMA_signal_6028), .Q (new_AGEMA_signal_6029) ) ;
    buf_clk new_AGEMA_reg_buffer_3261 ( .C (clk), .D (new_AGEMA_signal_6036), .Q (new_AGEMA_signal_6037) ) ;
    buf_clk new_AGEMA_reg_buffer_3269 ( .C (clk), .D (new_AGEMA_signal_6044), .Q (new_AGEMA_signal_6045) ) ;
    buf_clk new_AGEMA_reg_buffer_3277 ( .C (clk), .D (new_AGEMA_signal_6052), .Q (new_AGEMA_signal_6053) ) ;
    buf_clk new_AGEMA_reg_buffer_3285 ( .C (clk), .D (new_AGEMA_signal_6060), .Q (new_AGEMA_signal_6061) ) ;
    buf_clk new_AGEMA_reg_buffer_3293 ( .C (clk), .D (new_AGEMA_signal_6068), .Q (new_AGEMA_signal_6069) ) ;
    buf_clk new_AGEMA_reg_buffer_3301 ( .C (clk), .D (new_AGEMA_signal_6076), .Q (new_AGEMA_signal_6077) ) ;
    buf_clk new_AGEMA_reg_buffer_3309 ( .C (clk), .D (new_AGEMA_signal_6084), .Q (new_AGEMA_signal_6085) ) ;
    buf_clk new_AGEMA_reg_buffer_3317 ( .C (clk), .D (new_AGEMA_signal_6092), .Q (new_AGEMA_signal_6093) ) ;
    buf_clk new_AGEMA_reg_buffer_3325 ( .C (clk), .D (new_AGEMA_signal_6100), .Q (new_AGEMA_signal_6101) ) ;
    buf_clk new_AGEMA_reg_buffer_3333 ( .C (clk), .D (new_AGEMA_signal_6108), .Q (new_AGEMA_signal_6109) ) ;
    buf_clk new_AGEMA_reg_buffer_3341 ( .C (clk), .D (new_AGEMA_signal_6116), .Q (new_AGEMA_signal_6117) ) ;
    buf_clk new_AGEMA_reg_buffer_3349 ( .C (clk), .D (new_AGEMA_signal_6124), .Q (new_AGEMA_signal_6125) ) ;
    buf_clk new_AGEMA_reg_buffer_3357 ( .C (clk), .D (new_AGEMA_signal_6132), .Q (new_AGEMA_signal_6133) ) ;
    buf_clk new_AGEMA_reg_buffer_3365 ( .C (clk), .D (new_AGEMA_signal_6140), .Q (new_AGEMA_signal_6141) ) ;
    buf_clk new_AGEMA_reg_buffer_3373 ( .C (clk), .D (new_AGEMA_signal_6148), .Q (new_AGEMA_signal_6149) ) ;
    buf_clk new_AGEMA_reg_buffer_3381 ( .C (clk), .D (new_AGEMA_signal_6156), .Q (new_AGEMA_signal_6157) ) ;
    buf_clk new_AGEMA_reg_buffer_3389 ( .C (clk), .D (new_AGEMA_signal_6164), .Q (new_AGEMA_signal_6165) ) ;
    buf_clk new_AGEMA_reg_buffer_3397 ( .C (clk), .D (new_AGEMA_signal_6172), .Q (new_AGEMA_signal_6173) ) ;
    buf_clk new_AGEMA_reg_buffer_3405 ( .C (clk), .D (new_AGEMA_signal_6180), .Q (new_AGEMA_signal_6181) ) ;
    buf_clk new_AGEMA_reg_buffer_3413 ( .C (clk), .D (new_AGEMA_signal_6188), .Q (new_AGEMA_signal_6189) ) ;
    buf_clk new_AGEMA_reg_buffer_3421 ( .C (clk), .D (new_AGEMA_signal_6196), .Q (new_AGEMA_signal_6197) ) ;
    buf_clk new_AGEMA_reg_buffer_3429 ( .C (clk), .D (new_AGEMA_signal_6204), .Q (new_AGEMA_signal_6205) ) ;
    buf_clk new_AGEMA_reg_buffer_3437 ( .C (clk), .D (new_AGEMA_signal_6212), .Q (new_AGEMA_signal_6213) ) ;
    buf_clk new_AGEMA_reg_buffer_3445 ( .C (clk), .D (new_AGEMA_signal_6220), .Q (new_AGEMA_signal_6221) ) ;
    buf_clk new_AGEMA_reg_buffer_3453 ( .C (clk), .D (new_AGEMA_signal_6228), .Q (new_AGEMA_signal_6229) ) ;
    buf_clk new_AGEMA_reg_buffer_3461 ( .C (clk), .D (new_AGEMA_signal_6236), .Q (new_AGEMA_signal_6237) ) ;
    buf_clk new_AGEMA_reg_buffer_3469 ( .C (clk), .D (new_AGEMA_signal_6244), .Q (new_AGEMA_signal_6245) ) ;
    buf_clk new_AGEMA_reg_buffer_3477 ( .C (clk), .D (new_AGEMA_signal_6252), .Q (new_AGEMA_signal_6253) ) ;
    buf_clk new_AGEMA_reg_buffer_3485 ( .C (clk), .D (new_AGEMA_signal_6260), .Q (new_AGEMA_signal_6261) ) ;
    buf_clk new_AGEMA_reg_buffer_3493 ( .C (clk), .D (new_AGEMA_signal_6268), .Q (new_AGEMA_signal_6269) ) ;
    buf_clk new_AGEMA_reg_buffer_3501 ( .C (clk), .D (new_AGEMA_signal_6276), .Q (new_AGEMA_signal_6277) ) ;
    buf_clk new_AGEMA_reg_buffer_3509 ( .C (clk), .D (new_AGEMA_signal_6284), .Q (new_AGEMA_signal_6285) ) ;
    buf_clk new_AGEMA_reg_buffer_3517 ( .C (clk), .D (new_AGEMA_signal_6292), .Q (new_AGEMA_signal_6293) ) ;
    buf_clk new_AGEMA_reg_buffer_3525 ( .C (clk), .D (new_AGEMA_signal_6300), .Q (new_AGEMA_signal_6301) ) ;
    buf_clk new_AGEMA_reg_buffer_3533 ( .C (clk), .D (new_AGEMA_signal_6308), .Q (new_AGEMA_signal_6309) ) ;
    buf_clk new_AGEMA_reg_buffer_3541 ( .C (clk), .D (new_AGEMA_signal_6316), .Q (new_AGEMA_signal_6317) ) ;
    buf_clk new_AGEMA_reg_buffer_3549 ( .C (clk), .D (new_AGEMA_signal_6324), .Q (new_AGEMA_signal_6325) ) ;
    buf_clk new_AGEMA_reg_buffer_3557 ( .C (clk), .D (new_AGEMA_signal_6332), .Q (new_AGEMA_signal_6333) ) ;
    buf_clk new_AGEMA_reg_buffer_3565 ( .C (clk), .D (new_AGEMA_signal_6340), .Q (new_AGEMA_signal_6341) ) ;
    buf_clk new_AGEMA_reg_buffer_3573 ( .C (clk), .D (new_AGEMA_signal_6348), .Q (new_AGEMA_signal_6349) ) ;
    buf_clk new_AGEMA_reg_buffer_3581 ( .C (clk), .D (new_AGEMA_signal_6356), .Q (new_AGEMA_signal_6357) ) ;
    buf_clk new_AGEMA_reg_buffer_3589 ( .C (clk), .D (new_AGEMA_signal_6364), .Q (new_AGEMA_signal_6365) ) ;
    buf_clk new_AGEMA_reg_buffer_3597 ( .C (clk), .D (new_AGEMA_signal_6372), .Q (new_AGEMA_signal_6373) ) ;
    buf_clk new_AGEMA_reg_buffer_3605 ( .C (clk), .D (new_AGEMA_signal_6380), .Q (new_AGEMA_signal_6381) ) ;
    buf_clk new_AGEMA_reg_buffer_3613 ( .C (clk), .D (new_AGEMA_signal_6388), .Q (new_AGEMA_signal_6389) ) ;
    buf_clk new_AGEMA_reg_buffer_3621 ( .C (clk), .D (new_AGEMA_signal_6396), .Q (new_AGEMA_signal_6397) ) ;
    buf_clk new_AGEMA_reg_buffer_3629 ( .C (clk), .D (new_AGEMA_signal_6404), .Q (new_AGEMA_signal_6405) ) ;
    buf_clk new_AGEMA_reg_buffer_3637 ( .C (clk), .D (new_AGEMA_signal_6412), .Q (new_AGEMA_signal_6413) ) ;
    buf_clk new_AGEMA_reg_buffer_3645 ( .C (clk), .D (new_AGEMA_signal_6420), .Q (new_AGEMA_signal_6421) ) ;
    buf_clk new_AGEMA_reg_buffer_3653 ( .C (clk), .D (new_AGEMA_signal_6428), .Q (new_AGEMA_signal_6429) ) ;
    buf_clk new_AGEMA_reg_buffer_3661 ( .C (clk), .D (new_AGEMA_signal_6436), .Q (new_AGEMA_signal_6437) ) ;
    buf_clk new_AGEMA_reg_buffer_3669 ( .C (clk), .D (new_AGEMA_signal_6444), .Q (new_AGEMA_signal_6445) ) ;
    buf_clk new_AGEMA_reg_buffer_3677 ( .C (clk), .D (new_AGEMA_signal_6452), .Q (new_AGEMA_signal_6453) ) ;
    buf_clk new_AGEMA_reg_buffer_3685 ( .C (clk), .D (new_AGEMA_signal_6460), .Q (new_AGEMA_signal_6461) ) ;
    buf_clk new_AGEMA_reg_buffer_3693 ( .C (clk), .D (new_AGEMA_signal_6468), .Q (new_AGEMA_signal_6469) ) ;
    buf_clk new_AGEMA_reg_buffer_3701 ( .C (clk), .D (new_AGEMA_signal_6476), .Q (new_AGEMA_signal_6477) ) ;
    buf_clk new_AGEMA_reg_buffer_3709 ( .C (clk), .D (new_AGEMA_signal_6484), .Q (new_AGEMA_signal_6485) ) ;
    buf_clk new_AGEMA_reg_buffer_3717 ( .C (clk), .D (new_AGEMA_signal_6492), .Q (new_AGEMA_signal_6493) ) ;
    buf_clk new_AGEMA_reg_buffer_3725 ( .C (clk), .D (new_AGEMA_signal_6500), .Q (new_AGEMA_signal_6501) ) ;
    buf_clk new_AGEMA_reg_buffer_3733 ( .C (clk), .D (new_AGEMA_signal_6508), .Q (new_AGEMA_signal_6509) ) ;
    buf_clk new_AGEMA_reg_buffer_3741 ( .C (clk), .D (new_AGEMA_signal_6516), .Q (new_AGEMA_signal_6517) ) ;
    buf_clk new_AGEMA_reg_buffer_3749 ( .C (clk), .D (new_AGEMA_signal_6524), .Q (new_AGEMA_signal_6525) ) ;
    buf_clk new_AGEMA_reg_buffer_3757 ( .C (clk), .D (new_AGEMA_signal_6532), .Q (new_AGEMA_signal_6533) ) ;
    buf_clk new_AGEMA_reg_buffer_3765 ( .C (clk), .D (new_AGEMA_signal_6540), .Q (new_AGEMA_signal_6541) ) ;
    buf_clk new_AGEMA_reg_buffer_3773 ( .C (clk), .D (new_AGEMA_signal_6548), .Q (new_AGEMA_signal_6549) ) ;
    buf_clk new_AGEMA_reg_buffer_3781 ( .C (clk), .D (new_AGEMA_signal_6556), .Q (new_AGEMA_signal_6557) ) ;
    buf_clk new_AGEMA_reg_buffer_3789 ( .C (clk), .D (new_AGEMA_signal_6564), .Q (new_AGEMA_signal_6565) ) ;
    buf_clk new_AGEMA_reg_buffer_3797 ( .C (clk), .D (new_AGEMA_signal_6572), .Q (new_AGEMA_signal_6573) ) ;
    buf_clk new_AGEMA_reg_buffer_3805 ( .C (clk), .D (new_AGEMA_signal_6580), .Q (new_AGEMA_signal_6581) ) ;
    buf_clk new_AGEMA_reg_buffer_3813 ( .C (clk), .D (new_AGEMA_signal_6588), .Q (new_AGEMA_signal_6589) ) ;
    buf_clk new_AGEMA_reg_buffer_3821 ( .C (clk), .D (new_AGEMA_signal_6596), .Q (new_AGEMA_signal_6597) ) ;
    buf_clk new_AGEMA_reg_buffer_3829 ( .C (clk), .D (new_AGEMA_signal_6604), .Q (new_AGEMA_signal_6605) ) ;
    buf_clk new_AGEMA_reg_buffer_3837 ( .C (clk), .D (new_AGEMA_signal_6612), .Q (new_AGEMA_signal_6613) ) ;
    buf_clk new_AGEMA_reg_buffer_3845 ( .C (clk), .D (new_AGEMA_signal_6620), .Q (new_AGEMA_signal_6621) ) ;
    buf_clk new_AGEMA_reg_buffer_3853 ( .C (clk), .D (new_AGEMA_signal_6628), .Q (new_AGEMA_signal_6629) ) ;
    buf_clk new_AGEMA_reg_buffer_3861 ( .C (clk), .D (new_AGEMA_signal_6636), .Q (new_AGEMA_signal_6637) ) ;
    buf_clk new_AGEMA_reg_buffer_3869 ( .C (clk), .D (new_AGEMA_signal_6644), .Q (new_AGEMA_signal_6645) ) ;
    buf_clk new_AGEMA_reg_buffer_3877 ( .C (clk), .D (new_AGEMA_signal_6652), .Q (new_AGEMA_signal_6653) ) ;
    buf_clk new_AGEMA_reg_buffer_3885 ( .C (clk), .D (new_AGEMA_signal_6660), .Q (new_AGEMA_signal_6661) ) ;
    buf_clk new_AGEMA_reg_buffer_3893 ( .C (clk), .D (new_AGEMA_signal_6668), .Q (new_AGEMA_signal_6669) ) ;
    buf_clk new_AGEMA_reg_buffer_3901 ( .C (clk), .D (new_AGEMA_signal_6676), .Q (new_AGEMA_signal_6677) ) ;
    buf_clk new_AGEMA_reg_buffer_3909 ( .C (clk), .D (new_AGEMA_signal_6684), .Q (new_AGEMA_signal_6685) ) ;
    buf_clk new_AGEMA_reg_buffer_3917 ( .C (clk), .D (new_AGEMA_signal_6692), .Q (new_AGEMA_signal_6693) ) ;
    buf_clk new_AGEMA_reg_buffer_3925 ( .C (clk), .D (new_AGEMA_signal_6700), .Q (new_AGEMA_signal_6701) ) ;
    buf_clk new_AGEMA_reg_buffer_3933 ( .C (clk), .D (new_AGEMA_signal_6708), .Q (new_AGEMA_signal_6709) ) ;
    buf_clk new_AGEMA_reg_buffer_3941 ( .C (clk), .D (new_AGEMA_signal_6716), .Q (new_AGEMA_signal_6717) ) ;
    buf_clk new_AGEMA_reg_buffer_3949 ( .C (clk), .D (new_AGEMA_signal_6724), .Q (new_AGEMA_signal_6725) ) ;
    buf_clk new_AGEMA_reg_buffer_3957 ( .C (clk), .D (new_AGEMA_signal_6732), .Q (new_AGEMA_signal_6733) ) ;
    buf_clk new_AGEMA_reg_buffer_3965 ( .C (clk), .D (new_AGEMA_signal_6740), .Q (new_AGEMA_signal_6741) ) ;
    buf_clk new_AGEMA_reg_buffer_3973 ( .C (clk), .D (new_AGEMA_signal_6748), .Q (new_AGEMA_signal_6749) ) ;
    buf_clk new_AGEMA_reg_buffer_3981 ( .C (clk), .D (new_AGEMA_signal_6756), .Q (new_AGEMA_signal_6757) ) ;
    buf_clk new_AGEMA_reg_buffer_3989 ( .C (clk), .D (new_AGEMA_signal_6764), .Q (new_AGEMA_signal_6765) ) ;
    buf_clk new_AGEMA_reg_buffer_3997 ( .C (clk), .D (new_AGEMA_signal_6772), .Q (new_AGEMA_signal_6773) ) ;
    buf_clk new_AGEMA_reg_buffer_4005 ( .C (clk), .D (new_AGEMA_signal_6780), .Q (new_AGEMA_signal_6781) ) ;
    buf_clk new_AGEMA_reg_buffer_4013 ( .C (clk), .D (new_AGEMA_signal_6788), .Q (new_AGEMA_signal_6789) ) ;
    buf_clk new_AGEMA_reg_buffer_4021 ( .C (clk), .D (new_AGEMA_signal_6796), .Q (new_AGEMA_signal_6797) ) ;
    buf_clk new_AGEMA_reg_buffer_4029 ( .C (clk), .D (new_AGEMA_signal_6804), .Q (new_AGEMA_signal_6805) ) ;
    buf_clk new_AGEMA_reg_buffer_4037 ( .C (clk), .D (new_AGEMA_signal_6812), .Q (new_AGEMA_signal_6813) ) ;
    buf_clk new_AGEMA_reg_buffer_4045 ( .C (clk), .D (new_AGEMA_signal_6820), .Q (new_AGEMA_signal_6821) ) ;
    buf_clk new_AGEMA_reg_buffer_4053 ( .C (clk), .D (new_AGEMA_signal_6828), .Q (new_AGEMA_signal_6829) ) ;
    buf_clk new_AGEMA_reg_buffer_4061 ( .C (clk), .D (new_AGEMA_signal_6836), .Q (new_AGEMA_signal_6837) ) ;
    buf_clk new_AGEMA_reg_buffer_4069 ( .C (clk), .D (new_AGEMA_signal_6844), .Q (new_AGEMA_signal_6845) ) ;
    buf_clk new_AGEMA_reg_buffer_4077 ( .C (clk), .D (new_AGEMA_signal_6852), .Q (new_AGEMA_signal_6853) ) ;
    buf_clk new_AGEMA_reg_buffer_4085 ( .C (clk), .D (new_AGEMA_signal_6860), .Q (new_AGEMA_signal_6861) ) ;
    buf_clk new_AGEMA_reg_buffer_4093 ( .C (clk), .D (new_AGEMA_signal_6868), .Q (new_AGEMA_signal_6869) ) ;
    buf_clk new_AGEMA_reg_buffer_4101 ( .C (clk), .D (new_AGEMA_signal_6876), .Q (new_AGEMA_signal_6877) ) ;
    buf_clk new_AGEMA_reg_buffer_4109 ( .C (clk), .D (new_AGEMA_signal_6884), .Q (new_AGEMA_signal_6885) ) ;
    buf_clk new_AGEMA_reg_buffer_4117 ( .C (clk), .D (new_AGEMA_signal_6892), .Q (new_AGEMA_signal_6893) ) ;
    buf_clk new_AGEMA_reg_buffer_4125 ( .C (clk), .D (new_AGEMA_signal_6900), .Q (new_AGEMA_signal_6901) ) ;
    buf_clk new_AGEMA_reg_buffer_4133 ( .C (clk), .D (new_AGEMA_signal_6908), .Q (new_AGEMA_signal_6909) ) ;
    buf_clk new_AGEMA_reg_buffer_4141 ( .C (clk), .D (new_AGEMA_signal_6916), .Q (new_AGEMA_signal_6917) ) ;
    buf_clk new_AGEMA_reg_buffer_4149 ( .C (clk), .D (new_AGEMA_signal_6924), .Q (new_AGEMA_signal_6925) ) ;
    buf_clk new_AGEMA_reg_buffer_4157 ( .C (clk), .D (new_AGEMA_signal_6932), .Q (new_AGEMA_signal_6933) ) ;
    buf_clk new_AGEMA_reg_buffer_4165 ( .C (clk), .D (new_AGEMA_signal_6940), .Q (new_AGEMA_signal_6941) ) ;
    buf_clk new_AGEMA_reg_buffer_4173 ( .C (clk), .D (new_AGEMA_signal_6948), .Q (new_AGEMA_signal_6949) ) ;
    buf_clk new_AGEMA_reg_buffer_4181 ( .C (clk), .D (new_AGEMA_signal_6956), .Q (new_AGEMA_signal_6957) ) ;
    buf_clk new_AGEMA_reg_buffer_4193 ( .C (clk), .D (SubCellInst_SboxInst_0_n13), .Q (new_AGEMA_signal_6969) ) ;
    buf_clk new_AGEMA_reg_buffer_4197 ( .C (clk), .D (new_AGEMA_signal_1285), .Q (new_AGEMA_signal_6973) ) ;
    buf_clk new_AGEMA_reg_buffer_4201 ( .C (clk), .D (new_AGEMA_signal_1286), .Q (new_AGEMA_signal_6977) ) ;
    buf_clk new_AGEMA_reg_buffer_4211 ( .C (clk), .D (SubCellInst_SboxInst_1_n13), .Q (new_AGEMA_signal_6987) ) ;
    buf_clk new_AGEMA_reg_buffer_4215 ( .C (clk), .D (new_AGEMA_signal_1297), .Q (new_AGEMA_signal_6991) ) ;
    buf_clk new_AGEMA_reg_buffer_4219 ( .C (clk), .D (new_AGEMA_signal_1298), .Q (new_AGEMA_signal_6995) ) ;
    buf_clk new_AGEMA_reg_buffer_4229 ( .C (clk), .D (SubCellInst_SboxInst_2_n13), .Q (new_AGEMA_signal_7005) ) ;
    buf_clk new_AGEMA_reg_buffer_4233 ( .C (clk), .D (new_AGEMA_signal_1309), .Q (new_AGEMA_signal_7009) ) ;
    buf_clk new_AGEMA_reg_buffer_4237 ( .C (clk), .D (new_AGEMA_signal_1310), .Q (new_AGEMA_signal_7013) ) ;
    buf_clk new_AGEMA_reg_buffer_4247 ( .C (clk), .D (SubCellInst_SboxInst_3_n13), .Q (new_AGEMA_signal_7023) ) ;
    buf_clk new_AGEMA_reg_buffer_4251 ( .C (clk), .D (new_AGEMA_signal_1321), .Q (new_AGEMA_signal_7027) ) ;
    buf_clk new_AGEMA_reg_buffer_4255 ( .C (clk), .D (new_AGEMA_signal_1322), .Q (new_AGEMA_signal_7031) ) ;
    buf_clk new_AGEMA_reg_buffer_4265 ( .C (clk), .D (SubCellInst_SboxInst_4_n13), .Q (new_AGEMA_signal_7041) ) ;
    buf_clk new_AGEMA_reg_buffer_4269 ( .C (clk), .D (new_AGEMA_signal_1333), .Q (new_AGEMA_signal_7045) ) ;
    buf_clk new_AGEMA_reg_buffer_4273 ( .C (clk), .D (new_AGEMA_signal_1334), .Q (new_AGEMA_signal_7049) ) ;
    buf_clk new_AGEMA_reg_buffer_4283 ( .C (clk), .D (SubCellInst_SboxInst_5_n13), .Q (new_AGEMA_signal_7059) ) ;
    buf_clk new_AGEMA_reg_buffer_4287 ( .C (clk), .D (new_AGEMA_signal_1345), .Q (new_AGEMA_signal_7063) ) ;
    buf_clk new_AGEMA_reg_buffer_4291 ( .C (clk), .D (new_AGEMA_signal_1346), .Q (new_AGEMA_signal_7067) ) ;
    buf_clk new_AGEMA_reg_buffer_4301 ( .C (clk), .D (SubCellInst_SboxInst_6_n13), .Q (new_AGEMA_signal_7077) ) ;
    buf_clk new_AGEMA_reg_buffer_4305 ( .C (clk), .D (new_AGEMA_signal_1357), .Q (new_AGEMA_signal_7081) ) ;
    buf_clk new_AGEMA_reg_buffer_4309 ( .C (clk), .D (new_AGEMA_signal_1358), .Q (new_AGEMA_signal_7085) ) ;
    buf_clk new_AGEMA_reg_buffer_4319 ( .C (clk), .D (SubCellInst_SboxInst_7_n13), .Q (new_AGEMA_signal_7095) ) ;
    buf_clk new_AGEMA_reg_buffer_4323 ( .C (clk), .D (new_AGEMA_signal_1369), .Q (new_AGEMA_signal_7099) ) ;
    buf_clk new_AGEMA_reg_buffer_4327 ( .C (clk), .D (new_AGEMA_signal_1370), .Q (new_AGEMA_signal_7103) ) ;
    buf_clk new_AGEMA_reg_buffer_4337 ( .C (clk), .D (SubCellInst_SboxInst_8_n13), .Q (new_AGEMA_signal_7113) ) ;
    buf_clk new_AGEMA_reg_buffer_4341 ( .C (clk), .D (new_AGEMA_signal_1381), .Q (new_AGEMA_signal_7117) ) ;
    buf_clk new_AGEMA_reg_buffer_4345 ( .C (clk), .D (new_AGEMA_signal_1382), .Q (new_AGEMA_signal_7121) ) ;
    buf_clk new_AGEMA_reg_buffer_4355 ( .C (clk), .D (SubCellInst_SboxInst_9_n13), .Q (new_AGEMA_signal_7131) ) ;
    buf_clk new_AGEMA_reg_buffer_4359 ( .C (clk), .D (new_AGEMA_signal_1393), .Q (new_AGEMA_signal_7135) ) ;
    buf_clk new_AGEMA_reg_buffer_4363 ( .C (clk), .D (new_AGEMA_signal_1394), .Q (new_AGEMA_signal_7139) ) ;
    buf_clk new_AGEMA_reg_buffer_4373 ( .C (clk), .D (SubCellInst_SboxInst_10_n13), .Q (new_AGEMA_signal_7149) ) ;
    buf_clk new_AGEMA_reg_buffer_4377 ( .C (clk), .D (new_AGEMA_signal_1405), .Q (new_AGEMA_signal_7153) ) ;
    buf_clk new_AGEMA_reg_buffer_4381 ( .C (clk), .D (new_AGEMA_signal_1406), .Q (new_AGEMA_signal_7157) ) ;
    buf_clk new_AGEMA_reg_buffer_4391 ( .C (clk), .D (SubCellInst_SboxInst_11_n13), .Q (new_AGEMA_signal_7167) ) ;
    buf_clk new_AGEMA_reg_buffer_4395 ( .C (clk), .D (new_AGEMA_signal_1417), .Q (new_AGEMA_signal_7171) ) ;
    buf_clk new_AGEMA_reg_buffer_4399 ( .C (clk), .D (new_AGEMA_signal_1418), .Q (new_AGEMA_signal_7175) ) ;
    buf_clk new_AGEMA_reg_buffer_4409 ( .C (clk), .D (SubCellInst_SboxInst_12_n13), .Q (new_AGEMA_signal_7185) ) ;
    buf_clk new_AGEMA_reg_buffer_4413 ( .C (clk), .D (new_AGEMA_signal_1429), .Q (new_AGEMA_signal_7189) ) ;
    buf_clk new_AGEMA_reg_buffer_4417 ( .C (clk), .D (new_AGEMA_signal_1430), .Q (new_AGEMA_signal_7193) ) ;
    buf_clk new_AGEMA_reg_buffer_4427 ( .C (clk), .D (SubCellInst_SboxInst_13_n13), .Q (new_AGEMA_signal_7203) ) ;
    buf_clk new_AGEMA_reg_buffer_4431 ( .C (clk), .D (new_AGEMA_signal_1441), .Q (new_AGEMA_signal_7207) ) ;
    buf_clk new_AGEMA_reg_buffer_4435 ( .C (clk), .D (new_AGEMA_signal_1442), .Q (new_AGEMA_signal_7211) ) ;
    buf_clk new_AGEMA_reg_buffer_4445 ( .C (clk), .D (SubCellInst_SboxInst_14_n13), .Q (new_AGEMA_signal_7221) ) ;
    buf_clk new_AGEMA_reg_buffer_4449 ( .C (clk), .D (new_AGEMA_signal_1453), .Q (new_AGEMA_signal_7225) ) ;
    buf_clk new_AGEMA_reg_buffer_4453 ( .C (clk), .D (new_AGEMA_signal_1454), .Q (new_AGEMA_signal_7229) ) ;
    buf_clk new_AGEMA_reg_buffer_4463 ( .C (clk), .D (SubCellInst_SboxInst_15_n13), .Q (new_AGEMA_signal_7239) ) ;
    buf_clk new_AGEMA_reg_buffer_4467 ( .C (clk), .D (new_AGEMA_signal_1465), .Q (new_AGEMA_signal_7243) ) ;
    buf_clk new_AGEMA_reg_buffer_4471 ( .C (clk), .D (new_AGEMA_signal_1466), .Q (new_AGEMA_signal_7247) ) ;
    buf_clk new_AGEMA_reg_buffer_4669 ( .C (clk), .D (new_AGEMA_signal_7444), .Q (new_AGEMA_signal_7445) ) ;
    buf_clk new_AGEMA_reg_buffer_4677 ( .C (clk), .D (new_AGEMA_signal_7452), .Q (new_AGEMA_signal_7453) ) ;
    buf_clk new_AGEMA_reg_buffer_4685 ( .C (clk), .D (new_AGEMA_signal_7460), .Q (new_AGEMA_signal_7461) ) ;
    buf_clk new_AGEMA_reg_buffer_4693 ( .C (clk), .D (new_AGEMA_signal_7468), .Q (new_AGEMA_signal_7469) ) ;
    buf_clk new_AGEMA_reg_buffer_4701 ( .C (clk), .D (new_AGEMA_signal_7476), .Q (new_AGEMA_signal_7477) ) ;
    buf_clk new_AGEMA_reg_buffer_4709 ( .C (clk), .D (new_AGEMA_signal_7484), .Q (new_AGEMA_signal_7485) ) ;
    buf_clk new_AGEMA_reg_buffer_4717 ( .C (clk), .D (new_AGEMA_signal_7492), .Q (new_AGEMA_signal_7493) ) ;
    buf_clk new_AGEMA_reg_buffer_4725 ( .C (clk), .D (new_AGEMA_signal_7500), .Q (new_AGEMA_signal_7501) ) ;
    buf_clk new_AGEMA_reg_buffer_4733 ( .C (clk), .D (new_AGEMA_signal_7508), .Q (new_AGEMA_signal_7509) ) ;
    buf_clk new_AGEMA_reg_buffer_4741 ( .C (clk), .D (new_AGEMA_signal_7516), .Q (new_AGEMA_signal_7517) ) ;

    /* cells in depth 4 */
    or_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U18 ( .a ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, SubCellInst_SboxInst_0_n13}), .b ({new_AGEMA_signal_3600, new_AGEMA_signal_3598, new_AGEMA_signal_3596}), .clk (clk), .r ({Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_1566, new_AGEMA_signal_1565, SubCellInst_SboxInst_0_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U15 ( .a ({new_AGEMA_signal_1024, new_AGEMA_signal_1023, SubCellInst_SboxInst_0_n10}), .b ({new_AGEMA_signal_3606, new_AGEMA_signal_3604, new_AGEMA_signal_3602}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291]}), .c ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_0_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U11 ( .a ({new_AGEMA_signal_3612, new_AGEMA_signal_3610, new_AGEMA_signal_3608}), .b ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, SubCellInst_SboxInst_0_n4}), .clk (clk), .r ({Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_1570, new_AGEMA_signal_1569, SubCellInst_SboxInst_0_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U6 ( .a ({new_AGEMA_signal_3618, new_AGEMA_signal_3616, new_AGEMA_signal_3614}), .b ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, SubCellInst_SboxInst_0_n1}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297]}), .c ({new_AGEMA_signal_1284, new_AGEMA_signal_1283, SubCellInst_SboxInst_0_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U18 ( .a ({new_AGEMA_signal_1298, new_AGEMA_signal_1297, SubCellInst_SboxInst_1_n13}), .b ({new_AGEMA_signal_3624, new_AGEMA_signal_3622, new_AGEMA_signal_3620}), .clk (clk), .r ({Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_1576, new_AGEMA_signal_1575, SubCellInst_SboxInst_1_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U15 ( .a ({new_AGEMA_signal_1040, new_AGEMA_signal_1039, SubCellInst_SboxInst_1_n10}), .b ({new_AGEMA_signal_3630, new_AGEMA_signal_3628, new_AGEMA_signal_3626}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303]}), .c ({new_AGEMA_signal_1288, new_AGEMA_signal_1287, SubCellInst_SboxInst_1_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U11 ( .a ({new_AGEMA_signal_3636, new_AGEMA_signal_3634, new_AGEMA_signal_3632}), .b ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, SubCellInst_SboxInst_1_n4}), .clk (clk), .r ({Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_1580, new_AGEMA_signal_1579, SubCellInst_SboxInst_1_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U6 ( .a ({new_AGEMA_signal_3642, new_AGEMA_signal_3640, new_AGEMA_signal_3638}), .b ({new_AGEMA_signal_1044, new_AGEMA_signal_1043, SubCellInst_SboxInst_1_n1}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309]}), .c ({new_AGEMA_signal_1296, new_AGEMA_signal_1295, SubCellInst_SboxInst_1_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U18 ( .a ({new_AGEMA_signal_1310, new_AGEMA_signal_1309, SubCellInst_SboxInst_2_n13}), .b ({new_AGEMA_signal_3648, new_AGEMA_signal_3646, new_AGEMA_signal_3644}), .clk (clk), .r ({Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, SubCellInst_SboxInst_2_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U15 ( .a ({new_AGEMA_signal_1056, new_AGEMA_signal_1055, SubCellInst_SboxInst_2_n10}), .b ({new_AGEMA_signal_3654, new_AGEMA_signal_3652, new_AGEMA_signal_3650}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315]}), .c ({new_AGEMA_signal_1300, new_AGEMA_signal_1299, SubCellInst_SboxInst_2_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U11 ( .a ({new_AGEMA_signal_3660, new_AGEMA_signal_3658, new_AGEMA_signal_3656}), .b ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, SubCellInst_SboxInst_2_n4}), .clk (clk), .r ({Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_1590, new_AGEMA_signal_1589, SubCellInst_SboxInst_2_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U6 ( .a ({new_AGEMA_signal_3666, new_AGEMA_signal_3664, new_AGEMA_signal_3662}), .b ({new_AGEMA_signal_1060, new_AGEMA_signal_1059, SubCellInst_SboxInst_2_n1}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321]}), .c ({new_AGEMA_signal_1308, new_AGEMA_signal_1307, SubCellInst_SboxInst_2_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U18 ( .a ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, SubCellInst_SboxInst_3_n13}), .b ({new_AGEMA_signal_3672, new_AGEMA_signal_3670, new_AGEMA_signal_3668}), .clk (clk), .r ({Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_1596, new_AGEMA_signal_1595, SubCellInst_SboxInst_3_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U15 ( .a ({new_AGEMA_signal_1072, new_AGEMA_signal_1071, SubCellInst_SboxInst_3_n10}), .b ({new_AGEMA_signal_3678, new_AGEMA_signal_3676, new_AGEMA_signal_3674}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327]}), .c ({new_AGEMA_signal_1312, new_AGEMA_signal_1311, SubCellInst_SboxInst_3_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U11 ( .a ({new_AGEMA_signal_3684, new_AGEMA_signal_3682, new_AGEMA_signal_3680}), .b ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, SubCellInst_SboxInst_3_n4}), .clk (clk), .r ({Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_1600, new_AGEMA_signal_1599, SubCellInst_SboxInst_3_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U6 ( .a ({new_AGEMA_signal_3690, new_AGEMA_signal_3688, new_AGEMA_signal_3686}), .b ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, SubCellInst_SboxInst_3_n1}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333]}), .c ({new_AGEMA_signal_1320, new_AGEMA_signal_1319, SubCellInst_SboxInst_3_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U18 ( .a ({new_AGEMA_signal_1334, new_AGEMA_signal_1333, SubCellInst_SboxInst_4_n13}), .b ({new_AGEMA_signal_3696, new_AGEMA_signal_3694, new_AGEMA_signal_3692}), .clk (clk), .r ({Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_1606, new_AGEMA_signal_1605, SubCellInst_SboxInst_4_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U15 ( .a ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, SubCellInst_SboxInst_4_n10}), .b ({new_AGEMA_signal_3702, new_AGEMA_signal_3700, new_AGEMA_signal_3698}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339]}), .c ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, SubCellInst_SboxInst_4_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U11 ( .a ({new_AGEMA_signal_3708, new_AGEMA_signal_3706, new_AGEMA_signal_3704}), .b ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, SubCellInst_SboxInst_4_n4}), .clk (clk), .r ({Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_1610, new_AGEMA_signal_1609, SubCellInst_SboxInst_4_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U6 ( .a ({new_AGEMA_signal_3714, new_AGEMA_signal_3712, new_AGEMA_signal_3710}), .b ({new_AGEMA_signal_1092, new_AGEMA_signal_1091, SubCellInst_SboxInst_4_n1}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345]}), .c ({new_AGEMA_signal_1332, new_AGEMA_signal_1331, SubCellInst_SboxInst_4_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U18 ( .a ({new_AGEMA_signal_1346, new_AGEMA_signal_1345, SubCellInst_SboxInst_5_n13}), .b ({new_AGEMA_signal_3720, new_AGEMA_signal_3718, new_AGEMA_signal_3716}), .clk (clk), .r ({Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_1616, new_AGEMA_signal_1615, SubCellInst_SboxInst_5_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U15 ( .a ({new_AGEMA_signal_1104, new_AGEMA_signal_1103, SubCellInst_SboxInst_5_n10}), .b ({new_AGEMA_signal_3726, new_AGEMA_signal_3724, new_AGEMA_signal_3722}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351]}), .c ({new_AGEMA_signal_1336, new_AGEMA_signal_1335, SubCellInst_SboxInst_5_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U11 ( .a ({new_AGEMA_signal_3732, new_AGEMA_signal_3730, new_AGEMA_signal_3728}), .b ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, SubCellInst_SboxInst_5_n4}), .clk (clk), .r ({Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_1620, new_AGEMA_signal_1619, SubCellInst_SboxInst_5_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U6 ( .a ({new_AGEMA_signal_3738, new_AGEMA_signal_3736, new_AGEMA_signal_3734}), .b ({new_AGEMA_signal_1108, new_AGEMA_signal_1107, SubCellInst_SboxInst_5_n1}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357]}), .c ({new_AGEMA_signal_1344, new_AGEMA_signal_1343, SubCellInst_SboxInst_5_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U18 ( .a ({new_AGEMA_signal_1358, new_AGEMA_signal_1357, SubCellInst_SboxInst_6_n13}), .b ({new_AGEMA_signal_3744, new_AGEMA_signal_3742, new_AGEMA_signal_3740}), .clk (clk), .r ({Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_1626, new_AGEMA_signal_1625, SubCellInst_SboxInst_6_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U15 ( .a ({new_AGEMA_signal_1120, new_AGEMA_signal_1119, SubCellInst_SboxInst_6_n10}), .b ({new_AGEMA_signal_3750, new_AGEMA_signal_3748, new_AGEMA_signal_3746}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363]}), .c ({new_AGEMA_signal_1348, new_AGEMA_signal_1347, SubCellInst_SboxInst_6_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U11 ( .a ({new_AGEMA_signal_3756, new_AGEMA_signal_3754, new_AGEMA_signal_3752}), .b ({new_AGEMA_signal_1352, new_AGEMA_signal_1351, SubCellInst_SboxInst_6_n4}), .clk (clk), .r ({Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_1630, new_AGEMA_signal_1629, SubCellInst_SboxInst_6_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U6 ( .a ({new_AGEMA_signal_3762, new_AGEMA_signal_3760, new_AGEMA_signal_3758}), .b ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, SubCellInst_SboxInst_6_n1}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369]}), .c ({new_AGEMA_signal_1356, new_AGEMA_signal_1355, SubCellInst_SboxInst_6_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U18 ( .a ({new_AGEMA_signal_1370, new_AGEMA_signal_1369, SubCellInst_SboxInst_7_n13}), .b ({new_AGEMA_signal_3768, new_AGEMA_signal_3766, new_AGEMA_signal_3764}), .clk (clk), .r ({Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_1636, new_AGEMA_signal_1635, SubCellInst_SboxInst_7_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U15 ( .a ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, SubCellInst_SboxInst_7_n10}), .b ({new_AGEMA_signal_3774, new_AGEMA_signal_3772, new_AGEMA_signal_3770}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375]}), .c ({new_AGEMA_signal_1360, new_AGEMA_signal_1359, SubCellInst_SboxInst_7_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U11 ( .a ({new_AGEMA_signal_3780, new_AGEMA_signal_3778, new_AGEMA_signal_3776}), .b ({new_AGEMA_signal_1364, new_AGEMA_signal_1363, SubCellInst_SboxInst_7_n4}), .clk (clk), .r ({Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_1640, new_AGEMA_signal_1639, SubCellInst_SboxInst_7_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U6 ( .a ({new_AGEMA_signal_3786, new_AGEMA_signal_3784, new_AGEMA_signal_3782}), .b ({new_AGEMA_signal_1140, new_AGEMA_signal_1139, SubCellInst_SboxInst_7_n1}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381]}), .c ({new_AGEMA_signal_1368, new_AGEMA_signal_1367, SubCellInst_SboxInst_7_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U18 ( .a ({new_AGEMA_signal_1382, new_AGEMA_signal_1381, SubCellInst_SboxInst_8_n13}), .b ({new_AGEMA_signal_3792, new_AGEMA_signal_3790, new_AGEMA_signal_3788}), .clk (clk), .r ({Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_1646, new_AGEMA_signal_1645, SubCellInst_SboxInst_8_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U15 ( .a ({new_AGEMA_signal_1152, new_AGEMA_signal_1151, SubCellInst_SboxInst_8_n10}), .b ({new_AGEMA_signal_3798, new_AGEMA_signal_3796, new_AGEMA_signal_3794}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387]}), .c ({new_AGEMA_signal_1372, new_AGEMA_signal_1371, SubCellInst_SboxInst_8_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U11 ( .a ({new_AGEMA_signal_3804, new_AGEMA_signal_3802, new_AGEMA_signal_3800}), .b ({new_AGEMA_signal_1376, new_AGEMA_signal_1375, SubCellInst_SboxInst_8_n4}), .clk (clk), .r ({Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_1650, new_AGEMA_signal_1649, SubCellInst_SboxInst_8_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U6 ( .a ({new_AGEMA_signal_3810, new_AGEMA_signal_3808, new_AGEMA_signal_3806}), .b ({new_AGEMA_signal_1156, new_AGEMA_signal_1155, SubCellInst_SboxInst_8_n1}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393]}), .c ({new_AGEMA_signal_1380, new_AGEMA_signal_1379, SubCellInst_SboxInst_8_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U18 ( .a ({new_AGEMA_signal_1394, new_AGEMA_signal_1393, SubCellInst_SboxInst_9_n13}), .b ({new_AGEMA_signal_3816, new_AGEMA_signal_3814, new_AGEMA_signal_3812}), .clk (clk), .r ({Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_1656, new_AGEMA_signal_1655, SubCellInst_SboxInst_9_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U15 ( .a ({new_AGEMA_signal_1168, new_AGEMA_signal_1167, SubCellInst_SboxInst_9_n10}), .b ({new_AGEMA_signal_3822, new_AGEMA_signal_3820, new_AGEMA_signal_3818}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399]}), .c ({new_AGEMA_signal_1384, new_AGEMA_signal_1383, SubCellInst_SboxInst_9_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U11 ( .a ({new_AGEMA_signal_3828, new_AGEMA_signal_3826, new_AGEMA_signal_3824}), .b ({new_AGEMA_signal_1388, new_AGEMA_signal_1387, SubCellInst_SboxInst_9_n4}), .clk (clk), .r ({Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_1660, new_AGEMA_signal_1659, SubCellInst_SboxInst_9_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U6 ( .a ({new_AGEMA_signal_3834, new_AGEMA_signal_3832, new_AGEMA_signal_3830}), .b ({new_AGEMA_signal_1172, new_AGEMA_signal_1171, SubCellInst_SboxInst_9_n1}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405]}), .c ({new_AGEMA_signal_1392, new_AGEMA_signal_1391, SubCellInst_SboxInst_9_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U18 ( .a ({new_AGEMA_signal_1406, new_AGEMA_signal_1405, SubCellInst_SboxInst_10_n13}), .b ({new_AGEMA_signal_3840, new_AGEMA_signal_3838, new_AGEMA_signal_3836}), .clk (clk), .r ({Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_1666, new_AGEMA_signal_1665, SubCellInst_SboxInst_10_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U15 ( .a ({new_AGEMA_signal_1184, new_AGEMA_signal_1183, SubCellInst_SboxInst_10_n10}), .b ({new_AGEMA_signal_3846, new_AGEMA_signal_3844, new_AGEMA_signal_3842}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411]}), .c ({new_AGEMA_signal_1396, new_AGEMA_signal_1395, SubCellInst_SboxInst_10_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U11 ( .a ({new_AGEMA_signal_3852, new_AGEMA_signal_3850, new_AGEMA_signal_3848}), .b ({new_AGEMA_signal_1400, new_AGEMA_signal_1399, SubCellInst_SboxInst_10_n4}), .clk (clk), .r ({Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_1670, new_AGEMA_signal_1669, SubCellInst_SboxInst_10_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U6 ( .a ({new_AGEMA_signal_3858, new_AGEMA_signal_3856, new_AGEMA_signal_3854}), .b ({new_AGEMA_signal_1188, new_AGEMA_signal_1187, SubCellInst_SboxInst_10_n1}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417]}), .c ({new_AGEMA_signal_1404, new_AGEMA_signal_1403, SubCellInst_SboxInst_10_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U18 ( .a ({new_AGEMA_signal_1418, new_AGEMA_signal_1417, SubCellInst_SboxInst_11_n13}), .b ({new_AGEMA_signal_3864, new_AGEMA_signal_3862, new_AGEMA_signal_3860}), .clk (clk), .r ({Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, SubCellInst_SboxInst_11_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U15 ( .a ({new_AGEMA_signal_1200, new_AGEMA_signal_1199, SubCellInst_SboxInst_11_n10}), .b ({new_AGEMA_signal_3870, new_AGEMA_signal_3868, new_AGEMA_signal_3866}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423]}), .c ({new_AGEMA_signal_1408, new_AGEMA_signal_1407, SubCellInst_SboxInst_11_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U11 ( .a ({new_AGEMA_signal_3876, new_AGEMA_signal_3874, new_AGEMA_signal_3872}), .b ({new_AGEMA_signal_1412, new_AGEMA_signal_1411, SubCellInst_SboxInst_11_n4}), .clk (clk), .r ({Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_1680, new_AGEMA_signal_1679, SubCellInst_SboxInst_11_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U6 ( .a ({new_AGEMA_signal_3882, new_AGEMA_signal_3880, new_AGEMA_signal_3878}), .b ({new_AGEMA_signal_1204, new_AGEMA_signal_1203, SubCellInst_SboxInst_11_n1}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429]}), .c ({new_AGEMA_signal_1416, new_AGEMA_signal_1415, SubCellInst_SboxInst_11_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U18 ( .a ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, SubCellInst_SboxInst_12_n13}), .b ({new_AGEMA_signal_3888, new_AGEMA_signal_3886, new_AGEMA_signal_3884}), .clk (clk), .r ({Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_1686, new_AGEMA_signal_1685, SubCellInst_SboxInst_12_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U15 ( .a ({new_AGEMA_signal_1216, new_AGEMA_signal_1215, SubCellInst_SboxInst_12_n10}), .b ({new_AGEMA_signal_3894, new_AGEMA_signal_3892, new_AGEMA_signal_3890}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435]}), .c ({new_AGEMA_signal_1420, new_AGEMA_signal_1419, SubCellInst_SboxInst_12_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U11 ( .a ({new_AGEMA_signal_3900, new_AGEMA_signal_3898, new_AGEMA_signal_3896}), .b ({new_AGEMA_signal_1424, new_AGEMA_signal_1423, SubCellInst_SboxInst_12_n4}), .clk (clk), .r ({Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_1690, new_AGEMA_signal_1689, SubCellInst_SboxInst_12_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U6 ( .a ({new_AGEMA_signal_3906, new_AGEMA_signal_3904, new_AGEMA_signal_3902}), .b ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, SubCellInst_SboxInst_12_n1}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441]}), .c ({new_AGEMA_signal_1428, new_AGEMA_signal_1427, SubCellInst_SboxInst_12_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U18 ( .a ({new_AGEMA_signal_1442, new_AGEMA_signal_1441, SubCellInst_SboxInst_13_n13}), .b ({new_AGEMA_signal_3912, new_AGEMA_signal_3910, new_AGEMA_signal_3908}), .clk (clk), .r ({Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_1696, new_AGEMA_signal_1695, SubCellInst_SboxInst_13_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U15 ( .a ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, SubCellInst_SboxInst_13_n10}), .b ({new_AGEMA_signal_3918, new_AGEMA_signal_3916, new_AGEMA_signal_3914}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447]}), .c ({new_AGEMA_signal_1432, new_AGEMA_signal_1431, SubCellInst_SboxInst_13_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U11 ( .a ({new_AGEMA_signal_3924, new_AGEMA_signal_3922, new_AGEMA_signal_3920}), .b ({new_AGEMA_signal_1436, new_AGEMA_signal_1435, SubCellInst_SboxInst_13_n4}), .clk (clk), .r ({Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_1700, new_AGEMA_signal_1699, SubCellInst_SboxInst_13_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U6 ( .a ({new_AGEMA_signal_3930, new_AGEMA_signal_3928, new_AGEMA_signal_3926}), .b ({new_AGEMA_signal_1236, new_AGEMA_signal_1235, SubCellInst_SboxInst_13_n1}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453]}), .c ({new_AGEMA_signal_1440, new_AGEMA_signal_1439, SubCellInst_SboxInst_13_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U18 ( .a ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, SubCellInst_SboxInst_14_n13}), .b ({new_AGEMA_signal_3936, new_AGEMA_signal_3934, new_AGEMA_signal_3932}), .clk (clk), .r ({Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, SubCellInst_SboxInst_14_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U15 ( .a ({new_AGEMA_signal_1248, new_AGEMA_signal_1247, SubCellInst_SboxInst_14_n10}), .b ({new_AGEMA_signal_3942, new_AGEMA_signal_3940, new_AGEMA_signal_3938}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459]}), .c ({new_AGEMA_signal_1444, new_AGEMA_signal_1443, SubCellInst_SboxInst_14_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U11 ( .a ({new_AGEMA_signal_3948, new_AGEMA_signal_3946, new_AGEMA_signal_3944}), .b ({new_AGEMA_signal_1448, new_AGEMA_signal_1447, SubCellInst_SboxInst_14_n4}), .clk (clk), .r ({Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_1710, new_AGEMA_signal_1709, SubCellInst_SboxInst_14_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U6 ( .a ({new_AGEMA_signal_3954, new_AGEMA_signal_3952, new_AGEMA_signal_3950}), .b ({new_AGEMA_signal_1252, new_AGEMA_signal_1251, SubCellInst_SboxInst_14_n1}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465]}), .c ({new_AGEMA_signal_1452, new_AGEMA_signal_1451, SubCellInst_SboxInst_14_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U18 ( .a ({new_AGEMA_signal_1466, new_AGEMA_signal_1465, SubCellInst_SboxInst_15_n13}), .b ({new_AGEMA_signal_3960, new_AGEMA_signal_3958, new_AGEMA_signal_3956}), .clk (clk), .r ({Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_1716, new_AGEMA_signal_1715, SubCellInst_SboxInst_15_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U15 ( .a ({new_AGEMA_signal_1264, new_AGEMA_signal_1263, SubCellInst_SboxInst_15_n10}), .b ({new_AGEMA_signal_3966, new_AGEMA_signal_3964, new_AGEMA_signal_3962}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471]}), .c ({new_AGEMA_signal_1456, new_AGEMA_signal_1455, SubCellInst_SboxInst_15_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U11 ( .a ({new_AGEMA_signal_3972, new_AGEMA_signal_3970, new_AGEMA_signal_3968}), .b ({new_AGEMA_signal_1460, new_AGEMA_signal_1459, SubCellInst_SboxInst_15_n4}), .clk (clk), .r ({Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_1720, new_AGEMA_signal_1719, SubCellInst_SboxInst_15_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U6 ( .a ({new_AGEMA_signal_3978, new_AGEMA_signal_3976, new_AGEMA_signal_3974}), .b ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, SubCellInst_SboxInst_15_n1}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477]}), .c ({new_AGEMA_signal_1464, new_AGEMA_signal_1463, SubCellInst_SboxInst_15_n2}) ) ;
    buf_clk new_AGEMA_reg_buffer_1206 ( .C (clk), .D (new_AGEMA_signal_3981), .Q (new_AGEMA_signal_3982) ) ;
    buf_clk new_AGEMA_reg_buffer_1212 ( .C (clk), .D (new_AGEMA_signal_3987), .Q (new_AGEMA_signal_3988) ) ;
    buf_clk new_AGEMA_reg_buffer_1218 ( .C (clk), .D (new_AGEMA_signal_3993), .Q (new_AGEMA_signal_3994) ) ;
    buf_clk new_AGEMA_reg_buffer_1224 ( .C (clk), .D (new_AGEMA_signal_3999), .Q (new_AGEMA_signal_4000) ) ;
    buf_clk new_AGEMA_reg_buffer_1230 ( .C (clk), .D (new_AGEMA_signal_4005), .Q (new_AGEMA_signal_4006) ) ;
    buf_clk new_AGEMA_reg_buffer_1236 ( .C (clk), .D (new_AGEMA_signal_4011), .Q (new_AGEMA_signal_4012) ) ;
    buf_clk new_AGEMA_reg_buffer_1242 ( .C (clk), .D (new_AGEMA_signal_4017), .Q (new_AGEMA_signal_4018) ) ;
    buf_clk new_AGEMA_reg_buffer_1248 ( .C (clk), .D (new_AGEMA_signal_4023), .Q (new_AGEMA_signal_4024) ) ;
    buf_clk new_AGEMA_reg_buffer_1254 ( .C (clk), .D (new_AGEMA_signal_4029), .Q (new_AGEMA_signal_4030) ) ;
    buf_clk new_AGEMA_reg_buffer_1260 ( .C (clk), .D (new_AGEMA_signal_4035), .Q (new_AGEMA_signal_4036) ) ;
    buf_clk new_AGEMA_reg_buffer_1266 ( .C (clk), .D (new_AGEMA_signal_4041), .Q (new_AGEMA_signal_4042) ) ;
    buf_clk new_AGEMA_reg_buffer_1272 ( .C (clk), .D (new_AGEMA_signal_4047), .Q (new_AGEMA_signal_4048) ) ;
    buf_clk new_AGEMA_reg_buffer_1278 ( .C (clk), .D (new_AGEMA_signal_4053), .Q (new_AGEMA_signal_4054) ) ;
    buf_clk new_AGEMA_reg_buffer_1284 ( .C (clk), .D (new_AGEMA_signal_4059), .Q (new_AGEMA_signal_4060) ) ;
    buf_clk new_AGEMA_reg_buffer_1290 ( .C (clk), .D (new_AGEMA_signal_4065), .Q (new_AGEMA_signal_4066) ) ;
    buf_clk new_AGEMA_reg_buffer_1296 ( .C (clk), .D (new_AGEMA_signal_4071), .Q (new_AGEMA_signal_4072) ) ;
    buf_clk new_AGEMA_reg_buffer_1302 ( .C (clk), .D (new_AGEMA_signal_4077), .Q (new_AGEMA_signal_4078) ) ;
    buf_clk new_AGEMA_reg_buffer_1308 ( .C (clk), .D (new_AGEMA_signal_4083), .Q (new_AGEMA_signal_4084) ) ;
    buf_clk new_AGEMA_reg_buffer_1314 ( .C (clk), .D (new_AGEMA_signal_4089), .Q (new_AGEMA_signal_4090) ) ;
    buf_clk new_AGEMA_reg_buffer_1320 ( .C (clk), .D (new_AGEMA_signal_4095), .Q (new_AGEMA_signal_4096) ) ;
    buf_clk new_AGEMA_reg_buffer_1326 ( .C (clk), .D (new_AGEMA_signal_4101), .Q (new_AGEMA_signal_4102) ) ;
    buf_clk new_AGEMA_reg_buffer_1332 ( .C (clk), .D (new_AGEMA_signal_4107), .Q (new_AGEMA_signal_4108) ) ;
    buf_clk new_AGEMA_reg_buffer_1338 ( .C (clk), .D (new_AGEMA_signal_4113), .Q (new_AGEMA_signal_4114) ) ;
    buf_clk new_AGEMA_reg_buffer_1344 ( .C (clk), .D (new_AGEMA_signal_4119), .Q (new_AGEMA_signal_4120) ) ;
    buf_clk new_AGEMA_reg_buffer_1350 ( .C (clk), .D (new_AGEMA_signal_4125), .Q (new_AGEMA_signal_4126) ) ;
    buf_clk new_AGEMA_reg_buffer_1356 ( .C (clk), .D (new_AGEMA_signal_4131), .Q (new_AGEMA_signal_4132) ) ;
    buf_clk new_AGEMA_reg_buffer_1362 ( .C (clk), .D (new_AGEMA_signal_4137), .Q (new_AGEMA_signal_4138) ) ;
    buf_clk new_AGEMA_reg_buffer_1368 ( .C (clk), .D (new_AGEMA_signal_4143), .Q (new_AGEMA_signal_4144) ) ;
    buf_clk new_AGEMA_reg_buffer_1374 ( .C (clk), .D (new_AGEMA_signal_4149), .Q (new_AGEMA_signal_4150) ) ;
    buf_clk new_AGEMA_reg_buffer_1380 ( .C (clk), .D (new_AGEMA_signal_4155), .Q (new_AGEMA_signal_4156) ) ;
    buf_clk new_AGEMA_reg_buffer_1386 ( .C (clk), .D (new_AGEMA_signal_4161), .Q (new_AGEMA_signal_4162) ) ;
    buf_clk new_AGEMA_reg_buffer_1392 ( .C (clk), .D (new_AGEMA_signal_4167), .Q (new_AGEMA_signal_4168) ) ;
    buf_clk new_AGEMA_reg_buffer_1398 ( .C (clk), .D (new_AGEMA_signal_4173), .Q (new_AGEMA_signal_4174) ) ;
    buf_clk new_AGEMA_reg_buffer_1404 ( .C (clk), .D (new_AGEMA_signal_4179), .Q (new_AGEMA_signal_4180) ) ;
    buf_clk new_AGEMA_reg_buffer_1410 ( .C (clk), .D (new_AGEMA_signal_4185), .Q (new_AGEMA_signal_4186) ) ;
    buf_clk new_AGEMA_reg_buffer_1416 ( .C (clk), .D (new_AGEMA_signal_4191), .Q (new_AGEMA_signal_4192) ) ;
    buf_clk new_AGEMA_reg_buffer_1422 ( .C (clk), .D (new_AGEMA_signal_4197), .Q (new_AGEMA_signal_4198) ) ;
    buf_clk new_AGEMA_reg_buffer_1428 ( .C (clk), .D (new_AGEMA_signal_4203), .Q (new_AGEMA_signal_4204) ) ;
    buf_clk new_AGEMA_reg_buffer_1434 ( .C (clk), .D (new_AGEMA_signal_4209), .Q (new_AGEMA_signal_4210) ) ;
    buf_clk new_AGEMA_reg_buffer_1440 ( .C (clk), .D (new_AGEMA_signal_4215), .Q (new_AGEMA_signal_4216) ) ;
    buf_clk new_AGEMA_reg_buffer_1446 ( .C (clk), .D (new_AGEMA_signal_4221), .Q (new_AGEMA_signal_4222) ) ;
    buf_clk new_AGEMA_reg_buffer_1452 ( .C (clk), .D (new_AGEMA_signal_4227), .Q (new_AGEMA_signal_4228) ) ;
    buf_clk new_AGEMA_reg_buffer_1458 ( .C (clk), .D (new_AGEMA_signal_4233), .Q (new_AGEMA_signal_4234) ) ;
    buf_clk new_AGEMA_reg_buffer_1464 ( .C (clk), .D (new_AGEMA_signal_4239), .Q (new_AGEMA_signal_4240) ) ;
    buf_clk new_AGEMA_reg_buffer_1470 ( .C (clk), .D (new_AGEMA_signal_4245), .Q (new_AGEMA_signal_4246) ) ;
    buf_clk new_AGEMA_reg_buffer_1476 ( .C (clk), .D (new_AGEMA_signal_4251), .Q (new_AGEMA_signal_4252) ) ;
    buf_clk new_AGEMA_reg_buffer_1482 ( .C (clk), .D (new_AGEMA_signal_4257), .Q (new_AGEMA_signal_4258) ) ;
    buf_clk new_AGEMA_reg_buffer_1488 ( .C (clk), .D (new_AGEMA_signal_4263), .Q (new_AGEMA_signal_4264) ) ;
    buf_clk new_AGEMA_reg_buffer_1494 ( .C (clk), .D (new_AGEMA_signal_4269), .Q (new_AGEMA_signal_4270) ) ;
    buf_clk new_AGEMA_reg_buffer_1500 ( .C (clk), .D (new_AGEMA_signal_4275), .Q (new_AGEMA_signal_4276) ) ;
    buf_clk new_AGEMA_reg_buffer_1506 ( .C (clk), .D (new_AGEMA_signal_4281), .Q (new_AGEMA_signal_4282) ) ;
    buf_clk new_AGEMA_reg_buffer_1512 ( .C (clk), .D (new_AGEMA_signal_4287), .Q (new_AGEMA_signal_4288) ) ;
    buf_clk new_AGEMA_reg_buffer_1518 ( .C (clk), .D (new_AGEMA_signal_4293), .Q (new_AGEMA_signal_4294) ) ;
    buf_clk new_AGEMA_reg_buffer_1524 ( .C (clk), .D (new_AGEMA_signal_4299), .Q (new_AGEMA_signal_4300) ) ;
    buf_clk new_AGEMA_reg_buffer_1530 ( .C (clk), .D (new_AGEMA_signal_4305), .Q (new_AGEMA_signal_4306) ) ;
    buf_clk new_AGEMA_reg_buffer_1536 ( .C (clk), .D (new_AGEMA_signal_4311), .Q (new_AGEMA_signal_4312) ) ;
    buf_clk new_AGEMA_reg_buffer_1542 ( .C (clk), .D (new_AGEMA_signal_4317), .Q (new_AGEMA_signal_4318) ) ;
    buf_clk new_AGEMA_reg_buffer_1548 ( .C (clk), .D (new_AGEMA_signal_4323), .Q (new_AGEMA_signal_4324) ) ;
    buf_clk new_AGEMA_reg_buffer_1554 ( .C (clk), .D (new_AGEMA_signal_4329), .Q (new_AGEMA_signal_4330) ) ;
    buf_clk new_AGEMA_reg_buffer_1560 ( .C (clk), .D (new_AGEMA_signal_4335), .Q (new_AGEMA_signal_4336) ) ;
    buf_clk new_AGEMA_reg_buffer_1566 ( .C (clk), .D (new_AGEMA_signal_4341), .Q (new_AGEMA_signal_4342) ) ;
    buf_clk new_AGEMA_reg_buffer_1572 ( .C (clk), .D (new_AGEMA_signal_4347), .Q (new_AGEMA_signal_4348) ) ;
    buf_clk new_AGEMA_reg_buffer_1578 ( .C (clk), .D (new_AGEMA_signal_4353), .Q (new_AGEMA_signal_4354) ) ;
    buf_clk new_AGEMA_reg_buffer_1584 ( .C (clk), .D (new_AGEMA_signal_4359), .Q (new_AGEMA_signal_4360) ) ;
    buf_clk new_AGEMA_reg_buffer_1590 ( .C (clk), .D (new_AGEMA_signal_4365), .Q (new_AGEMA_signal_4366) ) ;
    buf_clk new_AGEMA_reg_buffer_1596 ( .C (clk), .D (new_AGEMA_signal_4371), .Q (new_AGEMA_signal_4372) ) ;
    buf_clk new_AGEMA_reg_buffer_1602 ( .C (clk), .D (new_AGEMA_signal_4377), .Q (new_AGEMA_signal_4378) ) ;
    buf_clk new_AGEMA_reg_buffer_1608 ( .C (clk), .D (new_AGEMA_signal_4383), .Q (new_AGEMA_signal_4384) ) ;
    buf_clk new_AGEMA_reg_buffer_1614 ( .C (clk), .D (new_AGEMA_signal_4389), .Q (new_AGEMA_signal_4390) ) ;
    buf_clk new_AGEMA_reg_buffer_1620 ( .C (clk), .D (new_AGEMA_signal_4395), .Q (new_AGEMA_signal_4396) ) ;
    buf_clk new_AGEMA_reg_buffer_1626 ( .C (clk), .D (new_AGEMA_signal_4401), .Q (new_AGEMA_signal_4402) ) ;
    buf_clk new_AGEMA_reg_buffer_1632 ( .C (clk), .D (new_AGEMA_signal_4407), .Q (new_AGEMA_signal_4408) ) ;
    buf_clk new_AGEMA_reg_buffer_1638 ( .C (clk), .D (new_AGEMA_signal_4413), .Q (new_AGEMA_signal_4414) ) ;
    buf_clk new_AGEMA_reg_buffer_1644 ( .C (clk), .D (new_AGEMA_signal_4419), .Q (new_AGEMA_signal_4420) ) ;
    buf_clk new_AGEMA_reg_buffer_1650 ( .C (clk), .D (new_AGEMA_signal_4425), .Q (new_AGEMA_signal_4426) ) ;
    buf_clk new_AGEMA_reg_buffer_1656 ( .C (clk), .D (new_AGEMA_signal_4431), .Q (new_AGEMA_signal_4432) ) ;
    buf_clk new_AGEMA_reg_buffer_1662 ( .C (clk), .D (new_AGEMA_signal_4437), .Q (new_AGEMA_signal_4438) ) ;
    buf_clk new_AGEMA_reg_buffer_1668 ( .C (clk), .D (new_AGEMA_signal_4443), .Q (new_AGEMA_signal_4444) ) ;
    buf_clk new_AGEMA_reg_buffer_1674 ( .C (clk), .D (new_AGEMA_signal_4449), .Q (new_AGEMA_signal_4450) ) ;
    buf_clk new_AGEMA_reg_buffer_1680 ( .C (clk), .D (new_AGEMA_signal_4455), .Q (new_AGEMA_signal_4456) ) ;
    buf_clk new_AGEMA_reg_buffer_1686 ( .C (clk), .D (new_AGEMA_signal_4461), .Q (new_AGEMA_signal_4462) ) ;
    buf_clk new_AGEMA_reg_buffer_1692 ( .C (clk), .D (new_AGEMA_signal_4467), .Q (new_AGEMA_signal_4468) ) ;
    buf_clk new_AGEMA_reg_buffer_1698 ( .C (clk), .D (new_AGEMA_signal_4473), .Q (new_AGEMA_signal_4474) ) ;
    buf_clk new_AGEMA_reg_buffer_1704 ( .C (clk), .D (new_AGEMA_signal_4479), .Q (new_AGEMA_signal_4480) ) ;
    buf_clk new_AGEMA_reg_buffer_1710 ( .C (clk), .D (new_AGEMA_signal_4485), .Q (new_AGEMA_signal_4486) ) ;
    buf_clk new_AGEMA_reg_buffer_1716 ( .C (clk), .D (new_AGEMA_signal_4491), .Q (new_AGEMA_signal_4492) ) ;
    buf_clk new_AGEMA_reg_buffer_1722 ( .C (clk), .D (new_AGEMA_signal_4497), .Q (new_AGEMA_signal_4498) ) ;
    buf_clk new_AGEMA_reg_buffer_1728 ( .C (clk), .D (new_AGEMA_signal_4503), .Q (new_AGEMA_signal_4504) ) ;
    buf_clk new_AGEMA_reg_buffer_1734 ( .C (clk), .D (new_AGEMA_signal_4509), .Q (new_AGEMA_signal_4510) ) ;
    buf_clk new_AGEMA_reg_buffer_1740 ( .C (clk), .D (new_AGEMA_signal_4515), .Q (new_AGEMA_signal_4516) ) ;
    buf_clk new_AGEMA_reg_buffer_1746 ( .C (clk), .D (new_AGEMA_signal_4521), .Q (new_AGEMA_signal_4522) ) ;
    buf_clk new_AGEMA_reg_buffer_1752 ( .C (clk), .D (new_AGEMA_signal_4527), .Q (new_AGEMA_signal_4528) ) ;
    buf_clk new_AGEMA_reg_buffer_1758 ( .C (clk), .D (new_AGEMA_signal_4533), .Q (new_AGEMA_signal_4534) ) ;
    buf_clk new_AGEMA_reg_buffer_1764 ( .C (clk), .D (new_AGEMA_signal_4539), .Q (new_AGEMA_signal_4540) ) ;
    buf_clk new_AGEMA_reg_buffer_1770 ( .C (clk), .D (new_AGEMA_signal_4545), .Q (new_AGEMA_signal_4546) ) ;
    buf_clk new_AGEMA_reg_buffer_1776 ( .C (clk), .D (new_AGEMA_signal_4551), .Q (new_AGEMA_signal_4552) ) ;
    buf_clk new_AGEMA_reg_buffer_1782 ( .C (clk), .D (new_AGEMA_signal_4557), .Q (new_AGEMA_signal_4558) ) ;
    buf_clk new_AGEMA_reg_buffer_1788 ( .C (clk), .D (new_AGEMA_signal_4563), .Q (new_AGEMA_signal_4564) ) ;
    buf_clk new_AGEMA_reg_buffer_1794 ( .C (clk), .D (new_AGEMA_signal_4569), .Q (new_AGEMA_signal_4570) ) ;
    buf_clk new_AGEMA_reg_buffer_1800 ( .C (clk), .D (new_AGEMA_signal_4575), .Q (new_AGEMA_signal_4576) ) ;
    buf_clk new_AGEMA_reg_buffer_1806 ( .C (clk), .D (new_AGEMA_signal_4581), .Q (new_AGEMA_signal_4582) ) ;
    buf_clk new_AGEMA_reg_buffer_1812 ( .C (clk), .D (new_AGEMA_signal_4587), .Q (new_AGEMA_signal_4588) ) ;
    buf_clk new_AGEMA_reg_buffer_1818 ( .C (clk), .D (new_AGEMA_signal_4593), .Q (new_AGEMA_signal_4594) ) ;
    buf_clk new_AGEMA_reg_buffer_1824 ( .C (clk), .D (new_AGEMA_signal_4599), .Q (new_AGEMA_signal_4600) ) ;
    buf_clk new_AGEMA_reg_buffer_1830 ( .C (clk), .D (new_AGEMA_signal_4605), .Q (new_AGEMA_signal_4606) ) ;
    buf_clk new_AGEMA_reg_buffer_1836 ( .C (clk), .D (new_AGEMA_signal_4611), .Q (new_AGEMA_signal_4612) ) ;
    buf_clk new_AGEMA_reg_buffer_1842 ( .C (clk), .D (new_AGEMA_signal_4617), .Q (new_AGEMA_signal_4618) ) ;
    buf_clk new_AGEMA_reg_buffer_1848 ( .C (clk), .D (new_AGEMA_signal_4623), .Q (new_AGEMA_signal_4624) ) ;
    buf_clk new_AGEMA_reg_buffer_1854 ( .C (clk), .D (new_AGEMA_signal_4629), .Q (new_AGEMA_signal_4630) ) ;
    buf_clk new_AGEMA_reg_buffer_1860 ( .C (clk), .D (new_AGEMA_signal_4635), .Q (new_AGEMA_signal_4636) ) ;
    buf_clk new_AGEMA_reg_buffer_1866 ( .C (clk), .D (new_AGEMA_signal_4641), .Q (new_AGEMA_signal_4642) ) ;
    buf_clk new_AGEMA_reg_buffer_1872 ( .C (clk), .D (new_AGEMA_signal_4647), .Q (new_AGEMA_signal_4648) ) ;
    buf_clk new_AGEMA_reg_buffer_1878 ( .C (clk), .D (new_AGEMA_signal_4653), .Q (new_AGEMA_signal_4654) ) ;
    buf_clk new_AGEMA_reg_buffer_1884 ( .C (clk), .D (new_AGEMA_signal_4659), .Q (new_AGEMA_signal_4660) ) ;
    buf_clk new_AGEMA_reg_buffer_1890 ( .C (clk), .D (new_AGEMA_signal_4665), .Q (new_AGEMA_signal_4666) ) ;
    buf_clk new_AGEMA_reg_buffer_1896 ( .C (clk), .D (new_AGEMA_signal_4671), .Q (new_AGEMA_signal_4672) ) ;
    buf_clk new_AGEMA_reg_buffer_1902 ( .C (clk), .D (new_AGEMA_signal_4677), .Q (new_AGEMA_signal_4678) ) ;
    buf_clk new_AGEMA_reg_buffer_1908 ( .C (clk), .D (new_AGEMA_signal_4683), .Q (new_AGEMA_signal_4684) ) ;
    buf_clk new_AGEMA_reg_buffer_1914 ( .C (clk), .D (new_AGEMA_signal_4689), .Q (new_AGEMA_signal_4690) ) ;
    buf_clk new_AGEMA_reg_buffer_1920 ( .C (clk), .D (new_AGEMA_signal_4695), .Q (new_AGEMA_signal_4696) ) ;
    buf_clk new_AGEMA_reg_buffer_1926 ( .C (clk), .D (new_AGEMA_signal_4701), .Q (new_AGEMA_signal_4702) ) ;
    buf_clk new_AGEMA_reg_buffer_1932 ( .C (clk), .D (new_AGEMA_signal_4707), .Q (new_AGEMA_signal_4708) ) ;
    buf_clk new_AGEMA_reg_buffer_1938 ( .C (clk), .D (new_AGEMA_signal_4713), .Q (new_AGEMA_signal_4714) ) ;
    buf_clk new_AGEMA_reg_buffer_1944 ( .C (clk), .D (new_AGEMA_signal_4719), .Q (new_AGEMA_signal_4720) ) ;
    buf_clk new_AGEMA_reg_buffer_1950 ( .C (clk), .D (new_AGEMA_signal_4725), .Q (new_AGEMA_signal_4726) ) ;
    buf_clk new_AGEMA_reg_buffer_1956 ( .C (clk), .D (new_AGEMA_signal_4731), .Q (new_AGEMA_signal_4732) ) ;
    buf_clk new_AGEMA_reg_buffer_1962 ( .C (clk), .D (new_AGEMA_signal_4737), .Q (new_AGEMA_signal_4738) ) ;
    buf_clk new_AGEMA_reg_buffer_1968 ( .C (clk), .D (new_AGEMA_signal_4743), .Q (new_AGEMA_signal_4744) ) ;
    buf_clk new_AGEMA_reg_buffer_1974 ( .C (clk), .D (new_AGEMA_signal_4749), .Q (new_AGEMA_signal_4750) ) ;
    buf_clk new_AGEMA_reg_buffer_1980 ( .C (clk), .D (new_AGEMA_signal_4755), .Q (new_AGEMA_signal_4756) ) ;
    buf_clk new_AGEMA_reg_buffer_1986 ( .C (clk), .D (new_AGEMA_signal_4761), .Q (new_AGEMA_signal_4762) ) ;
    buf_clk new_AGEMA_reg_buffer_1992 ( .C (clk), .D (new_AGEMA_signal_4767), .Q (new_AGEMA_signal_4768) ) ;
    buf_clk new_AGEMA_reg_buffer_1998 ( .C (clk), .D (new_AGEMA_signal_4773), .Q (new_AGEMA_signal_4774) ) ;
    buf_clk new_AGEMA_reg_buffer_2004 ( .C (clk), .D (new_AGEMA_signal_4779), .Q (new_AGEMA_signal_4780) ) ;
    buf_clk new_AGEMA_reg_buffer_2010 ( .C (clk), .D (new_AGEMA_signal_4785), .Q (new_AGEMA_signal_4786) ) ;
    buf_clk new_AGEMA_reg_buffer_2016 ( .C (clk), .D (new_AGEMA_signal_4791), .Q (new_AGEMA_signal_4792) ) ;
    buf_clk new_AGEMA_reg_buffer_2022 ( .C (clk), .D (new_AGEMA_signal_4797), .Q (new_AGEMA_signal_4798) ) ;
    buf_clk new_AGEMA_reg_buffer_2028 ( .C (clk), .D (new_AGEMA_signal_4803), .Q (new_AGEMA_signal_4804) ) ;
    buf_clk new_AGEMA_reg_buffer_2034 ( .C (clk), .D (new_AGEMA_signal_4809), .Q (new_AGEMA_signal_4810) ) ;
    buf_clk new_AGEMA_reg_buffer_2040 ( .C (clk), .D (new_AGEMA_signal_4815), .Q (new_AGEMA_signal_4816) ) ;
    buf_clk new_AGEMA_reg_buffer_2046 ( .C (clk), .D (new_AGEMA_signal_4821), .Q (new_AGEMA_signal_4822) ) ;
    buf_clk new_AGEMA_reg_buffer_2052 ( .C (clk), .D (new_AGEMA_signal_4827), .Q (new_AGEMA_signal_4828) ) ;
    buf_clk new_AGEMA_reg_buffer_2058 ( .C (clk), .D (new_AGEMA_signal_4833), .Q (new_AGEMA_signal_4834) ) ;
    buf_clk new_AGEMA_reg_buffer_2064 ( .C (clk), .D (new_AGEMA_signal_4839), .Q (new_AGEMA_signal_4840) ) ;
    buf_clk new_AGEMA_reg_buffer_2070 ( .C (clk), .D (new_AGEMA_signal_4845), .Q (new_AGEMA_signal_4846) ) ;
    buf_clk new_AGEMA_reg_buffer_2076 ( .C (clk), .D (new_AGEMA_signal_4851), .Q (new_AGEMA_signal_4852) ) ;
    buf_clk new_AGEMA_reg_buffer_2082 ( .C (clk), .D (new_AGEMA_signal_4857), .Q (new_AGEMA_signal_4858) ) ;
    buf_clk new_AGEMA_reg_buffer_2088 ( .C (clk), .D (new_AGEMA_signal_4863), .Q (new_AGEMA_signal_4864) ) ;
    buf_clk new_AGEMA_reg_buffer_2094 ( .C (clk), .D (new_AGEMA_signal_4869), .Q (new_AGEMA_signal_4870) ) ;
    buf_clk new_AGEMA_reg_buffer_2100 ( .C (clk), .D (new_AGEMA_signal_4875), .Q (new_AGEMA_signal_4876) ) ;
    buf_clk new_AGEMA_reg_buffer_2106 ( .C (clk), .D (new_AGEMA_signal_4881), .Q (new_AGEMA_signal_4882) ) ;
    buf_clk new_AGEMA_reg_buffer_2112 ( .C (clk), .D (new_AGEMA_signal_4887), .Q (new_AGEMA_signal_4888) ) ;
    buf_clk new_AGEMA_reg_buffer_2118 ( .C (clk), .D (new_AGEMA_signal_4893), .Q (new_AGEMA_signal_4894) ) ;
    buf_clk new_AGEMA_reg_buffer_2124 ( .C (clk), .D (new_AGEMA_signal_4899), .Q (new_AGEMA_signal_4900) ) ;
    buf_clk new_AGEMA_reg_buffer_2130 ( .C (clk), .D (new_AGEMA_signal_4905), .Q (new_AGEMA_signal_4906) ) ;
    buf_clk new_AGEMA_reg_buffer_2136 ( .C (clk), .D (new_AGEMA_signal_4911), .Q (new_AGEMA_signal_4912) ) ;
    buf_clk new_AGEMA_reg_buffer_2142 ( .C (clk), .D (new_AGEMA_signal_4917), .Q (new_AGEMA_signal_4918) ) ;
    buf_clk new_AGEMA_reg_buffer_2148 ( .C (clk), .D (new_AGEMA_signal_4923), .Q (new_AGEMA_signal_4924) ) ;
    buf_clk new_AGEMA_reg_buffer_2154 ( .C (clk), .D (new_AGEMA_signal_4929), .Q (new_AGEMA_signal_4930) ) ;
    buf_clk new_AGEMA_reg_buffer_2160 ( .C (clk), .D (new_AGEMA_signal_4935), .Q (new_AGEMA_signal_4936) ) ;
    buf_clk new_AGEMA_reg_buffer_2166 ( .C (clk), .D (new_AGEMA_signal_4941), .Q (new_AGEMA_signal_4942) ) ;
    buf_clk new_AGEMA_reg_buffer_2172 ( .C (clk), .D (new_AGEMA_signal_4947), .Q (new_AGEMA_signal_4948) ) ;
    buf_clk new_AGEMA_reg_buffer_2178 ( .C (clk), .D (new_AGEMA_signal_4953), .Q (new_AGEMA_signal_4954) ) ;
    buf_clk new_AGEMA_reg_buffer_2184 ( .C (clk), .D (new_AGEMA_signal_4959), .Q (new_AGEMA_signal_4960) ) ;
    buf_clk new_AGEMA_reg_buffer_2190 ( .C (clk), .D (new_AGEMA_signal_4965), .Q (new_AGEMA_signal_4966) ) ;
    buf_clk new_AGEMA_reg_buffer_2196 ( .C (clk), .D (new_AGEMA_signal_4971), .Q (new_AGEMA_signal_4972) ) ;
    buf_clk new_AGEMA_reg_buffer_2202 ( .C (clk), .D (new_AGEMA_signal_4977), .Q (new_AGEMA_signal_4978) ) ;
    buf_clk new_AGEMA_reg_buffer_2208 ( .C (clk), .D (new_AGEMA_signal_4983), .Q (new_AGEMA_signal_4984) ) ;
    buf_clk new_AGEMA_reg_buffer_2214 ( .C (clk), .D (new_AGEMA_signal_4989), .Q (new_AGEMA_signal_4990) ) ;
    buf_clk new_AGEMA_reg_buffer_2220 ( .C (clk), .D (new_AGEMA_signal_4995), .Q (new_AGEMA_signal_4996) ) ;
    buf_clk new_AGEMA_reg_buffer_2226 ( .C (clk), .D (new_AGEMA_signal_5001), .Q (new_AGEMA_signal_5002) ) ;
    buf_clk new_AGEMA_reg_buffer_2232 ( .C (clk), .D (new_AGEMA_signal_5007), .Q (new_AGEMA_signal_5008) ) ;
    buf_clk new_AGEMA_reg_buffer_2238 ( .C (clk), .D (new_AGEMA_signal_5013), .Q (new_AGEMA_signal_5014) ) ;
    buf_clk new_AGEMA_reg_buffer_2244 ( .C (clk), .D (new_AGEMA_signal_5019), .Q (new_AGEMA_signal_5020) ) ;
    buf_clk new_AGEMA_reg_buffer_2250 ( .C (clk), .D (new_AGEMA_signal_5025), .Q (new_AGEMA_signal_5026) ) ;
    buf_clk new_AGEMA_reg_buffer_2256 ( .C (clk), .D (new_AGEMA_signal_5031), .Q (new_AGEMA_signal_5032) ) ;
    buf_clk new_AGEMA_reg_buffer_2262 ( .C (clk), .D (new_AGEMA_signal_5037), .Q (new_AGEMA_signal_5038) ) ;
    buf_clk new_AGEMA_reg_buffer_2268 ( .C (clk), .D (new_AGEMA_signal_5043), .Q (new_AGEMA_signal_5044) ) ;
    buf_clk new_AGEMA_reg_buffer_2274 ( .C (clk), .D (new_AGEMA_signal_5049), .Q (new_AGEMA_signal_5050) ) ;
    buf_clk new_AGEMA_reg_buffer_2280 ( .C (clk), .D (new_AGEMA_signal_5055), .Q (new_AGEMA_signal_5056) ) ;
    buf_clk new_AGEMA_reg_buffer_2286 ( .C (clk), .D (new_AGEMA_signal_5061), .Q (new_AGEMA_signal_5062) ) ;
    buf_clk new_AGEMA_reg_buffer_2292 ( .C (clk), .D (new_AGEMA_signal_5067), .Q (new_AGEMA_signal_5068) ) ;
    buf_clk new_AGEMA_reg_buffer_2298 ( .C (clk), .D (new_AGEMA_signal_5073), .Q (new_AGEMA_signal_5074) ) ;
    buf_clk new_AGEMA_reg_buffer_2304 ( .C (clk), .D (new_AGEMA_signal_5079), .Q (new_AGEMA_signal_5080) ) ;
    buf_clk new_AGEMA_reg_buffer_2310 ( .C (clk), .D (new_AGEMA_signal_5085), .Q (new_AGEMA_signal_5086) ) ;
    buf_clk new_AGEMA_reg_buffer_2316 ( .C (clk), .D (new_AGEMA_signal_5091), .Q (new_AGEMA_signal_5092) ) ;
    buf_clk new_AGEMA_reg_buffer_2322 ( .C (clk), .D (new_AGEMA_signal_5097), .Q (new_AGEMA_signal_5098) ) ;
    buf_clk new_AGEMA_reg_buffer_2328 ( .C (clk), .D (new_AGEMA_signal_5103), .Q (new_AGEMA_signal_5104) ) ;
    buf_clk new_AGEMA_reg_buffer_2334 ( .C (clk), .D (new_AGEMA_signal_5109), .Q (new_AGEMA_signal_5110) ) ;
    buf_clk new_AGEMA_reg_buffer_2340 ( .C (clk), .D (new_AGEMA_signal_5115), .Q (new_AGEMA_signal_5116) ) ;
    buf_clk new_AGEMA_reg_buffer_2346 ( .C (clk), .D (new_AGEMA_signal_5121), .Q (new_AGEMA_signal_5122) ) ;
    buf_clk new_AGEMA_reg_buffer_2352 ( .C (clk), .D (new_AGEMA_signal_5127), .Q (new_AGEMA_signal_5128) ) ;
    buf_clk new_AGEMA_reg_buffer_2358 ( .C (clk), .D (new_AGEMA_signal_5133), .Q (new_AGEMA_signal_5134) ) ;
    buf_clk new_AGEMA_reg_buffer_2362 ( .C (clk), .D (new_AGEMA_signal_5137), .Q (new_AGEMA_signal_5138) ) ;
    buf_clk new_AGEMA_reg_buffer_2364 ( .C (clk), .D (new_AGEMA_signal_5139), .Q (new_AGEMA_signal_5140) ) ;
    buf_clk new_AGEMA_reg_buffer_2366 ( .C (clk), .D (new_AGEMA_signal_5141), .Q (new_AGEMA_signal_5142) ) ;
    buf_clk new_AGEMA_reg_buffer_2368 ( .C (clk), .D (new_AGEMA_signal_5143), .Q (new_AGEMA_signal_5144) ) ;
    buf_clk new_AGEMA_reg_buffer_2370 ( .C (clk), .D (new_AGEMA_signal_5145), .Q (new_AGEMA_signal_5146) ) ;
    buf_clk new_AGEMA_reg_buffer_2372 ( .C (clk), .D (new_AGEMA_signal_5147), .Q (new_AGEMA_signal_5148) ) ;
    buf_clk new_AGEMA_reg_buffer_2374 ( .C (clk), .D (new_AGEMA_signal_5149), .Q (new_AGEMA_signal_5150) ) ;
    buf_clk new_AGEMA_reg_buffer_2376 ( .C (clk), .D (new_AGEMA_signal_5151), .Q (new_AGEMA_signal_5152) ) ;
    buf_clk new_AGEMA_reg_buffer_2378 ( .C (clk), .D (new_AGEMA_signal_5153), .Q (new_AGEMA_signal_5154) ) ;
    buf_clk new_AGEMA_reg_buffer_2380 ( .C (clk), .D (new_AGEMA_signal_5155), .Q (new_AGEMA_signal_5156) ) ;
    buf_clk new_AGEMA_reg_buffer_2382 ( .C (clk), .D (new_AGEMA_signal_5157), .Q (new_AGEMA_signal_5158) ) ;
    buf_clk new_AGEMA_reg_buffer_2384 ( .C (clk), .D (new_AGEMA_signal_5159), .Q (new_AGEMA_signal_5160) ) ;
    buf_clk new_AGEMA_reg_buffer_2386 ( .C (clk), .D (new_AGEMA_signal_5161), .Q (new_AGEMA_signal_5162) ) ;
    buf_clk new_AGEMA_reg_buffer_2388 ( .C (clk), .D (new_AGEMA_signal_5163), .Q (new_AGEMA_signal_5164) ) ;
    buf_clk new_AGEMA_reg_buffer_2390 ( .C (clk), .D (new_AGEMA_signal_5165), .Q (new_AGEMA_signal_5166) ) ;
    buf_clk new_AGEMA_reg_buffer_2392 ( .C (clk), .D (new_AGEMA_signal_5167), .Q (new_AGEMA_signal_5168) ) ;
    buf_clk new_AGEMA_reg_buffer_2394 ( .C (clk), .D (new_AGEMA_signal_5169), .Q (new_AGEMA_signal_5170) ) ;
    buf_clk new_AGEMA_reg_buffer_2396 ( .C (clk), .D (new_AGEMA_signal_5171), .Q (new_AGEMA_signal_5172) ) ;
    buf_clk new_AGEMA_reg_buffer_2398 ( .C (clk), .D (new_AGEMA_signal_5173), .Q (new_AGEMA_signal_5174) ) ;
    buf_clk new_AGEMA_reg_buffer_2400 ( .C (clk), .D (new_AGEMA_signal_5175), .Q (new_AGEMA_signal_5176) ) ;
    buf_clk new_AGEMA_reg_buffer_2402 ( .C (clk), .D (new_AGEMA_signal_5177), .Q (new_AGEMA_signal_5178) ) ;
    buf_clk new_AGEMA_reg_buffer_2404 ( .C (clk), .D (new_AGEMA_signal_5179), .Q (new_AGEMA_signal_5180) ) ;
    buf_clk new_AGEMA_reg_buffer_2406 ( .C (clk), .D (new_AGEMA_signal_5181), .Q (new_AGEMA_signal_5182) ) ;
    buf_clk new_AGEMA_reg_buffer_2408 ( .C (clk), .D (new_AGEMA_signal_5183), .Q (new_AGEMA_signal_5184) ) ;
    buf_clk new_AGEMA_reg_buffer_2410 ( .C (clk), .D (new_AGEMA_signal_5185), .Q (new_AGEMA_signal_5186) ) ;
    buf_clk new_AGEMA_reg_buffer_2412 ( .C (clk), .D (new_AGEMA_signal_5187), .Q (new_AGEMA_signal_5188) ) ;
    buf_clk new_AGEMA_reg_buffer_2414 ( .C (clk), .D (new_AGEMA_signal_5189), .Q (new_AGEMA_signal_5190) ) ;
    buf_clk new_AGEMA_reg_buffer_2416 ( .C (clk), .D (new_AGEMA_signal_5191), .Q (new_AGEMA_signal_5192) ) ;
    buf_clk new_AGEMA_reg_buffer_2418 ( .C (clk), .D (new_AGEMA_signal_5193), .Q (new_AGEMA_signal_5194) ) ;
    buf_clk new_AGEMA_reg_buffer_2420 ( .C (clk), .D (new_AGEMA_signal_5195), .Q (new_AGEMA_signal_5196) ) ;
    buf_clk new_AGEMA_reg_buffer_2422 ( .C (clk), .D (new_AGEMA_signal_5197), .Q (new_AGEMA_signal_5198) ) ;
    buf_clk new_AGEMA_reg_buffer_2424 ( .C (clk), .D (new_AGEMA_signal_5199), .Q (new_AGEMA_signal_5200) ) ;
    buf_clk new_AGEMA_reg_buffer_2426 ( .C (clk), .D (new_AGEMA_signal_5201), .Q (new_AGEMA_signal_5202) ) ;
    buf_clk new_AGEMA_reg_buffer_2428 ( .C (clk), .D (new_AGEMA_signal_5203), .Q (new_AGEMA_signal_5204) ) ;
    buf_clk new_AGEMA_reg_buffer_2430 ( .C (clk), .D (new_AGEMA_signal_5205), .Q (new_AGEMA_signal_5206) ) ;
    buf_clk new_AGEMA_reg_buffer_2432 ( .C (clk), .D (new_AGEMA_signal_5207), .Q (new_AGEMA_signal_5208) ) ;
    buf_clk new_AGEMA_reg_buffer_2434 ( .C (clk), .D (new_AGEMA_signal_5209), .Q (new_AGEMA_signal_5210) ) ;
    buf_clk new_AGEMA_reg_buffer_2436 ( .C (clk), .D (new_AGEMA_signal_5211), .Q (new_AGEMA_signal_5212) ) ;
    buf_clk new_AGEMA_reg_buffer_2438 ( .C (clk), .D (new_AGEMA_signal_5213), .Q (new_AGEMA_signal_5214) ) ;
    buf_clk new_AGEMA_reg_buffer_2440 ( .C (clk), .D (new_AGEMA_signal_5215), .Q (new_AGEMA_signal_5216) ) ;
    buf_clk new_AGEMA_reg_buffer_2442 ( .C (clk), .D (new_AGEMA_signal_5217), .Q (new_AGEMA_signal_5218) ) ;
    buf_clk new_AGEMA_reg_buffer_2444 ( .C (clk), .D (new_AGEMA_signal_5219), .Q (new_AGEMA_signal_5220) ) ;
    buf_clk new_AGEMA_reg_buffer_2446 ( .C (clk), .D (new_AGEMA_signal_5221), .Q (new_AGEMA_signal_5222) ) ;
    buf_clk new_AGEMA_reg_buffer_2448 ( .C (clk), .D (new_AGEMA_signal_5223), .Q (new_AGEMA_signal_5224) ) ;
    buf_clk new_AGEMA_reg_buffer_2450 ( .C (clk), .D (new_AGEMA_signal_5225), .Q (new_AGEMA_signal_5226) ) ;
    buf_clk new_AGEMA_reg_buffer_2452 ( .C (clk), .D (new_AGEMA_signal_5227), .Q (new_AGEMA_signal_5228) ) ;
    buf_clk new_AGEMA_reg_buffer_2454 ( .C (clk), .D (new_AGEMA_signal_5229), .Q (new_AGEMA_signal_5230) ) ;
    buf_clk new_AGEMA_reg_buffer_2456 ( .C (clk), .D (new_AGEMA_signal_5231), .Q (new_AGEMA_signal_5232) ) ;
    buf_clk new_AGEMA_reg_buffer_2458 ( .C (clk), .D (new_AGEMA_signal_5233), .Q (new_AGEMA_signal_5234) ) ;
    buf_clk new_AGEMA_reg_buffer_2460 ( .C (clk), .D (new_AGEMA_signal_5235), .Q (new_AGEMA_signal_5236) ) ;
    buf_clk new_AGEMA_reg_buffer_2462 ( .C (clk), .D (new_AGEMA_signal_5237), .Q (new_AGEMA_signal_5238) ) ;
    buf_clk new_AGEMA_reg_buffer_2464 ( .C (clk), .D (new_AGEMA_signal_5239), .Q (new_AGEMA_signal_5240) ) ;
    buf_clk new_AGEMA_reg_buffer_2466 ( .C (clk), .D (new_AGEMA_signal_5241), .Q (new_AGEMA_signal_5242) ) ;
    buf_clk new_AGEMA_reg_buffer_2468 ( .C (clk), .D (new_AGEMA_signal_5243), .Q (new_AGEMA_signal_5244) ) ;
    buf_clk new_AGEMA_reg_buffer_2470 ( .C (clk), .D (new_AGEMA_signal_5245), .Q (new_AGEMA_signal_5246) ) ;
    buf_clk new_AGEMA_reg_buffer_2472 ( .C (clk), .D (new_AGEMA_signal_5247), .Q (new_AGEMA_signal_5248) ) ;
    buf_clk new_AGEMA_reg_buffer_2474 ( .C (clk), .D (new_AGEMA_signal_5249), .Q (new_AGEMA_signal_5250) ) ;
    buf_clk new_AGEMA_reg_buffer_2476 ( .C (clk), .D (new_AGEMA_signal_5251), .Q (new_AGEMA_signal_5252) ) ;
    buf_clk new_AGEMA_reg_buffer_2478 ( .C (clk), .D (new_AGEMA_signal_5253), .Q (new_AGEMA_signal_5254) ) ;
    buf_clk new_AGEMA_reg_buffer_2480 ( .C (clk), .D (new_AGEMA_signal_5255), .Q (new_AGEMA_signal_5256) ) ;
    buf_clk new_AGEMA_reg_buffer_2482 ( .C (clk), .D (new_AGEMA_signal_5257), .Q (new_AGEMA_signal_5258) ) ;
    buf_clk new_AGEMA_reg_buffer_2484 ( .C (clk), .D (new_AGEMA_signal_5259), .Q (new_AGEMA_signal_5260) ) ;
    buf_clk new_AGEMA_reg_buffer_2486 ( .C (clk), .D (new_AGEMA_signal_5261), .Q (new_AGEMA_signal_5262) ) ;
    buf_clk new_AGEMA_reg_buffer_2488 ( .C (clk), .D (new_AGEMA_signal_5263), .Q (new_AGEMA_signal_5264) ) ;
    buf_clk new_AGEMA_reg_buffer_2490 ( .C (clk), .D (new_AGEMA_signal_5265), .Q (new_AGEMA_signal_5266) ) ;
    buf_clk new_AGEMA_reg_buffer_2492 ( .C (clk), .D (new_AGEMA_signal_5267), .Q (new_AGEMA_signal_5268) ) ;
    buf_clk new_AGEMA_reg_buffer_2494 ( .C (clk), .D (new_AGEMA_signal_5269), .Q (new_AGEMA_signal_5270) ) ;
    buf_clk new_AGEMA_reg_buffer_2496 ( .C (clk), .D (new_AGEMA_signal_5271), .Q (new_AGEMA_signal_5272) ) ;
    buf_clk new_AGEMA_reg_buffer_2498 ( .C (clk), .D (new_AGEMA_signal_5273), .Q (new_AGEMA_signal_5274) ) ;
    buf_clk new_AGEMA_reg_buffer_2500 ( .C (clk), .D (new_AGEMA_signal_5275), .Q (new_AGEMA_signal_5276) ) ;
    buf_clk new_AGEMA_reg_buffer_2502 ( .C (clk), .D (new_AGEMA_signal_5277), .Q (new_AGEMA_signal_5278) ) ;
    buf_clk new_AGEMA_reg_buffer_2504 ( .C (clk), .D (new_AGEMA_signal_5279), .Q (new_AGEMA_signal_5280) ) ;
    buf_clk new_AGEMA_reg_buffer_2506 ( .C (clk), .D (new_AGEMA_signal_5281), .Q (new_AGEMA_signal_5282) ) ;
    buf_clk new_AGEMA_reg_buffer_2508 ( .C (clk), .D (new_AGEMA_signal_5283), .Q (new_AGEMA_signal_5284) ) ;
    buf_clk new_AGEMA_reg_buffer_2510 ( .C (clk), .D (new_AGEMA_signal_5285), .Q (new_AGEMA_signal_5286) ) ;
    buf_clk new_AGEMA_reg_buffer_2512 ( .C (clk), .D (new_AGEMA_signal_5287), .Q (new_AGEMA_signal_5288) ) ;
    buf_clk new_AGEMA_reg_buffer_2514 ( .C (clk), .D (new_AGEMA_signal_5289), .Q (new_AGEMA_signal_5290) ) ;
    buf_clk new_AGEMA_reg_buffer_2516 ( .C (clk), .D (new_AGEMA_signal_5291), .Q (new_AGEMA_signal_5292) ) ;
    buf_clk new_AGEMA_reg_buffer_2518 ( .C (clk), .D (new_AGEMA_signal_5293), .Q (new_AGEMA_signal_5294) ) ;
    buf_clk new_AGEMA_reg_buffer_2520 ( .C (clk), .D (new_AGEMA_signal_5295), .Q (new_AGEMA_signal_5296) ) ;
    buf_clk new_AGEMA_reg_buffer_2522 ( .C (clk), .D (new_AGEMA_signal_5297), .Q (new_AGEMA_signal_5298) ) ;
    buf_clk new_AGEMA_reg_buffer_2524 ( .C (clk), .D (new_AGEMA_signal_5299), .Q (new_AGEMA_signal_5300) ) ;
    buf_clk new_AGEMA_reg_buffer_2526 ( .C (clk), .D (new_AGEMA_signal_5301), .Q (new_AGEMA_signal_5302) ) ;
    buf_clk new_AGEMA_reg_buffer_2528 ( .C (clk), .D (new_AGEMA_signal_5303), .Q (new_AGEMA_signal_5304) ) ;
    buf_clk new_AGEMA_reg_buffer_2530 ( .C (clk), .D (new_AGEMA_signal_5305), .Q (new_AGEMA_signal_5306) ) ;
    buf_clk new_AGEMA_reg_buffer_2532 ( .C (clk), .D (new_AGEMA_signal_5307), .Q (new_AGEMA_signal_5308) ) ;
    buf_clk new_AGEMA_reg_buffer_2534 ( .C (clk), .D (new_AGEMA_signal_5309), .Q (new_AGEMA_signal_5310) ) ;
    buf_clk new_AGEMA_reg_buffer_2536 ( .C (clk), .D (new_AGEMA_signal_5311), .Q (new_AGEMA_signal_5312) ) ;
    buf_clk new_AGEMA_reg_buffer_2538 ( .C (clk), .D (new_AGEMA_signal_5313), .Q (new_AGEMA_signal_5314) ) ;
    buf_clk new_AGEMA_reg_buffer_2540 ( .C (clk), .D (new_AGEMA_signal_5315), .Q (new_AGEMA_signal_5316) ) ;
    buf_clk new_AGEMA_reg_buffer_2542 ( .C (clk), .D (new_AGEMA_signal_5317), .Q (new_AGEMA_signal_5318) ) ;
    buf_clk new_AGEMA_reg_buffer_2544 ( .C (clk), .D (new_AGEMA_signal_5319), .Q (new_AGEMA_signal_5320) ) ;
    buf_clk new_AGEMA_reg_buffer_2546 ( .C (clk), .D (new_AGEMA_signal_5321), .Q (new_AGEMA_signal_5322) ) ;
    buf_clk new_AGEMA_reg_buffer_2548 ( .C (clk), .D (new_AGEMA_signal_5323), .Q (new_AGEMA_signal_5324) ) ;
    buf_clk new_AGEMA_reg_buffer_2550 ( .C (clk), .D (new_AGEMA_signal_5325), .Q (new_AGEMA_signal_5326) ) ;
    buf_clk new_AGEMA_reg_buffer_2552 ( .C (clk), .D (new_AGEMA_signal_5327), .Q (new_AGEMA_signal_5328) ) ;
    buf_clk new_AGEMA_reg_buffer_2554 ( .C (clk), .D (new_AGEMA_signal_5329), .Q (new_AGEMA_signal_5330) ) ;
    buf_clk new_AGEMA_reg_buffer_2556 ( .C (clk), .D (new_AGEMA_signal_5331), .Q (new_AGEMA_signal_5332) ) ;
    buf_clk new_AGEMA_reg_buffer_2558 ( .C (clk), .D (new_AGEMA_signal_5333), .Q (new_AGEMA_signal_5334) ) ;
    buf_clk new_AGEMA_reg_buffer_2560 ( .C (clk), .D (new_AGEMA_signal_5335), .Q (new_AGEMA_signal_5336) ) ;
    buf_clk new_AGEMA_reg_buffer_2562 ( .C (clk), .D (new_AGEMA_signal_5337), .Q (new_AGEMA_signal_5338) ) ;
    buf_clk new_AGEMA_reg_buffer_2564 ( .C (clk), .D (new_AGEMA_signal_5339), .Q (new_AGEMA_signal_5340) ) ;
    buf_clk new_AGEMA_reg_buffer_2566 ( .C (clk), .D (new_AGEMA_signal_5341), .Q (new_AGEMA_signal_5342) ) ;
    buf_clk new_AGEMA_reg_buffer_2568 ( .C (clk), .D (new_AGEMA_signal_5343), .Q (new_AGEMA_signal_5344) ) ;
    buf_clk new_AGEMA_reg_buffer_2570 ( .C (clk), .D (new_AGEMA_signal_5345), .Q (new_AGEMA_signal_5346) ) ;
    buf_clk new_AGEMA_reg_buffer_2572 ( .C (clk), .D (new_AGEMA_signal_5347), .Q (new_AGEMA_signal_5348) ) ;
    buf_clk new_AGEMA_reg_buffer_2574 ( .C (clk), .D (new_AGEMA_signal_5349), .Q (new_AGEMA_signal_5350) ) ;
    buf_clk new_AGEMA_reg_buffer_2576 ( .C (clk), .D (new_AGEMA_signal_5351), .Q (new_AGEMA_signal_5352) ) ;
    buf_clk new_AGEMA_reg_buffer_2578 ( .C (clk), .D (new_AGEMA_signal_5353), .Q (new_AGEMA_signal_5354) ) ;
    buf_clk new_AGEMA_reg_buffer_2580 ( .C (clk), .D (new_AGEMA_signal_5355), .Q (new_AGEMA_signal_5356) ) ;
    buf_clk new_AGEMA_reg_buffer_2582 ( .C (clk), .D (new_AGEMA_signal_5357), .Q (new_AGEMA_signal_5358) ) ;
    buf_clk new_AGEMA_reg_buffer_2584 ( .C (clk), .D (new_AGEMA_signal_5359), .Q (new_AGEMA_signal_5360) ) ;
    buf_clk new_AGEMA_reg_buffer_2586 ( .C (clk), .D (new_AGEMA_signal_5361), .Q (new_AGEMA_signal_5362) ) ;
    buf_clk new_AGEMA_reg_buffer_2588 ( .C (clk), .D (new_AGEMA_signal_5363), .Q (new_AGEMA_signal_5364) ) ;
    buf_clk new_AGEMA_reg_buffer_2590 ( .C (clk), .D (new_AGEMA_signal_5365), .Q (new_AGEMA_signal_5366) ) ;
    buf_clk new_AGEMA_reg_buffer_2592 ( .C (clk), .D (new_AGEMA_signal_5367), .Q (new_AGEMA_signal_5368) ) ;
    buf_clk new_AGEMA_reg_buffer_2594 ( .C (clk), .D (new_AGEMA_signal_5369), .Q (new_AGEMA_signal_5370) ) ;
    buf_clk new_AGEMA_reg_buffer_2596 ( .C (clk), .D (new_AGEMA_signal_5371), .Q (new_AGEMA_signal_5372) ) ;
    buf_clk new_AGEMA_reg_buffer_2598 ( .C (clk), .D (new_AGEMA_signal_5373), .Q (new_AGEMA_signal_5374) ) ;
    buf_clk new_AGEMA_reg_buffer_2600 ( .C (clk), .D (new_AGEMA_signal_5375), .Q (new_AGEMA_signal_5376) ) ;
    buf_clk new_AGEMA_reg_buffer_2602 ( .C (clk), .D (new_AGEMA_signal_5377), .Q (new_AGEMA_signal_5378) ) ;
    buf_clk new_AGEMA_reg_buffer_2604 ( .C (clk), .D (new_AGEMA_signal_5379), .Q (new_AGEMA_signal_5380) ) ;
    buf_clk new_AGEMA_reg_buffer_2606 ( .C (clk), .D (new_AGEMA_signal_5381), .Q (new_AGEMA_signal_5382) ) ;
    buf_clk new_AGEMA_reg_buffer_2608 ( .C (clk), .D (new_AGEMA_signal_5383), .Q (new_AGEMA_signal_5384) ) ;
    buf_clk new_AGEMA_reg_buffer_2610 ( .C (clk), .D (new_AGEMA_signal_5385), .Q (new_AGEMA_signal_5386) ) ;
    buf_clk new_AGEMA_reg_buffer_2612 ( .C (clk), .D (new_AGEMA_signal_5387), .Q (new_AGEMA_signal_5388) ) ;
    buf_clk new_AGEMA_reg_buffer_2614 ( .C (clk), .D (new_AGEMA_signal_5389), .Q (new_AGEMA_signal_5390) ) ;
    buf_clk new_AGEMA_reg_buffer_2616 ( .C (clk), .D (new_AGEMA_signal_5391), .Q (new_AGEMA_signal_5392) ) ;
    buf_clk new_AGEMA_reg_buffer_2618 ( .C (clk), .D (new_AGEMA_signal_5393), .Q (new_AGEMA_signal_5394) ) ;
    buf_clk new_AGEMA_reg_buffer_2620 ( .C (clk), .D (new_AGEMA_signal_5395), .Q (new_AGEMA_signal_5396) ) ;
    buf_clk new_AGEMA_reg_buffer_2622 ( .C (clk), .D (new_AGEMA_signal_5397), .Q (new_AGEMA_signal_5398) ) ;
    buf_clk new_AGEMA_reg_buffer_2624 ( .C (clk), .D (new_AGEMA_signal_5399), .Q (new_AGEMA_signal_5400) ) ;
    buf_clk new_AGEMA_reg_buffer_2626 ( .C (clk), .D (new_AGEMA_signal_5401), .Q (new_AGEMA_signal_5402) ) ;
    buf_clk new_AGEMA_reg_buffer_2628 ( .C (clk), .D (new_AGEMA_signal_5403), .Q (new_AGEMA_signal_5404) ) ;
    buf_clk new_AGEMA_reg_buffer_2630 ( .C (clk), .D (new_AGEMA_signal_5405), .Q (new_AGEMA_signal_5406) ) ;
    buf_clk new_AGEMA_reg_buffer_2632 ( .C (clk), .D (new_AGEMA_signal_5407), .Q (new_AGEMA_signal_5408) ) ;
    buf_clk new_AGEMA_reg_buffer_2634 ( .C (clk), .D (new_AGEMA_signal_5409), .Q (new_AGEMA_signal_5410) ) ;
    buf_clk new_AGEMA_reg_buffer_2636 ( .C (clk), .D (new_AGEMA_signal_5411), .Q (new_AGEMA_signal_5412) ) ;
    buf_clk new_AGEMA_reg_buffer_2638 ( .C (clk), .D (new_AGEMA_signal_5413), .Q (new_AGEMA_signal_5414) ) ;
    buf_clk new_AGEMA_reg_buffer_2640 ( .C (clk), .D (new_AGEMA_signal_5415), .Q (new_AGEMA_signal_5416) ) ;
    buf_clk new_AGEMA_reg_buffer_2642 ( .C (clk), .D (new_AGEMA_signal_5417), .Q (new_AGEMA_signal_5418) ) ;
    buf_clk new_AGEMA_reg_buffer_2644 ( .C (clk), .D (new_AGEMA_signal_5419), .Q (new_AGEMA_signal_5420) ) ;
    buf_clk new_AGEMA_reg_buffer_2646 ( .C (clk), .D (new_AGEMA_signal_5421), .Q (new_AGEMA_signal_5422) ) ;
    buf_clk new_AGEMA_reg_buffer_2648 ( .C (clk), .D (new_AGEMA_signal_5423), .Q (new_AGEMA_signal_5424) ) ;
    buf_clk new_AGEMA_reg_buffer_2654 ( .C (clk), .D (new_AGEMA_signal_5429), .Q (new_AGEMA_signal_5430) ) ;
    buf_clk new_AGEMA_reg_buffer_2662 ( .C (clk), .D (new_AGEMA_signal_5437), .Q (new_AGEMA_signal_5438) ) ;
    buf_clk new_AGEMA_reg_buffer_2670 ( .C (clk), .D (new_AGEMA_signal_5445), .Q (new_AGEMA_signal_5446) ) ;
    buf_clk new_AGEMA_reg_buffer_2678 ( .C (clk), .D (new_AGEMA_signal_5453), .Q (new_AGEMA_signal_5454) ) ;
    buf_clk new_AGEMA_reg_buffer_2686 ( .C (clk), .D (new_AGEMA_signal_5461), .Q (new_AGEMA_signal_5462) ) ;
    buf_clk new_AGEMA_reg_buffer_2694 ( .C (clk), .D (new_AGEMA_signal_5469), .Q (new_AGEMA_signal_5470) ) ;
    buf_clk new_AGEMA_reg_buffer_2702 ( .C (clk), .D (new_AGEMA_signal_5477), .Q (new_AGEMA_signal_5478) ) ;
    buf_clk new_AGEMA_reg_buffer_2710 ( .C (clk), .D (new_AGEMA_signal_5485), .Q (new_AGEMA_signal_5486) ) ;
    buf_clk new_AGEMA_reg_buffer_2718 ( .C (clk), .D (new_AGEMA_signal_5493), .Q (new_AGEMA_signal_5494) ) ;
    buf_clk new_AGEMA_reg_buffer_2726 ( .C (clk), .D (new_AGEMA_signal_5501), .Q (new_AGEMA_signal_5502) ) ;
    buf_clk new_AGEMA_reg_buffer_2734 ( .C (clk), .D (new_AGEMA_signal_5509), .Q (new_AGEMA_signal_5510) ) ;
    buf_clk new_AGEMA_reg_buffer_2742 ( .C (clk), .D (new_AGEMA_signal_5517), .Q (new_AGEMA_signal_5518) ) ;
    buf_clk new_AGEMA_reg_buffer_2750 ( .C (clk), .D (new_AGEMA_signal_5525), .Q (new_AGEMA_signal_5526) ) ;
    buf_clk new_AGEMA_reg_buffer_2758 ( .C (clk), .D (new_AGEMA_signal_5533), .Q (new_AGEMA_signal_5534) ) ;
    buf_clk new_AGEMA_reg_buffer_2766 ( .C (clk), .D (new_AGEMA_signal_5541), .Q (new_AGEMA_signal_5542) ) ;
    buf_clk new_AGEMA_reg_buffer_2774 ( .C (clk), .D (new_AGEMA_signal_5549), .Q (new_AGEMA_signal_5550) ) ;
    buf_clk new_AGEMA_reg_buffer_2782 ( .C (clk), .D (new_AGEMA_signal_5557), .Q (new_AGEMA_signal_5558) ) ;
    buf_clk new_AGEMA_reg_buffer_2790 ( .C (clk), .D (new_AGEMA_signal_5565), .Q (new_AGEMA_signal_5566) ) ;
    buf_clk new_AGEMA_reg_buffer_2798 ( .C (clk), .D (new_AGEMA_signal_5573), .Q (new_AGEMA_signal_5574) ) ;
    buf_clk new_AGEMA_reg_buffer_2806 ( .C (clk), .D (new_AGEMA_signal_5581), .Q (new_AGEMA_signal_5582) ) ;
    buf_clk new_AGEMA_reg_buffer_2814 ( .C (clk), .D (new_AGEMA_signal_5589), .Q (new_AGEMA_signal_5590) ) ;
    buf_clk new_AGEMA_reg_buffer_2822 ( .C (clk), .D (new_AGEMA_signal_5597), .Q (new_AGEMA_signal_5598) ) ;
    buf_clk new_AGEMA_reg_buffer_2830 ( .C (clk), .D (new_AGEMA_signal_5605), .Q (new_AGEMA_signal_5606) ) ;
    buf_clk new_AGEMA_reg_buffer_2838 ( .C (clk), .D (new_AGEMA_signal_5613), .Q (new_AGEMA_signal_5614) ) ;
    buf_clk new_AGEMA_reg_buffer_2846 ( .C (clk), .D (new_AGEMA_signal_5621), .Q (new_AGEMA_signal_5622) ) ;
    buf_clk new_AGEMA_reg_buffer_2854 ( .C (clk), .D (new_AGEMA_signal_5629), .Q (new_AGEMA_signal_5630) ) ;
    buf_clk new_AGEMA_reg_buffer_2862 ( .C (clk), .D (new_AGEMA_signal_5637), .Q (new_AGEMA_signal_5638) ) ;
    buf_clk new_AGEMA_reg_buffer_2870 ( .C (clk), .D (new_AGEMA_signal_5645), .Q (new_AGEMA_signal_5646) ) ;
    buf_clk new_AGEMA_reg_buffer_2878 ( .C (clk), .D (new_AGEMA_signal_5653), .Q (new_AGEMA_signal_5654) ) ;
    buf_clk new_AGEMA_reg_buffer_2886 ( .C (clk), .D (new_AGEMA_signal_5661), .Q (new_AGEMA_signal_5662) ) ;
    buf_clk new_AGEMA_reg_buffer_2894 ( .C (clk), .D (new_AGEMA_signal_5669), .Q (new_AGEMA_signal_5670) ) ;
    buf_clk new_AGEMA_reg_buffer_2902 ( .C (clk), .D (new_AGEMA_signal_5677), .Q (new_AGEMA_signal_5678) ) ;
    buf_clk new_AGEMA_reg_buffer_2910 ( .C (clk), .D (new_AGEMA_signal_5685), .Q (new_AGEMA_signal_5686) ) ;
    buf_clk new_AGEMA_reg_buffer_2918 ( .C (clk), .D (new_AGEMA_signal_5693), .Q (new_AGEMA_signal_5694) ) ;
    buf_clk new_AGEMA_reg_buffer_2926 ( .C (clk), .D (new_AGEMA_signal_5701), .Q (new_AGEMA_signal_5702) ) ;
    buf_clk new_AGEMA_reg_buffer_2934 ( .C (clk), .D (new_AGEMA_signal_5709), .Q (new_AGEMA_signal_5710) ) ;
    buf_clk new_AGEMA_reg_buffer_2942 ( .C (clk), .D (new_AGEMA_signal_5717), .Q (new_AGEMA_signal_5718) ) ;
    buf_clk new_AGEMA_reg_buffer_2950 ( .C (clk), .D (new_AGEMA_signal_5725), .Q (new_AGEMA_signal_5726) ) ;
    buf_clk new_AGEMA_reg_buffer_2958 ( .C (clk), .D (new_AGEMA_signal_5733), .Q (new_AGEMA_signal_5734) ) ;
    buf_clk new_AGEMA_reg_buffer_2966 ( .C (clk), .D (new_AGEMA_signal_5741), .Q (new_AGEMA_signal_5742) ) ;
    buf_clk new_AGEMA_reg_buffer_2974 ( .C (clk), .D (new_AGEMA_signal_5749), .Q (new_AGEMA_signal_5750) ) ;
    buf_clk new_AGEMA_reg_buffer_2982 ( .C (clk), .D (new_AGEMA_signal_5757), .Q (new_AGEMA_signal_5758) ) ;
    buf_clk new_AGEMA_reg_buffer_2990 ( .C (clk), .D (new_AGEMA_signal_5765), .Q (new_AGEMA_signal_5766) ) ;
    buf_clk new_AGEMA_reg_buffer_2998 ( .C (clk), .D (new_AGEMA_signal_5773), .Q (new_AGEMA_signal_5774) ) ;
    buf_clk new_AGEMA_reg_buffer_3006 ( .C (clk), .D (new_AGEMA_signal_5781), .Q (new_AGEMA_signal_5782) ) ;
    buf_clk new_AGEMA_reg_buffer_3014 ( .C (clk), .D (new_AGEMA_signal_5789), .Q (new_AGEMA_signal_5790) ) ;
    buf_clk new_AGEMA_reg_buffer_3022 ( .C (clk), .D (new_AGEMA_signal_5797), .Q (new_AGEMA_signal_5798) ) ;
    buf_clk new_AGEMA_reg_buffer_3030 ( .C (clk), .D (new_AGEMA_signal_5805), .Q (new_AGEMA_signal_5806) ) ;
    buf_clk new_AGEMA_reg_buffer_3038 ( .C (clk), .D (new_AGEMA_signal_5813), .Q (new_AGEMA_signal_5814) ) ;
    buf_clk new_AGEMA_reg_buffer_3046 ( .C (clk), .D (new_AGEMA_signal_5821), .Q (new_AGEMA_signal_5822) ) ;
    buf_clk new_AGEMA_reg_buffer_3054 ( .C (clk), .D (new_AGEMA_signal_5829), .Q (new_AGEMA_signal_5830) ) ;
    buf_clk new_AGEMA_reg_buffer_3062 ( .C (clk), .D (new_AGEMA_signal_5837), .Q (new_AGEMA_signal_5838) ) ;
    buf_clk new_AGEMA_reg_buffer_3070 ( .C (clk), .D (new_AGEMA_signal_5845), .Q (new_AGEMA_signal_5846) ) ;
    buf_clk new_AGEMA_reg_buffer_3078 ( .C (clk), .D (new_AGEMA_signal_5853), .Q (new_AGEMA_signal_5854) ) ;
    buf_clk new_AGEMA_reg_buffer_3086 ( .C (clk), .D (new_AGEMA_signal_5861), .Q (new_AGEMA_signal_5862) ) ;
    buf_clk new_AGEMA_reg_buffer_3094 ( .C (clk), .D (new_AGEMA_signal_5869), .Q (new_AGEMA_signal_5870) ) ;
    buf_clk new_AGEMA_reg_buffer_3102 ( .C (clk), .D (new_AGEMA_signal_5877), .Q (new_AGEMA_signal_5878) ) ;
    buf_clk new_AGEMA_reg_buffer_3110 ( .C (clk), .D (new_AGEMA_signal_5885), .Q (new_AGEMA_signal_5886) ) ;
    buf_clk new_AGEMA_reg_buffer_3118 ( .C (clk), .D (new_AGEMA_signal_5893), .Q (new_AGEMA_signal_5894) ) ;
    buf_clk new_AGEMA_reg_buffer_3126 ( .C (clk), .D (new_AGEMA_signal_5901), .Q (new_AGEMA_signal_5902) ) ;
    buf_clk new_AGEMA_reg_buffer_3134 ( .C (clk), .D (new_AGEMA_signal_5909), .Q (new_AGEMA_signal_5910) ) ;
    buf_clk new_AGEMA_reg_buffer_3142 ( .C (clk), .D (new_AGEMA_signal_5917), .Q (new_AGEMA_signal_5918) ) ;
    buf_clk new_AGEMA_reg_buffer_3150 ( .C (clk), .D (new_AGEMA_signal_5925), .Q (new_AGEMA_signal_5926) ) ;
    buf_clk new_AGEMA_reg_buffer_3158 ( .C (clk), .D (new_AGEMA_signal_5933), .Q (new_AGEMA_signal_5934) ) ;
    buf_clk new_AGEMA_reg_buffer_3166 ( .C (clk), .D (new_AGEMA_signal_5941), .Q (new_AGEMA_signal_5942) ) ;
    buf_clk new_AGEMA_reg_buffer_3174 ( .C (clk), .D (new_AGEMA_signal_5949), .Q (new_AGEMA_signal_5950) ) ;
    buf_clk new_AGEMA_reg_buffer_3182 ( .C (clk), .D (new_AGEMA_signal_5957), .Q (new_AGEMA_signal_5958) ) ;
    buf_clk new_AGEMA_reg_buffer_3190 ( .C (clk), .D (new_AGEMA_signal_5965), .Q (new_AGEMA_signal_5966) ) ;
    buf_clk new_AGEMA_reg_buffer_3198 ( .C (clk), .D (new_AGEMA_signal_5973), .Q (new_AGEMA_signal_5974) ) ;
    buf_clk new_AGEMA_reg_buffer_3206 ( .C (clk), .D (new_AGEMA_signal_5981), .Q (new_AGEMA_signal_5982) ) ;
    buf_clk new_AGEMA_reg_buffer_3214 ( .C (clk), .D (new_AGEMA_signal_5989), .Q (new_AGEMA_signal_5990) ) ;
    buf_clk new_AGEMA_reg_buffer_3222 ( .C (clk), .D (new_AGEMA_signal_5997), .Q (new_AGEMA_signal_5998) ) ;
    buf_clk new_AGEMA_reg_buffer_3230 ( .C (clk), .D (new_AGEMA_signal_6005), .Q (new_AGEMA_signal_6006) ) ;
    buf_clk new_AGEMA_reg_buffer_3238 ( .C (clk), .D (new_AGEMA_signal_6013), .Q (new_AGEMA_signal_6014) ) ;
    buf_clk new_AGEMA_reg_buffer_3246 ( .C (clk), .D (new_AGEMA_signal_6021), .Q (new_AGEMA_signal_6022) ) ;
    buf_clk new_AGEMA_reg_buffer_3254 ( .C (clk), .D (new_AGEMA_signal_6029), .Q (new_AGEMA_signal_6030) ) ;
    buf_clk new_AGEMA_reg_buffer_3262 ( .C (clk), .D (new_AGEMA_signal_6037), .Q (new_AGEMA_signal_6038) ) ;
    buf_clk new_AGEMA_reg_buffer_3270 ( .C (clk), .D (new_AGEMA_signal_6045), .Q (new_AGEMA_signal_6046) ) ;
    buf_clk new_AGEMA_reg_buffer_3278 ( .C (clk), .D (new_AGEMA_signal_6053), .Q (new_AGEMA_signal_6054) ) ;
    buf_clk new_AGEMA_reg_buffer_3286 ( .C (clk), .D (new_AGEMA_signal_6061), .Q (new_AGEMA_signal_6062) ) ;
    buf_clk new_AGEMA_reg_buffer_3294 ( .C (clk), .D (new_AGEMA_signal_6069), .Q (new_AGEMA_signal_6070) ) ;
    buf_clk new_AGEMA_reg_buffer_3302 ( .C (clk), .D (new_AGEMA_signal_6077), .Q (new_AGEMA_signal_6078) ) ;
    buf_clk new_AGEMA_reg_buffer_3310 ( .C (clk), .D (new_AGEMA_signal_6085), .Q (new_AGEMA_signal_6086) ) ;
    buf_clk new_AGEMA_reg_buffer_3318 ( .C (clk), .D (new_AGEMA_signal_6093), .Q (new_AGEMA_signal_6094) ) ;
    buf_clk new_AGEMA_reg_buffer_3326 ( .C (clk), .D (new_AGEMA_signal_6101), .Q (new_AGEMA_signal_6102) ) ;
    buf_clk new_AGEMA_reg_buffer_3334 ( .C (clk), .D (new_AGEMA_signal_6109), .Q (new_AGEMA_signal_6110) ) ;
    buf_clk new_AGEMA_reg_buffer_3342 ( .C (clk), .D (new_AGEMA_signal_6117), .Q (new_AGEMA_signal_6118) ) ;
    buf_clk new_AGEMA_reg_buffer_3350 ( .C (clk), .D (new_AGEMA_signal_6125), .Q (new_AGEMA_signal_6126) ) ;
    buf_clk new_AGEMA_reg_buffer_3358 ( .C (clk), .D (new_AGEMA_signal_6133), .Q (new_AGEMA_signal_6134) ) ;
    buf_clk new_AGEMA_reg_buffer_3366 ( .C (clk), .D (new_AGEMA_signal_6141), .Q (new_AGEMA_signal_6142) ) ;
    buf_clk new_AGEMA_reg_buffer_3374 ( .C (clk), .D (new_AGEMA_signal_6149), .Q (new_AGEMA_signal_6150) ) ;
    buf_clk new_AGEMA_reg_buffer_3382 ( .C (clk), .D (new_AGEMA_signal_6157), .Q (new_AGEMA_signal_6158) ) ;
    buf_clk new_AGEMA_reg_buffer_3390 ( .C (clk), .D (new_AGEMA_signal_6165), .Q (new_AGEMA_signal_6166) ) ;
    buf_clk new_AGEMA_reg_buffer_3398 ( .C (clk), .D (new_AGEMA_signal_6173), .Q (new_AGEMA_signal_6174) ) ;
    buf_clk new_AGEMA_reg_buffer_3406 ( .C (clk), .D (new_AGEMA_signal_6181), .Q (new_AGEMA_signal_6182) ) ;
    buf_clk new_AGEMA_reg_buffer_3414 ( .C (clk), .D (new_AGEMA_signal_6189), .Q (new_AGEMA_signal_6190) ) ;
    buf_clk new_AGEMA_reg_buffer_3422 ( .C (clk), .D (new_AGEMA_signal_6197), .Q (new_AGEMA_signal_6198) ) ;
    buf_clk new_AGEMA_reg_buffer_3430 ( .C (clk), .D (new_AGEMA_signal_6205), .Q (new_AGEMA_signal_6206) ) ;
    buf_clk new_AGEMA_reg_buffer_3438 ( .C (clk), .D (new_AGEMA_signal_6213), .Q (new_AGEMA_signal_6214) ) ;
    buf_clk new_AGEMA_reg_buffer_3446 ( .C (clk), .D (new_AGEMA_signal_6221), .Q (new_AGEMA_signal_6222) ) ;
    buf_clk new_AGEMA_reg_buffer_3454 ( .C (clk), .D (new_AGEMA_signal_6229), .Q (new_AGEMA_signal_6230) ) ;
    buf_clk new_AGEMA_reg_buffer_3462 ( .C (clk), .D (new_AGEMA_signal_6237), .Q (new_AGEMA_signal_6238) ) ;
    buf_clk new_AGEMA_reg_buffer_3470 ( .C (clk), .D (new_AGEMA_signal_6245), .Q (new_AGEMA_signal_6246) ) ;
    buf_clk new_AGEMA_reg_buffer_3478 ( .C (clk), .D (new_AGEMA_signal_6253), .Q (new_AGEMA_signal_6254) ) ;
    buf_clk new_AGEMA_reg_buffer_3486 ( .C (clk), .D (new_AGEMA_signal_6261), .Q (new_AGEMA_signal_6262) ) ;
    buf_clk new_AGEMA_reg_buffer_3494 ( .C (clk), .D (new_AGEMA_signal_6269), .Q (new_AGEMA_signal_6270) ) ;
    buf_clk new_AGEMA_reg_buffer_3502 ( .C (clk), .D (new_AGEMA_signal_6277), .Q (new_AGEMA_signal_6278) ) ;
    buf_clk new_AGEMA_reg_buffer_3510 ( .C (clk), .D (new_AGEMA_signal_6285), .Q (new_AGEMA_signal_6286) ) ;
    buf_clk new_AGEMA_reg_buffer_3518 ( .C (clk), .D (new_AGEMA_signal_6293), .Q (new_AGEMA_signal_6294) ) ;
    buf_clk new_AGEMA_reg_buffer_3526 ( .C (clk), .D (new_AGEMA_signal_6301), .Q (new_AGEMA_signal_6302) ) ;
    buf_clk new_AGEMA_reg_buffer_3534 ( .C (clk), .D (new_AGEMA_signal_6309), .Q (new_AGEMA_signal_6310) ) ;
    buf_clk new_AGEMA_reg_buffer_3542 ( .C (clk), .D (new_AGEMA_signal_6317), .Q (new_AGEMA_signal_6318) ) ;
    buf_clk new_AGEMA_reg_buffer_3550 ( .C (clk), .D (new_AGEMA_signal_6325), .Q (new_AGEMA_signal_6326) ) ;
    buf_clk new_AGEMA_reg_buffer_3558 ( .C (clk), .D (new_AGEMA_signal_6333), .Q (new_AGEMA_signal_6334) ) ;
    buf_clk new_AGEMA_reg_buffer_3566 ( .C (clk), .D (new_AGEMA_signal_6341), .Q (new_AGEMA_signal_6342) ) ;
    buf_clk new_AGEMA_reg_buffer_3574 ( .C (clk), .D (new_AGEMA_signal_6349), .Q (new_AGEMA_signal_6350) ) ;
    buf_clk new_AGEMA_reg_buffer_3582 ( .C (clk), .D (new_AGEMA_signal_6357), .Q (new_AGEMA_signal_6358) ) ;
    buf_clk new_AGEMA_reg_buffer_3590 ( .C (clk), .D (new_AGEMA_signal_6365), .Q (new_AGEMA_signal_6366) ) ;
    buf_clk new_AGEMA_reg_buffer_3598 ( .C (clk), .D (new_AGEMA_signal_6373), .Q (new_AGEMA_signal_6374) ) ;
    buf_clk new_AGEMA_reg_buffer_3606 ( .C (clk), .D (new_AGEMA_signal_6381), .Q (new_AGEMA_signal_6382) ) ;
    buf_clk new_AGEMA_reg_buffer_3614 ( .C (clk), .D (new_AGEMA_signal_6389), .Q (new_AGEMA_signal_6390) ) ;
    buf_clk new_AGEMA_reg_buffer_3622 ( .C (clk), .D (new_AGEMA_signal_6397), .Q (new_AGEMA_signal_6398) ) ;
    buf_clk new_AGEMA_reg_buffer_3630 ( .C (clk), .D (new_AGEMA_signal_6405), .Q (new_AGEMA_signal_6406) ) ;
    buf_clk new_AGEMA_reg_buffer_3638 ( .C (clk), .D (new_AGEMA_signal_6413), .Q (new_AGEMA_signal_6414) ) ;
    buf_clk new_AGEMA_reg_buffer_3646 ( .C (clk), .D (new_AGEMA_signal_6421), .Q (new_AGEMA_signal_6422) ) ;
    buf_clk new_AGEMA_reg_buffer_3654 ( .C (clk), .D (new_AGEMA_signal_6429), .Q (new_AGEMA_signal_6430) ) ;
    buf_clk new_AGEMA_reg_buffer_3662 ( .C (clk), .D (new_AGEMA_signal_6437), .Q (new_AGEMA_signal_6438) ) ;
    buf_clk new_AGEMA_reg_buffer_3670 ( .C (clk), .D (new_AGEMA_signal_6445), .Q (new_AGEMA_signal_6446) ) ;
    buf_clk new_AGEMA_reg_buffer_3678 ( .C (clk), .D (new_AGEMA_signal_6453), .Q (new_AGEMA_signal_6454) ) ;
    buf_clk new_AGEMA_reg_buffer_3686 ( .C (clk), .D (new_AGEMA_signal_6461), .Q (new_AGEMA_signal_6462) ) ;
    buf_clk new_AGEMA_reg_buffer_3694 ( .C (clk), .D (new_AGEMA_signal_6469), .Q (new_AGEMA_signal_6470) ) ;
    buf_clk new_AGEMA_reg_buffer_3702 ( .C (clk), .D (new_AGEMA_signal_6477), .Q (new_AGEMA_signal_6478) ) ;
    buf_clk new_AGEMA_reg_buffer_3710 ( .C (clk), .D (new_AGEMA_signal_6485), .Q (new_AGEMA_signal_6486) ) ;
    buf_clk new_AGEMA_reg_buffer_3718 ( .C (clk), .D (new_AGEMA_signal_6493), .Q (new_AGEMA_signal_6494) ) ;
    buf_clk new_AGEMA_reg_buffer_3726 ( .C (clk), .D (new_AGEMA_signal_6501), .Q (new_AGEMA_signal_6502) ) ;
    buf_clk new_AGEMA_reg_buffer_3734 ( .C (clk), .D (new_AGEMA_signal_6509), .Q (new_AGEMA_signal_6510) ) ;
    buf_clk new_AGEMA_reg_buffer_3742 ( .C (clk), .D (new_AGEMA_signal_6517), .Q (new_AGEMA_signal_6518) ) ;
    buf_clk new_AGEMA_reg_buffer_3750 ( .C (clk), .D (new_AGEMA_signal_6525), .Q (new_AGEMA_signal_6526) ) ;
    buf_clk new_AGEMA_reg_buffer_3758 ( .C (clk), .D (new_AGEMA_signal_6533), .Q (new_AGEMA_signal_6534) ) ;
    buf_clk new_AGEMA_reg_buffer_3766 ( .C (clk), .D (new_AGEMA_signal_6541), .Q (new_AGEMA_signal_6542) ) ;
    buf_clk new_AGEMA_reg_buffer_3774 ( .C (clk), .D (new_AGEMA_signal_6549), .Q (new_AGEMA_signal_6550) ) ;
    buf_clk new_AGEMA_reg_buffer_3782 ( .C (clk), .D (new_AGEMA_signal_6557), .Q (new_AGEMA_signal_6558) ) ;
    buf_clk new_AGEMA_reg_buffer_3790 ( .C (clk), .D (new_AGEMA_signal_6565), .Q (new_AGEMA_signal_6566) ) ;
    buf_clk new_AGEMA_reg_buffer_3798 ( .C (clk), .D (new_AGEMA_signal_6573), .Q (new_AGEMA_signal_6574) ) ;
    buf_clk new_AGEMA_reg_buffer_3806 ( .C (clk), .D (new_AGEMA_signal_6581), .Q (new_AGEMA_signal_6582) ) ;
    buf_clk new_AGEMA_reg_buffer_3814 ( .C (clk), .D (new_AGEMA_signal_6589), .Q (new_AGEMA_signal_6590) ) ;
    buf_clk new_AGEMA_reg_buffer_3822 ( .C (clk), .D (new_AGEMA_signal_6597), .Q (new_AGEMA_signal_6598) ) ;
    buf_clk new_AGEMA_reg_buffer_3830 ( .C (clk), .D (new_AGEMA_signal_6605), .Q (new_AGEMA_signal_6606) ) ;
    buf_clk new_AGEMA_reg_buffer_3838 ( .C (clk), .D (new_AGEMA_signal_6613), .Q (new_AGEMA_signal_6614) ) ;
    buf_clk new_AGEMA_reg_buffer_3846 ( .C (clk), .D (new_AGEMA_signal_6621), .Q (new_AGEMA_signal_6622) ) ;
    buf_clk new_AGEMA_reg_buffer_3854 ( .C (clk), .D (new_AGEMA_signal_6629), .Q (new_AGEMA_signal_6630) ) ;
    buf_clk new_AGEMA_reg_buffer_3862 ( .C (clk), .D (new_AGEMA_signal_6637), .Q (new_AGEMA_signal_6638) ) ;
    buf_clk new_AGEMA_reg_buffer_3870 ( .C (clk), .D (new_AGEMA_signal_6645), .Q (new_AGEMA_signal_6646) ) ;
    buf_clk new_AGEMA_reg_buffer_3878 ( .C (clk), .D (new_AGEMA_signal_6653), .Q (new_AGEMA_signal_6654) ) ;
    buf_clk new_AGEMA_reg_buffer_3886 ( .C (clk), .D (new_AGEMA_signal_6661), .Q (new_AGEMA_signal_6662) ) ;
    buf_clk new_AGEMA_reg_buffer_3894 ( .C (clk), .D (new_AGEMA_signal_6669), .Q (new_AGEMA_signal_6670) ) ;
    buf_clk new_AGEMA_reg_buffer_3902 ( .C (clk), .D (new_AGEMA_signal_6677), .Q (new_AGEMA_signal_6678) ) ;
    buf_clk new_AGEMA_reg_buffer_3910 ( .C (clk), .D (new_AGEMA_signal_6685), .Q (new_AGEMA_signal_6686) ) ;
    buf_clk new_AGEMA_reg_buffer_3918 ( .C (clk), .D (new_AGEMA_signal_6693), .Q (new_AGEMA_signal_6694) ) ;
    buf_clk new_AGEMA_reg_buffer_3926 ( .C (clk), .D (new_AGEMA_signal_6701), .Q (new_AGEMA_signal_6702) ) ;
    buf_clk new_AGEMA_reg_buffer_3934 ( .C (clk), .D (new_AGEMA_signal_6709), .Q (new_AGEMA_signal_6710) ) ;
    buf_clk new_AGEMA_reg_buffer_3942 ( .C (clk), .D (new_AGEMA_signal_6717), .Q (new_AGEMA_signal_6718) ) ;
    buf_clk new_AGEMA_reg_buffer_3950 ( .C (clk), .D (new_AGEMA_signal_6725), .Q (new_AGEMA_signal_6726) ) ;
    buf_clk new_AGEMA_reg_buffer_3958 ( .C (clk), .D (new_AGEMA_signal_6733), .Q (new_AGEMA_signal_6734) ) ;
    buf_clk new_AGEMA_reg_buffer_3966 ( .C (clk), .D (new_AGEMA_signal_6741), .Q (new_AGEMA_signal_6742) ) ;
    buf_clk new_AGEMA_reg_buffer_3974 ( .C (clk), .D (new_AGEMA_signal_6749), .Q (new_AGEMA_signal_6750) ) ;
    buf_clk new_AGEMA_reg_buffer_3982 ( .C (clk), .D (new_AGEMA_signal_6757), .Q (new_AGEMA_signal_6758) ) ;
    buf_clk new_AGEMA_reg_buffer_3990 ( .C (clk), .D (new_AGEMA_signal_6765), .Q (new_AGEMA_signal_6766) ) ;
    buf_clk new_AGEMA_reg_buffer_3998 ( .C (clk), .D (new_AGEMA_signal_6773), .Q (new_AGEMA_signal_6774) ) ;
    buf_clk new_AGEMA_reg_buffer_4006 ( .C (clk), .D (new_AGEMA_signal_6781), .Q (new_AGEMA_signal_6782) ) ;
    buf_clk new_AGEMA_reg_buffer_4014 ( .C (clk), .D (new_AGEMA_signal_6789), .Q (new_AGEMA_signal_6790) ) ;
    buf_clk new_AGEMA_reg_buffer_4022 ( .C (clk), .D (new_AGEMA_signal_6797), .Q (new_AGEMA_signal_6798) ) ;
    buf_clk new_AGEMA_reg_buffer_4030 ( .C (clk), .D (new_AGEMA_signal_6805), .Q (new_AGEMA_signal_6806) ) ;
    buf_clk new_AGEMA_reg_buffer_4038 ( .C (clk), .D (new_AGEMA_signal_6813), .Q (new_AGEMA_signal_6814) ) ;
    buf_clk new_AGEMA_reg_buffer_4046 ( .C (clk), .D (new_AGEMA_signal_6821), .Q (new_AGEMA_signal_6822) ) ;
    buf_clk new_AGEMA_reg_buffer_4054 ( .C (clk), .D (new_AGEMA_signal_6829), .Q (new_AGEMA_signal_6830) ) ;
    buf_clk new_AGEMA_reg_buffer_4062 ( .C (clk), .D (new_AGEMA_signal_6837), .Q (new_AGEMA_signal_6838) ) ;
    buf_clk new_AGEMA_reg_buffer_4070 ( .C (clk), .D (new_AGEMA_signal_6845), .Q (new_AGEMA_signal_6846) ) ;
    buf_clk new_AGEMA_reg_buffer_4078 ( .C (clk), .D (new_AGEMA_signal_6853), .Q (new_AGEMA_signal_6854) ) ;
    buf_clk new_AGEMA_reg_buffer_4086 ( .C (clk), .D (new_AGEMA_signal_6861), .Q (new_AGEMA_signal_6862) ) ;
    buf_clk new_AGEMA_reg_buffer_4094 ( .C (clk), .D (new_AGEMA_signal_6869), .Q (new_AGEMA_signal_6870) ) ;
    buf_clk new_AGEMA_reg_buffer_4102 ( .C (clk), .D (new_AGEMA_signal_6877), .Q (new_AGEMA_signal_6878) ) ;
    buf_clk new_AGEMA_reg_buffer_4110 ( .C (clk), .D (new_AGEMA_signal_6885), .Q (new_AGEMA_signal_6886) ) ;
    buf_clk new_AGEMA_reg_buffer_4118 ( .C (clk), .D (new_AGEMA_signal_6893), .Q (new_AGEMA_signal_6894) ) ;
    buf_clk new_AGEMA_reg_buffer_4126 ( .C (clk), .D (new_AGEMA_signal_6901), .Q (new_AGEMA_signal_6902) ) ;
    buf_clk new_AGEMA_reg_buffer_4134 ( .C (clk), .D (new_AGEMA_signal_6909), .Q (new_AGEMA_signal_6910) ) ;
    buf_clk new_AGEMA_reg_buffer_4142 ( .C (clk), .D (new_AGEMA_signal_6917), .Q (new_AGEMA_signal_6918) ) ;
    buf_clk new_AGEMA_reg_buffer_4150 ( .C (clk), .D (new_AGEMA_signal_6925), .Q (new_AGEMA_signal_6926) ) ;
    buf_clk new_AGEMA_reg_buffer_4158 ( .C (clk), .D (new_AGEMA_signal_6933), .Q (new_AGEMA_signal_6934) ) ;
    buf_clk new_AGEMA_reg_buffer_4166 ( .C (clk), .D (new_AGEMA_signal_6941), .Q (new_AGEMA_signal_6942) ) ;
    buf_clk new_AGEMA_reg_buffer_4174 ( .C (clk), .D (new_AGEMA_signal_6949), .Q (new_AGEMA_signal_6950) ) ;
    buf_clk new_AGEMA_reg_buffer_4182 ( .C (clk), .D (new_AGEMA_signal_6957), .Q (new_AGEMA_signal_6958) ) ;
    buf_clk new_AGEMA_reg_buffer_4194 ( .C (clk), .D (new_AGEMA_signal_6969), .Q (new_AGEMA_signal_6970) ) ;
    buf_clk new_AGEMA_reg_buffer_4198 ( .C (clk), .D (new_AGEMA_signal_6973), .Q (new_AGEMA_signal_6974) ) ;
    buf_clk new_AGEMA_reg_buffer_4202 ( .C (clk), .D (new_AGEMA_signal_6977), .Q (new_AGEMA_signal_6978) ) ;
    buf_clk new_AGEMA_reg_buffer_4212 ( .C (clk), .D (new_AGEMA_signal_6987), .Q (new_AGEMA_signal_6988) ) ;
    buf_clk new_AGEMA_reg_buffer_4216 ( .C (clk), .D (new_AGEMA_signal_6991), .Q (new_AGEMA_signal_6992) ) ;
    buf_clk new_AGEMA_reg_buffer_4220 ( .C (clk), .D (new_AGEMA_signal_6995), .Q (new_AGEMA_signal_6996) ) ;
    buf_clk new_AGEMA_reg_buffer_4230 ( .C (clk), .D (new_AGEMA_signal_7005), .Q (new_AGEMA_signal_7006) ) ;
    buf_clk new_AGEMA_reg_buffer_4234 ( .C (clk), .D (new_AGEMA_signal_7009), .Q (new_AGEMA_signal_7010) ) ;
    buf_clk new_AGEMA_reg_buffer_4238 ( .C (clk), .D (new_AGEMA_signal_7013), .Q (new_AGEMA_signal_7014) ) ;
    buf_clk new_AGEMA_reg_buffer_4248 ( .C (clk), .D (new_AGEMA_signal_7023), .Q (new_AGEMA_signal_7024) ) ;
    buf_clk new_AGEMA_reg_buffer_4252 ( .C (clk), .D (new_AGEMA_signal_7027), .Q (new_AGEMA_signal_7028) ) ;
    buf_clk new_AGEMA_reg_buffer_4256 ( .C (clk), .D (new_AGEMA_signal_7031), .Q (new_AGEMA_signal_7032) ) ;
    buf_clk new_AGEMA_reg_buffer_4266 ( .C (clk), .D (new_AGEMA_signal_7041), .Q (new_AGEMA_signal_7042) ) ;
    buf_clk new_AGEMA_reg_buffer_4270 ( .C (clk), .D (new_AGEMA_signal_7045), .Q (new_AGEMA_signal_7046) ) ;
    buf_clk new_AGEMA_reg_buffer_4274 ( .C (clk), .D (new_AGEMA_signal_7049), .Q (new_AGEMA_signal_7050) ) ;
    buf_clk new_AGEMA_reg_buffer_4284 ( .C (clk), .D (new_AGEMA_signal_7059), .Q (new_AGEMA_signal_7060) ) ;
    buf_clk new_AGEMA_reg_buffer_4288 ( .C (clk), .D (new_AGEMA_signal_7063), .Q (new_AGEMA_signal_7064) ) ;
    buf_clk new_AGEMA_reg_buffer_4292 ( .C (clk), .D (new_AGEMA_signal_7067), .Q (new_AGEMA_signal_7068) ) ;
    buf_clk new_AGEMA_reg_buffer_4302 ( .C (clk), .D (new_AGEMA_signal_7077), .Q (new_AGEMA_signal_7078) ) ;
    buf_clk new_AGEMA_reg_buffer_4306 ( .C (clk), .D (new_AGEMA_signal_7081), .Q (new_AGEMA_signal_7082) ) ;
    buf_clk new_AGEMA_reg_buffer_4310 ( .C (clk), .D (new_AGEMA_signal_7085), .Q (new_AGEMA_signal_7086) ) ;
    buf_clk new_AGEMA_reg_buffer_4320 ( .C (clk), .D (new_AGEMA_signal_7095), .Q (new_AGEMA_signal_7096) ) ;
    buf_clk new_AGEMA_reg_buffer_4324 ( .C (clk), .D (new_AGEMA_signal_7099), .Q (new_AGEMA_signal_7100) ) ;
    buf_clk new_AGEMA_reg_buffer_4328 ( .C (clk), .D (new_AGEMA_signal_7103), .Q (new_AGEMA_signal_7104) ) ;
    buf_clk new_AGEMA_reg_buffer_4338 ( .C (clk), .D (new_AGEMA_signal_7113), .Q (new_AGEMA_signal_7114) ) ;
    buf_clk new_AGEMA_reg_buffer_4342 ( .C (clk), .D (new_AGEMA_signal_7117), .Q (new_AGEMA_signal_7118) ) ;
    buf_clk new_AGEMA_reg_buffer_4346 ( .C (clk), .D (new_AGEMA_signal_7121), .Q (new_AGEMA_signal_7122) ) ;
    buf_clk new_AGEMA_reg_buffer_4356 ( .C (clk), .D (new_AGEMA_signal_7131), .Q (new_AGEMA_signal_7132) ) ;
    buf_clk new_AGEMA_reg_buffer_4360 ( .C (clk), .D (new_AGEMA_signal_7135), .Q (new_AGEMA_signal_7136) ) ;
    buf_clk new_AGEMA_reg_buffer_4364 ( .C (clk), .D (new_AGEMA_signal_7139), .Q (new_AGEMA_signal_7140) ) ;
    buf_clk new_AGEMA_reg_buffer_4374 ( .C (clk), .D (new_AGEMA_signal_7149), .Q (new_AGEMA_signal_7150) ) ;
    buf_clk new_AGEMA_reg_buffer_4378 ( .C (clk), .D (new_AGEMA_signal_7153), .Q (new_AGEMA_signal_7154) ) ;
    buf_clk new_AGEMA_reg_buffer_4382 ( .C (clk), .D (new_AGEMA_signal_7157), .Q (new_AGEMA_signal_7158) ) ;
    buf_clk new_AGEMA_reg_buffer_4392 ( .C (clk), .D (new_AGEMA_signal_7167), .Q (new_AGEMA_signal_7168) ) ;
    buf_clk new_AGEMA_reg_buffer_4396 ( .C (clk), .D (new_AGEMA_signal_7171), .Q (new_AGEMA_signal_7172) ) ;
    buf_clk new_AGEMA_reg_buffer_4400 ( .C (clk), .D (new_AGEMA_signal_7175), .Q (new_AGEMA_signal_7176) ) ;
    buf_clk new_AGEMA_reg_buffer_4410 ( .C (clk), .D (new_AGEMA_signal_7185), .Q (new_AGEMA_signal_7186) ) ;
    buf_clk new_AGEMA_reg_buffer_4414 ( .C (clk), .D (new_AGEMA_signal_7189), .Q (new_AGEMA_signal_7190) ) ;
    buf_clk new_AGEMA_reg_buffer_4418 ( .C (clk), .D (new_AGEMA_signal_7193), .Q (new_AGEMA_signal_7194) ) ;
    buf_clk new_AGEMA_reg_buffer_4428 ( .C (clk), .D (new_AGEMA_signal_7203), .Q (new_AGEMA_signal_7204) ) ;
    buf_clk new_AGEMA_reg_buffer_4432 ( .C (clk), .D (new_AGEMA_signal_7207), .Q (new_AGEMA_signal_7208) ) ;
    buf_clk new_AGEMA_reg_buffer_4436 ( .C (clk), .D (new_AGEMA_signal_7211), .Q (new_AGEMA_signal_7212) ) ;
    buf_clk new_AGEMA_reg_buffer_4446 ( .C (clk), .D (new_AGEMA_signal_7221), .Q (new_AGEMA_signal_7222) ) ;
    buf_clk new_AGEMA_reg_buffer_4450 ( .C (clk), .D (new_AGEMA_signal_7225), .Q (new_AGEMA_signal_7226) ) ;
    buf_clk new_AGEMA_reg_buffer_4454 ( .C (clk), .D (new_AGEMA_signal_7229), .Q (new_AGEMA_signal_7230) ) ;
    buf_clk new_AGEMA_reg_buffer_4464 ( .C (clk), .D (new_AGEMA_signal_7239), .Q (new_AGEMA_signal_7240) ) ;
    buf_clk new_AGEMA_reg_buffer_4468 ( .C (clk), .D (new_AGEMA_signal_7243), .Q (new_AGEMA_signal_7244) ) ;
    buf_clk new_AGEMA_reg_buffer_4472 ( .C (clk), .D (new_AGEMA_signal_7247), .Q (new_AGEMA_signal_7248) ) ;
    buf_clk new_AGEMA_reg_buffer_4670 ( .C (clk), .D (new_AGEMA_signal_7445), .Q (new_AGEMA_signal_7446) ) ;
    buf_clk new_AGEMA_reg_buffer_4678 ( .C (clk), .D (new_AGEMA_signal_7453), .Q (new_AGEMA_signal_7454) ) ;
    buf_clk new_AGEMA_reg_buffer_4686 ( .C (clk), .D (new_AGEMA_signal_7461), .Q (new_AGEMA_signal_7462) ) ;
    buf_clk new_AGEMA_reg_buffer_4694 ( .C (clk), .D (new_AGEMA_signal_7469), .Q (new_AGEMA_signal_7470) ) ;
    buf_clk new_AGEMA_reg_buffer_4702 ( .C (clk), .D (new_AGEMA_signal_7477), .Q (new_AGEMA_signal_7478) ) ;
    buf_clk new_AGEMA_reg_buffer_4710 ( .C (clk), .D (new_AGEMA_signal_7485), .Q (new_AGEMA_signal_7486) ) ;
    buf_clk new_AGEMA_reg_buffer_4718 ( .C (clk), .D (new_AGEMA_signal_7493), .Q (new_AGEMA_signal_7494) ) ;
    buf_clk new_AGEMA_reg_buffer_4726 ( .C (clk), .D (new_AGEMA_signal_7501), .Q (new_AGEMA_signal_7502) ) ;
    buf_clk new_AGEMA_reg_buffer_4734 ( .C (clk), .D (new_AGEMA_signal_7509), .Q (new_AGEMA_signal_7510) ) ;
    buf_clk new_AGEMA_reg_buffer_4742 ( .C (clk), .D (new_AGEMA_signal_7517), .Q (new_AGEMA_signal_7518) ) ;

    /* cells in depth 5 */
    buf_clk new_AGEMA_reg_buffer_1207 ( .C (clk), .D (new_AGEMA_signal_3982), .Q (new_AGEMA_signal_3983) ) ;
    buf_clk new_AGEMA_reg_buffer_1213 ( .C (clk), .D (new_AGEMA_signal_3988), .Q (new_AGEMA_signal_3989) ) ;
    buf_clk new_AGEMA_reg_buffer_1219 ( .C (clk), .D (new_AGEMA_signal_3994), .Q (new_AGEMA_signal_3995) ) ;
    buf_clk new_AGEMA_reg_buffer_1225 ( .C (clk), .D (new_AGEMA_signal_4000), .Q (new_AGEMA_signal_4001) ) ;
    buf_clk new_AGEMA_reg_buffer_1231 ( .C (clk), .D (new_AGEMA_signal_4006), .Q (new_AGEMA_signal_4007) ) ;
    buf_clk new_AGEMA_reg_buffer_1237 ( .C (clk), .D (new_AGEMA_signal_4012), .Q (new_AGEMA_signal_4013) ) ;
    buf_clk new_AGEMA_reg_buffer_1243 ( .C (clk), .D (new_AGEMA_signal_4018), .Q (new_AGEMA_signal_4019) ) ;
    buf_clk new_AGEMA_reg_buffer_1249 ( .C (clk), .D (new_AGEMA_signal_4024), .Q (new_AGEMA_signal_4025) ) ;
    buf_clk new_AGEMA_reg_buffer_1255 ( .C (clk), .D (new_AGEMA_signal_4030), .Q (new_AGEMA_signal_4031) ) ;
    buf_clk new_AGEMA_reg_buffer_1261 ( .C (clk), .D (new_AGEMA_signal_4036), .Q (new_AGEMA_signal_4037) ) ;
    buf_clk new_AGEMA_reg_buffer_1267 ( .C (clk), .D (new_AGEMA_signal_4042), .Q (new_AGEMA_signal_4043) ) ;
    buf_clk new_AGEMA_reg_buffer_1273 ( .C (clk), .D (new_AGEMA_signal_4048), .Q (new_AGEMA_signal_4049) ) ;
    buf_clk new_AGEMA_reg_buffer_1279 ( .C (clk), .D (new_AGEMA_signal_4054), .Q (new_AGEMA_signal_4055) ) ;
    buf_clk new_AGEMA_reg_buffer_1285 ( .C (clk), .D (new_AGEMA_signal_4060), .Q (new_AGEMA_signal_4061) ) ;
    buf_clk new_AGEMA_reg_buffer_1291 ( .C (clk), .D (new_AGEMA_signal_4066), .Q (new_AGEMA_signal_4067) ) ;
    buf_clk new_AGEMA_reg_buffer_1297 ( .C (clk), .D (new_AGEMA_signal_4072), .Q (new_AGEMA_signal_4073) ) ;
    buf_clk new_AGEMA_reg_buffer_1303 ( .C (clk), .D (new_AGEMA_signal_4078), .Q (new_AGEMA_signal_4079) ) ;
    buf_clk new_AGEMA_reg_buffer_1309 ( .C (clk), .D (new_AGEMA_signal_4084), .Q (new_AGEMA_signal_4085) ) ;
    buf_clk new_AGEMA_reg_buffer_1315 ( .C (clk), .D (new_AGEMA_signal_4090), .Q (new_AGEMA_signal_4091) ) ;
    buf_clk new_AGEMA_reg_buffer_1321 ( .C (clk), .D (new_AGEMA_signal_4096), .Q (new_AGEMA_signal_4097) ) ;
    buf_clk new_AGEMA_reg_buffer_1327 ( .C (clk), .D (new_AGEMA_signal_4102), .Q (new_AGEMA_signal_4103) ) ;
    buf_clk new_AGEMA_reg_buffer_1333 ( .C (clk), .D (new_AGEMA_signal_4108), .Q (new_AGEMA_signal_4109) ) ;
    buf_clk new_AGEMA_reg_buffer_1339 ( .C (clk), .D (new_AGEMA_signal_4114), .Q (new_AGEMA_signal_4115) ) ;
    buf_clk new_AGEMA_reg_buffer_1345 ( .C (clk), .D (new_AGEMA_signal_4120), .Q (new_AGEMA_signal_4121) ) ;
    buf_clk new_AGEMA_reg_buffer_1351 ( .C (clk), .D (new_AGEMA_signal_4126), .Q (new_AGEMA_signal_4127) ) ;
    buf_clk new_AGEMA_reg_buffer_1357 ( .C (clk), .D (new_AGEMA_signal_4132), .Q (new_AGEMA_signal_4133) ) ;
    buf_clk new_AGEMA_reg_buffer_1363 ( .C (clk), .D (new_AGEMA_signal_4138), .Q (new_AGEMA_signal_4139) ) ;
    buf_clk new_AGEMA_reg_buffer_1369 ( .C (clk), .D (new_AGEMA_signal_4144), .Q (new_AGEMA_signal_4145) ) ;
    buf_clk new_AGEMA_reg_buffer_1375 ( .C (clk), .D (new_AGEMA_signal_4150), .Q (new_AGEMA_signal_4151) ) ;
    buf_clk new_AGEMA_reg_buffer_1381 ( .C (clk), .D (new_AGEMA_signal_4156), .Q (new_AGEMA_signal_4157) ) ;
    buf_clk new_AGEMA_reg_buffer_1387 ( .C (clk), .D (new_AGEMA_signal_4162), .Q (new_AGEMA_signal_4163) ) ;
    buf_clk new_AGEMA_reg_buffer_1393 ( .C (clk), .D (new_AGEMA_signal_4168), .Q (new_AGEMA_signal_4169) ) ;
    buf_clk new_AGEMA_reg_buffer_1399 ( .C (clk), .D (new_AGEMA_signal_4174), .Q (new_AGEMA_signal_4175) ) ;
    buf_clk new_AGEMA_reg_buffer_1405 ( .C (clk), .D (new_AGEMA_signal_4180), .Q (new_AGEMA_signal_4181) ) ;
    buf_clk new_AGEMA_reg_buffer_1411 ( .C (clk), .D (new_AGEMA_signal_4186), .Q (new_AGEMA_signal_4187) ) ;
    buf_clk new_AGEMA_reg_buffer_1417 ( .C (clk), .D (new_AGEMA_signal_4192), .Q (new_AGEMA_signal_4193) ) ;
    buf_clk new_AGEMA_reg_buffer_1423 ( .C (clk), .D (new_AGEMA_signal_4198), .Q (new_AGEMA_signal_4199) ) ;
    buf_clk new_AGEMA_reg_buffer_1429 ( .C (clk), .D (new_AGEMA_signal_4204), .Q (new_AGEMA_signal_4205) ) ;
    buf_clk new_AGEMA_reg_buffer_1435 ( .C (clk), .D (new_AGEMA_signal_4210), .Q (new_AGEMA_signal_4211) ) ;
    buf_clk new_AGEMA_reg_buffer_1441 ( .C (clk), .D (new_AGEMA_signal_4216), .Q (new_AGEMA_signal_4217) ) ;
    buf_clk new_AGEMA_reg_buffer_1447 ( .C (clk), .D (new_AGEMA_signal_4222), .Q (new_AGEMA_signal_4223) ) ;
    buf_clk new_AGEMA_reg_buffer_1453 ( .C (clk), .D (new_AGEMA_signal_4228), .Q (new_AGEMA_signal_4229) ) ;
    buf_clk new_AGEMA_reg_buffer_1459 ( .C (clk), .D (new_AGEMA_signal_4234), .Q (new_AGEMA_signal_4235) ) ;
    buf_clk new_AGEMA_reg_buffer_1465 ( .C (clk), .D (new_AGEMA_signal_4240), .Q (new_AGEMA_signal_4241) ) ;
    buf_clk new_AGEMA_reg_buffer_1471 ( .C (clk), .D (new_AGEMA_signal_4246), .Q (new_AGEMA_signal_4247) ) ;
    buf_clk new_AGEMA_reg_buffer_1477 ( .C (clk), .D (new_AGEMA_signal_4252), .Q (new_AGEMA_signal_4253) ) ;
    buf_clk new_AGEMA_reg_buffer_1483 ( .C (clk), .D (new_AGEMA_signal_4258), .Q (new_AGEMA_signal_4259) ) ;
    buf_clk new_AGEMA_reg_buffer_1489 ( .C (clk), .D (new_AGEMA_signal_4264), .Q (new_AGEMA_signal_4265) ) ;
    buf_clk new_AGEMA_reg_buffer_1495 ( .C (clk), .D (new_AGEMA_signal_4270), .Q (new_AGEMA_signal_4271) ) ;
    buf_clk new_AGEMA_reg_buffer_1501 ( .C (clk), .D (new_AGEMA_signal_4276), .Q (new_AGEMA_signal_4277) ) ;
    buf_clk new_AGEMA_reg_buffer_1507 ( .C (clk), .D (new_AGEMA_signal_4282), .Q (new_AGEMA_signal_4283) ) ;
    buf_clk new_AGEMA_reg_buffer_1513 ( .C (clk), .D (new_AGEMA_signal_4288), .Q (new_AGEMA_signal_4289) ) ;
    buf_clk new_AGEMA_reg_buffer_1519 ( .C (clk), .D (new_AGEMA_signal_4294), .Q (new_AGEMA_signal_4295) ) ;
    buf_clk new_AGEMA_reg_buffer_1525 ( .C (clk), .D (new_AGEMA_signal_4300), .Q (new_AGEMA_signal_4301) ) ;
    buf_clk new_AGEMA_reg_buffer_1531 ( .C (clk), .D (new_AGEMA_signal_4306), .Q (new_AGEMA_signal_4307) ) ;
    buf_clk new_AGEMA_reg_buffer_1537 ( .C (clk), .D (new_AGEMA_signal_4312), .Q (new_AGEMA_signal_4313) ) ;
    buf_clk new_AGEMA_reg_buffer_1543 ( .C (clk), .D (new_AGEMA_signal_4318), .Q (new_AGEMA_signal_4319) ) ;
    buf_clk new_AGEMA_reg_buffer_1549 ( .C (clk), .D (new_AGEMA_signal_4324), .Q (new_AGEMA_signal_4325) ) ;
    buf_clk new_AGEMA_reg_buffer_1555 ( .C (clk), .D (new_AGEMA_signal_4330), .Q (new_AGEMA_signal_4331) ) ;
    buf_clk new_AGEMA_reg_buffer_1561 ( .C (clk), .D (new_AGEMA_signal_4336), .Q (new_AGEMA_signal_4337) ) ;
    buf_clk new_AGEMA_reg_buffer_1567 ( .C (clk), .D (new_AGEMA_signal_4342), .Q (new_AGEMA_signal_4343) ) ;
    buf_clk new_AGEMA_reg_buffer_1573 ( .C (clk), .D (new_AGEMA_signal_4348), .Q (new_AGEMA_signal_4349) ) ;
    buf_clk new_AGEMA_reg_buffer_1579 ( .C (clk), .D (new_AGEMA_signal_4354), .Q (new_AGEMA_signal_4355) ) ;
    buf_clk new_AGEMA_reg_buffer_1585 ( .C (clk), .D (new_AGEMA_signal_4360), .Q (new_AGEMA_signal_4361) ) ;
    buf_clk new_AGEMA_reg_buffer_1591 ( .C (clk), .D (new_AGEMA_signal_4366), .Q (new_AGEMA_signal_4367) ) ;
    buf_clk new_AGEMA_reg_buffer_1597 ( .C (clk), .D (new_AGEMA_signal_4372), .Q (new_AGEMA_signal_4373) ) ;
    buf_clk new_AGEMA_reg_buffer_1603 ( .C (clk), .D (new_AGEMA_signal_4378), .Q (new_AGEMA_signal_4379) ) ;
    buf_clk new_AGEMA_reg_buffer_1609 ( .C (clk), .D (new_AGEMA_signal_4384), .Q (new_AGEMA_signal_4385) ) ;
    buf_clk new_AGEMA_reg_buffer_1615 ( .C (clk), .D (new_AGEMA_signal_4390), .Q (new_AGEMA_signal_4391) ) ;
    buf_clk new_AGEMA_reg_buffer_1621 ( .C (clk), .D (new_AGEMA_signal_4396), .Q (new_AGEMA_signal_4397) ) ;
    buf_clk new_AGEMA_reg_buffer_1627 ( .C (clk), .D (new_AGEMA_signal_4402), .Q (new_AGEMA_signal_4403) ) ;
    buf_clk new_AGEMA_reg_buffer_1633 ( .C (clk), .D (new_AGEMA_signal_4408), .Q (new_AGEMA_signal_4409) ) ;
    buf_clk new_AGEMA_reg_buffer_1639 ( .C (clk), .D (new_AGEMA_signal_4414), .Q (new_AGEMA_signal_4415) ) ;
    buf_clk new_AGEMA_reg_buffer_1645 ( .C (clk), .D (new_AGEMA_signal_4420), .Q (new_AGEMA_signal_4421) ) ;
    buf_clk new_AGEMA_reg_buffer_1651 ( .C (clk), .D (new_AGEMA_signal_4426), .Q (new_AGEMA_signal_4427) ) ;
    buf_clk new_AGEMA_reg_buffer_1657 ( .C (clk), .D (new_AGEMA_signal_4432), .Q (new_AGEMA_signal_4433) ) ;
    buf_clk new_AGEMA_reg_buffer_1663 ( .C (clk), .D (new_AGEMA_signal_4438), .Q (new_AGEMA_signal_4439) ) ;
    buf_clk new_AGEMA_reg_buffer_1669 ( .C (clk), .D (new_AGEMA_signal_4444), .Q (new_AGEMA_signal_4445) ) ;
    buf_clk new_AGEMA_reg_buffer_1675 ( .C (clk), .D (new_AGEMA_signal_4450), .Q (new_AGEMA_signal_4451) ) ;
    buf_clk new_AGEMA_reg_buffer_1681 ( .C (clk), .D (new_AGEMA_signal_4456), .Q (new_AGEMA_signal_4457) ) ;
    buf_clk new_AGEMA_reg_buffer_1687 ( .C (clk), .D (new_AGEMA_signal_4462), .Q (new_AGEMA_signal_4463) ) ;
    buf_clk new_AGEMA_reg_buffer_1693 ( .C (clk), .D (new_AGEMA_signal_4468), .Q (new_AGEMA_signal_4469) ) ;
    buf_clk new_AGEMA_reg_buffer_1699 ( .C (clk), .D (new_AGEMA_signal_4474), .Q (new_AGEMA_signal_4475) ) ;
    buf_clk new_AGEMA_reg_buffer_1705 ( .C (clk), .D (new_AGEMA_signal_4480), .Q (new_AGEMA_signal_4481) ) ;
    buf_clk new_AGEMA_reg_buffer_1711 ( .C (clk), .D (new_AGEMA_signal_4486), .Q (new_AGEMA_signal_4487) ) ;
    buf_clk new_AGEMA_reg_buffer_1717 ( .C (clk), .D (new_AGEMA_signal_4492), .Q (new_AGEMA_signal_4493) ) ;
    buf_clk new_AGEMA_reg_buffer_1723 ( .C (clk), .D (new_AGEMA_signal_4498), .Q (new_AGEMA_signal_4499) ) ;
    buf_clk new_AGEMA_reg_buffer_1729 ( .C (clk), .D (new_AGEMA_signal_4504), .Q (new_AGEMA_signal_4505) ) ;
    buf_clk new_AGEMA_reg_buffer_1735 ( .C (clk), .D (new_AGEMA_signal_4510), .Q (new_AGEMA_signal_4511) ) ;
    buf_clk new_AGEMA_reg_buffer_1741 ( .C (clk), .D (new_AGEMA_signal_4516), .Q (new_AGEMA_signal_4517) ) ;
    buf_clk new_AGEMA_reg_buffer_1747 ( .C (clk), .D (new_AGEMA_signal_4522), .Q (new_AGEMA_signal_4523) ) ;
    buf_clk new_AGEMA_reg_buffer_1753 ( .C (clk), .D (new_AGEMA_signal_4528), .Q (new_AGEMA_signal_4529) ) ;
    buf_clk new_AGEMA_reg_buffer_1759 ( .C (clk), .D (new_AGEMA_signal_4534), .Q (new_AGEMA_signal_4535) ) ;
    buf_clk new_AGEMA_reg_buffer_1765 ( .C (clk), .D (new_AGEMA_signal_4540), .Q (new_AGEMA_signal_4541) ) ;
    buf_clk new_AGEMA_reg_buffer_1771 ( .C (clk), .D (new_AGEMA_signal_4546), .Q (new_AGEMA_signal_4547) ) ;
    buf_clk new_AGEMA_reg_buffer_1777 ( .C (clk), .D (new_AGEMA_signal_4552), .Q (new_AGEMA_signal_4553) ) ;
    buf_clk new_AGEMA_reg_buffer_1783 ( .C (clk), .D (new_AGEMA_signal_4558), .Q (new_AGEMA_signal_4559) ) ;
    buf_clk new_AGEMA_reg_buffer_1789 ( .C (clk), .D (new_AGEMA_signal_4564), .Q (new_AGEMA_signal_4565) ) ;
    buf_clk new_AGEMA_reg_buffer_1795 ( .C (clk), .D (new_AGEMA_signal_4570), .Q (new_AGEMA_signal_4571) ) ;
    buf_clk new_AGEMA_reg_buffer_1801 ( .C (clk), .D (new_AGEMA_signal_4576), .Q (new_AGEMA_signal_4577) ) ;
    buf_clk new_AGEMA_reg_buffer_1807 ( .C (clk), .D (new_AGEMA_signal_4582), .Q (new_AGEMA_signal_4583) ) ;
    buf_clk new_AGEMA_reg_buffer_1813 ( .C (clk), .D (new_AGEMA_signal_4588), .Q (new_AGEMA_signal_4589) ) ;
    buf_clk new_AGEMA_reg_buffer_1819 ( .C (clk), .D (new_AGEMA_signal_4594), .Q (new_AGEMA_signal_4595) ) ;
    buf_clk new_AGEMA_reg_buffer_1825 ( .C (clk), .D (new_AGEMA_signal_4600), .Q (new_AGEMA_signal_4601) ) ;
    buf_clk new_AGEMA_reg_buffer_1831 ( .C (clk), .D (new_AGEMA_signal_4606), .Q (new_AGEMA_signal_4607) ) ;
    buf_clk new_AGEMA_reg_buffer_1837 ( .C (clk), .D (new_AGEMA_signal_4612), .Q (new_AGEMA_signal_4613) ) ;
    buf_clk new_AGEMA_reg_buffer_1843 ( .C (clk), .D (new_AGEMA_signal_4618), .Q (new_AGEMA_signal_4619) ) ;
    buf_clk new_AGEMA_reg_buffer_1849 ( .C (clk), .D (new_AGEMA_signal_4624), .Q (new_AGEMA_signal_4625) ) ;
    buf_clk new_AGEMA_reg_buffer_1855 ( .C (clk), .D (new_AGEMA_signal_4630), .Q (new_AGEMA_signal_4631) ) ;
    buf_clk new_AGEMA_reg_buffer_1861 ( .C (clk), .D (new_AGEMA_signal_4636), .Q (new_AGEMA_signal_4637) ) ;
    buf_clk new_AGEMA_reg_buffer_1867 ( .C (clk), .D (new_AGEMA_signal_4642), .Q (new_AGEMA_signal_4643) ) ;
    buf_clk new_AGEMA_reg_buffer_1873 ( .C (clk), .D (new_AGEMA_signal_4648), .Q (new_AGEMA_signal_4649) ) ;
    buf_clk new_AGEMA_reg_buffer_1879 ( .C (clk), .D (new_AGEMA_signal_4654), .Q (new_AGEMA_signal_4655) ) ;
    buf_clk new_AGEMA_reg_buffer_1885 ( .C (clk), .D (new_AGEMA_signal_4660), .Q (new_AGEMA_signal_4661) ) ;
    buf_clk new_AGEMA_reg_buffer_1891 ( .C (clk), .D (new_AGEMA_signal_4666), .Q (new_AGEMA_signal_4667) ) ;
    buf_clk new_AGEMA_reg_buffer_1897 ( .C (clk), .D (new_AGEMA_signal_4672), .Q (new_AGEMA_signal_4673) ) ;
    buf_clk new_AGEMA_reg_buffer_1903 ( .C (clk), .D (new_AGEMA_signal_4678), .Q (new_AGEMA_signal_4679) ) ;
    buf_clk new_AGEMA_reg_buffer_1909 ( .C (clk), .D (new_AGEMA_signal_4684), .Q (new_AGEMA_signal_4685) ) ;
    buf_clk new_AGEMA_reg_buffer_1915 ( .C (clk), .D (new_AGEMA_signal_4690), .Q (new_AGEMA_signal_4691) ) ;
    buf_clk new_AGEMA_reg_buffer_1921 ( .C (clk), .D (new_AGEMA_signal_4696), .Q (new_AGEMA_signal_4697) ) ;
    buf_clk new_AGEMA_reg_buffer_1927 ( .C (clk), .D (new_AGEMA_signal_4702), .Q (new_AGEMA_signal_4703) ) ;
    buf_clk new_AGEMA_reg_buffer_1933 ( .C (clk), .D (new_AGEMA_signal_4708), .Q (new_AGEMA_signal_4709) ) ;
    buf_clk new_AGEMA_reg_buffer_1939 ( .C (clk), .D (new_AGEMA_signal_4714), .Q (new_AGEMA_signal_4715) ) ;
    buf_clk new_AGEMA_reg_buffer_1945 ( .C (clk), .D (new_AGEMA_signal_4720), .Q (new_AGEMA_signal_4721) ) ;
    buf_clk new_AGEMA_reg_buffer_1951 ( .C (clk), .D (new_AGEMA_signal_4726), .Q (new_AGEMA_signal_4727) ) ;
    buf_clk new_AGEMA_reg_buffer_1957 ( .C (clk), .D (new_AGEMA_signal_4732), .Q (new_AGEMA_signal_4733) ) ;
    buf_clk new_AGEMA_reg_buffer_1963 ( .C (clk), .D (new_AGEMA_signal_4738), .Q (new_AGEMA_signal_4739) ) ;
    buf_clk new_AGEMA_reg_buffer_1969 ( .C (clk), .D (new_AGEMA_signal_4744), .Q (new_AGEMA_signal_4745) ) ;
    buf_clk new_AGEMA_reg_buffer_1975 ( .C (clk), .D (new_AGEMA_signal_4750), .Q (new_AGEMA_signal_4751) ) ;
    buf_clk new_AGEMA_reg_buffer_1981 ( .C (clk), .D (new_AGEMA_signal_4756), .Q (new_AGEMA_signal_4757) ) ;
    buf_clk new_AGEMA_reg_buffer_1987 ( .C (clk), .D (new_AGEMA_signal_4762), .Q (new_AGEMA_signal_4763) ) ;
    buf_clk new_AGEMA_reg_buffer_1993 ( .C (clk), .D (new_AGEMA_signal_4768), .Q (new_AGEMA_signal_4769) ) ;
    buf_clk new_AGEMA_reg_buffer_1999 ( .C (clk), .D (new_AGEMA_signal_4774), .Q (new_AGEMA_signal_4775) ) ;
    buf_clk new_AGEMA_reg_buffer_2005 ( .C (clk), .D (new_AGEMA_signal_4780), .Q (new_AGEMA_signal_4781) ) ;
    buf_clk new_AGEMA_reg_buffer_2011 ( .C (clk), .D (new_AGEMA_signal_4786), .Q (new_AGEMA_signal_4787) ) ;
    buf_clk new_AGEMA_reg_buffer_2017 ( .C (clk), .D (new_AGEMA_signal_4792), .Q (new_AGEMA_signal_4793) ) ;
    buf_clk new_AGEMA_reg_buffer_2023 ( .C (clk), .D (new_AGEMA_signal_4798), .Q (new_AGEMA_signal_4799) ) ;
    buf_clk new_AGEMA_reg_buffer_2029 ( .C (clk), .D (new_AGEMA_signal_4804), .Q (new_AGEMA_signal_4805) ) ;
    buf_clk new_AGEMA_reg_buffer_2035 ( .C (clk), .D (new_AGEMA_signal_4810), .Q (new_AGEMA_signal_4811) ) ;
    buf_clk new_AGEMA_reg_buffer_2041 ( .C (clk), .D (new_AGEMA_signal_4816), .Q (new_AGEMA_signal_4817) ) ;
    buf_clk new_AGEMA_reg_buffer_2047 ( .C (clk), .D (new_AGEMA_signal_4822), .Q (new_AGEMA_signal_4823) ) ;
    buf_clk new_AGEMA_reg_buffer_2053 ( .C (clk), .D (new_AGEMA_signal_4828), .Q (new_AGEMA_signal_4829) ) ;
    buf_clk new_AGEMA_reg_buffer_2059 ( .C (clk), .D (new_AGEMA_signal_4834), .Q (new_AGEMA_signal_4835) ) ;
    buf_clk new_AGEMA_reg_buffer_2065 ( .C (clk), .D (new_AGEMA_signal_4840), .Q (new_AGEMA_signal_4841) ) ;
    buf_clk new_AGEMA_reg_buffer_2071 ( .C (clk), .D (new_AGEMA_signal_4846), .Q (new_AGEMA_signal_4847) ) ;
    buf_clk new_AGEMA_reg_buffer_2077 ( .C (clk), .D (new_AGEMA_signal_4852), .Q (new_AGEMA_signal_4853) ) ;
    buf_clk new_AGEMA_reg_buffer_2083 ( .C (clk), .D (new_AGEMA_signal_4858), .Q (new_AGEMA_signal_4859) ) ;
    buf_clk new_AGEMA_reg_buffer_2089 ( .C (clk), .D (new_AGEMA_signal_4864), .Q (new_AGEMA_signal_4865) ) ;
    buf_clk new_AGEMA_reg_buffer_2095 ( .C (clk), .D (new_AGEMA_signal_4870), .Q (new_AGEMA_signal_4871) ) ;
    buf_clk new_AGEMA_reg_buffer_2101 ( .C (clk), .D (new_AGEMA_signal_4876), .Q (new_AGEMA_signal_4877) ) ;
    buf_clk new_AGEMA_reg_buffer_2107 ( .C (clk), .D (new_AGEMA_signal_4882), .Q (new_AGEMA_signal_4883) ) ;
    buf_clk new_AGEMA_reg_buffer_2113 ( .C (clk), .D (new_AGEMA_signal_4888), .Q (new_AGEMA_signal_4889) ) ;
    buf_clk new_AGEMA_reg_buffer_2119 ( .C (clk), .D (new_AGEMA_signal_4894), .Q (new_AGEMA_signal_4895) ) ;
    buf_clk new_AGEMA_reg_buffer_2125 ( .C (clk), .D (new_AGEMA_signal_4900), .Q (new_AGEMA_signal_4901) ) ;
    buf_clk new_AGEMA_reg_buffer_2131 ( .C (clk), .D (new_AGEMA_signal_4906), .Q (new_AGEMA_signal_4907) ) ;
    buf_clk new_AGEMA_reg_buffer_2137 ( .C (clk), .D (new_AGEMA_signal_4912), .Q (new_AGEMA_signal_4913) ) ;
    buf_clk new_AGEMA_reg_buffer_2143 ( .C (clk), .D (new_AGEMA_signal_4918), .Q (new_AGEMA_signal_4919) ) ;
    buf_clk new_AGEMA_reg_buffer_2149 ( .C (clk), .D (new_AGEMA_signal_4924), .Q (new_AGEMA_signal_4925) ) ;
    buf_clk new_AGEMA_reg_buffer_2155 ( .C (clk), .D (new_AGEMA_signal_4930), .Q (new_AGEMA_signal_4931) ) ;
    buf_clk new_AGEMA_reg_buffer_2161 ( .C (clk), .D (new_AGEMA_signal_4936), .Q (new_AGEMA_signal_4937) ) ;
    buf_clk new_AGEMA_reg_buffer_2167 ( .C (clk), .D (new_AGEMA_signal_4942), .Q (new_AGEMA_signal_4943) ) ;
    buf_clk new_AGEMA_reg_buffer_2173 ( .C (clk), .D (new_AGEMA_signal_4948), .Q (new_AGEMA_signal_4949) ) ;
    buf_clk new_AGEMA_reg_buffer_2179 ( .C (clk), .D (new_AGEMA_signal_4954), .Q (new_AGEMA_signal_4955) ) ;
    buf_clk new_AGEMA_reg_buffer_2185 ( .C (clk), .D (new_AGEMA_signal_4960), .Q (new_AGEMA_signal_4961) ) ;
    buf_clk new_AGEMA_reg_buffer_2191 ( .C (clk), .D (new_AGEMA_signal_4966), .Q (new_AGEMA_signal_4967) ) ;
    buf_clk new_AGEMA_reg_buffer_2197 ( .C (clk), .D (new_AGEMA_signal_4972), .Q (new_AGEMA_signal_4973) ) ;
    buf_clk new_AGEMA_reg_buffer_2203 ( .C (clk), .D (new_AGEMA_signal_4978), .Q (new_AGEMA_signal_4979) ) ;
    buf_clk new_AGEMA_reg_buffer_2209 ( .C (clk), .D (new_AGEMA_signal_4984), .Q (new_AGEMA_signal_4985) ) ;
    buf_clk new_AGEMA_reg_buffer_2215 ( .C (clk), .D (new_AGEMA_signal_4990), .Q (new_AGEMA_signal_4991) ) ;
    buf_clk new_AGEMA_reg_buffer_2221 ( .C (clk), .D (new_AGEMA_signal_4996), .Q (new_AGEMA_signal_4997) ) ;
    buf_clk new_AGEMA_reg_buffer_2227 ( .C (clk), .D (new_AGEMA_signal_5002), .Q (new_AGEMA_signal_5003) ) ;
    buf_clk new_AGEMA_reg_buffer_2233 ( .C (clk), .D (new_AGEMA_signal_5008), .Q (new_AGEMA_signal_5009) ) ;
    buf_clk new_AGEMA_reg_buffer_2239 ( .C (clk), .D (new_AGEMA_signal_5014), .Q (new_AGEMA_signal_5015) ) ;
    buf_clk new_AGEMA_reg_buffer_2245 ( .C (clk), .D (new_AGEMA_signal_5020), .Q (new_AGEMA_signal_5021) ) ;
    buf_clk new_AGEMA_reg_buffer_2251 ( .C (clk), .D (new_AGEMA_signal_5026), .Q (new_AGEMA_signal_5027) ) ;
    buf_clk new_AGEMA_reg_buffer_2257 ( .C (clk), .D (new_AGEMA_signal_5032), .Q (new_AGEMA_signal_5033) ) ;
    buf_clk new_AGEMA_reg_buffer_2263 ( .C (clk), .D (new_AGEMA_signal_5038), .Q (new_AGEMA_signal_5039) ) ;
    buf_clk new_AGEMA_reg_buffer_2269 ( .C (clk), .D (new_AGEMA_signal_5044), .Q (new_AGEMA_signal_5045) ) ;
    buf_clk new_AGEMA_reg_buffer_2275 ( .C (clk), .D (new_AGEMA_signal_5050), .Q (new_AGEMA_signal_5051) ) ;
    buf_clk new_AGEMA_reg_buffer_2281 ( .C (clk), .D (new_AGEMA_signal_5056), .Q (new_AGEMA_signal_5057) ) ;
    buf_clk new_AGEMA_reg_buffer_2287 ( .C (clk), .D (new_AGEMA_signal_5062), .Q (new_AGEMA_signal_5063) ) ;
    buf_clk new_AGEMA_reg_buffer_2293 ( .C (clk), .D (new_AGEMA_signal_5068), .Q (new_AGEMA_signal_5069) ) ;
    buf_clk new_AGEMA_reg_buffer_2299 ( .C (clk), .D (new_AGEMA_signal_5074), .Q (new_AGEMA_signal_5075) ) ;
    buf_clk new_AGEMA_reg_buffer_2305 ( .C (clk), .D (new_AGEMA_signal_5080), .Q (new_AGEMA_signal_5081) ) ;
    buf_clk new_AGEMA_reg_buffer_2311 ( .C (clk), .D (new_AGEMA_signal_5086), .Q (new_AGEMA_signal_5087) ) ;
    buf_clk new_AGEMA_reg_buffer_2317 ( .C (clk), .D (new_AGEMA_signal_5092), .Q (new_AGEMA_signal_5093) ) ;
    buf_clk new_AGEMA_reg_buffer_2323 ( .C (clk), .D (new_AGEMA_signal_5098), .Q (new_AGEMA_signal_5099) ) ;
    buf_clk new_AGEMA_reg_buffer_2329 ( .C (clk), .D (new_AGEMA_signal_5104), .Q (new_AGEMA_signal_5105) ) ;
    buf_clk new_AGEMA_reg_buffer_2335 ( .C (clk), .D (new_AGEMA_signal_5110), .Q (new_AGEMA_signal_5111) ) ;
    buf_clk new_AGEMA_reg_buffer_2341 ( .C (clk), .D (new_AGEMA_signal_5116), .Q (new_AGEMA_signal_5117) ) ;
    buf_clk new_AGEMA_reg_buffer_2347 ( .C (clk), .D (new_AGEMA_signal_5122), .Q (new_AGEMA_signal_5123) ) ;
    buf_clk new_AGEMA_reg_buffer_2353 ( .C (clk), .D (new_AGEMA_signal_5128), .Q (new_AGEMA_signal_5129) ) ;
    buf_clk new_AGEMA_reg_buffer_2359 ( .C (clk), .D (new_AGEMA_signal_5134), .Q (new_AGEMA_signal_5135) ) ;
    buf_clk new_AGEMA_reg_buffer_2655 ( .C (clk), .D (new_AGEMA_signal_5430), .Q (new_AGEMA_signal_5431) ) ;
    buf_clk new_AGEMA_reg_buffer_2663 ( .C (clk), .D (new_AGEMA_signal_5438), .Q (new_AGEMA_signal_5439) ) ;
    buf_clk new_AGEMA_reg_buffer_2671 ( .C (clk), .D (new_AGEMA_signal_5446), .Q (new_AGEMA_signal_5447) ) ;
    buf_clk new_AGEMA_reg_buffer_2679 ( .C (clk), .D (new_AGEMA_signal_5454), .Q (new_AGEMA_signal_5455) ) ;
    buf_clk new_AGEMA_reg_buffer_2687 ( .C (clk), .D (new_AGEMA_signal_5462), .Q (new_AGEMA_signal_5463) ) ;
    buf_clk new_AGEMA_reg_buffer_2695 ( .C (clk), .D (new_AGEMA_signal_5470), .Q (new_AGEMA_signal_5471) ) ;
    buf_clk new_AGEMA_reg_buffer_2703 ( .C (clk), .D (new_AGEMA_signal_5478), .Q (new_AGEMA_signal_5479) ) ;
    buf_clk new_AGEMA_reg_buffer_2711 ( .C (clk), .D (new_AGEMA_signal_5486), .Q (new_AGEMA_signal_5487) ) ;
    buf_clk new_AGEMA_reg_buffer_2719 ( .C (clk), .D (new_AGEMA_signal_5494), .Q (new_AGEMA_signal_5495) ) ;
    buf_clk new_AGEMA_reg_buffer_2727 ( .C (clk), .D (new_AGEMA_signal_5502), .Q (new_AGEMA_signal_5503) ) ;
    buf_clk new_AGEMA_reg_buffer_2735 ( .C (clk), .D (new_AGEMA_signal_5510), .Q (new_AGEMA_signal_5511) ) ;
    buf_clk new_AGEMA_reg_buffer_2743 ( .C (clk), .D (new_AGEMA_signal_5518), .Q (new_AGEMA_signal_5519) ) ;
    buf_clk new_AGEMA_reg_buffer_2751 ( .C (clk), .D (new_AGEMA_signal_5526), .Q (new_AGEMA_signal_5527) ) ;
    buf_clk new_AGEMA_reg_buffer_2759 ( .C (clk), .D (new_AGEMA_signal_5534), .Q (new_AGEMA_signal_5535) ) ;
    buf_clk new_AGEMA_reg_buffer_2767 ( .C (clk), .D (new_AGEMA_signal_5542), .Q (new_AGEMA_signal_5543) ) ;
    buf_clk new_AGEMA_reg_buffer_2775 ( .C (clk), .D (new_AGEMA_signal_5550), .Q (new_AGEMA_signal_5551) ) ;
    buf_clk new_AGEMA_reg_buffer_2783 ( .C (clk), .D (new_AGEMA_signal_5558), .Q (new_AGEMA_signal_5559) ) ;
    buf_clk new_AGEMA_reg_buffer_2791 ( .C (clk), .D (new_AGEMA_signal_5566), .Q (new_AGEMA_signal_5567) ) ;
    buf_clk new_AGEMA_reg_buffer_2799 ( .C (clk), .D (new_AGEMA_signal_5574), .Q (new_AGEMA_signal_5575) ) ;
    buf_clk new_AGEMA_reg_buffer_2807 ( .C (clk), .D (new_AGEMA_signal_5582), .Q (new_AGEMA_signal_5583) ) ;
    buf_clk new_AGEMA_reg_buffer_2815 ( .C (clk), .D (new_AGEMA_signal_5590), .Q (new_AGEMA_signal_5591) ) ;
    buf_clk new_AGEMA_reg_buffer_2823 ( .C (clk), .D (new_AGEMA_signal_5598), .Q (new_AGEMA_signal_5599) ) ;
    buf_clk new_AGEMA_reg_buffer_2831 ( .C (clk), .D (new_AGEMA_signal_5606), .Q (new_AGEMA_signal_5607) ) ;
    buf_clk new_AGEMA_reg_buffer_2839 ( .C (clk), .D (new_AGEMA_signal_5614), .Q (new_AGEMA_signal_5615) ) ;
    buf_clk new_AGEMA_reg_buffer_2847 ( .C (clk), .D (new_AGEMA_signal_5622), .Q (new_AGEMA_signal_5623) ) ;
    buf_clk new_AGEMA_reg_buffer_2855 ( .C (clk), .D (new_AGEMA_signal_5630), .Q (new_AGEMA_signal_5631) ) ;
    buf_clk new_AGEMA_reg_buffer_2863 ( .C (clk), .D (new_AGEMA_signal_5638), .Q (new_AGEMA_signal_5639) ) ;
    buf_clk new_AGEMA_reg_buffer_2871 ( .C (clk), .D (new_AGEMA_signal_5646), .Q (new_AGEMA_signal_5647) ) ;
    buf_clk new_AGEMA_reg_buffer_2879 ( .C (clk), .D (new_AGEMA_signal_5654), .Q (new_AGEMA_signal_5655) ) ;
    buf_clk new_AGEMA_reg_buffer_2887 ( .C (clk), .D (new_AGEMA_signal_5662), .Q (new_AGEMA_signal_5663) ) ;
    buf_clk new_AGEMA_reg_buffer_2895 ( .C (clk), .D (new_AGEMA_signal_5670), .Q (new_AGEMA_signal_5671) ) ;
    buf_clk new_AGEMA_reg_buffer_2903 ( .C (clk), .D (new_AGEMA_signal_5678), .Q (new_AGEMA_signal_5679) ) ;
    buf_clk new_AGEMA_reg_buffer_2911 ( .C (clk), .D (new_AGEMA_signal_5686), .Q (new_AGEMA_signal_5687) ) ;
    buf_clk new_AGEMA_reg_buffer_2919 ( .C (clk), .D (new_AGEMA_signal_5694), .Q (new_AGEMA_signal_5695) ) ;
    buf_clk new_AGEMA_reg_buffer_2927 ( .C (clk), .D (new_AGEMA_signal_5702), .Q (new_AGEMA_signal_5703) ) ;
    buf_clk new_AGEMA_reg_buffer_2935 ( .C (clk), .D (new_AGEMA_signal_5710), .Q (new_AGEMA_signal_5711) ) ;
    buf_clk new_AGEMA_reg_buffer_2943 ( .C (clk), .D (new_AGEMA_signal_5718), .Q (new_AGEMA_signal_5719) ) ;
    buf_clk new_AGEMA_reg_buffer_2951 ( .C (clk), .D (new_AGEMA_signal_5726), .Q (new_AGEMA_signal_5727) ) ;
    buf_clk new_AGEMA_reg_buffer_2959 ( .C (clk), .D (new_AGEMA_signal_5734), .Q (new_AGEMA_signal_5735) ) ;
    buf_clk new_AGEMA_reg_buffer_2967 ( .C (clk), .D (new_AGEMA_signal_5742), .Q (new_AGEMA_signal_5743) ) ;
    buf_clk new_AGEMA_reg_buffer_2975 ( .C (clk), .D (new_AGEMA_signal_5750), .Q (new_AGEMA_signal_5751) ) ;
    buf_clk new_AGEMA_reg_buffer_2983 ( .C (clk), .D (new_AGEMA_signal_5758), .Q (new_AGEMA_signal_5759) ) ;
    buf_clk new_AGEMA_reg_buffer_2991 ( .C (clk), .D (new_AGEMA_signal_5766), .Q (new_AGEMA_signal_5767) ) ;
    buf_clk new_AGEMA_reg_buffer_2999 ( .C (clk), .D (new_AGEMA_signal_5774), .Q (new_AGEMA_signal_5775) ) ;
    buf_clk new_AGEMA_reg_buffer_3007 ( .C (clk), .D (new_AGEMA_signal_5782), .Q (new_AGEMA_signal_5783) ) ;
    buf_clk new_AGEMA_reg_buffer_3015 ( .C (clk), .D (new_AGEMA_signal_5790), .Q (new_AGEMA_signal_5791) ) ;
    buf_clk new_AGEMA_reg_buffer_3023 ( .C (clk), .D (new_AGEMA_signal_5798), .Q (new_AGEMA_signal_5799) ) ;
    buf_clk new_AGEMA_reg_buffer_3031 ( .C (clk), .D (new_AGEMA_signal_5806), .Q (new_AGEMA_signal_5807) ) ;
    buf_clk new_AGEMA_reg_buffer_3039 ( .C (clk), .D (new_AGEMA_signal_5814), .Q (new_AGEMA_signal_5815) ) ;
    buf_clk new_AGEMA_reg_buffer_3047 ( .C (clk), .D (new_AGEMA_signal_5822), .Q (new_AGEMA_signal_5823) ) ;
    buf_clk new_AGEMA_reg_buffer_3055 ( .C (clk), .D (new_AGEMA_signal_5830), .Q (new_AGEMA_signal_5831) ) ;
    buf_clk new_AGEMA_reg_buffer_3063 ( .C (clk), .D (new_AGEMA_signal_5838), .Q (new_AGEMA_signal_5839) ) ;
    buf_clk new_AGEMA_reg_buffer_3071 ( .C (clk), .D (new_AGEMA_signal_5846), .Q (new_AGEMA_signal_5847) ) ;
    buf_clk new_AGEMA_reg_buffer_3079 ( .C (clk), .D (new_AGEMA_signal_5854), .Q (new_AGEMA_signal_5855) ) ;
    buf_clk new_AGEMA_reg_buffer_3087 ( .C (clk), .D (new_AGEMA_signal_5862), .Q (new_AGEMA_signal_5863) ) ;
    buf_clk new_AGEMA_reg_buffer_3095 ( .C (clk), .D (new_AGEMA_signal_5870), .Q (new_AGEMA_signal_5871) ) ;
    buf_clk new_AGEMA_reg_buffer_3103 ( .C (clk), .D (new_AGEMA_signal_5878), .Q (new_AGEMA_signal_5879) ) ;
    buf_clk new_AGEMA_reg_buffer_3111 ( .C (clk), .D (new_AGEMA_signal_5886), .Q (new_AGEMA_signal_5887) ) ;
    buf_clk new_AGEMA_reg_buffer_3119 ( .C (clk), .D (new_AGEMA_signal_5894), .Q (new_AGEMA_signal_5895) ) ;
    buf_clk new_AGEMA_reg_buffer_3127 ( .C (clk), .D (new_AGEMA_signal_5902), .Q (new_AGEMA_signal_5903) ) ;
    buf_clk new_AGEMA_reg_buffer_3135 ( .C (clk), .D (new_AGEMA_signal_5910), .Q (new_AGEMA_signal_5911) ) ;
    buf_clk new_AGEMA_reg_buffer_3143 ( .C (clk), .D (new_AGEMA_signal_5918), .Q (new_AGEMA_signal_5919) ) ;
    buf_clk new_AGEMA_reg_buffer_3151 ( .C (clk), .D (new_AGEMA_signal_5926), .Q (new_AGEMA_signal_5927) ) ;
    buf_clk new_AGEMA_reg_buffer_3159 ( .C (clk), .D (new_AGEMA_signal_5934), .Q (new_AGEMA_signal_5935) ) ;
    buf_clk new_AGEMA_reg_buffer_3167 ( .C (clk), .D (new_AGEMA_signal_5942), .Q (new_AGEMA_signal_5943) ) ;
    buf_clk new_AGEMA_reg_buffer_3175 ( .C (clk), .D (new_AGEMA_signal_5950), .Q (new_AGEMA_signal_5951) ) ;
    buf_clk new_AGEMA_reg_buffer_3183 ( .C (clk), .D (new_AGEMA_signal_5958), .Q (new_AGEMA_signal_5959) ) ;
    buf_clk new_AGEMA_reg_buffer_3191 ( .C (clk), .D (new_AGEMA_signal_5966), .Q (new_AGEMA_signal_5967) ) ;
    buf_clk new_AGEMA_reg_buffer_3199 ( .C (clk), .D (new_AGEMA_signal_5974), .Q (new_AGEMA_signal_5975) ) ;
    buf_clk new_AGEMA_reg_buffer_3207 ( .C (clk), .D (new_AGEMA_signal_5982), .Q (new_AGEMA_signal_5983) ) ;
    buf_clk new_AGEMA_reg_buffer_3215 ( .C (clk), .D (new_AGEMA_signal_5990), .Q (new_AGEMA_signal_5991) ) ;
    buf_clk new_AGEMA_reg_buffer_3223 ( .C (clk), .D (new_AGEMA_signal_5998), .Q (new_AGEMA_signal_5999) ) ;
    buf_clk new_AGEMA_reg_buffer_3231 ( .C (clk), .D (new_AGEMA_signal_6006), .Q (new_AGEMA_signal_6007) ) ;
    buf_clk new_AGEMA_reg_buffer_3239 ( .C (clk), .D (new_AGEMA_signal_6014), .Q (new_AGEMA_signal_6015) ) ;
    buf_clk new_AGEMA_reg_buffer_3247 ( .C (clk), .D (new_AGEMA_signal_6022), .Q (new_AGEMA_signal_6023) ) ;
    buf_clk new_AGEMA_reg_buffer_3255 ( .C (clk), .D (new_AGEMA_signal_6030), .Q (new_AGEMA_signal_6031) ) ;
    buf_clk new_AGEMA_reg_buffer_3263 ( .C (clk), .D (new_AGEMA_signal_6038), .Q (new_AGEMA_signal_6039) ) ;
    buf_clk new_AGEMA_reg_buffer_3271 ( .C (clk), .D (new_AGEMA_signal_6046), .Q (new_AGEMA_signal_6047) ) ;
    buf_clk new_AGEMA_reg_buffer_3279 ( .C (clk), .D (new_AGEMA_signal_6054), .Q (new_AGEMA_signal_6055) ) ;
    buf_clk new_AGEMA_reg_buffer_3287 ( .C (clk), .D (new_AGEMA_signal_6062), .Q (new_AGEMA_signal_6063) ) ;
    buf_clk new_AGEMA_reg_buffer_3295 ( .C (clk), .D (new_AGEMA_signal_6070), .Q (new_AGEMA_signal_6071) ) ;
    buf_clk new_AGEMA_reg_buffer_3303 ( .C (clk), .D (new_AGEMA_signal_6078), .Q (new_AGEMA_signal_6079) ) ;
    buf_clk new_AGEMA_reg_buffer_3311 ( .C (clk), .D (new_AGEMA_signal_6086), .Q (new_AGEMA_signal_6087) ) ;
    buf_clk new_AGEMA_reg_buffer_3319 ( .C (clk), .D (new_AGEMA_signal_6094), .Q (new_AGEMA_signal_6095) ) ;
    buf_clk new_AGEMA_reg_buffer_3327 ( .C (clk), .D (new_AGEMA_signal_6102), .Q (new_AGEMA_signal_6103) ) ;
    buf_clk new_AGEMA_reg_buffer_3335 ( .C (clk), .D (new_AGEMA_signal_6110), .Q (new_AGEMA_signal_6111) ) ;
    buf_clk new_AGEMA_reg_buffer_3343 ( .C (clk), .D (new_AGEMA_signal_6118), .Q (new_AGEMA_signal_6119) ) ;
    buf_clk new_AGEMA_reg_buffer_3351 ( .C (clk), .D (new_AGEMA_signal_6126), .Q (new_AGEMA_signal_6127) ) ;
    buf_clk new_AGEMA_reg_buffer_3359 ( .C (clk), .D (new_AGEMA_signal_6134), .Q (new_AGEMA_signal_6135) ) ;
    buf_clk new_AGEMA_reg_buffer_3367 ( .C (clk), .D (new_AGEMA_signal_6142), .Q (new_AGEMA_signal_6143) ) ;
    buf_clk new_AGEMA_reg_buffer_3375 ( .C (clk), .D (new_AGEMA_signal_6150), .Q (new_AGEMA_signal_6151) ) ;
    buf_clk new_AGEMA_reg_buffer_3383 ( .C (clk), .D (new_AGEMA_signal_6158), .Q (new_AGEMA_signal_6159) ) ;
    buf_clk new_AGEMA_reg_buffer_3391 ( .C (clk), .D (new_AGEMA_signal_6166), .Q (new_AGEMA_signal_6167) ) ;
    buf_clk new_AGEMA_reg_buffer_3399 ( .C (clk), .D (new_AGEMA_signal_6174), .Q (new_AGEMA_signal_6175) ) ;
    buf_clk new_AGEMA_reg_buffer_3407 ( .C (clk), .D (new_AGEMA_signal_6182), .Q (new_AGEMA_signal_6183) ) ;
    buf_clk new_AGEMA_reg_buffer_3415 ( .C (clk), .D (new_AGEMA_signal_6190), .Q (new_AGEMA_signal_6191) ) ;
    buf_clk new_AGEMA_reg_buffer_3423 ( .C (clk), .D (new_AGEMA_signal_6198), .Q (new_AGEMA_signal_6199) ) ;
    buf_clk new_AGEMA_reg_buffer_3431 ( .C (clk), .D (new_AGEMA_signal_6206), .Q (new_AGEMA_signal_6207) ) ;
    buf_clk new_AGEMA_reg_buffer_3439 ( .C (clk), .D (new_AGEMA_signal_6214), .Q (new_AGEMA_signal_6215) ) ;
    buf_clk new_AGEMA_reg_buffer_3447 ( .C (clk), .D (new_AGEMA_signal_6222), .Q (new_AGEMA_signal_6223) ) ;
    buf_clk new_AGEMA_reg_buffer_3455 ( .C (clk), .D (new_AGEMA_signal_6230), .Q (new_AGEMA_signal_6231) ) ;
    buf_clk new_AGEMA_reg_buffer_3463 ( .C (clk), .D (new_AGEMA_signal_6238), .Q (new_AGEMA_signal_6239) ) ;
    buf_clk new_AGEMA_reg_buffer_3471 ( .C (clk), .D (new_AGEMA_signal_6246), .Q (new_AGEMA_signal_6247) ) ;
    buf_clk new_AGEMA_reg_buffer_3479 ( .C (clk), .D (new_AGEMA_signal_6254), .Q (new_AGEMA_signal_6255) ) ;
    buf_clk new_AGEMA_reg_buffer_3487 ( .C (clk), .D (new_AGEMA_signal_6262), .Q (new_AGEMA_signal_6263) ) ;
    buf_clk new_AGEMA_reg_buffer_3495 ( .C (clk), .D (new_AGEMA_signal_6270), .Q (new_AGEMA_signal_6271) ) ;
    buf_clk new_AGEMA_reg_buffer_3503 ( .C (clk), .D (new_AGEMA_signal_6278), .Q (new_AGEMA_signal_6279) ) ;
    buf_clk new_AGEMA_reg_buffer_3511 ( .C (clk), .D (new_AGEMA_signal_6286), .Q (new_AGEMA_signal_6287) ) ;
    buf_clk new_AGEMA_reg_buffer_3519 ( .C (clk), .D (new_AGEMA_signal_6294), .Q (new_AGEMA_signal_6295) ) ;
    buf_clk new_AGEMA_reg_buffer_3527 ( .C (clk), .D (new_AGEMA_signal_6302), .Q (new_AGEMA_signal_6303) ) ;
    buf_clk new_AGEMA_reg_buffer_3535 ( .C (clk), .D (new_AGEMA_signal_6310), .Q (new_AGEMA_signal_6311) ) ;
    buf_clk new_AGEMA_reg_buffer_3543 ( .C (clk), .D (new_AGEMA_signal_6318), .Q (new_AGEMA_signal_6319) ) ;
    buf_clk new_AGEMA_reg_buffer_3551 ( .C (clk), .D (new_AGEMA_signal_6326), .Q (new_AGEMA_signal_6327) ) ;
    buf_clk new_AGEMA_reg_buffer_3559 ( .C (clk), .D (new_AGEMA_signal_6334), .Q (new_AGEMA_signal_6335) ) ;
    buf_clk new_AGEMA_reg_buffer_3567 ( .C (clk), .D (new_AGEMA_signal_6342), .Q (new_AGEMA_signal_6343) ) ;
    buf_clk new_AGEMA_reg_buffer_3575 ( .C (clk), .D (new_AGEMA_signal_6350), .Q (new_AGEMA_signal_6351) ) ;
    buf_clk new_AGEMA_reg_buffer_3583 ( .C (clk), .D (new_AGEMA_signal_6358), .Q (new_AGEMA_signal_6359) ) ;
    buf_clk new_AGEMA_reg_buffer_3591 ( .C (clk), .D (new_AGEMA_signal_6366), .Q (new_AGEMA_signal_6367) ) ;
    buf_clk new_AGEMA_reg_buffer_3599 ( .C (clk), .D (new_AGEMA_signal_6374), .Q (new_AGEMA_signal_6375) ) ;
    buf_clk new_AGEMA_reg_buffer_3607 ( .C (clk), .D (new_AGEMA_signal_6382), .Q (new_AGEMA_signal_6383) ) ;
    buf_clk new_AGEMA_reg_buffer_3615 ( .C (clk), .D (new_AGEMA_signal_6390), .Q (new_AGEMA_signal_6391) ) ;
    buf_clk new_AGEMA_reg_buffer_3623 ( .C (clk), .D (new_AGEMA_signal_6398), .Q (new_AGEMA_signal_6399) ) ;
    buf_clk new_AGEMA_reg_buffer_3631 ( .C (clk), .D (new_AGEMA_signal_6406), .Q (new_AGEMA_signal_6407) ) ;
    buf_clk new_AGEMA_reg_buffer_3639 ( .C (clk), .D (new_AGEMA_signal_6414), .Q (new_AGEMA_signal_6415) ) ;
    buf_clk new_AGEMA_reg_buffer_3647 ( .C (clk), .D (new_AGEMA_signal_6422), .Q (new_AGEMA_signal_6423) ) ;
    buf_clk new_AGEMA_reg_buffer_3655 ( .C (clk), .D (new_AGEMA_signal_6430), .Q (new_AGEMA_signal_6431) ) ;
    buf_clk new_AGEMA_reg_buffer_3663 ( .C (clk), .D (new_AGEMA_signal_6438), .Q (new_AGEMA_signal_6439) ) ;
    buf_clk new_AGEMA_reg_buffer_3671 ( .C (clk), .D (new_AGEMA_signal_6446), .Q (new_AGEMA_signal_6447) ) ;
    buf_clk new_AGEMA_reg_buffer_3679 ( .C (clk), .D (new_AGEMA_signal_6454), .Q (new_AGEMA_signal_6455) ) ;
    buf_clk new_AGEMA_reg_buffer_3687 ( .C (clk), .D (new_AGEMA_signal_6462), .Q (new_AGEMA_signal_6463) ) ;
    buf_clk new_AGEMA_reg_buffer_3695 ( .C (clk), .D (new_AGEMA_signal_6470), .Q (new_AGEMA_signal_6471) ) ;
    buf_clk new_AGEMA_reg_buffer_3703 ( .C (clk), .D (new_AGEMA_signal_6478), .Q (new_AGEMA_signal_6479) ) ;
    buf_clk new_AGEMA_reg_buffer_3711 ( .C (clk), .D (new_AGEMA_signal_6486), .Q (new_AGEMA_signal_6487) ) ;
    buf_clk new_AGEMA_reg_buffer_3719 ( .C (clk), .D (new_AGEMA_signal_6494), .Q (new_AGEMA_signal_6495) ) ;
    buf_clk new_AGEMA_reg_buffer_3727 ( .C (clk), .D (new_AGEMA_signal_6502), .Q (new_AGEMA_signal_6503) ) ;
    buf_clk new_AGEMA_reg_buffer_3735 ( .C (clk), .D (new_AGEMA_signal_6510), .Q (new_AGEMA_signal_6511) ) ;
    buf_clk new_AGEMA_reg_buffer_3743 ( .C (clk), .D (new_AGEMA_signal_6518), .Q (new_AGEMA_signal_6519) ) ;
    buf_clk new_AGEMA_reg_buffer_3751 ( .C (clk), .D (new_AGEMA_signal_6526), .Q (new_AGEMA_signal_6527) ) ;
    buf_clk new_AGEMA_reg_buffer_3759 ( .C (clk), .D (new_AGEMA_signal_6534), .Q (new_AGEMA_signal_6535) ) ;
    buf_clk new_AGEMA_reg_buffer_3767 ( .C (clk), .D (new_AGEMA_signal_6542), .Q (new_AGEMA_signal_6543) ) ;
    buf_clk new_AGEMA_reg_buffer_3775 ( .C (clk), .D (new_AGEMA_signal_6550), .Q (new_AGEMA_signal_6551) ) ;
    buf_clk new_AGEMA_reg_buffer_3783 ( .C (clk), .D (new_AGEMA_signal_6558), .Q (new_AGEMA_signal_6559) ) ;
    buf_clk new_AGEMA_reg_buffer_3791 ( .C (clk), .D (new_AGEMA_signal_6566), .Q (new_AGEMA_signal_6567) ) ;
    buf_clk new_AGEMA_reg_buffer_3799 ( .C (clk), .D (new_AGEMA_signal_6574), .Q (new_AGEMA_signal_6575) ) ;
    buf_clk new_AGEMA_reg_buffer_3807 ( .C (clk), .D (new_AGEMA_signal_6582), .Q (new_AGEMA_signal_6583) ) ;
    buf_clk new_AGEMA_reg_buffer_3815 ( .C (clk), .D (new_AGEMA_signal_6590), .Q (new_AGEMA_signal_6591) ) ;
    buf_clk new_AGEMA_reg_buffer_3823 ( .C (clk), .D (new_AGEMA_signal_6598), .Q (new_AGEMA_signal_6599) ) ;
    buf_clk new_AGEMA_reg_buffer_3831 ( .C (clk), .D (new_AGEMA_signal_6606), .Q (new_AGEMA_signal_6607) ) ;
    buf_clk new_AGEMA_reg_buffer_3839 ( .C (clk), .D (new_AGEMA_signal_6614), .Q (new_AGEMA_signal_6615) ) ;
    buf_clk new_AGEMA_reg_buffer_3847 ( .C (clk), .D (new_AGEMA_signal_6622), .Q (new_AGEMA_signal_6623) ) ;
    buf_clk new_AGEMA_reg_buffer_3855 ( .C (clk), .D (new_AGEMA_signal_6630), .Q (new_AGEMA_signal_6631) ) ;
    buf_clk new_AGEMA_reg_buffer_3863 ( .C (clk), .D (new_AGEMA_signal_6638), .Q (new_AGEMA_signal_6639) ) ;
    buf_clk new_AGEMA_reg_buffer_3871 ( .C (clk), .D (new_AGEMA_signal_6646), .Q (new_AGEMA_signal_6647) ) ;
    buf_clk new_AGEMA_reg_buffer_3879 ( .C (clk), .D (new_AGEMA_signal_6654), .Q (new_AGEMA_signal_6655) ) ;
    buf_clk new_AGEMA_reg_buffer_3887 ( .C (clk), .D (new_AGEMA_signal_6662), .Q (new_AGEMA_signal_6663) ) ;
    buf_clk new_AGEMA_reg_buffer_3895 ( .C (clk), .D (new_AGEMA_signal_6670), .Q (new_AGEMA_signal_6671) ) ;
    buf_clk new_AGEMA_reg_buffer_3903 ( .C (clk), .D (new_AGEMA_signal_6678), .Q (new_AGEMA_signal_6679) ) ;
    buf_clk new_AGEMA_reg_buffer_3911 ( .C (clk), .D (new_AGEMA_signal_6686), .Q (new_AGEMA_signal_6687) ) ;
    buf_clk new_AGEMA_reg_buffer_3919 ( .C (clk), .D (new_AGEMA_signal_6694), .Q (new_AGEMA_signal_6695) ) ;
    buf_clk new_AGEMA_reg_buffer_3927 ( .C (clk), .D (new_AGEMA_signal_6702), .Q (new_AGEMA_signal_6703) ) ;
    buf_clk new_AGEMA_reg_buffer_3935 ( .C (clk), .D (new_AGEMA_signal_6710), .Q (new_AGEMA_signal_6711) ) ;
    buf_clk new_AGEMA_reg_buffer_3943 ( .C (clk), .D (new_AGEMA_signal_6718), .Q (new_AGEMA_signal_6719) ) ;
    buf_clk new_AGEMA_reg_buffer_3951 ( .C (clk), .D (new_AGEMA_signal_6726), .Q (new_AGEMA_signal_6727) ) ;
    buf_clk new_AGEMA_reg_buffer_3959 ( .C (clk), .D (new_AGEMA_signal_6734), .Q (new_AGEMA_signal_6735) ) ;
    buf_clk new_AGEMA_reg_buffer_3967 ( .C (clk), .D (new_AGEMA_signal_6742), .Q (new_AGEMA_signal_6743) ) ;
    buf_clk new_AGEMA_reg_buffer_3975 ( .C (clk), .D (new_AGEMA_signal_6750), .Q (new_AGEMA_signal_6751) ) ;
    buf_clk new_AGEMA_reg_buffer_3983 ( .C (clk), .D (new_AGEMA_signal_6758), .Q (new_AGEMA_signal_6759) ) ;
    buf_clk new_AGEMA_reg_buffer_3991 ( .C (clk), .D (new_AGEMA_signal_6766), .Q (new_AGEMA_signal_6767) ) ;
    buf_clk new_AGEMA_reg_buffer_3999 ( .C (clk), .D (new_AGEMA_signal_6774), .Q (new_AGEMA_signal_6775) ) ;
    buf_clk new_AGEMA_reg_buffer_4007 ( .C (clk), .D (new_AGEMA_signal_6782), .Q (new_AGEMA_signal_6783) ) ;
    buf_clk new_AGEMA_reg_buffer_4015 ( .C (clk), .D (new_AGEMA_signal_6790), .Q (new_AGEMA_signal_6791) ) ;
    buf_clk new_AGEMA_reg_buffer_4023 ( .C (clk), .D (new_AGEMA_signal_6798), .Q (new_AGEMA_signal_6799) ) ;
    buf_clk new_AGEMA_reg_buffer_4031 ( .C (clk), .D (new_AGEMA_signal_6806), .Q (new_AGEMA_signal_6807) ) ;
    buf_clk new_AGEMA_reg_buffer_4039 ( .C (clk), .D (new_AGEMA_signal_6814), .Q (new_AGEMA_signal_6815) ) ;
    buf_clk new_AGEMA_reg_buffer_4047 ( .C (clk), .D (new_AGEMA_signal_6822), .Q (new_AGEMA_signal_6823) ) ;
    buf_clk new_AGEMA_reg_buffer_4055 ( .C (clk), .D (new_AGEMA_signal_6830), .Q (new_AGEMA_signal_6831) ) ;
    buf_clk new_AGEMA_reg_buffer_4063 ( .C (clk), .D (new_AGEMA_signal_6838), .Q (new_AGEMA_signal_6839) ) ;
    buf_clk new_AGEMA_reg_buffer_4071 ( .C (clk), .D (new_AGEMA_signal_6846), .Q (new_AGEMA_signal_6847) ) ;
    buf_clk new_AGEMA_reg_buffer_4079 ( .C (clk), .D (new_AGEMA_signal_6854), .Q (new_AGEMA_signal_6855) ) ;
    buf_clk new_AGEMA_reg_buffer_4087 ( .C (clk), .D (new_AGEMA_signal_6862), .Q (new_AGEMA_signal_6863) ) ;
    buf_clk new_AGEMA_reg_buffer_4095 ( .C (clk), .D (new_AGEMA_signal_6870), .Q (new_AGEMA_signal_6871) ) ;
    buf_clk new_AGEMA_reg_buffer_4103 ( .C (clk), .D (new_AGEMA_signal_6878), .Q (new_AGEMA_signal_6879) ) ;
    buf_clk new_AGEMA_reg_buffer_4111 ( .C (clk), .D (new_AGEMA_signal_6886), .Q (new_AGEMA_signal_6887) ) ;
    buf_clk new_AGEMA_reg_buffer_4119 ( .C (clk), .D (new_AGEMA_signal_6894), .Q (new_AGEMA_signal_6895) ) ;
    buf_clk new_AGEMA_reg_buffer_4127 ( .C (clk), .D (new_AGEMA_signal_6902), .Q (new_AGEMA_signal_6903) ) ;
    buf_clk new_AGEMA_reg_buffer_4135 ( .C (clk), .D (new_AGEMA_signal_6910), .Q (new_AGEMA_signal_6911) ) ;
    buf_clk new_AGEMA_reg_buffer_4143 ( .C (clk), .D (new_AGEMA_signal_6918), .Q (new_AGEMA_signal_6919) ) ;
    buf_clk new_AGEMA_reg_buffer_4151 ( .C (clk), .D (new_AGEMA_signal_6926), .Q (new_AGEMA_signal_6927) ) ;
    buf_clk new_AGEMA_reg_buffer_4159 ( .C (clk), .D (new_AGEMA_signal_6934), .Q (new_AGEMA_signal_6935) ) ;
    buf_clk new_AGEMA_reg_buffer_4167 ( .C (clk), .D (new_AGEMA_signal_6942), .Q (new_AGEMA_signal_6943) ) ;
    buf_clk new_AGEMA_reg_buffer_4175 ( .C (clk), .D (new_AGEMA_signal_6950), .Q (new_AGEMA_signal_6951) ) ;
    buf_clk new_AGEMA_reg_buffer_4183 ( .C (clk), .D (new_AGEMA_signal_6958), .Q (new_AGEMA_signal_6959) ) ;
    buf_clk new_AGEMA_reg_buffer_4187 ( .C (clk), .D (new_AGEMA_signal_5138), .Q (new_AGEMA_signal_6963) ) ;
    buf_clk new_AGEMA_reg_buffer_4189 ( .C (clk), .D (new_AGEMA_signal_5140), .Q (new_AGEMA_signal_6965) ) ;
    buf_clk new_AGEMA_reg_buffer_4191 ( .C (clk), .D (new_AGEMA_signal_5142), .Q (new_AGEMA_signal_6967) ) ;
    buf_clk new_AGEMA_reg_buffer_4195 ( .C (clk), .D (new_AGEMA_signal_6970), .Q (new_AGEMA_signal_6971) ) ;
    buf_clk new_AGEMA_reg_buffer_4199 ( .C (clk), .D (new_AGEMA_signal_6974), .Q (new_AGEMA_signal_6975) ) ;
    buf_clk new_AGEMA_reg_buffer_4203 ( .C (clk), .D (new_AGEMA_signal_6978), .Q (new_AGEMA_signal_6979) ) ;
    buf_clk new_AGEMA_reg_buffer_4205 ( .C (clk), .D (new_AGEMA_signal_5156), .Q (new_AGEMA_signal_6981) ) ;
    buf_clk new_AGEMA_reg_buffer_4207 ( .C (clk), .D (new_AGEMA_signal_5158), .Q (new_AGEMA_signal_6983) ) ;
    buf_clk new_AGEMA_reg_buffer_4209 ( .C (clk), .D (new_AGEMA_signal_5160), .Q (new_AGEMA_signal_6985) ) ;
    buf_clk new_AGEMA_reg_buffer_4213 ( .C (clk), .D (new_AGEMA_signal_6988), .Q (new_AGEMA_signal_6989) ) ;
    buf_clk new_AGEMA_reg_buffer_4217 ( .C (clk), .D (new_AGEMA_signal_6992), .Q (new_AGEMA_signal_6993) ) ;
    buf_clk new_AGEMA_reg_buffer_4221 ( .C (clk), .D (new_AGEMA_signal_6996), .Q (new_AGEMA_signal_6997) ) ;
    buf_clk new_AGEMA_reg_buffer_4223 ( .C (clk), .D (new_AGEMA_signal_5174), .Q (new_AGEMA_signal_6999) ) ;
    buf_clk new_AGEMA_reg_buffer_4225 ( .C (clk), .D (new_AGEMA_signal_5176), .Q (new_AGEMA_signal_7001) ) ;
    buf_clk new_AGEMA_reg_buffer_4227 ( .C (clk), .D (new_AGEMA_signal_5178), .Q (new_AGEMA_signal_7003) ) ;
    buf_clk new_AGEMA_reg_buffer_4231 ( .C (clk), .D (new_AGEMA_signal_7006), .Q (new_AGEMA_signal_7007) ) ;
    buf_clk new_AGEMA_reg_buffer_4235 ( .C (clk), .D (new_AGEMA_signal_7010), .Q (new_AGEMA_signal_7011) ) ;
    buf_clk new_AGEMA_reg_buffer_4239 ( .C (clk), .D (new_AGEMA_signal_7014), .Q (new_AGEMA_signal_7015) ) ;
    buf_clk new_AGEMA_reg_buffer_4241 ( .C (clk), .D (new_AGEMA_signal_5192), .Q (new_AGEMA_signal_7017) ) ;
    buf_clk new_AGEMA_reg_buffer_4243 ( .C (clk), .D (new_AGEMA_signal_5194), .Q (new_AGEMA_signal_7019) ) ;
    buf_clk new_AGEMA_reg_buffer_4245 ( .C (clk), .D (new_AGEMA_signal_5196), .Q (new_AGEMA_signal_7021) ) ;
    buf_clk new_AGEMA_reg_buffer_4249 ( .C (clk), .D (new_AGEMA_signal_7024), .Q (new_AGEMA_signal_7025) ) ;
    buf_clk new_AGEMA_reg_buffer_4253 ( .C (clk), .D (new_AGEMA_signal_7028), .Q (new_AGEMA_signal_7029) ) ;
    buf_clk new_AGEMA_reg_buffer_4257 ( .C (clk), .D (new_AGEMA_signal_7032), .Q (new_AGEMA_signal_7033) ) ;
    buf_clk new_AGEMA_reg_buffer_4259 ( .C (clk), .D (new_AGEMA_signal_5210), .Q (new_AGEMA_signal_7035) ) ;
    buf_clk new_AGEMA_reg_buffer_4261 ( .C (clk), .D (new_AGEMA_signal_5212), .Q (new_AGEMA_signal_7037) ) ;
    buf_clk new_AGEMA_reg_buffer_4263 ( .C (clk), .D (new_AGEMA_signal_5214), .Q (new_AGEMA_signal_7039) ) ;
    buf_clk new_AGEMA_reg_buffer_4267 ( .C (clk), .D (new_AGEMA_signal_7042), .Q (new_AGEMA_signal_7043) ) ;
    buf_clk new_AGEMA_reg_buffer_4271 ( .C (clk), .D (new_AGEMA_signal_7046), .Q (new_AGEMA_signal_7047) ) ;
    buf_clk new_AGEMA_reg_buffer_4275 ( .C (clk), .D (new_AGEMA_signal_7050), .Q (new_AGEMA_signal_7051) ) ;
    buf_clk new_AGEMA_reg_buffer_4277 ( .C (clk), .D (new_AGEMA_signal_5228), .Q (new_AGEMA_signal_7053) ) ;
    buf_clk new_AGEMA_reg_buffer_4279 ( .C (clk), .D (new_AGEMA_signal_5230), .Q (new_AGEMA_signal_7055) ) ;
    buf_clk new_AGEMA_reg_buffer_4281 ( .C (clk), .D (new_AGEMA_signal_5232), .Q (new_AGEMA_signal_7057) ) ;
    buf_clk new_AGEMA_reg_buffer_4285 ( .C (clk), .D (new_AGEMA_signal_7060), .Q (new_AGEMA_signal_7061) ) ;
    buf_clk new_AGEMA_reg_buffer_4289 ( .C (clk), .D (new_AGEMA_signal_7064), .Q (new_AGEMA_signal_7065) ) ;
    buf_clk new_AGEMA_reg_buffer_4293 ( .C (clk), .D (new_AGEMA_signal_7068), .Q (new_AGEMA_signal_7069) ) ;
    buf_clk new_AGEMA_reg_buffer_4295 ( .C (clk), .D (new_AGEMA_signal_5246), .Q (new_AGEMA_signal_7071) ) ;
    buf_clk new_AGEMA_reg_buffer_4297 ( .C (clk), .D (new_AGEMA_signal_5248), .Q (new_AGEMA_signal_7073) ) ;
    buf_clk new_AGEMA_reg_buffer_4299 ( .C (clk), .D (new_AGEMA_signal_5250), .Q (new_AGEMA_signal_7075) ) ;
    buf_clk new_AGEMA_reg_buffer_4303 ( .C (clk), .D (new_AGEMA_signal_7078), .Q (new_AGEMA_signal_7079) ) ;
    buf_clk new_AGEMA_reg_buffer_4307 ( .C (clk), .D (new_AGEMA_signal_7082), .Q (new_AGEMA_signal_7083) ) ;
    buf_clk new_AGEMA_reg_buffer_4311 ( .C (clk), .D (new_AGEMA_signal_7086), .Q (new_AGEMA_signal_7087) ) ;
    buf_clk new_AGEMA_reg_buffer_4313 ( .C (clk), .D (new_AGEMA_signal_5264), .Q (new_AGEMA_signal_7089) ) ;
    buf_clk new_AGEMA_reg_buffer_4315 ( .C (clk), .D (new_AGEMA_signal_5266), .Q (new_AGEMA_signal_7091) ) ;
    buf_clk new_AGEMA_reg_buffer_4317 ( .C (clk), .D (new_AGEMA_signal_5268), .Q (new_AGEMA_signal_7093) ) ;
    buf_clk new_AGEMA_reg_buffer_4321 ( .C (clk), .D (new_AGEMA_signal_7096), .Q (new_AGEMA_signal_7097) ) ;
    buf_clk new_AGEMA_reg_buffer_4325 ( .C (clk), .D (new_AGEMA_signal_7100), .Q (new_AGEMA_signal_7101) ) ;
    buf_clk new_AGEMA_reg_buffer_4329 ( .C (clk), .D (new_AGEMA_signal_7104), .Q (new_AGEMA_signal_7105) ) ;
    buf_clk new_AGEMA_reg_buffer_4331 ( .C (clk), .D (new_AGEMA_signal_5282), .Q (new_AGEMA_signal_7107) ) ;
    buf_clk new_AGEMA_reg_buffer_4333 ( .C (clk), .D (new_AGEMA_signal_5284), .Q (new_AGEMA_signal_7109) ) ;
    buf_clk new_AGEMA_reg_buffer_4335 ( .C (clk), .D (new_AGEMA_signal_5286), .Q (new_AGEMA_signal_7111) ) ;
    buf_clk new_AGEMA_reg_buffer_4339 ( .C (clk), .D (new_AGEMA_signal_7114), .Q (new_AGEMA_signal_7115) ) ;
    buf_clk new_AGEMA_reg_buffer_4343 ( .C (clk), .D (new_AGEMA_signal_7118), .Q (new_AGEMA_signal_7119) ) ;
    buf_clk new_AGEMA_reg_buffer_4347 ( .C (clk), .D (new_AGEMA_signal_7122), .Q (new_AGEMA_signal_7123) ) ;
    buf_clk new_AGEMA_reg_buffer_4349 ( .C (clk), .D (new_AGEMA_signal_5300), .Q (new_AGEMA_signal_7125) ) ;
    buf_clk new_AGEMA_reg_buffer_4351 ( .C (clk), .D (new_AGEMA_signal_5302), .Q (new_AGEMA_signal_7127) ) ;
    buf_clk new_AGEMA_reg_buffer_4353 ( .C (clk), .D (new_AGEMA_signal_5304), .Q (new_AGEMA_signal_7129) ) ;
    buf_clk new_AGEMA_reg_buffer_4357 ( .C (clk), .D (new_AGEMA_signal_7132), .Q (new_AGEMA_signal_7133) ) ;
    buf_clk new_AGEMA_reg_buffer_4361 ( .C (clk), .D (new_AGEMA_signal_7136), .Q (new_AGEMA_signal_7137) ) ;
    buf_clk new_AGEMA_reg_buffer_4365 ( .C (clk), .D (new_AGEMA_signal_7140), .Q (new_AGEMA_signal_7141) ) ;
    buf_clk new_AGEMA_reg_buffer_4367 ( .C (clk), .D (new_AGEMA_signal_5318), .Q (new_AGEMA_signal_7143) ) ;
    buf_clk new_AGEMA_reg_buffer_4369 ( .C (clk), .D (new_AGEMA_signal_5320), .Q (new_AGEMA_signal_7145) ) ;
    buf_clk new_AGEMA_reg_buffer_4371 ( .C (clk), .D (new_AGEMA_signal_5322), .Q (new_AGEMA_signal_7147) ) ;
    buf_clk new_AGEMA_reg_buffer_4375 ( .C (clk), .D (new_AGEMA_signal_7150), .Q (new_AGEMA_signal_7151) ) ;
    buf_clk new_AGEMA_reg_buffer_4379 ( .C (clk), .D (new_AGEMA_signal_7154), .Q (new_AGEMA_signal_7155) ) ;
    buf_clk new_AGEMA_reg_buffer_4383 ( .C (clk), .D (new_AGEMA_signal_7158), .Q (new_AGEMA_signal_7159) ) ;
    buf_clk new_AGEMA_reg_buffer_4385 ( .C (clk), .D (new_AGEMA_signal_5336), .Q (new_AGEMA_signal_7161) ) ;
    buf_clk new_AGEMA_reg_buffer_4387 ( .C (clk), .D (new_AGEMA_signal_5338), .Q (new_AGEMA_signal_7163) ) ;
    buf_clk new_AGEMA_reg_buffer_4389 ( .C (clk), .D (new_AGEMA_signal_5340), .Q (new_AGEMA_signal_7165) ) ;
    buf_clk new_AGEMA_reg_buffer_4393 ( .C (clk), .D (new_AGEMA_signal_7168), .Q (new_AGEMA_signal_7169) ) ;
    buf_clk new_AGEMA_reg_buffer_4397 ( .C (clk), .D (new_AGEMA_signal_7172), .Q (new_AGEMA_signal_7173) ) ;
    buf_clk new_AGEMA_reg_buffer_4401 ( .C (clk), .D (new_AGEMA_signal_7176), .Q (new_AGEMA_signal_7177) ) ;
    buf_clk new_AGEMA_reg_buffer_4403 ( .C (clk), .D (new_AGEMA_signal_5354), .Q (new_AGEMA_signal_7179) ) ;
    buf_clk new_AGEMA_reg_buffer_4405 ( .C (clk), .D (new_AGEMA_signal_5356), .Q (new_AGEMA_signal_7181) ) ;
    buf_clk new_AGEMA_reg_buffer_4407 ( .C (clk), .D (new_AGEMA_signal_5358), .Q (new_AGEMA_signal_7183) ) ;
    buf_clk new_AGEMA_reg_buffer_4411 ( .C (clk), .D (new_AGEMA_signal_7186), .Q (new_AGEMA_signal_7187) ) ;
    buf_clk new_AGEMA_reg_buffer_4415 ( .C (clk), .D (new_AGEMA_signal_7190), .Q (new_AGEMA_signal_7191) ) ;
    buf_clk new_AGEMA_reg_buffer_4419 ( .C (clk), .D (new_AGEMA_signal_7194), .Q (new_AGEMA_signal_7195) ) ;
    buf_clk new_AGEMA_reg_buffer_4421 ( .C (clk), .D (new_AGEMA_signal_5372), .Q (new_AGEMA_signal_7197) ) ;
    buf_clk new_AGEMA_reg_buffer_4423 ( .C (clk), .D (new_AGEMA_signal_5374), .Q (new_AGEMA_signal_7199) ) ;
    buf_clk new_AGEMA_reg_buffer_4425 ( .C (clk), .D (new_AGEMA_signal_5376), .Q (new_AGEMA_signal_7201) ) ;
    buf_clk new_AGEMA_reg_buffer_4429 ( .C (clk), .D (new_AGEMA_signal_7204), .Q (new_AGEMA_signal_7205) ) ;
    buf_clk new_AGEMA_reg_buffer_4433 ( .C (clk), .D (new_AGEMA_signal_7208), .Q (new_AGEMA_signal_7209) ) ;
    buf_clk new_AGEMA_reg_buffer_4437 ( .C (clk), .D (new_AGEMA_signal_7212), .Q (new_AGEMA_signal_7213) ) ;
    buf_clk new_AGEMA_reg_buffer_4439 ( .C (clk), .D (new_AGEMA_signal_5390), .Q (new_AGEMA_signal_7215) ) ;
    buf_clk new_AGEMA_reg_buffer_4441 ( .C (clk), .D (new_AGEMA_signal_5392), .Q (new_AGEMA_signal_7217) ) ;
    buf_clk new_AGEMA_reg_buffer_4443 ( .C (clk), .D (new_AGEMA_signal_5394), .Q (new_AGEMA_signal_7219) ) ;
    buf_clk new_AGEMA_reg_buffer_4447 ( .C (clk), .D (new_AGEMA_signal_7222), .Q (new_AGEMA_signal_7223) ) ;
    buf_clk new_AGEMA_reg_buffer_4451 ( .C (clk), .D (new_AGEMA_signal_7226), .Q (new_AGEMA_signal_7227) ) ;
    buf_clk new_AGEMA_reg_buffer_4455 ( .C (clk), .D (new_AGEMA_signal_7230), .Q (new_AGEMA_signal_7231) ) ;
    buf_clk new_AGEMA_reg_buffer_4457 ( .C (clk), .D (new_AGEMA_signal_5408), .Q (new_AGEMA_signal_7233) ) ;
    buf_clk new_AGEMA_reg_buffer_4459 ( .C (clk), .D (new_AGEMA_signal_5410), .Q (new_AGEMA_signal_7235) ) ;
    buf_clk new_AGEMA_reg_buffer_4461 ( .C (clk), .D (new_AGEMA_signal_5412), .Q (new_AGEMA_signal_7237) ) ;
    buf_clk new_AGEMA_reg_buffer_4465 ( .C (clk), .D (new_AGEMA_signal_7240), .Q (new_AGEMA_signal_7241) ) ;
    buf_clk new_AGEMA_reg_buffer_4469 ( .C (clk), .D (new_AGEMA_signal_7244), .Q (new_AGEMA_signal_7245) ) ;
    buf_clk new_AGEMA_reg_buffer_4473 ( .C (clk), .D (new_AGEMA_signal_7248), .Q (new_AGEMA_signal_7249) ) ;
    buf_clk new_AGEMA_reg_buffer_4671 ( .C (clk), .D (new_AGEMA_signal_7446), .Q (new_AGEMA_signal_7447) ) ;
    buf_clk new_AGEMA_reg_buffer_4679 ( .C (clk), .D (new_AGEMA_signal_7454), .Q (new_AGEMA_signal_7455) ) ;
    buf_clk new_AGEMA_reg_buffer_4687 ( .C (clk), .D (new_AGEMA_signal_7462), .Q (new_AGEMA_signal_7463) ) ;
    buf_clk new_AGEMA_reg_buffer_4695 ( .C (clk), .D (new_AGEMA_signal_7470), .Q (new_AGEMA_signal_7471) ) ;
    buf_clk new_AGEMA_reg_buffer_4703 ( .C (clk), .D (new_AGEMA_signal_7478), .Q (new_AGEMA_signal_7479) ) ;
    buf_clk new_AGEMA_reg_buffer_4711 ( .C (clk), .D (new_AGEMA_signal_7486), .Q (new_AGEMA_signal_7487) ) ;
    buf_clk new_AGEMA_reg_buffer_4719 ( .C (clk), .D (new_AGEMA_signal_7494), .Q (new_AGEMA_signal_7495) ) ;
    buf_clk new_AGEMA_reg_buffer_4727 ( .C (clk), .D (new_AGEMA_signal_7502), .Q (new_AGEMA_signal_7503) ) ;
    buf_clk new_AGEMA_reg_buffer_4735 ( .C (clk), .D (new_AGEMA_signal_7510), .Q (new_AGEMA_signal_7511) ) ;
    buf_clk new_AGEMA_reg_buffer_4743 ( .C (clk), .D (new_AGEMA_signal_7518), .Q (new_AGEMA_signal_7519) ) ;

    /* cells in depth 6 */
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_1_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1728, new_AGEMA_signal_1727, Feedback[1]}), .a ({new_AGEMA_signal_4002, new_AGEMA_signal_3996, new_AGEMA_signal_3990}), .c ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, MCOutput[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_3_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, Feedback[3]}), .a ({new_AGEMA_signal_4020, new_AGEMA_signal_4014, new_AGEMA_signal_4008}), .c ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, MCOutput[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_5_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1736, new_AGEMA_signal_1735, Feedback[5]}), .a ({new_AGEMA_signal_4038, new_AGEMA_signal_4032, new_AGEMA_signal_4026}), .c ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, MCOutput[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_7_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1732, new_AGEMA_signal_1731, Feedback[7]}), .a ({new_AGEMA_signal_4056, new_AGEMA_signal_4050, new_AGEMA_signal_4044}), .c ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, MCOutput[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_9_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1744, new_AGEMA_signal_1743, Feedback[9]}), .a ({new_AGEMA_signal_4074, new_AGEMA_signal_4068, new_AGEMA_signal_4062}), .c ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, MCOutput[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_11_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1740, new_AGEMA_signal_1739, Feedback[11]}), .a ({new_AGEMA_signal_4092, new_AGEMA_signal_4086, new_AGEMA_signal_4080}), .c ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, MCOutput[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_13_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1752, new_AGEMA_signal_1751, Feedback[13]}), .a ({new_AGEMA_signal_4110, new_AGEMA_signal_4104, new_AGEMA_signal_4098}), .c ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, MCOutput[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_15_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, Feedback[15]}), .a ({new_AGEMA_signal_4128, new_AGEMA_signal_4122, new_AGEMA_signal_4116}), .c ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, MCOutput[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_17_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1760, new_AGEMA_signal_1759, Feedback[17]}), .a ({new_AGEMA_signal_4146, new_AGEMA_signal_4140, new_AGEMA_signal_4134}), .c ({new_AGEMA_signal_2210, new_AGEMA_signal_2209, MCOutput[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_19_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1756, new_AGEMA_signal_1755, Feedback[19]}), .a ({new_AGEMA_signal_4164, new_AGEMA_signal_4158, new_AGEMA_signal_4152}), .c ({new_AGEMA_signal_2218, new_AGEMA_signal_2217, MCOutput[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_21_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1768, new_AGEMA_signal_1767, Feedback[21]}), .a ({new_AGEMA_signal_4182, new_AGEMA_signal_4176, new_AGEMA_signal_4170}), .c ({new_AGEMA_signal_2226, new_AGEMA_signal_2225, MCOutput[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_23_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1764, new_AGEMA_signal_1763, Feedback[23]}), .a ({new_AGEMA_signal_4200, new_AGEMA_signal_4194, new_AGEMA_signal_4188}), .c ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, MCOutput[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_25_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1776, new_AGEMA_signal_1775, Feedback[25]}), .a ({new_AGEMA_signal_4218, new_AGEMA_signal_4212, new_AGEMA_signal_4206}), .c ({new_AGEMA_signal_2242, new_AGEMA_signal_2241, MCOutput[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_27_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1772, new_AGEMA_signal_1771, Feedback[27]}), .a ({new_AGEMA_signal_4236, new_AGEMA_signal_4230, new_AGEMA_signal_4224}), .c ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, MCOutput[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_29_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1784, new_AGEMA_signal_1783, Feedback[29]}), .a ({new_AGEMA_signal_4254, new_AGEMA_signal_4248, new_AGEMA_signal_4242}), .c ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, MCOutput[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_31_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1780, new_AGEMA_signal_1779, Feedback[31]}), .a ({new_AGEMA_signal_4272, new_AGEMA_signal_4266, new_AGEMA_signal_4260}), .c ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, MCOutput[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_33_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1792, new_AGEMA_signal_1791, Feedback[33]}), .a ({new_AGEMA_signal_4290, new_AGEMA_signal_4284, new_AGEMA_signal_4278}), .c ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, MCInput[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_35_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, Feedback[35]}), .a ({new_AGEMA_signal_4308, new_AGEMA_signal_4302, new_AGEMA_signal_4296}), .c ({new_AGEMA_signal_2282, new_AGEMA_signal_2281, MCInput[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_37_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1800, new_AGEMA_signal_1799, Feedback[37]}), .a ({new_AGEMA_signal_4326, new_AGEMA_signal_4320, new_AGEMA_signal_4314}), .c ({new_AGEMA_signal_2290, new_AGEMA_signal_2289, MCInput[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_39_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, Feedback[39]}), .a ({new_AGEMA_signal_4344, new_AGEMA_signal_4338, new_AGEMA_signal_4332}), .c ({new_AGEMA_signal_2298, new_AGEMA_signal_2297, MCInput[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_41_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1808, new_AGEMA_signal_1807, Feedback[41]}), .a ({new_AGEMA_signal_4362, new_AGEMA_signal_4356, new_AGEMA_signal_4350}), .c ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, MCInput[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_43_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1804, new_AGEMA_signal_1803, Feedback[43]}), .a ({new_AGEMA_signal_4380, new_AGEMA_signal_4374, new_AGEMA_signal_4368}), .c ({new_AGEMA_signal_2314, new_AGEMA_signal_2313, MCInput[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_45_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1816, new_AGEMA_signal_1815, Feedback[45]}), .a ({new_AGEMA_signal_4398, new_AGEMA_signal_4392, new_AGEMA_signal_4386}), .c ({new_AGEMA_signal_2322, new_AGEMA_signal_2321, MCInput[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_47_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1812, new_AGEMA_signal_1811, Feedback[47]}), .a ({new_AGEMA_signal_4416, new_AGEMA_signal_4410, new_AGEMA_signal_4404}), .c ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, MCInput[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_49_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1824, new_AGEMA_signal_1823, Feedback[49]}), .a ({new_AGEMA_signal_4434, new_AGEMA_signal_4428, new_AGEMA_signal_4422}), .c ({new_AGEMA_signal_2338, new_AGEMA_signal_2337, MCInput[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_51_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1820, new_AGEMA_signal_1819, Feedback[51]}), .a ({new_AGEMA_signal_4452, new_AGEMA_signal_4446, new_AGEMA_signal_4440}), .c ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, MCInput[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_53_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1832, new_AGEMA_signal_1831, Feedback[53]}), .a ({new_AGEMA_signal_4470, new_AGEMA_signal_4464, new_AGEMA_signal_4458}), .c ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, MCInput[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_55_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1828, new_AGEMA_signal_1827, Feedback[55]}), .a ({new_AGEMA_signal_4488, new_AGEMA_signal_4482, new_AGEMA_signal_4476}), .c ({new_AGEMA_signal_2362, new_AGEMA_signal_2361, MCInput[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_57_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1840, new_AGEMA_signal_1839, Feedback[57]}), .a ({new_AGEMA_signal_4506, new_AGEMA_signal_4500, new_AGEMA_signal_4494}), .c ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, MCInput[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_59_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1836, new_AGEMA_signal_1835, Feedback[59]}), .a ({new_AGEMA_signal_4524, new_AGEMA_signal_4518, new_AGEMA_signal_4512}), .c ({new_AGEMA_signal_2378, new_AGEMA_signal_2377, MCInput[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_61_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1848, new_AGEMA_signal_1847, Feedback[61]}), .a ({new_AGEMA_signal_4542, new_AGEMA_signal_4536, new_AGEMA_signal_4530}), .c ({new_AGEMA_signal_2386, new_AGEMA_signal_2385, MCInput[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_63_U1 ( .s (new_AGEMA_signal_3984), .b ({new_AGEMA_signal_1844, new_AGEMA_signal_1843, Feedback[63]}), .a ({new_AGEMA_signal_4560, new_AGEMA_signal_4554, new_AGEMA_signal_4548}), .c ({new_AGEMA_signal_2394, new_AGEMA_signal_2393, MCInput[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_1_U3 ( .a ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, MCInst_XOR_r0_Inst_1_n2}), .b ({new_AGEMA_signal_2418, new_AGEMA_signal_2417, MCInst_XOR_r0_Inst_1_n1}), .c ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, MCOutput[49]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_1_U2 ( .a ({new_AGEMA_signal_2210, new_AGEMA_signal_2209, MCOutput[17]}), .b ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, MCOutput[1]}), .c ({new_AGEMA_signal_2418, new_AGEMA_signal_2417, MCInst_XOR_r0_Inst_1_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2338, new_AGEMA_signal_2337, MCInput[49]}), .c ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, MCInst_XOR_r0_Inst_1_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_1_U2 ( .a ({new_AGEMA_signal_2422, new_AGEMA_signal_2421, MCInst_XOR_r1_Inst_1_n1}), .b ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, MCOutput[1]}), .c ({new_AGEMA_signal_2578, new_AGEMA_signal_2577, MCOutput[33]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, MCInput[33]}), .c ({new_AGEMA_signal_2422, new_AGEMA_signal_2421, MCInst_XOR_r1_Inst_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_3_U3 ( .a ({new_AGEMA_signal_2432, new_AGEMA_signal_2431, MCInst_XOR_r0_Inst_3_n2}), .b ({new_AGEMA_signal_2430, new_AGEMA_signal_2429, MCInst_XOR_r0_Inst_3_n1}), .c ({new_AGEMA_signal_2584, new_AGEMA_signal_2583, MCOutput[51]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_3_U2 ( .a ({new_AGEMA_signal_2218, new_AGEMA_signal_2217, MCOutput[19]}), .b ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, MCOutput[3]}), .c ({new_AGEMA_signal_2430, new_AGEMA_signal_2429, MCInst_XOR_r0_Inst_3_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, MCInput[51]}), .c ({new_AGEMA_signal_2432, new_AGEMA_signal_2431, MCInst_XOR_r0_Inst_3_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_3_U2 ( .a ({new_AGEMA_signal_2434, new_AGEMA_signal_2433, MCInst_XOR_r1_Inst_3_n1}), .b ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, MCOutput[3]}), .c ({new_AGEMA_signal_2586, new_AGEMA_signal_2585, MCOutput[35]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2282, new_AGEMA_signal_2281, MCInput[35]}), .c ({new_AGEMA_signal_2434, new_AGEMA_signal_2433, MCInst_XOR_r1_Inst_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_5_U3 ( .a ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, MCInst_XOR_r0_Inst_5_n2}), .b ({new_AGEMA_signal_2442, new_AGEMA_signal_2441, MCInst_XOR_r0_Inst_5_n1}), .c ({new_AGEMA_signal_2592, new_AGEMA_signal_2591, MCOutput[53]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_5_U2 ( .a ({new_AGEMA_signal_2226, new_AGEMA_signal_2225, MCOutput[21]}), .b ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, MCOutput[5]}), .c ({new_AGEMA_signal_2442, new_AGEMA_signal_2441, MCInst_XOR_r0_Inst_5_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_5_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, MCInput[53]}), .c ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, MCInst_XOR_r0_Inst_5_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_5_U2 ( .a ({new_AGEMA_signal_2446, new_AGEMA_signal_2445, MCInst_XOR_r1_Inst_5_n1}), .b ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, MCOutput[5]}), .c ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, MCOutput[37]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_5_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2290, new_AGEMA_signal_2289, MCInput[37]}), .c ({new_AGEMA_signal_2446, new_AGEMA_signal_2445, MCInst_XOR_r1_Inst_5_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_7_U3 ( .a ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, MCInst_XOR_r0_Inst_7_n2}), .b ({new_AGEMA_signal_2454, new_AGEMA_signal_2453, MCInst_XOR_r0_Inst_7_n1}), .c ({new_AGEMA_signal_2600, new_AGEMA_signal_2599, MCOutput[55]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_7_U2 ( .a ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, MCOutput[23]}), .b ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, MCOutput[7]}), .c ({new_AGEMA_signal_2454, new_AGEMA_signal_2453, MCInst_XOR_r0_Inst_7_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_7_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2362, new_AGEMA_signal_2361, MCInput[55]}), .c ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, MCInst_XOR_r0_Inst_7_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_7_U2 ( .a ({new_AGEMA_signal_2458, new_AGEMA_signal_2457, MCInst_XOR_r1_Inst_7_n1}), .b ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, MCOutput[7]}), .c ({new_AGEMA_signal_2602, new_AGEMA_signal_2601, MCOutput[39]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_7_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2298, new_AGEMA_signal_2297, MCInput[39]}), .c ({new_AGEMA_signal_2458, new_AGEMA_signal_2457, MCInst_XOR_r1_Inst_7_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_9_U3 ( .a ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, MCInst_XOR_r0_Inst_9_n2}), .b ({new_AGEMA_signal_2466, new_AGEMA_signal_2465, MCInst_XOR_r0_Inst_9_n1}), .c ({new_AGEMA_signal_2608, new_AGEMA_signal_2607, MCOutput[57]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_9_U2 ( .a ({new_AGEMA_signal_2242, new_AGEMA_signal_2241, MCOutput[25]}), .b ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, MCOutput[9]}), .c ({new_AGEMA_signal_2466, new_AGEMA_signal_2465, MCInst_XOR_r0_Inst_9_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_9_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, MCInput[57]}), .c ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, MCInst_XOR_r0_Inst_9_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_9_U2 ( .a ({new_AGEMA_signal_2470, new_AGEMA_signal_2469, MCInst_XOR_r1_Inst_9_n1}), .b ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, MCOutput[9]}), .c ({new_AGEMA_signal_2610, new_AGEMA_signal_2609, MCOutput[41]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_9_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, MCInput[41]}), .c ({new_AGEMA_signal_2470, new_AGEMA_signal_2469, MCInst_XOR_r1_Inst_9_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_11_U3 ( .a ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, MCInst_XOR_r0_Inst_11_n2}), .b ({new_AGEMA_signal_2478, new_AGEMA_signal_2477, MCInst_XOR_r0_Inst_11_n1}), .c ({new_AGEMA_signal_2616, new_AGEMA_signal_2615, MCOutput[59]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_11_U2 ( .a ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, MCOutput[27]}), .b ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, MCOutput[11]}), .c ({new_AGEMA_signal_2478, new_AGEMA_signal_2477, MCInst_XOR_r0_Inst_11_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_11_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2378, new_AGEMA_signal_2377, MCInput[59]}), .c ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, MCInst_XOR_r0_Inst_11_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_11_U2 ( .a ({new_AGEMA_signal_2482, new_AGEMA_signal_2481, MCInst_XOR_r1_Inst_11_n1}), .b ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, MCOutput[11]}), .c ({new_AGEMA_signal_2618, new_AGEMA_signal_2617, MCOutput[43]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_11_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2314, new_AGEMA_signal_2313, MCInput[43]}), .c ({new_AGEMA_signal_2482, new_AGEMA_signal_2481, MCInst_XOR_r1_Inst_11_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_13_U3 ( .a ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, MCInst_XOR_r0_Inst_13_n2}), .b ({new_AGEMA_signal_2490, new_AGEMA_signal_2489, MCInst_XOR_r0_Inst_13_n1}), .c ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, MCOutput[61]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_13_U2 ( .a ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, MCOutput[29]}), .b ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, MCOutput[13]}), .c ({new_AGEMA_signal_2490, new_AGEMA_signal_2489, MCInst_XOR_r0_Inst_13_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_13_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2386, new_AGEMA_signal_2385, MCInput[61]}), .c ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, MCInst_XOR_r0_Inst_13_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_13_U2 ( .a ({new_AGEMA_signal_2494, new_AGEMA_signal_2493, MCInst_XOR_r1_Inst_13_n1}), .b ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, MCOutput[13]}), .c ({new_AGEMA_signal_2626, new_AGEMA_signal_2625, MCOutput[45]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_13_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2322, new_AGEMA_signal_2321, MCInput[45]}), .c ({new_AGEMA_signal_2494, new_AGEMA_signal_2493, MCInst_XOR_r1_Inst_13_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_15_U3 ( .a ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, MCInst_XOR_r0_Inst_15_n2}), .b ({new_AGEMA_signal_2502, new_AGEMA_signal_2501, MCInst_XOR_r0_Inst_15_n1}), .c ({new_AGEMA_signal_2632, new_AGEMA_signal_2631, MCOutput[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_15_U2 ( .a ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, MCOutput[31]}), .b ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, MCOutput[15]}), .c ({new_AGEMA_signal_2502, new_AGEMA_signal_2501, MCInst_XOR_r0_Inst_15_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_15_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2394, new_AGEMA_signal_2393, MCInput[63]}), .c ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, MCInst_XOR_r0_Inst_15_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_15_U2 ( .a ({new_AGEMA_signal_2506, new_AGEMA_signal_2505, MCInst_XOR_r1_Inst_15_n1}), .b ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, MCOutput[15]}), .c ({new_AGEMA_signal_2634, new_AGEMA_signal_2633, MCOutput[47]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_15_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, MCInput[47]}), .c ({new_AGEMA_signal_2506, new_AGEMA_signal_2505, MCInst_XOR_r1_Inst_15_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2702, new_AGEMA_signal_2701, AddKeyXOR1_XORInst_0_1_n1}), .b ({new_AGEMA_signal_4578, new_AGEMA_signal_4572, new_AGEMA_signal_4566}), .c ({new_AGEMA_signal_2766, new_AGEMA_signal_2765, AddRoundKeyOutput[49]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, MCOutput[49]}), .c ({new_AGEMA_signal_2702, new_AGEMA_signal_2701, AddKeyXOR1_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2706, new_AGEMA_signal_2705, AddKeyXOR1_XORInst_0_3_n1}), .b ({new_AGEMA_signal_4596, new_AGEMA_signal_4590, new_AGEMA_signal_4584}), .c ({new_AGEMA_signal_2770, new_AGEMA_signal_2769, AddRoundKeyOutput[51]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2584, new_AGEMA_signal_2583, MCOutput[51]}), .c ({new_AGEMA_signal_2706, new_AGEMA_signal_2705, AddKeyXOR1_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, AddKeyXOR1_XORInst_1_1_n1}), .b ({new_AGEMA_signal_4614, new_AGEMA_signal_4608, new_AGEMA_signal_4602}), .c ({new_AGEMA_signal_2774, new_AGEMA_signal_2773, AddRoundKeyOutput[53]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2592, new_AGEMA_signal_2591, MCOutput[53]}), .c ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, AddKeyXOR1_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, AddKeyXOR1_XORInst_1_3_n1}), .b ({new_AGEMA_signal_4632, new_AGEMA_signal_4626, new_AGEMA_signal_4620}), .c ({new_AGEMA_signal_2778, new_AGEMA_signal_2777, AddRoundKeyOutput[55]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2600, new_AGEMA_signal_2599, MCOutput[55]}), .c ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, AddKeyXOR1_XORInst_1_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_2718, new_AGEMA_signal_2717, AddKeyXOR1_XORInst_2_1_n1}), .b ({new_AGEMA_signal_4650, new_AGEMA_signal_4644, new_AGEMA_signal_4638}), .c ({new_AGEMA_signal_2782, new_AGEMA_signal_2781, AddRoundKeyOutput[57]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2608, new_AGEMA_signal_2607, MCOutput[57]}), .c ({new_AGEMA_signal_2718, new_AGEMA_signal_2717, AddKeyXOR1_XORInst_2_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_2722, new_AGEMA_signal_2721, AddKeyXOR1_XORInst_2_3_n1}), .b ({new_AGEMA_signal_4668, new_AGEMA_signal_4662, new_AGEMA_signal_4656}), .c ({new_AGEMA_signal_2786, new_AGEMA_signal_2785, AddRoundKeyOutput[59]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2616, new_AGEMA_signal_2615, MCOutput[59]}), .c ({new_AGEMA_signal_2722, new_AGEMA_signal_2721, AddKeyXOR1_XORInst_2_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, AddKeyXOR1_XORInst_3_1_n1}), .b ({new_AGEMA_signal_4686, new_AGEMA_signal_4680, new_AGEMA_signal_4674}), .c ({new_AGEMA_signal_2790, new_AGEMA_signal_2789, AddRoundKeyOutput[61]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, MCOutput[61]}), .c ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, AddKeyXOR1_XORInst_3_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_2730, new_AGEMA_signal_2729, AddKeyXOR1_XORInst_3_3_n1}), .b ({new_AGEMA_signal_4704, new_AGEMA_signal_4698, new_AGEMA_signal_4692}), .c ({new_AGEMA_signal_2794, new_AGEMA_signal_2793, AddRoundKeyOutput[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2632, new_AGEMA_signal_2631, MCOutput[63]}), .c ({new_AGEMA_signal_2730, new_AGEMA_signal_2729, AddKeyXOR1_XORInst_3_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_0_1_U3 ( .a ({new_AGEMA_signal_2734, new_AGEMA_signal_2733, AddKeyConstXOR_XORInst_0_1_n2}), .b ({new_AGEMA_signal_4722, new_AGEMA_signal_4716, new_AGEMA_signal_4710}), .c ({new_AGEMA_signal_2798, new_AGEMA_signal_2797, AddRoundKeyOutput[41]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2610, new_AGEMA_signal_2609, MCOutput[41]}), .c ({new_AGEMA_signal_2734, new_AGEMA_signal_2733, AddKeyConstXOR_XORInst_0_1_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_0_3_U3 ( .a ({new_AGEMA_signal_2738, new_AGEMA_signal_2737, AddKeyConstXOR_XORInst_0_3_n2}), .b ({new_AGEMA_signal_4740, new_AGEMA_signal_4734, new_AGEMA_signal_4728}), .c ({new_AGEMA_signal_2802, new_AGEMA_signal_2801, AddRoundKeyOutput[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2618, new_AGEMA_signal_2617, MCOutput[43]}), .c ({new_AGEMA_signal_2738, new_AGEMA_signal_2737, AddKeyConstXOR_XORInst_0_3_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_1_1_U3 ( .a ({new_AGEMA_signal_2742, new_AGEMA_signal_2741, AddKeyConstXOR_XORInst_1_1_n2}), .b ({new_AGEMA_signal_4758, new_AGEMA_signal_4752, new_AGEMA_signal_4746}), .c ({new_AGEMA_signal_2806, new_AGEMA_signal_2805, AddRoundKeyOutput[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2626, new_AGEMA_signal_2625, MCOutput[45]}), .c ({new_AGEMA_signal_2742, new_AGEMA_signal_2741, AddKeyConstXOR_XORInst_1_1_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_1_3_U3 ( .a ({new_AGEMA_signal_2746, new_AGEMA_signal_2745, AddKeyConstXOR_XORInst_1_3_n2}), .b ({new_AGEMA_signal_4776, new_AGEMA_signal_4770, new_AGEMA_signal_4764}), .c ({new_AGEMA_signal_2810, new_AGEMA_signal_2809, AddRoundKeyOutput[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2634, new_AGEMA_signal_2633, MCOutput[47]}), .c ({new_AGEMA_signal_2746, new_AGEMA_signal_2745, AddKeyConstXOR_XORInst_1_3_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, AddKeyXOR2_XORInst_0_1_n1}), .b ({new_AGEMA_signal_4794, new_AGEMA_signal_4788, new_AGEMA_signal_4782}), .c ({new_AGEMA_signal_2638, new_AGEMA_signal_2637, AddRoundKeyOutput[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, MCOutput[1]}), .c ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, AddKeyXOR2_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2514, new_AGEMA_signal_2513, AddKeyXOR2_XORInst_0_3_n1}), .b ({new_AGEMA_signal_4812, new_AGEMA_signal_4806, new_AGEMA_signal_4800}), .c ({new_AGEMA_signal_2642, new_AGEMA_signal_2641, AddRoundKeyOutput[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, MCOutput[3]}), .c ({new_AGEMA_signal_2514, new_AGEMA_signal_2513, AddKeyXOR2_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2518, new_AGEMA_signal_2517, AddKeyXOR2_XORInst_1_1_n1}), .b ({new_AGEMA_signal_4830, new_AGEMA_signal_4824, new_AGEMA_signal_4818}), .c ({new_AGEMA_signal_2646, new_AGEMA_signal_2645, AddRoundKeyOutput[5]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, MCOutput[5]}), .c ({new_AGEMA_signal_2518, new_AGEMA_signal_2517, AddKeyXOR2_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, AddKeyXOR2_XORInst_1_3_n1}), .b ({new_AGEMA_signal_4848, new_AGEMA_signal_4842, new_AGEMA_signal_4836}), .c ({new_AGEMA_signal_2650, new_AGEMA_signal_2649, AddRoundKeyOutput[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, MCOutput[7]}), .c ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, AddKeyXOR2_XORInst_1_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_2526, new_AGEMA_signal_2525, AddKeyXOR2_XORInst_2_1_n1}), .b ({new_AGEMA_signal_4866, new_AGEMA_signal_4860, new_AGEMA_signal_4854}), .c ({new_AGEMA_signal_2654, new_AGEMA_signal_2653, AddRoundKeyOutput[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, MCOutput[9]}), .c ({new_AGEMA_signal_2526, new_AGEMA_signal_2525, AddKeyXOR2_XORInst_2_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_2530, new_AGEMA_signal_2529, AddKeyXOR2_XORInst_2_3_n1}), .b ({new_AGEMA_signal_4884, new_AGEMA_signal_4878, new_AGEMA_signal_4872}), .c ({new_AGEMA_signal_2658, new_AGEMA_signal_2657, AddRoundKeyOutput[11]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, MCOutput[11]}), .c ({new_AGEMA_signal_2530, new_AGEMA_signal_2529, AddKeyXOR2_XORInst_2_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, AddKeyXOR2_XORInst_3_1_n1}), .b ({new_AGEMA_signal_4902, new_AGEMA_signal_4896, new_AGEMA_signal_4890}), .c ({new_AGEMA_signal_2662, new_AGEMA_signal_2661, AddRoundKeyOutput[13]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, MCOutput[13]}), .c ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, AddKeyXOR2_XORInst_3_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_2538, new_AGEMA_signal_2537, AddKeyXOR2_XORInst_3_3_n1}), .b ({new_AGEMA_signal_4920, new_AGEMA_signal_4914, new_AGEMA_signal_4908}), .c ({new_AGEMA_signal_2666, new_AGEMA_signal_2665, AddRoundKeyOutput[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, MCOutput[15]}), .c ({new_AGEMA_signal_2538, new_AGEMA_signal_2537, AddKeyXOR2_XORInst_3_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_4_1_U2 ( .a ({new_AGEMA_signal_2542, new_AGEMA_signal_2541, AddKeyXOR2_XORInst_4_1_n1}), .b ({new_AGEMA_signal_4938, new_AGEMA_signal_4932, new_AGEMA_signal_4926}), .c ({new_AGEMA_signal_2670, new_AGEMA_signal_2669, AddRoundKeyOutput[17]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_4_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2210, new_AGEMA_signal_2209, MCOutput[17]}), .c ({new_AGEMA_signal_2542, new_AGEMA_signal_2541, AddKeyXOR2_XORInst_4_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_4_3_U2 ( .a ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, AddKeyXOR2_XORInst_4_3_n1}), .b ({new_AGEMA_signal_4956, new_AGEMA_signal_4950, new_AGEMA_signal_4944}), .c ({new_AGEMA_signal_2674, new_AGEMA_signal_2673, AddRoundKeyOutput[19]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_4_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2218, new_AGEMA_signal_2217, MCOutput[19]}), .c ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, AddKeyXOR2_XORInst_4_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_5_1_U2 ( .a ({new_AGEMA_signal_2550, new_AGEMA_signal_2549, AddKeyXOR2_XORInst_5_1_n1}), .b ({new_AGEMA_signal_4974, new_AGEMA_signal_4968, new_AGEMA_signal_4962}), .c ({new_AGEMA_signal_2678, new_AGEMA_signal_2677, AddRoundKeyOutput[21]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_5_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2226, new_AGEMA_signal_2225, MCOutput[21]}), .c ({new_AGEMA_signal_2550, new_AGEMA_signal_2549, AddKeyXOR2_XORInst_5_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_5_3_U2 ( .a ({new_AGEMA_signal_2554, new_AGEMA_signal_2553, AddKeyXOR2_XORInst_5_3_n1}), .b ({new_AGEMA_signal_4992, new_AGEMA_signal_4986, new_AGEMA_signal_4980}), .c ({new_AGEMA_signal_2682, new_AGEMA_signal_2681, AddRoundKeyOutput[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_5_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, MCOutput[23]}), .c ({new_AGEMA_signal_2554, new_AGEMA_signal_2553, AddKeyXOR2_XORInst_5_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_6_1_U2 ( .a ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, AddKeyXOR2_XORInst_6_1_n1}), .b ({new_AGEMA_signal_5010, new_AGEMA_signal_5004, new_AGEMA_signal_4998}), .c ({new_AGEMA_signal_2686, new_AGEMA_signal_2685, AddRoundKeyOutput[25]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_6_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2242, new_AGEMA_signal_2241, MCOutput[25]}), .c ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, AddKeyXOR2_XORInst_6_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_6_3_U2 ( .a ({new_AGEMA_signal_2562, new_AGEMA_signal_2561, AddKeyXOR2_XORInst_6_3_n1}), .b ({new_AGEMA_signal_5028, new_AGEMA_signal_5022, new_AGEMA_signal_5016}), .c ({new_AGEMA_signal_2690, new_AGEMA_signal_2689, AddRoundKeyOutput[27]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_6_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, MCOutput[27]}), .c ({new_AGEMA_signal_2562, new_AGEMA_signal_2561, AddKeyXOR2_XORInst_6_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_7_1_U2 ( .a ({new_AGEMA_signal_2566, new_AGEMA_signal_2565, AddKeyXOR2_XORInst_7_1_n1}), .b ({new_AGEMA_signal_5046, new_AGEMA_signal_5040, new_AGEMA_signal_5034}), .c ({new_AGEMA_signal_2694, new_AGEMA_signal_2693, AddRoundKeyOutput[29]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_7_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, MCOutput[29]}), .c ({new_AGEMA_signal_2566, new_AGEMA_signal_2565, AddKeyXOR2_XORInst_7_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_7_3_U2 ( .a ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, AddKeyXOR2_XORInst_7_3_n1}), .b ({new_AGEMA_signal_5064, new_AGEMA_signal_5058, new_AGEMA_signal_5052}), .c ({new_AGEMA_signal_2698, new_AGEMA_signal_2697, AddRoundKeyOutput[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_7_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, MCOutput[31]}), .c ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, AddKeyXOR2_XORInst_7_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_8_1_U2 ( .a ({new_AGEMA_signal_2750, new_AGEMA_signal_2749, AddKeyXOR2_XORInst_8_1_n1}), .b ({new_AGEMA_signal_5082, new_AGEMA_signal_5076, new_AGEMA_signal_5070}), .c ({new_AGEMA_signal_2814, new_AGEMA_signal_2813, AddRoundKeyOutput[33]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_8_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2578, new_AGEMA_signal_2577, MCOutput[33]}), .c ({new_AGEMA_signal_2750, new_AGEMA_signal_2749, AddKeyXOR2_XORInst_8_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_8_3_U2 ( .a ({new_AGEMA_signal_2754, new_AGEMA_signal_2753, AddKeyXOR2_XORInst_8_3_n1}), .b ({new_AGEMA_signal_5100, new_AGEMA_signal_5094, new_AGEMA_signal_5088}), .c ({new_AGEMA_signal_2818, new_AGEMA_signal_2817, AddRoundKeyOutput[35]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_8_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2586, new_AGEMA_signal_2585, MCOutput[35]}), .c ({new_AGEMA_signal_2754, new_AGEMA_signal_2753, AddKeyXOR2_XORInst_8_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_9_1_U2 ( .a ({new_AGEMA_signal_2758, new_AGEMA_signal_2757, AddKeyXOR2_XORInst_9_1_n1}), .b ({new_AGEMA_signal_5118, new_AGEMA_signal_5112, new_AGEMA_signal_5106}), .c ({new_AGEMA_signal_2822, new_AGEMA_signal_2821, AddRoundKeyOutput[37]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_9_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, MCOutput[37]}), .c ({new_AGEMA_signal_2758, new_AGEMA_signal_2757, AddKeyXOR2_XORInst_9_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_9_3_U2 ( .a ({new_AGEMA_signal_2762, new_AGEMA_signal_2761, AddKeyXOR2_XORInst_9_3_n1}), .b ({new_AGEMA_signal_5136, new_AGEMA_signal_5130, new_AGEMA_signal_5124}), .c ({new_AGEMA_signal_2826, new_AGEMA_signal_2825, AddRoundKeyOutput[39]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_9_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2602, new_AGEMA_signal_2601, MCOutput[39]}), .c ({new_AGEMA_signal_2762, new_AGEMA_signal_2761, AddKeyXOR2_XORInst_9_3_n1}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U19 ( .a ({new_AGEMA_signal_5142, new_AGEMA_signal_5140, new_AGEMA_signal_5138}), .b ({new_AGEMA_signal_1566, new_AGEMA_signal_1565, SubCellInst_SboxInst_0_n14}), .clk (clk), .r ({Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, Feedback[3]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U16 ( .a ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_0_n11}), .b ({new_AGEMA_signal_5148, new_AGEMA_signal_5146, new_AGEMA_signal_5144}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483]}), .c ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, SubCellInst_SboxInst_0_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U12 ( .a ({new_AGEMA_signal_5154, new_AGEMA_signal_5152, new_AGEMA_signal_5150}), .b ({new_AGEMA_signal_1570, new_AGEMA_signal_1569, SubCellInst_SboxInst_0_n5}), .clk (clk), .r ({Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_1728, new_AGEMA_signal_1727, Feedback[1]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U7 ( .a ({new_AGEMA_signal_5148, new_AGEMA_signal_5146, new_AGEMA_signal_5144}), .b ({new_AGEMA_signal_1284, new_AGEMA_signal_1283, SubCellInst_SboxInst_0_n2}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489]}), .c ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, SubCellInst_SboxInst_0_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U19 ( .a ({new_AGEMA_signal_5160, new_AGEMA_signal_5158, new_AGEMA_signal_5156}), .b ({new_AGEMA_signal_1576, new_AGEMA_signal_1575, SubCellInst_SboxInst_1_n14}), .clk (clk), .r ({Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_1732, new_AGEMA_signal_1731, Feedback[7]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U16 ( .a ({new_AGEMA_signal_1288, new_AGEMA_signal_1287, SubCellInst_SboxInst_1_n11}), .b ({new_AGEMA_signal_5166, new_AGEMA_signal_5164, new_AGEMA_signal_5162}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495]}), .c ({new_AGEMA_signal_1578, new_AGEMA_signal_1577, SubCellInst_SboxInst_1_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U12 ( .a ({new_AGEMA_signal_5172, new_AGEMA_signal_5170, new_AGEMA_signal_5168}), .b ({new_AGEMA_signal_1580, new_AGEMA_signal_1579, SubCellInst_SboxInst_1_n5}), .clk (clk), .r ({Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_1736, new_AGEMA_signal_1735, Feedback[5]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U7 ( .a ({new_AGEMA_signal_5166, new_AGEMA_signal_5164, new_AGEMA_signal_5162}), .b ({new_AGEMA_signal_1296, new_AGEMA_signal_1295, SubCellInst_SboxInst_1_n2}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501]}), .c ({new_AGEMA_signal_1582, new_AGEMA_signal_1581, SubCellInst_SboxInst_1_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U19 ( .a ({new_AGEMA_signal_5178, new_AGEMA_signal_5176, new_AGEMA_signal_5174}), .b ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, SubCellInst_SboxInst_2_n14}), .clk (clk), .r ({Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_1740, new_AGEMA_signal_1739, Feedback[11]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U16 ( .a ({new_AGEMA_signal_1300, new_AGEMA_signal_1299, SubCellInst_SboxInst_2_n11}), .b ({new_AGEMA_signal_5184, new_AGEMA_signal_5182, new_AGEMA_signal_5180}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507]}), .c ({new_AGEMA_signal_1588, new_AGEMA_signal_1587, SubCellInst_SboxInst_2_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U12 ( .a ({new_AGEMA_signal_5190, new_AGEMA_signal_5188, new_AGEMA_signal_5186}), .b ({new_AGEMA_signal_1590, new_AGEMA_signal_1589, SubCellInst_SboxInst_2_n5}), .clk (clk), .r ({Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_1744, new_AGEMA_signal_1743, Feedback[9]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U7 ( .a ({new_AGEMA_signal_5184, new_AGEMA_signal_5182, new_AGEMA_signal_5180}), .b ({new_AGEMA_signal_1308, new_AGEMA_signal_1307, SubCellInst_SboxInst_2_n2}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513]}), .c ({new_AGEMA_signal_1592, new_AGEMA_signal_1591, SubCellInst_SboxInst_2_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U19 ( .a ({new_AGEMA_signal_5196, new_AGEMA_signal_5194, new_AGEMA_signal_5192}), .b ({new_AGEMA_signal_1596, new_AGEMA_signal_1595, SubCellInst_SboxInst_3_n14}), .clk (clk), .r ({Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, Feedback[15]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U16 ( .a ({new_AGEMA_signal_1312, new_AGEMA_signal_1311, SubCellInst_SboxInst_3_n11}), .b ({new_AGEMA_signal_5202, new_AGEMA_signal_5200, new_AGEMA_signal_5198}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519]}), .c ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, SubCellInst_SboxInst_3_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U12 ( .a ({new_AGEMA_signal_5208, new_AGEMA_signal_5206, new_AGEMA_signal_5204}), .b ({new_AGEMA_signal_1600, new_AGEMA_signal_1599, SubCellInst_SboxInst_3_n5}), .clk (clk), .r ({Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_1752, new_AGEMA_signal_1751, Feedback[13]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U7 ( .a ({new_AGEMA_signal_5202, new_AGEMA_signal_5200, new_AGEMA_signal_5198}), .b ({new_AGEMA_signal_1320, new_AGEMA_signal_1319, SubCellInst_SboxInst_3_n2}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525]}), .c ({new_AGEMA_signal_1602, new_AGEMA_signal_1601, SubCellInst_SboxInst_3_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U19 ( .a ({new_AGEMA_signal_5214, new_AGEMA_signal_5212, new_AGEMA_signal_5210}), .b ({new_AGEMA_signal_1606, new_AGEMA_signal_1605, SubCellInst_SboxInst_4_n14}), .clk (clk), .r ({Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_1756, new_AGEMA_signal_1755, Feedback[19]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U16 ( .a ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, SubCellInst_SboxInst_4_n11}), .b ({new_AGEMA_signal_5220, new_AGEMA_signal_5218, new_AGEMA_signal_5216}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531]}), .c ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, SubCellInst_SboxInst_4_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U12 ( .a ({new_AGEMA_signal_5226, new_AGEMA_signal_5224, new_AGEMA_signal_5222}), .b ({new_AGEMA_signal_1610, new_AGEMA_signal_1609, SubCellInst_SboxInst_4_n5}), .clk (clk), .r ({Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_1760, new_AGEMA_signal_1759, Feedback[17]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U7 ( .a ({new_AGEMA_signal_5220, new_AGEMA_signal_5218, new_AGEMA_signal_5216}), .b ({new_AGEMA_signal_1332, new_AGEMA_signal_1331, SubCellInst_SboxInst_4_n2}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537]}), .c ({new_AGEMA_signal_1612, new_AGEMA_signal_1611, SubCellInst_SboxInst_4_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U19 ( .a ({new_AGEMA_signal_5232, new_AGEMA_signal_5230, new_AGEMA_signal_5228}), .b ({new_AGEMA_signal_1616, new_AGEMA_signal_1615, SubCellInst_SboxInst_5_n14}), .clk (clk), .r ({Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_1764, new_AGEMA_signal_1763, Feedback[23]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U16 ( .a ({new_AGEMA_signal_1336, new_AGEMA_signal_1335, SubCellInst_SboxInst_5_n11}), .b ({new_AGEMA_signal_5238, new_AGEMA_signal_5236, new_AGEMA_signal_5234}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543]}), .c ({new_AGEMA_signal_1618, new_AGEMA_signal_1617, SubCellInst_SboxInst_5_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U12 ( .a ({new_AGEMA_signal_5244, new_AGEMA_signal_5242, new_AGEMA_signal_5240}), .b ({new_AGEMA_signal_1620, new_AGEMA_signal_1619, SubCellInst_SboxInst_5_n5}), .clk (clk), .r ({Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_1768, new_AGEMA_signal_1767, Feedback[21]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U7 ( .a ({new_AGEMA_signal_5238, new_AGEMA_signal_5236, new_AGEMA_signal_5234}), .b ({new_AGEMA_signal_1344, new_AGEMA_signal_1343, SubCellInst_SboxInst_5_n2}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549]}), .c ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, SubCellInst_SboxInst_5_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U19 ( .a ({new_AGEMA_signal_5250, new_AGEMA_signal_5248, new_AGEMA_signal_5246}), .b ({new_AGEMA_signal_1626, new_AGEMA_signal_1625, SubCellInst_SboxInst_6_n14}), .clk (clk), .r ({Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_1772, new_AGEMA_signal_1771, Feedback[27]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U16 ( .a ({new_AGEMA_signal_1348, new_AGEMA_signal_1347, SubCellInst_SboxInst_6_n11}), .b ({new_AGEMA_signal_5256, new_AGEMA_signal_5254, new_AGEMA_signal_5252}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555]}), .c ({new_AGEMA_signal_1628, new_AGEMA_signal_1627, SubCellInst_SboxInst_6_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U12 ( .a ({new_AGEMA_signal_5262, new_AGEMA_signal_5260, new_AGEMA_signal_5258}), .b ({new_AGEMA_signal_1630, new_AGEMA_signal_1629, SubCellInst_SboxInst_6_n5}), .clk (clk), .r ({Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_1776, new_AGEMA_signal_1775, Feedback[25]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U7 ( .a ({new_AGEMA_signal_5256, new_AGEMA_signal_5254, new_AGEMA_signal_5252}), .b ({new_AGEMA_signal_1356, new_AGEMA_signal_1355, SubCellInst_SboxInst_6_n2}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561]}), .c ({new_AGEMA_signal_1632, new_AGEMA_signal_1631, SubCellInst_SboxInst_6_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U19 ( .a ({new_AGEMA_signal_5268, new_AGEMA_signal_5266, new_AGEMA_signal_5264}), .b ({new_AGEMA_signal_1636, new_AGEMA_signal_1635, SubCellInst_SboxInst_7_n14}), .clk (clk), .r ({Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_1780, new_AGEMA_signal_1779, Feedback[31]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U16 ( .a ({new_AGEMA_signal_1360, new_AGEMA_signal_1359, SubCellInst_SboxInst_7_n11}), .b ({new_AGEMA_signal_5274, new_AGEMA_signal_5272, new_AGEMA_signal_5270}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567]}), .c ({new_AGEMA_signal_1638, new_AGEMA_signal_1637, SubCellInst_SboxInst_7_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U12 ( .a ({new_AGEMA_signal_5280, new_AGEMA_signal_5278, new_AGEMA_signal_5276}), .b ({new_AGEMA_signal_1640, new_AGEMA_signal_1639, SubCellInst_SboxInst_7_n5}), .clk (clk), .r ({Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_1784, new_AGEMA_signal_1783, Feedback[29]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U7 ( .a ({new_AGEMA_signal_5274, new_AGEMA_signal_5272, new_AGEMA_signal_5270}), .b ({new_AGEMA_signal_1368, new_AGEMA_signal_1367, SubCellInst_SboxInst_7_n2}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573]}), .c ({new_AGEMA_signal_1642, new_AGEMA_signal_1641, SubCellInst_SboxInst_7_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U19 ( .a ({new_AGEMA_signal_5286, new_AGEMA_signal_5284, new_AGEMA_signal_5282}), .b ({new_AGEMA_signal_1646, new_AGEMA_signal_1645, SubCellInst_SboxInst_8_n14}), .clk (clk), .r ({Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, Feedback[35]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U16 ( .a ({new_AGEMA_signal_1372, new_AGEMA_signal_1371, SubCellInst_SboxInst_8_n11}), .b ({new_AGEMA_signal_5292, new_AGEMA_signal_5290, new_AGEMA_signal_5288}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579]}), .c ({new_AGEMA_signal_1648, new_AGEMA_signal_1647, SubCellInst_SboxInst_8_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U12 ( .a ({new_AGEMA_signal_5298, new_AGEMA_signal_5296, new_AGEMA_signal_5294}), .b ({new_AGEMA_signal_1650, new_AGEMA_signal_1649, SubCellInst_SboxInst_8_n5}), .clk (clk), .r ({Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_1792, new_AGEMA_signal_1791, Feedback[33]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U7 ( .a ({new_AGEMA_signal_5292, new_AGEMA_signal_5290, new_AGEMA_signal_5288}), .b ({new_AGEMA_signal_1380, new_AGEMA_signal_1379, SubCellInst_SboxInst_8_n2}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585]}), .c ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, SubCellInst_SboxInst_8_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U19 ( .a ({new_AGEMA_signal_5304, new_AGEMA_signal_5302, new_AGEMA_signal_5300}), .b ({new_AGEMA_signal_1656, new_AGEMA_signal_1655, SubCellInst_SboxInst_9_n14}), .clk (clk), .r ({Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, Feedback[39]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U16 ( .a ({new_AGEMA_signal_1384, new_AGEMA_signal_1383, SubCellInst_SboxInst_9_n11}), .b ({new_AGEMA_signal_5310, new_AGEMA_signal_5308, new_AGEMA_signal_5306}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591]}), .c ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, SubCellInst_SboxInst_9_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U12 ( .a ({new_AGEMA_signal_5316, new_AGEMA_signal_5314, new_AGEMA_signal_5312}), .b ({new_AGEMA_signal_1660, new_AGEMA_signal_1659, SubCellInst_SboxInst_9_n5}), .clk (clk), .r ({Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_1800, new_AGEMA_signal_1799, Feedback[37]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U7 ( .a ({new_AGEMA_signal_5310, new_AGEMA_signal_5308, new_AGEMA_signal_5306}), .b ({new_AGEMA_signal_1392, new_AGEMA_signal_1391, SubCellInst_SboxInst_9_n2}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597]}), .c ({new_AGEMA_signal_1662, new_AGEMA_signal_1661, SubCellInst_SboxInst_9_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U19 ( .a ({new_AGEMA_signal_5322, new_AGEMA_signal_5320, new_AGEMA_signal_5318}), .b ({new_AGEMA_signal_1666, new_AGEMA_signal_1665, SubCellInst_SboxInst_10_n14}), .clk (clk), .r ({Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_1804, new_AGEMA_signal_1803, Feedback[43]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U16 ( .a ({new_AGEMA_signal_1396, new_AGEMA_signal_1395, SubCellInst_SboxInst_10_n11}), .b ({new_AGEMA_signal_5328, new_AGEMA_signal_5326, new_AGEMA_signal_5324}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603]}), .c ({new_AGEMA_signal_1668, new_AGEMA_signal_1667, SubCellInst_SboxInst_10_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U12 ( .a ({new_AGEMA_signal_5334, new_AGEMA_signal_5332, new_AGEMA_signal_5330}), .b ({new_AGEMA_signal_1670, new_AGEMA_signal_1669, SubCellInst_SboxInst_10_n5}), .clk (clk), .r ({Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_1808, new_AGEMA_signal_1807, Feedback[41]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U7 ( .a ({new_AGEMA_signal_5328, new_AGEMA_signal_5326, new_AGEMA_signal_5324}), .b ({new_AGEMA_signal_1404, new_AGEMA_signal_1403, SubCellInst_SboxInst_10_n2}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609]}), .c ({new_AGEMA_signal_1672, new_AGEMA_signal_1671, SubCellInst_SboxInst_10_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U19 ( .a ({new_AGEMA_signal_5340, new_AGEMA_signal_5338, new_AGEMA_signal_5336}), .b ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, SubCellInst_SboxInst_11_n14}), .clk (clk), .r ({Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_1812, new_AGEMA_signal_1811, Feedback[47]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U16 ( .a ({new_AGEMA_signal_1408, new_AGEMA_signal_1407, SubCellInst_SboxInst_11_n11}), .b ({new_AGEMA_signal_5346, new_AGEMA_signal_5344, new_AGEMA_signal_5342}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615]}), .c ({new_AGEMA_signal_1678, new_AGEMA_signal_1677, SubCellInst_SboxInst_11_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U12 ( .a ({new_AGEMA_signal_5352, new_AGEMA_signal_5350, new_AGEMA_signal_5348}), .b ({new_AGEMA_signal_1680, new_AGEMA_signal_1679, SubCellInst_SboxInst_11_n5}), .clk (clk), .r ({Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_1816, new_AGEMA_signal_1815, Feedback[45]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U7 ( .a ({new_AGEMA_signal_5346, new_AGEMA_signal_5344, new_AGEMA_signal_5342}), .b ({new_AGEMA_signal_1416, new_AGEMA_signal_1415, SubCellInst_SboxInst_11_n2}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621]}), .c ({new_AGEMA_signal_1682, new_AGEMA_signal_1681, SubCellInst_SboxInst_11_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U19 ( .a ({new_AGEMA_signal_5358, new_AGEMA_signal_5356, new_AGEMA_signal_5354}), .b ({new_AGEMA_signal_1686, new_AGEMA_signal_1685, SubCellInst_SboxInst_12_n14}), .clk (clk), .r ({Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_1820, new_AGEMA_signal_1819, Feedback[51]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U16 ( .a ({new_AGEMA_signal_1420, new_AGEMA_signal_1419, SubCellInst_SboxInst_12_n11}), .b ({new_AGEMA_signal_5364, new_AGEMA_signal_5362, new_AGEMA_signal_5360}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627]}), .c ({new_AGEMA_signal_1688, new_AGEMA_signal_1687, SubCellInst_SboxInst_12_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U12 ( .a ({new_AGEMA_signal_5370, new_AGEMA_signal_5368, new_AGEMA_signal_5366}), .b ({new_AGEMA_signal_1690, new_AGEMA_signal_1689, SubCellInst_SboxInst_12_n5}), .clk (clk), .r ({Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_1824, new_AGEMA_signal_1823, Feedback[49]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U7 ( .a ({new_AGEMA_signal_5364, new_AGEMA_signal_5362, new_AGEMA_signal_5360}), .b ({new_AGEMA_signal_1428, new_AGEMA_signal_1427, SubCellInst_SboxInst_12_n2}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633]}), .c ({new_AGEMA_signal_1692, new_AGEMA_signal_1691, SubCellInst_SboxInst_12_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U19 ( .a ({new_AGEMA_signal_5376, new_AGEMA_signal_5374, new_AGEMA_signal_5372}), .b ({new_AGEMA_signal_1696, new_AGEMA_signal_1695, SubCellInst_SboxInst_13_n14}), .clk (clk), .r ({Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_1828, new_AGEMA_signal_1827, Feedback[55]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U16 ( .a ({new_AGEMA_signal_1432, new_AGEMA_signal_1431, SubCellInst_SboxInst_13_n11}), .b ({new_AGEMA_signal_5382, new_AGEMA_signal_5380, new_AGEMA_signal_5378}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639]}), .c ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, SubCellInst_SboxInst_13_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U12 ( .a ({new_AGEMA_signal_5388, new_AGEMA_signal_5386, new_AGEMA_signal_5384}), .b ({new_AGEMA_signal_1700, new_AGEMA_signal_1699, SubCellInst_SboxInst_13_n5}), .clk (clk), .r ({Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_1832, new_AGEMA_signal_1831, Feedback[53]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U7 ( .a ({new_AGEMA_signal_5382, new_AGEMA_signal_5380, new_AGEMA_signal_5378}), .b ({new_AGEMA_signal_1440, new_AGEMA_signal_1439, SubCellInst_SboxInst_13_n2}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645]}), .c ({new_AGEMA_signal_1702, new_AGEMA_signal_1701, SubCellInst_SboxInst_13_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U19 ( .a ({new_AGEMA_signal_5394, new_AGEMA_signal_5392, new_AGEMA_signal_5390}), .b ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, SubCellInst_SboxInst_14_n14}), .clk (clk), .r ({Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_1836, new_AGEMA_signal_1835, Feedback[59]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U16 ( .a ({new_AGEMA_signal_1444, new_AGEMA_signal_1443, SubCellInst_SboxInst_14_n11}), .b ({new_AGEMA_signal_5400, new_AGEMA_signal_5398, new_AGEMA_signal_5396}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651]}), .c ({new_AGEMA_signal_1708, new_AGEMA_signal_1707, SubCellInst_SboxInst_14_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U12 ( .a ({new_AGEMA_signal_5406, new_AGEMA_signal_5404, new_AGEMA_signal_5402}), .b ({new_AGEMA_signal_1710, new_AGEMA_signal_1709, SubCellInst_SboxInst_14_n5}), .clk (clk), .r ({Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_1840, new_AGEMA_signal_1839, Feedback[57]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U7 ( .a ({new_AGEMA_signal_5400, new_AGEMA_signal_5398, new_AGEMA_signal_5396}), .b ({new_AGEMA_signal_1452, new_AGEMA_signal_1451, SubCellInst_SboxInst_14_n2}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657]}), .c ({new_AGEMA_signal_1712, new_AGEMA_signal_1711, SubCellInst_SboxInst_14_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U19 ( .a ({new_AGEMA_signal_5412, new_AGEMA_signal_5410, new_AGEMA_signal_5408}), .b ({new_AGEMA_signal_1716, new_AGEMA_signal_1715, SubCellInst_SboxInst_15_n14}), .clk (clk), .r ({Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_1844, new_AGEMA_signal_1843, Feedback[63]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U16 ( .a ({new_AGEMA_signal_1456, new_AGEMA_signal_1455, SubCellInst_SboxInst_15_n11}), .b ({new_AGEMA_signal_5418, new_AGEMA_signal_5416, new_AGEMA_signal_5414}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663]}), .c ({new_AGEMA_signal_1718, new_AGEMA_signal_1717, SubCellInst_SboxInst_15_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U12 ( .a ({new_AGEMA_signal_5424, new_AGEMA_signal_5422, new_AGEMA_signal_5420}), .b ({new_AGEMA_signal_1720, new_AGEMA_signal_1719, SubCellInst_SboxInst_15_n5}), .clk (clk), .r ({Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_1848, new_AGEMA_signal_1847, Feedback[61]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U7 ( .a ({new_AGEMA_signal_5418, new_AGEMA_signal_5416, new_AGEMA_signal_5414}), .b ({new_AGEMA_signal_1464, new_AGEMA_signal_1463, SubCellInst_SboxInst_15_n2}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669]}), .c ({new_AGEMA_signal_1722, new_AGEMA_signal_1721, SubCellInst_SboxInst_15_n3}) ) ;
    buf_clk new_AGEMA_reg_buffer_1208 ( .C (clk), .D (new_AGEMA_signal_3983), .Q (new_AGEMA_signal_3984) ) ;
    buf_clk new_AGEMA_reg_buffer_1214 ( .C (clk), .D (new_AGEMA_signal_3989), .Q (new_AGEMA_signal_3990) ) ;
    buf_clk new_AGEMA_reg_buffer_1220 ( .C (clk), .D (new_AGEMA_signal_3995), .Q (new_AGEMA_signal_3996) ) ;
    buf_clk new_AGEMA_reg_buffer_1226 ( .C (clk), .D (new_AGEMA_signal_4001), .Q (new_AGEMA_signal_4002) ) ;
    buf_clk new_AGEMA_reg_buffer_1232 ( .C (clk), .D (new_AGEMA_signal_4007), .Q (new_AGEMA_signal_4008) ) ;
    buf_clk new_AGEMA_reg_buffer_1238 ( .C (clk), .D (new_AGEMA_signal_4013), .Q (new_AGEMA_signal_4014) ) ;
    buf_clk new_AGEMA_reg_buffer_1244 ( .C (clk), .D (new_AGEMA_signal_4019), .Q (new_AGEMA_signal_4020) ) ;
    buf_clk new_AGEMA_reg_buffer_1250 ( .C (clk), .D (new_AGEMA_signal_4025), .Q (new_AGEMA_signal_4026) ) ;
    buf_clk new_AGEMA_reg_buffer_1256 ( .C (clk), .D (new_AGEMA_signal_4031), .Q (new_AGEMA_signal_4032) ) ;
    buf_clk new_AGEMA_reg_buffer_1262 ( .C (clk), .D (new_AGEMA_signal_4037), .Q (new_AGEMA_signal_4038) ) ;
    buf_clk new_AGEMA_reg_buffer_1268 ( .C (clk), .D (new_AGEMA_signal_4043), .Q (new_AGEMA_signal_4044) ) ;
    buf_clk new_AGEMA_reg_buffer_1274 ( .C (clk), .D (new_AGEMA_signal_4049), .Q (new_AGEMA_signal_4050) ) ;
    buf_clk new_AGEMA_reg_buffer_1280 ( .C (clk), .D (new_AGEMA_signal_4055), .Q (new_AGEMA_signal_4056) ) ;
    buf_clk new_AGEMA_reg_buffer_1286 ( .C (clk), .D (new_AGEMA_signal_4061), .Q (new_AGEMA_signal_4062) ) ;
    buf_clk new_AGEMA_reg_buffer_1292 ( .C (clk), .D (new_AGEMA_signal_4067), .Q (new_AGEMA_signal_4068) ) ;
    buf_clk new_AGEMA_reg_buffer_1298 ( .C (clk), .D (new_AGEMA_signal_4073), .Q (new_AGEMA_signal_4074) ) ;
    buf_clk new_AGEMA_reg_buffer_1304 ( .C (clk), .D (new_AGEMA_signal_4079), .Q (new_AGEMA_signal_4080) ) ;
    buf_clk new_AGEMA_reg_buffer_1310 ( .C (clk), .D (new_AGEMA_signal_4085), .Q (new_AGEMA_signal_4086) ) ;
    buf_clk new_AGEMA_reg_buffer_1316 ( .C (clk), .D (new_AGEMA_signal_4091), .Q (new_AGEMA_signal_4092) ) ;
    buf_clk new_AGEMA_reg_buffer_1322 ( .C (clk), .D (new_AGEMA_signal_4097), .Q (new_AGEMA_signal_4098) ) ;
    buf_clk new_AGEMA_reg_buffer_1328 ( .C (clk), .D (new_AGEMA_signal_4103), .Q (new_AGEMA_signal_4104) ) ;
    buf_clk new_AGEMA_reg_buffer_1334 ( .C (clk), .D (new_AGEMA_signal_4109), .Q (new_AGEMA_signal_4110) ) ;
    buf_clk new_AGEMA_reg_buffer_1340 ( .C (clk), .D (new_AGEMA_signal_4115), .Q (new_AGEMA_signal_4116) ) ;
    buf_clk new_AGEMA_reg_buffer_1346 ( .C (clk), .D (new_AGEMA_signal_4121), .Q (new_AGEMA_signal_4122) ) ;
    buf_clk new_AGEMA_reg_buffer_1352 ( .C (clk), .D (new_AGEMA_signal_4127), .Q (new_AGEMA_signal_4128) ) ;
    buf_clk new_AGEMA_reg_buffer_1358 ( .C (clk), .D (new_AGEMA_signal_4133), .Q (new_AGEMA_signal_4134) ) ;
    buf_clk new_AGEMA_reg_buffer_1364 ( .C (clk), .D (new_AGEMA_signal_4139), .Q (new_AGEMA_signal_4140) ) ;
    buf_clk new_AGEMA_reg_buffer_1370 ( .C (clk), .D (new_AGEMA_signal_4145), .Q (new_AGEMA_signal_4146) ) ;
    buf_clk new_AGEMA_reg_buffer_1376 ( .C (clk), .D (new_AGEMA_signal_4151), .Q (new_AGEMA_signal_4152) ) ;
    buf_clk new_AGEMA_reg_buffer_1382 ( .C (clk), .D (new_AGEMA_signal_4157), .Q (new_AGEMA_signal_4158) ) ;
    buf_clk new_AGEMA_reg_buffer_1388 ( .C (clk), .D (new_AGEMA_signal_4163), .Q (new_AGEMA_signal_4164) ) ;
    buf_clk new_AGEMA_reg_buffer_1394 ( .C (clk), .D (new_AGEMA_signal_4169), .Q (new_AGEMA_signal_4170) ) ;
    buf_clk new_AGEMA_reg_buffer_1400 ( .C (clk), .D (new_AGEMA_signal_4175), .Q (new_AGEMA_signal_4176) ) ;
    buf_clk new_AGEMA_reg_buffer_1406 ( .C (clk), .D (new_AGEMA_signal_4181), .Q (new_AGEMA_signal_4182) ) ;
    buf_clk new_AGEMA_reg_buffer_1412 ( .C (clk), .D (new_AGEMA_signal_4187), .Q (new_AGEMA_signal_4188) ) ;
    buf_clk new_AGEMA_reg_buffer_1418 ( .C (clk), .D (new_AGEMA_signal_4193), .Q (new_AGEMA_signal_4194) ) ;
    buf_clk new_AGEMA_reg_buffer_1424 ( .C (clk), .D (new_AGEMA_signal_4199), .Q (new_AGEMA_signal_4200) ) ;
    buf_clk new_AGEMA_reg_buffer_1430 ( .C (clk), .D (new_AGEMA_signal_4205), .Q (new_AGEMA_signal_4206) ) ;
    buf_clk new_AGEMA_reg_buffer_1436 ( .C (clk), .D (new_AGEMA_signal_4211), .Q (new_AGEMA_signal_4212) ) ;
    buf_clk new_AGEMA_reg_buffer_1442 ( .C (clk), .D (new_AGEMA_signal_4217), .Q (new_AGEMA_signal_4218) ) ;
    buf_clk new_AGEMA_reg_buffer_1448 ( .C (clk), .D (new_AGEMA_signal_4223), .Q (new_AGEMA_signal_4224) ) ;
    buf_clk new_AGEMA_reg_buffer_1454 ( .C (clk), .D (new_AGEMA_signal_4229), .Q (new_AGEMA_signal_4230) ) ;
    buf_clk new_AGEMA_reg_buffer_1460 ( .C (clk), .D (new_AGEMA_signal_4235), .Q (new_AGEMA_signal_4236) ) ;
    buf_clk new_AGEMA_reg_buffer_1466 ( .C (clk), .D (new_AGEMA_signal_4241), .Q (new_AGEMA_signal_4242) ) ;
    buf_clk new_AGEMA_reg_buffer_1472 ( .C (clk), .D (new_AGEMA_signal_4247), .Q (new_AGEMA_signal_4248) ) ;
    buf_clk new_AGEMA_reg_buffer_1478 ( .C (clk), .D (new_AGEMA_signal_4253), .Q (new_AGEMA_signal_4254) ) ;
    buf_clk new_AGEMA_reg_buffer_1484 ( .C (clk), .D (new_AGEMA_signal_4259), .Q (new_AGEMA_signal_4260) ) ;
    buf_clk new_AGEMA_reg_buffer_1490 ( .C (clk), .D (new_AGEMA_signal_4265), .Q (new_AGEMA_signal_4266) ) ;
    buf_clk new_AGEMA_reg_buffer_1496 ( .C (clk), .D (new_AGEMA_signal_4271), .Q (new_AGEMA_signal_4272) ) ;
    buf_clk new_AGEMA_reg_buffer_1502 ( .C (clk), .D (new_AGEMA_signal_4277), .Q (new_AGEMA_signal_4278) ) ;
    buf_clk new_AGEMA_reg_buffer_1508 ( .C (clk), .D (new_AGEMA_signal_4283), .Q (new_AGEMA_signal_4284) ) ;
    buf_clk new_AGEMA_reg_buffer_1514 ( .C (clk), .D (new_AGEMA_signal_4289), .Q (new_AGEMA_signal_4290) ) ;
    buf_clk new_AGEMA_reg_buffer_1520 ( .C (clk), .D (new_AGEMA_signal_4295), .Q (new_AGEMA_signal_4296) ) ;
    buf_clk new_AGEMA_reg_buffer_1526 ( .C (clk), .D (new_AGEMA_signal_4301), .Q (new_AGEMA_signal_4302) ) ;
    buf_clk new_AGEMA_reg_buffer_1532 ( .C (clk), .D (new_AGEMA_signal_4307), .Q (new_AGEMA_signal_4308) ) ;
    buf_clk new_AGEMA_reg_buffer_1538 ( .C (clk), .D (new_AGEMA_signal_4313), .Q (new_AGEMA_signal_4314) ) ;
    buf_clk new_AGEMA_reg_buffer_1544 ( .C (clk), .D (new_AGEMA_signal_4319), .Q (new_AGEMA_signal_4320) ) ;
    buf_clk new_AGEMA_reg_buffer_1550 ( .C (clk), .D (new_AGEMA_signal_4325), .Q (new_AGEMA_signal_4326) ) ;
    buf_clk new_AGEMA_reg_buffer_1556 ( .C (clk), .D (new_AGEMA_signal_4331), .Q (new_AGEMA_signal_4332) ) ;
    buf_clk new_AGEMA_reg_buffer_1562 ( .C (clk), .D (new_AGEMA_signal_4337), .Q (new_AGEMA_signal_4338) ) ;
    buf_clk new_AGEMA_reg_buffer_1568 ( .C (clk), .D (new_AGEMA_signal_4343), .Q (new_AGEMA_signal_4344) ) ;
    buf_clk new_AGEMA_reg_buffer_1574 ( .C (clk), .D (new_AGEMA_signal_4349), .Q (new_AGEMA_signal_4350) ) ;
    buf_clk new_AGEMA_reg_buffer_1580 ( .C (clk), .D (new_AGEMA_signal_4355), .Q (new_AGEMA_signal_4356) ) ;
    buf_clk new_AGEMA_reg_buffer_1586 ( .C (clk), .D (new_AGEMA_signal_4361), .Q (new_AGEMA_signal_4362) ) ;
    buf_clk new_AGEMA_reg_buffer_1592 ( .C (clk), .D (new_AGEMA_signal_4367), .Q (new_AGEMA_signal_4368) ) ;
    buf_clk new_AGEMA_reg_buffer_1598 ( .C (clk), .D (new_AGEMA_signal_4373), .Q (new_AGEMA_signal_4374) ) ;
    buf_clk new_AGEMA_reg_buffer_1604 ( .C (clk), .D (new_AGEMA_signal_4379), .Q (new_AGEMA_signal_4380) ) ;
    buf_clk new_AGEMA_reg_buffer_1610 ( .C (clk), .D (new_AGEMA_signal_4385), .Q (new_AGEMA_signal_4386) ) ;
    buf_clk new_AGEMA_reg_buffer_1616 ( .C (clk), .D (new_AGEMA_signal_4391), .Q (new_AGEMA_signal_4392) ) ;
    buf_clk new_AGEMA_reg_buffer_1622 ( .C (clk), .D (new_AGEMA_signal_4397), .Q (new_AGEMA_signal_4398) ) ;
    buf_clk new_AGEMA_reg_buffer_1628 ( .C (clk), .D (new_AGEMA_signal_4403), .Q (new_AGEMA_signal_4404) ) ;
    buf_clk new_AGEMA_reg_buffer_1634 ( .C (clk), .D (new_AGEMA_signal_4409), .Q (new_AGEMA_signal_4410) ) ;
    buf_clk new_AGEMA_reg_buffer_1640 ( .C (clk), .D (new_AGEMA_signal_4415), .Q (new_AGEMA_signal_4416) ) ;
    buf_clk new_AGEMA_reg_buffer_1646 ( .C (clk), .D (new_AGEMA_signal_4421), .Q (new_AGEMA_signal_4422) ) ;
    buf_clk new_AGEMA_reg_buffer_1652 ( .C (clk), .D (new_AGEMA_signal_4427), .Q (new_AGEMA_signal_4428) ) ;
    buf_clk new_AGEMA_reg_buffer_1658 ( .C (clk), .D (new_AGEMA_signal_4433), .Q (new_AGEMA_signal_4434) ) ;
    buf_clk new_AGEMA_reg_buffer_1664 ( .C (clk), .D (new_AGEMA_signal_4439), .Q (new_AGEMA_signal_4440) ) ;
    buf_clk new_AGEMA_reg_buffer_1670 ( .C (clk), .D (new_AGEMA_signal_4445), .Q (new_AGEMA_signal_4446) ) ;
    buf_clk new_AGEMA_reg_buffer_1676 ( .C (clk), .D (new_AGEMA_signal_4451), .Q (new_AGEMA_signal_4452) ) ;
    buf_clk new_AGEMA_reg_buffer_1682 ( .C (clk), .D (new_AGEMA_signal_4457), .Q (new_AGEMA_signal_4458) ) ;
    buf_clk new_AGEMA_reg_buffer_1688 ( .C (clk), .D (new_AGEMA_signal_4463), .Q (new_AGEMA_signal_4464) ) ;
    buf_clk new_AGEMA_reg_buffer_1694 ( .C (clk), .D (new_AGEMA_signal_4469), .Q (new_AGEMA_signal_4470) ) ;
    buf_clk new_AGEMA_reg_buffer_1700 ( .C (clk), .D (new_AGEMA_signal_4475), .Q (new_AGEMA_signal_4476) ) ;
    buf_clk new_AGEMA_reg_buffer_1706 ( .C (clk), .D (new_AGEMA_signal_4481), .Q (new_AGEMA_signal_4482) ) ;
    buf_clk new_AGEMA_reg_buffer_1712 ( .C (clk), .D (new_AGEMA_signal_4487), .Q (new_AGEMA_signal_4488) ) ;
    buf_clk new_AGEMA_reg_buffer_1718 ( .C (clk), .D (new_AGEMA_signal_4493), .Q (new_AGEMA_signal_4494) ) ;
    buf_clk new_AGEMA_reg_buffer_1724 ( .C (clk), .D (new_AGEMA_signal_4499), .Q (new_AGEMA_signal_4500) ) ;
    buf_clk new_AGEMA_reg_buffer_1730 ( .C (clk), .D (new_AGEMA_signal_4505), .Q (new_AGEMA_signal_4506) ) ;
    buf_clk new_AGEMA_reg_buffer_1736 ( .C (clk), .D (new_AGEMA_signal_4511), .Q (new_AGEMA_signal_4512) ) ;
    buf_clk new_AGEMA_reg_buffer_1742 ( .C (clk), .D (new_AGEMA_signal_4517), .Q (new_AGEMA_signal_4518) ) ;
    buf_clk new_AGEMA_reg_buffer_1748 ( .C (clk), .D (new_AGEMA_signal_4523), .Q (new_AGEMA_signal_4524) ) ;
    buf_clk new_AGEMA_reg_buffer_1754 ( .C (clk), .D (new_AGEMA_signal_4529), .Q (new_AGEMA_signal_4530) ) ;
    buf_clk new_AGEMA_reg_buffer_1760 ( .C (clk), .D (new_AGEMA_signal_4535), .Q (new_AGEMA_signal_4536) ) ;
    buf_clk new_AGEMA_reg_buffer_1766 ( .C (clk), .D (new_AGEMA_signal_4541), .Q (new_AGEMA_signal_4542) ) ;
    buf_clk new_AGEMA_reg_buffer_1772 ( .C (clk), .D (new_AGEMA_signal_4547), .Q (new_AGEMA_signal_4548) ) ;
    buf_clk new_AGEMA_reg_buffer_1778 ( .C (clk), .D (new_AGEMA_signal_4553), .Q (new_AGEMA_signal_4554) ) ;
    buf_clk new_AGEMA_reg_buffer_1784 ( .C (clk), .D (new_AGEMA_signal_4559), .Q (new_AGEMA_signal_4560) ) ;
    buf_clk new_AGEMA_reg_buffer_1790 ( .C (clk), .D (new_AGEMA_signal_4565), .Q (new_AGEMA_signal_4566) ) ;
    buf_clk new_AGEMA_reg_buffer_1796 ( .C (clk), .D (new_AGEMA_signal_4571), .Q (new_AGEMA_signal_4572) ) ;
    buf_clk new_AGEMA_reg_buffer_1802 ( .C (clk), .D (new_AGEMA_signal_4577), .Q (new_AGEMA_signal_4578) ) ;
    buf_clk new_AGEMA_reg_buffer_1808 ( .C (clk), .D (new_AGEMA_signal_4583), .Q (new_AGEMA_signal_4584) ) ;
    buf_clk new_AGEMA_reg_buffer_1814 ( .C (clk), .D (new_AGEMA_signal_4589), .Q (new_AGEMA_signal_4590) ) ;
    buf_clk new_AGEMA_reg_buffer_1820 ( .C (clk), .D (new_AGEMA_signal_4595), .Q (new_AGEMA_signal_4596) ) ;
    buf_clk new_AGEMA_reg_buffer_1826 ( .C (clk), .D (new_AGEMA_signal_4601), .Q (new_AGEMA_signal_4602) ) ;
    buf_clk new_AGEMA_reg_buffer_1832 ( .C (clk), .D (new_AGEMA_signal_4607), .Q (new_AGEMA_signal_4608) ) ;
    buf_clk new_AGEMA_reg_buffer_1838 ( .C (clk), .D (new_AGEMA_signal_4613), .Q (new_AGEMA_signal_4614) ) ;
    buf_clk new_AGEMA_reg_buffer_1844 ( .C (clk), .D (new_AGEMA_signal_4619), .Q (new_AGEMA_signal_4620) ) ;
    buf_clk new_AGEMA_reg_buffer_1850 ( .C (clk), .D (new_AGEMA_signal_4625), .Q (new_AGEMA_signal_4626) ) ;
    buf_clk new_AGEMA_reg_buffer_1856 ( .C (clk), .D (new_AGEMA_signal_4631), .Q (new_AGEMA_signal_4632) ) ;
    buf_clk new_AGEMA_reg_buffer_1862 ( .C (clk), .D (new_AGEMA_signal_4637), .Q (new_AGEMA_signal_4638) ) ;
    buf_clk new_AGEMA_reg_buffer_1868 ( .C (clk), .D (new_AGEMA_signal_4643), .Q (new_AGEMA_signal_4644) ) ;
    buf_clk new_AGEMA_reg_buffer_1874 ( .C (clk), .D (new_AGEMA_signal_4649), .Q (new_AGEMA_signal_4650) ) ;
    buf_clk new_AGEMA_reg_buffer_1880 ( .C (clk), .D (new_AGEMA_signal_4655), .Q (new_AGEMA_signal_4656) ) ;
    buf_clk new_AGEMA_reg_buffer_1886 ( .C (clk), .D (new_AGEMA_signal_4661), .Q (new_AGEMA_signal_4662) ) ;
    buf_clk new_AGEMA_reg_buffer_1892 ( .C (clk), .D (new_AGEMA_signal_4667), .Q (new_AGEMA_signal_4668) ) ;
    buf_clk new_AGEMA_reg_buffer_1898 ( .C (clk), .D (new_AGEMA_signal_4673), .Q (new_AGEMA_signal_4674) ) ;
    buf_clk new_AGEMA_reg_buffer_1904 ( .C (clk), .D (new_AGEMA_signal_4679), .Q (new_AGEMA_signal_4680) ) ;
    buf_clk new_AGEMA_reg_buffer_1910 ( .C (clk), .D (new_AGEMA_signal_4685), .Q (new_AGEMA_signal_4686) ) ;
    buf_clk new_AGEMA_reg_buffer_1916 ( .C (clk), .D (new_AGEMA_signal_4691), .Q (new_AGEMA_signal_4692) ) ;
    buf_clk new_AGEMA_reg_buffer_1922 ( .C (clk), .D (new_AGEMA_signal_4697), .Q (new_AGEMA_signal_4698) ) ;
    buf_clk new_AGEMA_reg_buffer_1928 ( .C (clk), .D (new_AGEMA_signal_4703), .Q (new_AGEMA_signal_4704) ) ;
    buf_clk new_AGEMA_reg_buffer_1934 ( .C (clk), .D (new_AGEMA_signal_4709), .Q (new_AGEMA_signal_4710) ) ;
    buf_clk new_AGEMA_reg_buffer_1940 ( .C (clk), .D (new_AGEMA_signal_4715), .Q (new_AGEMA_signal_4716) ) ;
    buf_clk new_AGEMA_reg_buffer_1946 ( .C (clk), .D (new_AGEMA_signal_4721), .Q (new_AGEMA_signal_4722) ) ;
    buf_clk new_AGEMA_reg_buffer_1952 ( .C (clk), .D (new_AGEMA_signal_4727), .Q (new_AGEMA_signal_4728) ) ;
    buf_clk new_AGEMA_reg_buffer_1958 ( .C (clk), .D (new_AGEMA_signal_4733), .Q (new_AGEMA_signal_4734) ) ;
    buf_clk new_AGEMA_reg_buffer_1964 ( .C (clk), .D (new_AGEMA_signal_4739), .Q (new_AGEMA_signal_4740) ) ;
    buf_clk new_AGEMA_reg_buffer_1970 ( .C (clk), .D (new_AGEMA_signal_4745), .Q (new_AGEMA_signal_4746) ) ;
    buf_clk new_AGEMA_reg_buffer_1976 ( .C (clk), .D (new_AGEMA_signal_4751), .Q (new_AGEMA_signal_4752) ) ;
    buf_clk new_AGEMA_reg_buffer_1982 ( .C (clk), .D (new_AGEMA_signal_4757), .Q (new_AGEMA_signal_4758) ) ;
    buf_clk new_AGEMA_reg_buffer_1988 ( .C (clk), .D (new_AGEMA_signal_4763), .Q (new_AGEMA_signal_4764) ) ;
    buf_clk new_AGEMA_reg_buffer_1994 ( .C (clk), .D (new_AGEMA_signal_4769), .Q (new_AGEMA_signal_4770) ) ;
    buf_clk new_AGEMA_reg_buffer_2000 ( .C (clk), .D (new_AGEMA_signal_4775), .Q (new_AGEMA_signal_4776) ) ;
    buf_clk new_AGEMA_reg_buffer_2006 ( .C (clk), .D (new_AGEMA_signal_4781), .Q (new_AGEMA_signal_4782) ) ;
    buf_clk new_AGEMA_reg_buffer_2012 ( .C (clk), .D (new_AGEMA_signal_4787), .Q (new_AGEMA_signal_4788) ) ;
    buf_clk new_AGEMA_reg_buffer_2018 ( .C (clk), .D (new_AGEMA_signal_4793), .Q (new_AGEMA_signal_4794) ) ;
    buf_clk new_AGEMA_reg_buffer_2024 ( .C (clk), .D (new_AGEMA_signal_4799), .Q (new_AGEMA_signal_4800) ) ;
    buf_clk new_AGEMA_reg_buffer_2030 ( .C (clk), .D (new_AGEMA_signal_4805), .Q (new_AGEMA_signal_4806) ) ;
    buf_clk new_AGEMA_reg_buffer_2036 ( .C (clk), .D (new_AGEMA_signal_4811), .Q (new_AGEMA_signal_4812) ) ;
    buf_clk new_AGEMA_reg_buffer_2042 ( .C (clk), .D (new_AGEMA_signal_4817), .Q (new_AGEMA_signal_4818) ) ;
    buf_clk new_AGEMA_reg_buffer_2048 ( .C (clk), .D (new_AGEMA_signal_4823), .Q (new_AGEMA_signal_4824) ) ;
    buf_clk new_AGEMA_reg_buffer_2054 ( .C (clk), .D (new_AGEMA_signal_4829), .Q (new_AGEMA_signal_4830) ) ;
    buf_clk new_AGEMA_reg_buffer_2060 ( .C (clk), .D (new_AGEMA_signal_4835), .Q (new_AGEMA_signal_4836) ) ;
    buf_clk new_AGEMA_reg_buffer_2066 ( .C (clk), .D (new_AGEMA_signal_4841), .Q (new_AGEMA_signal_4842) ) ;
    buf_clk new_AGEMA_reg_buffer_2072 ( .C (clk), .D (new_AGEMA_signal_4847), .Q (new_AGEMA_signal_4848) ) ;
    buf_clk new_AGEMA_reg_buffer_2078 ( .C (clk), .D (new_AGEMA_signal_4853), .Q (new_AGEMA_signal_4854) ) ;
    buf_clk new_AGEMA_reg_buffer_2084 ( .C (clk), .D (new_AGEMA_signal_4859), .Q (new_AGEMA_signal_4860) ) ;
    buf_clk new_AGEMA_reg_buffer_2090 ( .C (clk), .D (new_AGEMA_signal_4865), .Q (new_AGEMA_signal_4866) ) ;
    buf_clk new_AGEMA_reg_buffer_2096 ( .C (clk), .D (new_AGEMA_signal_4871), .Q (new_AGEMA_signal_4872) ) ;
    buf_clk new_AGEMA_reg_buffer_2102 ( .C (clk), .D (new_AGEMA_signal_4877), .Q (new_AGEMA_signal_4878) ) ;
    buf_clk new_AGEMA_reg_buffer_2108 ( .C (clk), .D (new_AGEMA_signal_4883), .Q (new_AGEMA_signal_4884) ) ;
    buf_clk new_AGEMA_reg_buffer_2114 ( .C (clk), .D (new_AGEMA_signal_4889), .Q (new_AGEMA_signal_4890) ) ;
    buf_clk new_AGEMA_reg_buffer_2120 ( .C (clk), .D (new_AGEMA_signal_4895), .Q (new_AGEMA_signal_4896) ) ;
    buf_clk new_AGEMA_reg_buffer_2126 ( .C (clk), .D (new_AGEMA_signal_4901), .Q (new_AGEMA_signal_4902) ) ;
    buf_clk new_AGEMA_reg_buffer_2132 ( .C (clk), .D (new_AGEMA_signal_4907), .Q (new_AGEMA_signal_4908) ) ;
    buf_clk new_AGEMA_reg_buffer_2138 ( .C (clk), .D (new_AGEMA_signal_4913), .Q (new_AGEMA_signal_4914) ) ;
    buf_clk new_AGEMA_reg_buffer_2144 ( .C (clk), .D (new_AGEMA_signal_4919), .Q (new_AGEMA_signal_4920) ) ;
    buf_clk new_AGEMA_reg_buffer_2150 ( .C (clk), .D (new_AGEMA_signal_4925), .Q (new_AGEMA_signal_4926) ) ;
    buf_clk new_AGEMA_reg_buffer_2156 ( .C (clk), .D (new_AGEMA_signal_4931), .Q (new_AGEMA_signal_4932) ) ;
    buf_clk new_AGEMA_reg_buffer_2162 ( .C (clk), .D (new_AGEMA_signal_4937), .Q (new_AGEMA_signal_4938) ) ;
    buf_clk new_AGEMA_reg_buffer_2168 ( .C (clk), .D (new_AGEMA_signal_4943), .Q (new_AGEMA_signal_4944) ) ;
    buf_clk new_AGEMA_reg_buffer_2174 ( .C (clk), .D (new_AGEMA_signal_4949), .Q (new_AGEMA_signal_4950) ) ;
    buf_clk new_AGEMA_reg_buffer_2180 ( .C (clk), .D (new_AGEMA_signal_4955), .Q (new_AGEMA_signal_4956) ) ;
    buf_clk new_AGEMA_reg_buffer_2186 ( .C (clk), .D (new_AGEMA_signal_4961), .Q (new_AGEMA_signal_4962) ) ;
    buf_clk new_AGEMA_reg_buffer_2192 ( .C (clk), .D (new_AGEMA_signal_4967), .Q (new_AGEMA_signal_4968) ) ;
    buf_clk new_AGEMA_reg_buffer_2198 ( .C (clk), .D (new_AGEMA_signal_4973), .Q (new_AGEMA_signal_4974) ) ;
    buf_clk new_AGEMA_reg_buffer_2204 ( .C (clk), .D (new_AGEMA_signal_4979), .Q (new_AGEMA_signal_4980) ) ;
    buf_clk new_AGEMA_reg_buffer_2210 ( .C (clk), .D (new_AGEMA_signal_4985), .Q (new_AGEMA_signal_4986) ) ;
    buf_clk new_AGEMA_reg_buffer_2216 ( .C (clk), .D (new_AGEMA_signal_4991), .Q (new_AGEMA_signal_4992) ) ;
    buf_clk new_AGEMA_reg_buffer_2222 ( .C (clk), .D (new_AGEMA_signal_4997), .Q (new_AGEMA_signal_4998) ) ;
    buf_clk new_AGEMA_reg_buffer_2228 ( .C (clk), .D (new_AGEMA_signal_5003), .Q (new_AGEMA_signal_5004) ) ;
    buf_clk new_AGEMA_reg_buffer_2234 ( .C (clk), .D (new_AGEMA_signal_5009), .Q (new_AGEMA_signal_5010) ) ;
    buf_clk new_AGEMA_reg_buffer_2240 ( .C (clk), .D (new_AGEMA_signal_5015), .Q (new_AGEMA_signal_5016) ) ;
    buf_clk new_AGEMA_reg_buffer_2246 ( .C (clk), .D (new_AGEMA_signal_5021), .Q (new_AGEMA_signal_5022) ) ;
    buf_clk new_AGEMA_reg_buffer_2252 ( .C (clk), .D (new_AGEMA_signal_5027), .Q (new_AGEMA_signal_5028) ) ;
    buf_clk new_AGEMA_reg_buffer_2258 ( .C (clk), .D (new_AGEMA_signal_5033), .Q (new_AGEMA_signal_5034) ) ;
    buf_clk new_AGEMA_reg_buffer_2264 ( .C (clk), .D (new_AGEMA_signal_5039), .Q (new_AGEMA_signal_5040) ) ;
    buf_clk new_AGEMA_reg_buffer_2270 ( .C (clk), .D (new_AGEMA_signal_5045), .Q (new_AGEMA_signal_5046) ) ;
    buf_clk new_AGEMA_reg_buffer_2276 ( .C (clk), .D (new_AGEMA_signal_5051), .Q (new_AGEMA_signal_5052) ) ;
    buf_clk new_AGEMA_reg_buffer_2282 ( .C (clk), .D (new_AGEMA_signal_5057), .Q (new_AGEMA_signal_5058) ) ;
    buf_clk new_AGEMA_reg_buffer_2288 ( .C (clk), .D (new_AGEMA_signal_5063), .Q (new_AGEMA_signal_5064) ) ;
    buf_clk new_AGEMA_reg_buffer_2294 ( .C (clk), .D (new_AGEMA_signal_5069), .Q (new_AGEMA_signal_5070) ) ;
    buf_clk new_AGEMA_reg_buffer_2300 ( .C (clk), .D (new_AGEMA_signal_5075), .Q (new_AGEMA_signal_5076) ) ;
    buf_clk new_AGEMA_reg_buffer_2306 ( .C (clk), .D (new_AGEMA_signal_5081), .Q (new_AGEMA_signal_5082) ) ;
    buf_clk new_AGEMA_reg_buffer_2312 ( .C (clk), .D (new_AGEMA_signal_5087), .Q (new_AGEMA_signal_5088) ) ;
    buf_clk new_AGEMA_reg_buffer_2318 ( .C (clk), .D (new_AGEMA_signal_5093), .Q (new_AGEMA_signal_5094) ) ;
    buf_clk new_AGEMA_reg_buffer_2324 ( .C (clk), .D (new_AGEMA_signal_5099), .Q (new_AGEMA_signal_5100) ) ;
    buf_clk new_AGEMA_reg_buffer_2330 ( .C (clk), .D (new_AGEMA_signal_5105), .Q (new_AGEMA_signal_5106) ) ;
    buf_clk new_AGEMA_reg_buffer_2336 ( .C (clk), .D (new_AGEMA_signal_5111), .Q (new_AGEMA_signal_5112) ) ;
    buf_clk new_AGEMA_reg_buffer_2342 ( .C (clk), .D (new_AGEMA_signal_5117), .Q (new_AGEMA_signal_5118) ) ;
    buf_clk new_AGEMA_reg_buffer_2348 ( .C (clk), .D (new_AGEMA_signal_5123), .Q (new_AGEMA_signal_5124) ) ;
    buf_clk new_AGEMA_reg_buffer_2354 ( .C (clk), .D (new_AGEMA_signal_5129), .Q (new_AGEMA_signal_5130) ) ;
    buf_clk new_AGEMA_reg_buffer_2360 ( .C (clk), .D (new_AGEMA_signal_5135), .Q (new_AGEMA_signal_5136) ) ;
    buf_clk new_AGEMA_reg_buffer_2656 ( .C (clk), .D (new_AGEMA_signal_5431), .Q (new_AGEMA_signal_5432) ) ;
    buf_clk new_AGEMA_reg_buffer_2664 ( .C (clk), .D (new_AGEMA_signal_5439), .Q (new_AGEMA_signal_5440) ) ;
    buf_clk new_AGEMA_reg_buffer_2672 ( .C (clk), .D (new_AGEMA_signal_5447), .Q (new_AGEMA_signal_5448) ) ;
    buf_clk new_AGEMA_reg_buffer_2680 ( .C (clk), .D (new_AGEMA_signal_5455), .Q (new_AGEMA_signal_5456) ) ;
    buf_clk new_AGEMA_reg_buffer_2688 ( .C (clk), .D (new_AGEMA_signal_5463), .Q (new_AGEMA_signal_5464) ) ;
    buf_clk new_AGEMA_reg_buffer_2696 ( .C (clk), .D (new_AGEMA_signal_5471), .Q (new_AGEMA_signal_5472) ) ;
    buf_clk new_AGEMA_reg_buffer_2704 ( .C (clk), .D (new_AGEMA_signal_5479), .Q (new_AGEMA_signal_5480) ) ;
    buf_clk new_AGEMA_reg_buffer_2712 ( .C (clk), .D (new_AGEMA_signal_5487), .Q (new_AGEMA_signal_5488) ) ;
    buf_clk new_AGEMA_reg_buffer_2720 ( .C (clk), .D (new_AGEMA_signal_5495), .Q (new_AGEMA_signal_5496) ) ;
    buf_clk new_AGEMA_reg_buffer_2728 ( .C (clk), .D (new_AGEMA_signal_5503), .Q (new_AGEMA_signal_5504) ) ;
    buf_clk new_AGEMA_reg_buffer_2736 ( .C (clk), .D (new_AGEMA_signal_5511), .Q (new_AGEMA_signal_5512) ) ;
    buf_clk new_AGEMA_reg_buffer_2744 ( .C (clk), .D (new_AGEMA_signal_5519), .Q (new_AGEMA_signal_5520) ) ;
    buf_clk new_AGEMA_reg_buffer_2752 ( .C (clk), .D (new_AGEMA_signal_5527), .Q (new_AGEMA_signal_5528) ) ;
    buf_clk new_AGEMA_reg_buffer_2760 ( .C (clk), .D (new_AGEMA_signal_5535), .Q (new_AGEMA_signal_5536) ) ;
    buf_clk new_AGEMA_reg_buffer_2768 ( .C (clk), .D (new_AGEMA_signal_5543), .Q (new_AGEMA_signal_5544) ) ;
    buf_clk new_AGEMA_reg_buffer_2776 ( .C (clk), .D (new_AGEMA_signal_5551), .Q (new_AGEMA_signal_5552) ) ;
    buf_clk new_AGEMA_reg_buffer_2784 ( .C (clk), .D (new_AGEMA_signal_5559), .Q (new_AGEMA_signal_5560) ) ;
    buf_clk new_AGEMA_reg_buffer_2792 ( .C (clk), .D (new_AGEMA_signal_5567), .Q (new_AGEMA_signal_5568) ) ;
    buf_clk new_AGEMA_reg_buffer_2800 ( .C (clk), .D (new_AGEMA_signal_5575), .Q (new_AGEMA_signal_5576) ) ;
    buf_clk new_AGEMA_reg_buffer_2808 ( .C (clk), .D (new_AGEMA_signal_5583), .Q (new_AGEMA_signal_5584) ) ;
    buf_clk new_AGEMA_reg_buffer_2816 ( .C (clk), .D (new_AGEMA_signal_5591), .Q (new_AGEMA_signal_5592) ) ;
    buf_clk new_AGEMA_reg_buffer_2824 ( .C (clk), .D (new_AGEMA_signal_5599), .Q (new_AGEMA_signal_5600) ) ;
    buf_clk new_AGEMA_reg_buffer_2832 ( .C (clk), .D (new_AGEMA_signal_5607), .Q (new_AGEMA_signal_5608) ) ;
    buf_clk new_AGEMA_reg_buffer_2840 ( .C (clk), .D (new_AGEMA_signal_5615), .Q (new_AGEMA_signal_5616) ) ;
    buf_clk new_AGEMA_reg_buffer_2848 ( .C (clk), .D (new_AGEMA_signal_5623), .Q (new_AGEMA_signal_5624) ) ;
    buf_clk new_AGEMA_reg_buffer_2856 ( .C (clk), .D (new_AGEMA_signal_5631), .Q (new_AGEMA_signal_5632) ) ;
    buf_clk new_AGEMA_reg_buffer_2864 ( .C (clk), .D (new_AGEMA_signal_5639), .Q (new_AGEMA_signal_5640) ) ;
    buf_clk new_AGEMA_reg_buffer_2872 ( .C (clk), .D (new_AGEMA_signal_5647), .Q (new_AGEMA_signal_5648) ) ;
    buf_clk new_AGEMA_reg_buffer_2880 ( .C (clk), .D (new_AGEMA_signal_5655), .Q (new_AGEMA_signal_5656) ) ;
    buf_clk new_AGEMA_reg_buffer_2888 ( .C (clk), .D (new_AGEMA_signal_5663), .Q (new_AGEMA_signal_5664) ) ;
    buf_clk new_AGEMA_reg_buffer_2896 ( .C (clk), .D (new_AGEMA_signal_5671), .Q (new_AGEMA_signal_5672) ) ;
    buf_clk new_AGEMA_reg_buffer_2904 ( .C (clk), .D (new_AGEMA_signal_5679), .Q (new_AGEMA_signal_5680) ) ;
    buf_clk new_AGEMA_reg_buffer_2912 ( .C (clk), .D (new_AGEMA_signal_5687), .Q (new_AGEMA_signal_5688) ) ;
    buf_clk new_AGEMA_reg_buffer_2920 ( .C (clk), .D (new_AGEMA_signal_5695), .Q (new_AGEMA_signal_5696) ) ;
    buf_clk new_AGEMA_reg_buffer_2928 ( .C (clk), .D (new_AGEMA_signal_5703), .Q (new_AGEMA_signal_5704) ) ;
    buf_clk new_AGEMA_reg_buffer_2936 ( .C (clk), .D (new_AGEMA_signal_5711), .Q (new_AGEMA_signal_5712) ) ;
    buf_clk new_AGEMA_reg_buffer_2944 ( .C (clk), .D (new_AGEMA_signal_5719), .Q (new_AGEMA_signal_5720) ) ;
    buf_clk new_AGEMA_reg_buffer_2952 ( .C (clk), .D (new_AGEMA_signal_5727), .Q (new_AGEMA_signal_5728) ) ;
    buf_clk new_AGEMA_reg_buffer_2960 ( .C (clk), .D (new_AGEMA_signal_5735), .Q (new_AGEMA_signal_5736) ) ;
    buf_clk new_AGEMA_reg_buffer_2968 ( .C (clk), .D (new_AGEMA_signal_5743), .Q (new_AGEMA_signal_5744) ) ;
    buf_clk new_AGEMA_reg_buffer_2976 ( .C (clk), .D (new_AGEMA_signal_5751), .Q (new_AGEMA_signal_5752) ) ;
    buf_clk new_AGEMA_reg_buffer_2984 ( .C (clk), .D (new_AGEMA_signal_5759), .Q (new_AGEMA_signal_5760) ) ;
    buf_clk new_AGEMA_reg_buffer_2992 ( .C (clk), .D (new_AGEMA_signal_5767), .Q (new_AGEMA_signal_5768) ) ;
    buf_clk new_AGEMA_reg_buffer_3000 ( .C (clk), .D (new_AGEMA_signal_5775), .Q (new_AGEMA_signal_5776) ) ;
    buf_clk new_AGEMA_reg_buffer_3008 ( .C (clk), .D (new_AGEMA_signal_5783), .Q (new_AGEMA_signal_5784) ) ;
    buf_clk new_AGEMA_reg_buffer_3016 ( .C (clk), .D (new_AGEMA_signal_5791), .Q (new_AGEMA_signal_5792) ) ;
    buf_clk new_AGEMA_reg_buffer_3024 ( .C (clk), .D (new_AGEMA_signal_5799), .Q (new_AGEMA_signal_5800) ) ;
    buf_clk new_AGEMA_reg_buffer_3032 ( .C (clk), .D (new_AGEMA_signal_5807), .Q (new_AGEMA_signal_5808) ) ;
    buf_clk new_AGEMA_reg_buffer_3040 ( .C (clk), .D (new_AGEMA_signal_5815), .Q (new_AGEMA_signal_5816) ) ;
    buf_clk new_AGEMA_reg_buffer_3048 ( .C (clk), .D (new_AGEMA_signal_5823), .Q (new_AGEMA_signal_5824) ) ;
    buf_clk new_AGEMA_reg_buffer_3056 ( .C (clk), .D (new_AGEMA_signal_5831), .Q (new_AGEMA_signal_5832) ) ;
    buf_clk new_AGEMA_reg_buffer_3064 ( .C (clk), .D (new_AGEMA_signal_5839), .Q (new_AGEMA_signal_5840) ) ;
    buf_clk new_AGEMA_reg_buffer_3072 ( .C (clk), .D (new_AGEMA_signal_5847), .Q (new_AGEMA_signal_5848) ) ;
    buf_clk new_AGEMA_reg_buffer_3080 ( .C (clk), .D (new_AGEMA_signal_5855), .Q (new_AGEMA_signal_5856) ) ;
    buf_clk new_AGEMA_reg_buffer_3088 ( .C (clk), .D (new_AGEMA_signal_5863), .Q (new_AGEMA_signal_5864) ) ;
    buf_clk new_AGEMA_reg_buffer_3096 ( .C (clk), .D (new_AGEMA_signal_5871), .Q (new_AGEMA_signal_5872) ) ;
    buf_clk new_AGEMA_reg_buffer_3104 ( .C (clk), .D (new_AGEMA_signal_5879), .Q (new_AGEMA_signal_5880) ) ;
    buf_clk new_AGEMA_reg_buffer_3112 ( .C (clk), .D (new_AGEMA_signal_5887), .Q (new_AGEMA_signal_5888) ) ;
    buf_clk new_AGEMA_reg_buffer_3120 ( .C (clk), .D (new_AGEMA_signal_5895), .Q (new_AGEMA_signal_5896) ) ;
    buf_clk new_AGEMA_reg_buffer_3128 ( .C (clk), .D (new_AGEMA_signal_5903), .Q (new_AGEMA_signal_5904) ) ;
    buf_clk new_AGEMA_reg_buffer_3136 ( .C (clk), .D (new_AGEMA_signal_5911), .Q (new_AGEMA_signal_5912) ) ;
    buf_clk new_AGEMA_reg_buffer_3144 ( .C (clk), .D (new_AGEMA_signal_5919), .Q (new_AGEMA_signal_5920) ) ;
    buf_clk new_AGEMA_reg_buffer_3152 ( .C (clk), .D (new_AGEMA_signal_5927), .Q (new_AGEMA_signal_5928) ) ;
    buf_clk new_AGEMA_reg_buffer_3160 ( .C (clk), .D (new_AGEMA_signal_5935), .Q (new_AGEMA_signal_5936) ) ;
    buf_clk new_AGEMA_reg_buffer_3168 ( .C (clk), .D (new_AGEMA_signal_5943), .Q (new_AGEMA_signal_5944) ) ;
    buf_clk new_AGEMA_reg_buffer_3176 ( .C (clk), .D (new_AGEMA_signal_5951), .Q (new_AGEMA_signal_5952) ) ;
    buf_clk new_AGEMA_reg_buffer_3184 ( .C (clk), .D (new_AGEMA_signal_5959), .Q (new_AGEMA_signal_5960) ) ;
    buf_clk new_AGEMA_reg_buffer_3192 ( .C (clk), .D (new_AGEMA_signal_5967), .Q (new_AGEMA_signal_5968) ) ;
    buf_clk new_AGEMA_reg_buffer_3200 ( .C (clk), .D (new_AGEMA_signal_5975), .Q (new_AGEMA_signal_5976) ) ;
    buf_clk new_AGEMA_reg_buffer_3208 ( .C (clk), .D (new_AGEMA_signal_5983), .Q (new_AGEMA_signal_5984) ) ;
    buf_clk new_AGEMA_reg_buffer_3216 ( .C (clk), .D (new_AGEMA_signal_5991), .Q (new_AGEMA_signal_5992) ) ;
    buf_clk new_AGEMA_reg_buffer_3224 ( .C (clk), .D (new_AGEMA_signal_5999), .Q (new_AGEMA_signal_6000) ) ;
    buf_clk new_AGEMA_reg_buffer_3232 ( .C (clk), .D (new_AGEMA_signal_6007), .Q (new_AGEMA_signal_6008) ) ;
    buf_clk new_AGEMA_reg_buffer_3240 ( .C (clk), .D (new_AGEMA_signal_6015), .Q (new_AGEMA_signal_6016) ) ;
    buf_clk new_AGEMA_reg_buffer_3248 ( .C (clk), .D (new_AGEMA_signal_6023), .Q (new_AGEMA_signal_6024) ) ;
    buf_clk new_AGEMA_reg_buffer_3256 ( .C (clk), .D (new_AGEMA_signal_6031), .Q (new_AGEMA_signal_6032) ) ;
    buf_clk new_AGEMA_reg_buffer_3264 ( .C (clk), .D (new_AGEMA_signal_6039), .Q (new_AGEMA_signal_6040) ) ;
    buf_clk new_AGEMA_reg_buffer_3272 ( .C (clk), .D (new_AGEMA_signal_6047), .Q (new_AGEMA_signal_6048) ) ;
    buf_clk new_AGEMA_reg_buffer_3280 ( .C (clk), .D (new_AGEMA_signal_6055), .Q (new_AGEMA_signal_6056) ) ;
    buf_clk new_AGEMA_reg_buffer_3288 ( .C (clk), .D (new_AGEMA_signal_6063), .Q (new_AGEMA_signal_6064) ) ;
    buf_clk new_AGEMA_reg_buffer_3296 ( .C (clk), .D (new_AGEMA_signal_6071), .Q (new_AGEMA_signal_6072) ) ;
    buf_clk new_AGEMA_reg_buffer_3304 ( .C (clk), .D (new_AGEMA_signal_6079), .Q (new_AGEMA_signal_6080) ) ;
    buf_clk new_AGEMA_reg_buffer_3312 ( .C (clk), .D (new_AGEMA_signal_6087), .Q (new_AGEMA_signal_6088) ) ;
    buf_clk new_AGEMA_reg_buffer_3320 ( .C (clk), .D (new_AGEMA_signal_6095), .Q (new_AGEMA_signal_6096) ) ;
    buf_clk new_AGEMA_reg_buffer_3328 ( .C (clk), .D (new_AGEMA_signal_6103), .Q (new_AGEMA_signal_6104) ) ;
    buf_clk new_AGEMA_reg_buffer_3336 ( .C (clk), .D (new_AGEMA_signal_6111), .Q (new_AGEMA_signal_6112) ) ;
    buf_clk new_AGEMA_reg_buffer_3344 ( .C (clk), .D (new_AGEMA_signal_6119), .Q (new_AGEMA_signal_6120) ) ;
    buf_clk new_AGEMA_reg_buffer_3352 ( .C (clk), .D (new_AGEMA_signal_6127), .Q (new_AGEMA_signal_6128) ) ;
    buf_clk new_AGEMA_reg_buffer_3360 ( .C (clk), .D (new_AGEMA_signal_6135), .Q (new_AGEMA_signal_6136) ) ;
    buf_clk new_AGEMA_reg_buffer_3368 ( .C (clk), .D (new_AGEMA_signal_6143), .Q (new_AGEMA_signal_6144) ) ;
    buf_clk new_AGEMA_reg_buffer_3376 ( .C (clk), .D (new_AGEMA_signal_6151), .Q (new_AGEMA_signal_6152) ) ;
    buf_clk new_AGEMA_reg_buffer_3384 ( .C (clk), .D (new_AGEMA_signal_6159), .Q (new_AGEMA_signal_6160) ) ;
    buf_clk new_AGEMA_reg_buffer_3392 ( .C (clk), .D (new_AGEMA_signal_6167), .Q (new_AGEMA_signal_6168) ) ;
    buf_clk new_AGEMA_reg_buffer_3400 ( .C (clk), .D (new_AGEMA_signal_6175), .Q (new_AGEMA_signal_6176) ) ;
    buf_clk new_AGEMA_reg_buffer_3408 ( .C (clk), .D (new_AGEMA_signal_6183), .Q (new_AGEMA_signal_6184) ) ;
    buf_clk new_AGEMA_reg_buffer_3416 ( .C (clk), .D (new_AGEMA_signal_6191), .Q (new_AGEMA_signal_6192) ) ;
    buf_clk new_AGEMA_reg_buffer_3424 ( .C (clk), .D (new_AGEMA_signal_6199), .Q (new_AGEMA_signal_6200) ) ;
    buf_clk new_AGEMA_reg_buffer_3432 ( .C (clk), .D (new_AGEMA_signal_6207), .Q (new_AGEMA_signal_6208) ) ;
    buf_clk new_AGEMA_reg_buffer_3440 ( .C (clk), .D (new_AGEMA_signal_6215), .Q (new_AGEMA_signal_6216) ) ;
    buf_clk new_AGEMA_reg_buffer_3448 ( .C (clk), .D (new_AGEMA_signal_6223), .Q (new_AGEMA_signal_6224) ) ;
    buf_clk new_AGEMA_reg_buffer_3456 ( .C (clk), .D (new_AGEMA_signal_6231), .Q (new_AGEMA_signal_6232) ) ;
    buf_clk new_AGEMA_reg_buffer_3464 ( .C (clk), .D (new_AGEMA_signal_6239), .Q (new_AGEMA_signal_6240) ) ;
    buf_clk new_AGEMA_reg_buffer_3472 ( .C (clk), .D (new_AGEMA_signal_6247), .Q (new_AGEMA_signal_6248) ) ;
    buf_clk new_AGEMA_reg_buffer_3480 ( .C (clk), .D (new_AGEMA_signal_6255), .Q (new_AGEMA_signal_6256) ) ;
    buf_clk new_AGEMA_reg_buffer_3488 ( .C (clk), .D (new_AGEMA_signal_6263), .Q (new_AGEMA_signal_6264) ) ;
    buf_clk new_AGEMA_reg_buffer_3496 ( .C (clk), .D (new_AGEMA_signal_6271), .Q (new_AGEMA_signal_6272) ) ;
    buf_clk new_AGEMA_reg_buffer_3504 ( .C (clk), .D (new_AGEMA_signal_6279), .Q (new_AGEMA_signal_6280) ) ;
    buf_clk new_AGEMA_reg_buffer_3512 ( .C (clk), .D (new_AGEMA_signal_6287), .Q (new_AGEMA_signal_6288) ) ;
    buf_clk new_AGEMA_reg_buffer_3520 ( .C (clk), .D (new_AGEMA_signal_6295), .Q (new_AGEMA_signal_6296) ) ;
    buf_clk new_AGEMA_reg_buffer_3528 ( .C (clk), .D (new_AGEMA_signal_6303), .Q (new_AGEMA_signal_6304) ) ;
    buf_clk new_AGEMA_reg_buffer_3536 ( .C (clk), .D (new_AGEMA_signal_6311), .Q (new_AGEMA_signal_6312) ) ;
    buf_clk new_AGEMA_reg_buffer_3544 ( .C (clk), .D (new_AGEMA_signal_6319), .Q (new_AGEMA_signal_6320) ) ;
    buf_clk new_AGEMA_reg_buffer_3552 ( .C (clk), .D (new_AGEMA_signal_6327), .Q (new_AGEMA_signal_6328) ) ;
    buf_clk new_AGEMA_reg_buffer_3560 ( .C (clk), .D (new_AGEMA_signal_6335), .Q (new_AGEMA_signal_6336) ) ;
    buf_clk new_AGEMA_reg_buffer_3568 ( .C (clk), .D (new_AGEMA_signal_6343), .Q (new_AGEMA_signal_6344) ) ;
    buf_clk new_AGEMA_reg_buffer_3576 ( .C (clk), .D (new_AGEMA_signal_6351), .Q (new_AGEMA_signal_6352) ) ;
    buf_clk new_AGEMA_reg_buffer_3584 ( .C (clk), .D (new_AGEMA_signal_6359), .Q (new_AGEMA_signal_6360) ) ;
    buf_clk new_AGEMA_reg_buffer_3592 ( .C (clk), .D (new_AGEMA_signal_6367), .Q (new_AGEMA_signal_6368) ) ;
    buf_clk new_AGEMA_reg_buffer_3600 ( .C (clk), .D (new_AGEMA_signal_6375), .Q (new_AGEMA_signal_6376) ) ;
    buf_clk new_AGEMA_reg_buffer_3608 ( .C (clk), .D (new_AGEMA_signal_6383), .Q (new_AGEMA_signal_6384) ) ;
    buf_clk new_AGEMA_reg_buffer_3616 ( .C (clk), .D (new_AGEMA_signal_6391), .Q (new_AGEMA_signal_6392) ) ;
    buf_clk new_AGEMA_reg_buffer_3624 ( .C (clk), .D (new_AGEMA_signal_6399), .Q (new_AGEMA_signal_6400) ) ;
    buf_clk new_AGEMA_reg_buffer_3632 ( .C (clk), .D (new_AGEMA_signal_6407), .Q (new_AGEMA_signal_6408) ) ;
    buf_clk new_AGEMA_reg_buffer_3640 ( .C (clk), .D (new_AGEMA_signal_6415), .Q (new_AGEMA_signal_6416) ) ;
    buf_clk new_AGEMA_reg_buffer_3648 ( .C (clk), .D (new_AGEMA_signal_6423), .Q (new_AGEMA_signal_6424) ) ;
    buf_clk new_AGEMA_reg_buffer_3656 ( .C (clk), .D (new_AGEMA_signal_6431), .Q (new_AGEMA_signal_6432) ) ;
    buf_clk new_AGEMA_reg_buffer_3664 ( .C (clk), .D (new_AGEMA_signal_6439), .Q (new_AGEMA_signal_6440) ) ;
    buf_clk new_AGEMA_reg_buffer_3672 ( .C (clk), .D (new_AGEMA_signal_6447), .Q (new_AGEMA_signal_6448) ) ;
    buf_clk new_AGEMA_reg_buffer_3680 ( .C (clk), .D (new_AGEMA_signal_6455), .Q (new_AGEMA_signal_6456) ) ;
    buf_clk new_AGEMA_reg_buffer_3688 ( .C (clk), .D (new_AGEMA_signal_6463), .Q (new_AGEMA_signal_6464) ) ;
    buf_clk new_AGEMA_reg_buffer_3696 ( .C (clk), .D (new_AGEMA_signal_6471), .Q (new_AGEMA_signal_6472) ) ;
    buf_clk new_AGEMA_reg_buffer_3704 ( .C (clk), .D (new_AGEMA_signal_6479), .Q (new_AGEMA_signal_6480) ) ;
    buf_clk new_AGEMA_reg_buffer_3712 ( .C (clk), .D (new_AGEMA_signal_6487), .Q (new_AGEMA_signal_6488) ) ;
    buf_clk new_AGEMA_reg_buffer_3720 ( .C (clk), .D (new_AGEMA_signal_6495), .Q (new_AGEMA_signal_6496) ) ;
    buf_clk new_AGEMA_reg_buffer_3728 ( .C (clk), .D (new_AGEMA_signal_6503), .Q (new_AGEMA_signal_6504) ) ;
    buf_clk new_AGEMA_reg_buffer_3736 ( .C (clk), .D (new_AGEMA_signal_6511), .Q (new_AGEMA_signal_6512) ) ;
    buf_clk new_AGEMA_reg_buffer_3744 ( .C (clk), .D (new_AGEMA_signal_6519), .Q (new_AGEMA_signal_6520) ) ;
    buf_clk new_AGEMA_reg_buffer_3752 ( .C (clk), .D (new_AGEMA_signal_6527), .Q (new_AGEMA_signal_6528) ) ;
    buf_clk new_AGEMA_reg_buffer_3760 ( .C (clk), .D (new_AGEMA_signal_6535), .Q (new_AGEMA_signal_6536) ) ;
    buf_clk new_AGEMA_reg_buffer_3768 ( .C (clk), .D (new_AGEMA_signal_6543), .Q (new_AGEMA_signal_6544) ) ;
    buf_clk new_AGEMA_reg_buffer_3776 ( .C (clk), .D (new_AGEMA_signal_6551), .Q (new_AGEMA_signal_6552) ) ;
    buf_clk new_AGEMA_reg_buffer_3784 ( .C (clk), .D (new_AGEMA_signal_6559), .Q (new_AGEMA_signal_6560) ) ;
    buf_clk new_AGEMA_reg_buffer_3792 ( .C (clk), .D (new_AGEMA_signal_6567), .Q (new_AGEMA_signal_6568) ) ;
    buf_clk new_AGEMA_reg_buffer_3800 ( .C (clk), .D (new_AGEMA_signal_6575), .Q (new_AGEMA_signal_6576) ) ;
    buf_clk new_AGEMA_reg_buffer_3808 ( .C (clk), .D (new_AGEMA_signal_6583), .Q (new_AGEMA_signal_6584) ) ;
    buf_clk new_AGEMA_reg_buffer_3816 ( .C (clk), .D (new_AGEMA_signal_6591), .Q (new_AGEMA_signal_6592) ) ;
    buf_clk new_AGEMA_reg_buffer_3824 ( .C (clk), .D (new_AGEMA_signal_6599), .Q (new_AGEMA_signal_6600) ) ;
    buf_clk new_AGEMA_reg_buffer_3832 ( .C (clk), .D (new_AGEMA_signal_6607), .Q (new_AGEMA_signal_6608) ) ;
    buf_clk new_AGEMA_reg_buffer_3840 ( .C (clk), .D (new_AGEMA_signal_6615), .Q (new_AGEMA_signal_6616) ) ;
    buf_clk new_AGEMA_reg_buffer_3848 ( .C (clk), .D (new_AGEMA_signal_6623), .Q (new_AGEMA_signal_6624) ) ;
    buf_clk new_AGEMA_reg_buffer_3856 ( .C (clk), .D (new_AGEMA_signal_6631), .Q (new_AGEMA_signal_6632) ) ;
    buf_clk new_AGEMA_reg_buffer_3864 ( .C (clk), .D (new_AGEMA_signal_6639), .Q (new_AGEMA_signal_6640) ) ;
    buf_clk new_AGEMA_reg_buffer_3872 ( .C (clk), .D (new_AGEMA_signal_6647), .Q (new_AGEMA_signal_6648) ) ;
    buf_clk new_AGEMA_reg_buffer_3880 ( .C (clk), .D (new_AGEMA_signal_6655), .Q (new_AGEMA_signal_6656) ) ;
    buf_clk new_AGEMA_reg_buffer_3888 ( .C (clk), .D (new_AGEMA_signal_6663), .Q (new_AGEMA_signal_6664) ) ;
    buf_clk new_AGEMA_reg_buffer_3896 ( .C (clk), .D (new_AGEMA_signal_6671), .Q (new_AGEMA_signal_6672) ) ;
    buf_clk new_AGEMA_reg_buffer_3904 ( .C (clk), .D (new_AGEMA_signal_6679), .Q (new_AGEMA_signal_6680) ) ;
    buf_clk new_AGEMA_reg_buffer_3912 ( .C (clk), .D (new_AGEMA_signal_6687), .Q (new_AGEMA_signal_6688) ) ;
    buf_clk new_AGEMA_reg_buffer_3920 ( .C (clk), .D (new_AGEMA_signal_6695), .Q (new_AGEMA_signal_6696) ) ;
    buf_clk new_AGEMA_reg_buffer_3928 ( .C (clk), .D (new_AGEMA_signal_6703), .Q (new_AGEMA_signal_6704) ) ;
    buf_clk new_AGEMA_reg_buffer_3936 ( .C (clk), .D (new_AGEMA_signal_6711), .Q (new_AGEMA_signal_6712) ) ;
    buf_clk new_AGEMA_reg_buffer_3944 ( .C (clk), .D (new_AGEMA_signal_6719), .Q (new_AGEMA_signal_6720) ) ;
    buf_clk new_AGEMA_reg_buffer_3952 ( .C (clk), .D (new_AGEMA_signal_6727), .Q (new_AGEMA_signal_6728) ) ;
    buf_clk new_AGEMA_reg_buffer_3960 ( .C (clk), .D (new_AGEMA_signal_6735), .Q (new_AGEMA_signal_6736) ) ;
    buf_clk new_AGEMA_reg_buffer_3968 ( .C (clk), .D (new_AGEMA_signal_6743), .Q (new_AGEMA_signal_6744) ) ;
    buf_clk new_AGEMA_reg_buffer_3976 ( .C (clk), .D (new_AGEMA_signal_6751), .Q (new_AGEMA_signal_6752) ) ;
    buf_clk new_AGEMA_reg_buffer_3984 ( .C (clk), .D (new_AGEMA_signal_6759), .Q (new_AGEMA_signal_6760) ) ;
    buf_clk new_AGEMA_reg_buffer_3992 ( .C (clk), .D (new_AGEMA_signal_6767), .Q (new_AGEMA_signal_6768) ) ;
    buf_clk new_AGEMA_reg_buffer_4000 ( .C (clk), .D (new_AGEMA_signal_6775), .Q (new_AGEMA_signal_6776) ) ;
    buf_clk new_AGEMA_reg_buffer_4008 ( .C (clk), .D (new_AGEMA_signal_6783), .Q (new_AGEMA_signal_6784) ) ;
    buf_clk new_AGEMA_reg_buffer_4016 ( .C (clk), .D (new_AGEMA_signal_6791), .Q (new_AGEMA_signal_6792) ) ;
    buf_clk new_AGEMA_reg_buffer_4024 ( .C (clk), .D (new_AGEMA_signal_6799), .Q (new_AGEMA_signal_6800) ) ;
    buf_clk new_AGEMA_reg_buffer_4032 ( .C (clk), .D (new_AGEMA_signal_6807), .Q (new_AGEMA_signal_6808) ) ;
    buf_clk new_AGEMA_reg_buffer_4040 ( .C (clk), .D (new_AGEMA_signal_6815), .Q (new_AGEMA_signal_6816) ) ;
    buf_clk new_AGEMA_reg_buffer_4048 ( .C (clk), .D (new_AGEMA_signal_6823), .Q (new_AGEMA_signal_6824) ) ;
    buf_clk new_AGEMA_reg_buffer_4056 ( .C (clk), .D (new_AGEMA_signal_6831), .Q (new_AGEMA_signal_6832) ) ;
    buf_clk new_AGEMA_reg_buffer_4064 ( .C (clk), .D (new_AGEMA_signal_6839), .Q (new_AGEMA_signal_6840) ) ;
    buf_clk new_AGEMA_reg_buffer_4072 ( .C (clk), .D (new_AGEMA_signal_6847), .Q (new_AGEMA_signal_6848) ) ;
    buf_clk new_AGEMA_reg_buffer_4080 ( .C (clk), .D (new_AGEMA_signal_6855), .Q (new_AGEMA_signal_6856) ) ;
    buf_clk new_AGEMA_reg_buffer_4088 ( .C (clk), .D (new_AGEMA_signal_6863), .Q (new_AGEMA_signal_6864) ) ;
    buf_clk new_AGEMA_reg_buffer_4096 ( .C (clk), .D (new_AGEMA_signal_6871), .Q (new_AGEMA_signal_6872) ) ;
    buf_clk new_AGEMA_reg_buffer_4104 ( .C (clk), .D (new_AGEMA_signal_6879), .Q (new_AGEMA_signal_6880) ) ;
    buf_clk new_AGEMA_reg_buffer_4112 ( .C (clk), .D (new_AGEMA_signal_6887), .Q (new_AGEMA_signal_6888) ) ;
    buf_clk new_AGEMA_reg_buffer_4120 ( .C (clk), .D (new_AGEMA_signal_6895), .Q (new_AGEMA_signal_6896) ) ;
    buf_clk new_AGEMA_reg_buffer_4128 ( .C (clk), .D (new_AGEMA_signal_6903), .Q (new_AGEMA_signal_6904) ) ;
    buf_clk new_AGEMA_reg_buffer_4136 ( .C (clk), .D (new_AGEMA_signal_6911), .Q (new_AGEMA_signal_6912) ) ;
    buf_clk new_AGEMA_reg_buffer_4144 ( .C (clk), .D (new_AGEMA_signal_6919), .Q (new_AGEMA_signal_6920) ) ;
    buf_clk new_AGEMA_reg_buffer_4152 ( .C (clk), .D (new_AGEMA_signal_6927), .Q (new_AGEMA_signal_6928) ) ;
    buf_clk new_AGEMA_reg_buffer_4160 ( .C (clk), .D (new_AGEMA_signal_6935), .Q (new_AGEMA_signal_6936) ) ;
    buf_clk new_AGEMA_reg_buffer_4168 ( .C (clk), .D (new_AGEMA_signal_6943), .Q (new_AGEMA_signal_6944) ) ;
    buf_clk new_AGEMA_reg_buffer_4176 ( .C (clk), .D (new_AGEMA_signal_6951), .Q (new_AGEMA_signal_6952) ) ;
    buf_clk new_AGEMA_reg_buffer_4184 ( .C (clk), .D (new_AGEMA_signal_6959), .Q (new_AGEMA_signal_6960) ) ;
    buf_clk new_AGEMA_reg_buffer_4188 ( .C (clk), .D (new_AGEMA_signal_6963), .Q (new_AGEMA_signal_6964) ) ;
    buf_clk new_AGEMA_reg_buffer_4190 ( .C (clk), .D (new_AGEMA_signal_6965), .Q (new_AGEMA_signal_6966) ) ;
    buf_clk new_AGEMA_reg_buffer_4192 ( .C (clk), .D (new_AGEMA_signal_6967), .Q (new_AGEMA_signal_6968) ) ;
    buf_clk new_AGEMA_reg_buffer_4196 ( .C (clk), .D (new_AGEMA_signal_6971), .Q (new_AGEMA_signal_6972) ) ;
    buf_clk new_AGEMA_reg_buffer_4200 ( .C (clk), .D (new_AGEMA_signal_6975), .Q (new_AGEMA_signal_6976) ) ;
    buf_clk new_AGEMA_reg_buffer_4204 ( .C (clk), .D (new_AGEMA_signal_6979), .Q (new_AGEMA_signal_6980) ) ;
    buf_clk new_AGEMA_reg_buffer_4206 ( .C (clk), .D (new_AGEMA_signal_6981), .Q (new_AGEMA_signal_6982) ) ;
    buf_clk new_AGEMA_reg_buffer_4208 ( .C (clk), .D (new_AGEMA_signal_6983), .Q (new_AGEMA_signal_6984) ) ;
    buf_clk new_AGEMA_reg_buffer_4210 ( .C (clk), .D (new_AGEMA_signal_6985), .Q (new_AGEMA_signal_6986) ) ;
    buf_clk new_AGEMA_reg_buffer_4214 ( .C (clk), .D (new_AGEMA_signal_6989), .Q (new_AGEMA_signal_6990) ) ;
    buf_clk new_AGEMA_reg_buffer_4218 ( .C (clk), .D (new_AGEMA_signal_6993), .Q (new_AGEMA_signal_6994) ) ;
    buf_clk new_AGEMA_reg_buffer_4222 ( .C (clk), .D (new_AGEMA_signal_6997), .Q (new_AGEMA_signal_6998) ) ;
    buf_clk new_AGEMA_reg_buffer_4224 ( .C (clk), .D (new_AGEMA_signal_6999), .Q (new_AGEMA_signal_7000) ) ;
    buf_clk new_AGEMA_reg_buffer_4226 ( .C (clk), .D (new_AGEMA_signal_7001), .Q (new_AGEMA_signal_7002) ) ;
    buf_clk new_AGEMA_reg_buffer_4228 ( .C (clk), .D (new_AGEMA_signal_7003), .Q (new_AGEMA_signal_7004) ) ;
    buf_clk new_AGEMA_reg_buffer_4232 ( .C (clk), .D (new_AGEMA_signal_7007), .Q (new_AGEMA_signal_7008) ) ;
    buf_clk new_AGEMA_reg_buffer_4236 ( .C (clk), .D (new_AGEMA_signal_7011), .Q (new_AGEMA_signal_7012) ) ;
    buf_clk new_AGEMA_reg_buffer_4240 ( .C (clk), .D (new_AGEMA_signal_7015), .Q (new_AGEMA_signal_7016) ) ;
    buf_clk new_AGEMA_reg_buffer_4242 ( .C (clk), .D (new_AGEMA_signal_7017), .Q (new_AGEMA_signal_7018) ) ;
    buf_clk new_AGEMA_reg_buffer_4244 ( .C (clk), .D (new_AGEMA_signal_7019), .Q (new_AGEMA_signal_7020) ) ;
    buf_clk new_AGEMA_reg_buffer_4246 ( .C (clk), .D (new_AGEMA_signal_7021), .Q (new_AGEMA_signal_7022) ) ;
    buf_clk new_AGEMA_reg_buffer_4250 ( .C (clk), .D (new_AGEMA_signal_7025), .Q (new_AGEMA_signal_7026) ) ;
    buf_clk new_AGEMA_reg_buffer_4254 ( .C (clk), .D (new_AGEMA_signal_7029), .Q (new_AGEMA_signal_7030) ) ;
    buf_clk new_AGEMA_reg_buffer_4258 ( .C (clk), .D (new_AGEMA_signal_7033), .Q (new_AGEMA_signal_7034) ) ;
    buf_clk new_AGEMA_reg_buffer_4260 ( .C (clk), .D (new_AGEMA_signal_7035), .Q (new_AGEMA_signal_7036) ) ;
    buf_clk new_AGEMA_reg_buffer_4262 ( .C (clk), .D (new_AGEMA_signal_7037), .Q (new_AGEMA_signal_7038) ) ;
    buf_clk new_AGEMA_reg_buffer_4264 ( .C (clk), .D (new_AGEMA_signal_7039), .Q (new_AGEMA_signal_7040) ) ;
    buf_clk new_AGEMA_reg_buffer_4268 ( .C (clk), .D (new_AGEMA_signal_7043), .Q (new_AGEMA_signal_7044) ) ;
    buf_clk new_AGEMA_reg_buffer_4272 ( .C (clk), .D (new_AGEMA_signal_7047), .Q (new_AGEMA_signal_7048) ) ;
    buf_clk new_AGEMA_reg_buffer_4276 ( .C (clk), .D (new_AGEMA_signal_7051), .Q (new_AGEMA_signal_7052) ) ;
    buf_clk new_AGEMA_reg_buffer_4278 ( .C (clk), .D (new_AGEMA_signal_7053), .Q (new_AGEMA_signal_7054) ) ;
    buf_clk new_AGEMA_reg_buffer_4280 ( .C (clk), .D (new_AGEMA_signal_7055), .Q (new_AGEMA_signal_7056) ) ;
    buf_clk new_AGEMA_reg_buffer_4282 ( .C (clk), .D (new_AGEMA_signal_7057), .Q (new_AGEMA_signal_7058) ) ;
    buf_clk new_AGEMA_reg_buffer_4286 ( .C (clk), .D (new_AGEMA_signal_7061), .Q (new_AGEMA_signal_7062) ) ;
    buf_clk new_AGEMA_reg_buffer_4290 ( .C (clk), .D (new_AGEMA_signal_7065), .Q (new_AGEMA_signal_7066) ) ;
    buf_clk new_AGEMA_reg_buffer_4294 ( .C (clk), .D (new_AGEMA_signal_7069), .Q (new_AGEMA_signal_7070) ) ;
    buf_clk new_AGEMA_reg_buffer_4296 ( .C (clk), .D (new_AGEMA_signal_7071), .Q (new_AGEMA_signal_7072) ) ;
    buf_clk new_AGEMA_reg_buffer_4298 ( .C (clk), .D (new_AGEMA_signal_7073), .Q (new_AGEMA_signal_7074) ) ;
    buf_clk new_AGEMA_reg_buffer_4300 ( .C (clk), .D (new_AGEMA_signal_7075), .Q (new_AGEMA_signal_7076) ) ;
    buf_clk new_AGEMA_reg_buffer_4304 ( .C (clk), .D (new_AGEMA_signal_7079), .Q (new_AGEMA_signal_7080) ) ;
    buf_clk new_AGEMA_reg_buffer_4308 ( .C (clk), .D (new_AGEMA_signal_7083), .Q (new_AGEMA_signal_7084) ) ;
    buf_clk new_AGEMA_reg_buffer_4312 ( .C (clk), .D (new_AGEMA_signal_7087), .Q (new_AGEMA_signal_7088) ) ;
    buf_clk new_AGEMA_reg_buffer_4314 ( .C (clk), .D (new_AGEMA_signal_7089), .Q (new_AGEMA_signal_7090) ) ;
    buf_clk new_AGEMA_reg_buffer_4316 ( .C (clk), .D (new_AGEMA_signal_7091), .Q (new_AGEMA_signal_7092) ) ;
    buf_clk new_AGEMA_reg_buffer_4318 ( .C (clk), .D (new_AGEMA_signal_7093), .Q (new_AGEMA_signal_7094) ) ;
    buf_clk new_AGEMA_reg_buffer_4322 ( .C (clk), .D (new_AGEMA_signal_7097), .Q (new_AGEMA_signal_7098) ) ;
    buf_clk new_AGEMA_reg_buffer_4326 ( .C (clk), .D (new_AGEMA_signal_7101), .Q (new_AGEMA_signal_7102) ) ;
    buf_clk new_AGEMA_reg_buffer_4330 ( .C (clk), .D (new_AGEMA_signal_7105), .Q (new_AGEMA_signal_7106) ) ;
    buf_clk new_AGEMA_reg_buffer_4332 ( .C (clk), .D (new_AGEMA_signal_7107), .Q (new_AGEMA_signal_7108) ) ;
    buf_clk new_AGEMA_reg_buffer_4334 ( .C (clk), .D (new_AGEMA_signal_7109), .Q (new_AGEMA_signal_7110) ) ;
    buf_clk new_AGEMA_reg_buffer_4336 ( .C (clk), .D (new_AGEMA_signal_7111), .Q (new_AGEMA_signal_7112) ) ;
    buf_clk new_AGEMA_reg_buffer_4340 ( .C (clk), .D (new_AGEMA_signal_7115), .Q (new_AGEMA_signal_7116) ) ;
    buf_clk new_AGEMA_reg_buffer_4344 ( .C (clk), .D (new_AGEMA_signal_7119), .Q (new_AGEMA_signal_7120) ) ;
    buf_clk new_AGEMA_reg_buffer_4348 ( .C (clk), .D (new_AGEMA_signal_7123), .Q (new_AGEMA_signal_7124) ) ;
    buf_clk new_AGEMA_reg_buffer_4350 ( .C (clk), .D (new_AGEMA_signal_7125), .Q (new_AGEMA_signal_7126) ) ;
    buf_clk new_AGEMA_reg_buffer_4352 ( .C (clk), .D (new_AGEMA_signal_7127), .Q (new_AGEMA_signal_7128) ) ;
    buf_clk new_AGEMA_reg_buffer_4354 ( .C (clk), .D (new_AGEMA_signal_7129), .Q (new_AGEMA_signal_7130) ) ;
    buf_clk new_AGEMA_reg_buffer_4358 ( .C (clk), .D (new_AGEMA_signal_7133), .Q (new_AGEMA_signal_7134) ) ;
    buf_clk new_AGEMA_reg_buffer_4362 ( .C (clk), .D (new_AGEMA_signal_7137), .Q (new_AGEMA_signal_7138) ) ;
    buf_clk new_AGEMA_reg_buffer_4366 ( .C (clk), .D (new_AGEMA_signal_7141), .Q (new_AGEMA_signal_7142) ) ;
    buf_clk new_AGEMA_reg_buffer_4368 ( .C (clk), .D (new_AGEMA_signal_7143), .Q (new_AGEMA_signal_7144) ) ;
    buf_clk new_AGEMA_reg_buffer_4370 ( .C (clk), .D (new_AGEMA_signal_7145), .Q (new_AGEMA_signal_7146) ) ;
    buf_clk new_AGEMA_reg_buffer_4372 ( .C (clk), .D (new_AGEMA_signal_7147), .Q (new_AGEMA_signal_7148) ) ;
    buf_clk new_AGEMA_reg_buffer_4376 ( .C (clk), .D (new_AGEMA_signal_7151), .Q (new_AGEMA_signal_7152) ) ;
    buf_clk new_AGEMA_reg_buffer_4380 ( .C (clk), .D (new_AGEMA_signal_7155), .Q (new_AGEMA_signal_7156) ) ;
    buf_clk new_AGEMA_reg_buffer_4384 ( .C (clk), .D (new_AGEMA_signal_7159), .Q (new_AGEMA_signal_7160) ) ;
    buf_clk new_AGEMA_reg_buffer_4386 ( .C (clk), .D (new_AGEMA_signal_7161), .Q (new_AGEMA_signal_7162) ) ;
    buf_clk new_AGEMA_reg_buffer_4388 ( .C (clk), .D (new_AGEMA_signal_7163), .Q (new_AGEMA_signal_7164) ) ;
    buf_clk new_AGEMA_reg_buffer_4390 ( .C (clk), .D (new_AGEMA_signal_7165), .Q (new_AGEMA_signal_7166) ) ;
    buf_clk new_AGEMA_reg_buffer_4394 ( .C (clk), .D (new_AGEMA_signal_7169), .Q (new_AGEMA_signal_7170) ) ;
    buf_clk new_AGEMA_reg_buffer_4398 ( .C (clk), .D (new_AGEMA_signal_7173), .Q (new_AGEMA_signal_7174) ) ;
    buf_clk new_AGEMA_reg_buffer_4402 ( .C (clk), .D (new_AGEMA_signal_7177), .Q (new_AGEMA_signal_7178) ) ;
    buf_clk new_AGEMA_reg_buffer_4404 ( .C (clk), .D (new_AGEMA_signal_7179), .Q (new_AGEMA_signal_7180) ) ;
    buf_clk new_AGEMA_reg_buffer_4406 ( .C (clk), .D (new_AGEMA_signal_7181), .Q (new_AGEMA_signal_7182) ) ;
    buf_clk new_AGEMA_reg_buffer_4408 ( .C (clk), .D (new_AGEMA_signal_7183), .Q (new_AGEMA_signal_7184) ) ;
    buf_clk new_AGEMA_reg_buffer_4412 ( .C (clk), .D (new_AGEMA_signal_7187), .Q (new_AGEMA_signal_7188) ) ;
    buf_clk new_AGEMA_reg_buffer_4416 ( .C (clk), .D (new_AGEMA_signal_7191), .Q (new_AGEMA_signal_7192) ) ;
    buf_clk new_AGEMA_reg_buffer_4420 ( .C (clk), .D (new_AGEMA_signal_7195), .Q (new_AGEMA_signal_7196) ) ;
    buf_clk new_AGEMA_reg_buffer_4422 ( .C (clk), .D (new_AGEMA_signal_7197), .Q (new_AGEMA_signal_7198) ) ;
    buf_clk new_AGEMA_reg_buffer_4424 ( .C (clk), .D (new_AGEMA_signal_7199), .Q (new_AGEMA_signal_7200) ) ;
    buf_clk new_AGEMA_reg_buffer_4426 ( .C (clk), .D (new_AGEMA_signal_7201), .Q (new_AGEMA_signal_7202) ) ;
    buf_clk new_AGEMA_reg_buffer_4430 ( .C (clk), .D (new_AGEMA_signal_7205), .Q (new_AGEMA_signal_7206) ) ;
    buf_clk new_AGEMA_reg_buffer_4434 ( .C (clk), .D (new_AGEMA_signal_7209), .Q (new_AGEMA_signal_7210) ) ;
    buf_clk new_AGEMA_reg_buffer_4438 ( .C (clk), .D (new_AGEMA_signal_7213), .Q (new_AGEMA_signal_7214) ) ;
    buf_clk new_AGEMA_reg_buffer_4440 ( .C (clk), .D (new_AGEMA_signal_7215), .Q (new_AGEMA_signal_7216) ) ;
    buf_clk new_AGEMA_reg_buffer_4442 ( .C (clk), .D (new_AGEMA_signal_7217), .Q (new_AGEMA_signal_7218) ) ;
    buf_clk new_AGEMA_reg_buffer_4444 ( .C (clk), .D (new_AGEMA_signal_7219), .Q (new_AGEMA_signal_7220) ) ;
    buf_clk new_AGEMA_reg_buffer_4448 ( .C (clk), .D (new_AGEMA_signal_7223), .Q (new_AGEMA_signal_7224) ) ;
    buf_clk new_AGEMA_reg_buffer_4452 ( .C (clk), .D (new_AGEMA_signal_7227), .Q (new_AGEMA_signal_7228) ) ;
    buf_clk new_AGEMA_reg_buffer_4456 ( .C (clk), .D (new_AGEMA_signal_7231), .Q (new_AGEMA_signal_7232) ) ;
    buf_clk new_AGEMA_reg_buffer_4458 ( .C (clk), .D (new_AGEMA_signal_7233), .Q (new_AGEMA_signal_7234) ) ;
    buf_clk new_AGEMA_reg_buffer_4460 ( .C (clk), .D (new_AGEMA_signal_7235), .Q (new_AGEMA_signal_7236) ) ;
    buf_clk new_AGEMA_reg_buffer_4462 ( .C (clk), .D (new_AGEMA_signal_7237), .Q (new_AGEMA_signal_7238) ) ;
    buf_clk new_AGEMA_reg_buffer_4466 ( .C (clk), .D (new_AGEMA_signal_7241), .Q (new_AGEMA_signal_7242) ) ;
    buf_clk new_AGEMA_reg_buffer_4470 ( .C (clk), .D (new_AGEMA_signal_7245), .Q (new_AGEMA_signal_7246) ) ;
    buf_clk new_AGEMA_reg_buffer_4474 ( .C (clk), .D (new_AGEMA_signal_7249), .Q (new_AGEMA_signal_7250) ) ;
    buf_clk new_AGEMA_reg_buffer_4672 ( .C (clk), .D (new_AGEMA_signal_7447), .Q (new_AGEMA_signal_7448) ) ;
    buf_clk new_AGEMA_reg_buffer_4680 ( .C (clk), .D (new_AGEMA_signal_7455), .Q (new_AGEMA_signal_7456) ) ;
    buf_clk new_AGEMA_reg_buffer_4688 ( .C (clk), .D (new_AGEMA_signal_7463), .Q (new_AGEMA_signal_7464) ) ;
    buf_clk new_AGEMA_reg_buffer_4696 ( .C (clk), .D (new_AGEMA_signal_7471), .Q (new_AGEMA_signal_7472) ) ;
    buf_clk new_AGEMA_reg_buffer_4704 ( .C (clk), .D (new_AGEMA_signal_7479), .Q (new_AGEMA_signal_7480) ) ;
    buf_clk new_AGEMA_reg_buffer_4712 ( .C (clk), .D (new_AGEMA_signal_7487), .Q (new_AGEMA_signal_7488) ) ;
    buf_clk new_AGEMA_reg_buffer_4720 ( .C (clk), .D (new_AGEMA_signal_7495), .Q (new_AGEMA_signal_7496) ) ;
    buf_clk new_AGEMA_reg_buffer_4728 ( .C (clk), .D (new_AGEMA_signal_7503), .Q (new_AGEMA_signal_7504) ) ;
    buf_clk new_AGEMA_reg_buffer_4736 ( .C (clk), .D (new_AGEMA_signal_7511), .Q (new_AGEMA_signal_7512) ) ;
    buf_clk new_AGEMA_reg_buffer_4744 ( .C (clk), .D (new_AGEMA_signal_7519), .Q (new_AGEMA_signal_7520) ) ;

    /* cells in depth 7 */
    buf_clk new_AGEMA_reg_buffer_2649 ( .C (clk), .D (new_AGEMA_signal_3984), .Q (new_AGEMA_signal_5425) ) ;
    buf_clk new_AGEMA_reg_buffer_2657 ( .C (clk), .D (new_AGEMA_signal_5432), .Q (new_AGEMA_signal_5433) ) ;
    buf_clk new_AGEMA_reg_buffer_2665 ( .C (clk), .D (new_AGEMA_signal_5440), .Q (new_AGEMA_signal_5441) ) ;
    buf_clk new_AGEMA_reg_buffer_2673 ( .C (clk), .D (new_AGEMA_signal_5448), .Q (new_AGEMA_signal_5449) ) ;
    buf_clk new_AGEMA_reg_buffer_2681 ( .C (clk), .D (new_AGEMA_signal_5456), .Q (new_AGEMA_signal_5457) ) ;
    buf_clk new_AGEMA_reg_buffer_2689 ( .C (clk), .D (new_AGEMA_signal_5464), .Q (new_AGEMA_signal_5465) ) ;
    buf_clk new_AGEMA_reg_buffer_2697 ( .C (clk), .D (new_AGEMA_signal_5472), .Q (new_AGEMA_signal_5473) ) ;
    buf_clk new_AGEMA_reg_buffer_2705 ( .C (clk), .D (new_AGEMA_signal_5480), .Q (new_AGEMA_signal_5481) ) ;
    buf_clk new_AGEMA_reg_buffer_2713 ( .C (clk), .D (new_AGEMA_signal_5488), .Q (new_AGEMA_signal_5489) ) ;
    buf_clk new_AGEMA_reg_buffer_2721 ( .C (clk), .D (new_AGEMA_signal_5496), .Q (new_AGEMA_signal_5497) ) ;
    buf_clk new_AGEMA_reg_buffer_2729 ( .C (clk), .D (new_AGEMA_signal_5504), .Q (new_AGEMA_signal_5505) ) ;
    buf_clk new_AGEMA_reg_buffer_2737 ( .C (clk), .D (new_AGEMA_signal_5512), .Q (new_AGEMA_signal_5513) ) ;
    buf_clk new_AGEMA_reg_buffer_2745 ( .C (clk), .D (new_AGEMA_signal_5520), .Q (new_AGEMA_signal_5521) ) ;
    buf_clk new_AGEMA_reg_buffer_2753 ( .C (clk), .D (new_AGEMA_signal_5528), .Q (new_AGEMA_signal_5529) ) ;
    buf_clk new_AGEMA_reg_buffer_2761 ( .C (clk), .D (new_AGEMA_signal_5536), .Q (new_AGEMA_signal_5537) ) ;
    buf_clk new_AGEMA_reg_buffer_2769 ( .C (clk), .D (new_AGEMA_signal_5544), .Q (new_AGEMA_signal_5545) ) ;
    buf_clk new_AGEMA_reg_buffer_2777 ( .C (clk), .D (new_AGEMA_signal_5552), .Q (new_AGEMA_signal_5553) ) ;
    buf_clk new_AGEMA_reg_buffer_2785 ( .C (clk), .D (new_AGEMA_signal_5560), .Q (new_AGEMA_signal_5561) ) ;
    buf_clk new_AGEMA_reg_buffer_2793 ( .C (clk), .D (new_AGEMA_signal_5568), .Q (new_AGEMA_signal_5569) ) ;
    buf_clk new_AGEMA_reg_buffer_2801 ( .C (clk), .D (new_AGEMA_signal_5576), .Q (new_AGEMA_signal_5577) ) ;
    buf_clk new_AGEMA_reg_buffer_2809 ( .C (clk), .D (new_AGEMA_signal_5584), .Q (new_AGEMA_signal_5585) ) ;
    buf_clk new_AGEMA_reg_buffer_2817 ( .C (clk), .D (new_AGEMA_signal_5592), .Q (new_AGEMA_signal_5593) ) ;
    buf_clk new_AGEMA_reg_buffer_2825 ( .C (clk), .D (new_AGEMA_signal_5600), .Q (new_AGEMA_signal_5601) ) ;
    buf_clk new_AGEMA_reg_buffer_2833 ( .C (clk), .D (new_AGEMA_signal_5608), .Q (new_AGEMA_signal_5609) ) ;
    buf_clk new_AGEMA_reg_buffer_2841 ( .C (clk), .D (new_AGEMA_signal_5616), .Q (new_AGEMA_signal_5617) ) ;
    buf_clk new_AGEMA_reg_buffer_2849 ( .C (clk), .D (new_AGEMA_signal_5624), .Q (new_AGEMA_signal_5625) ) ;
    buf_clk new_AGEMA_reg_buffer_2857 ( .C (clk), .D (new_AGEMA_signal_5632), .Q (new_AGEMA_signal_5633) ) ;
    buf_clk new_AGEMA_reg_buffer_2865 ( .C (clk), .D (new_AGEMA_signal_5640), .Q (new_AGEMA_signal_5641) ) ;
    buf_clk new_AGEMA_reg_buffer_2873 ( .C (clk), .D (new_AGEMA_signal_5648), .Q (new_AGEMA_signal_5649) ) ;
    buf_clk new_AGEMA_reg_buffer_2881 ( .C (clk), .D (new_AGEMA_signal_5656), .Q (new_AGEMA_signal_5657) ) ;
    buf_clk new_AGEMA_reg_buffer_2889 ( .C (clk), .D (new_AGEMA_signal_5664), .Q (new_AGEMA_signal_5665) ) ;
    buf_clk new_AGEMA_reg_buffer_2897 ( .C (clk), .D (new_AGEMA_signal_5672), .Q (new_AGEMA_signal_5673) ) ;
    buf_clk new_AGEMA_reg_buffer_2905 ( .C (clk), .D (new_AGEMA_signal_5680), .Q (new_AGEMA_signal_5681) ) ;
    buf_clk new_AGEMA_reg_buffer_2913 ( .C (clk), .D (new_AGEMA_signal_5688), .Q (new_AGEMA_signal_5689) ) ;
    buf_clk new_AGEMA_reg_buffer_2921 ( .C (clk), .D (new_AGEMA_signal_5696), .Q (new_AGEMA_signal_5697) ) ;
    buf_clk new_AGEMA_reg_buffer_2929 ( .C (clk), .D (new_AGEMA_signal_5704), .Q (new_AGEMA_signal_5705) ) ;
    buf_clk new_AGEMA_reg_buffer_2937 ( .C (clk), .D (new_AGEMA_signal_5712), .Q (new_AGEMA_signal_5713) ) ;
    buf_clk new_AGEMA_reg_buffer_2945 ( .C (clk), .D (new_AGEMA_signal_5720), .Q (new_AGEMA_signal_5721) ) ;
    buf_clk new_AGEMA_reg_buffer_2953 ( .C (clk), .D (new_AGEMA_signal_5728), .Q (new_AGEMA_signal_5729) ) ;
    buf_clk new_AGEMA_reg_buffer_2961 ( .C (clk), .D (new_AGEMA_signal_5736), .Q (new_AGEMA_signal_5737) ) ;
    buf_clk new_AGEMA_reg_buffer_2969 ( .C (clk), .D (new_AGEMA_signal_5744), .Q (new_AGEMA_signal_5745) ) ;
    buf_clk new_AGEMA_reg_buffer_2977 ( .C (clk), .D (new_AGEMA_signal_5752), .Q (new_AGEMA_signal_5753) ) ;
    buf_clk new_AGEMA_reg_buffer_2985 ( .C (clk), .D (new_AGEMA_signal_5760), .Q (new_AGEMA_signal_5761) ) ;
    buf_clk new_AGEMA_reg_buffer_2993 ( .C (clk), .D (new_AGEMA_signal_5768), .Q (new_AGEMA_signal_5769) ) ;
    buf_clk new_AGEMA_reg_buffer_3001 ( .C (clk), .D (new_AGEMA_signal_5776), .Q (new_AGEMA_signal_5777) ) ;
    buf_clk new_AGEMA_reg_buffer_3009 ( .C (clk), .D (new_AGEMA_signal_5784), .Q (new_AGEMA_signal_5785) ) ;
    buf_clk new_AGEMA_reg_buffer_3017 ( .C (clk), .D (new_AGEMA_signal_5792), .Q (new_AGEMA_signal_5793) ) ;
    buf_clk new_AGEMA_reg_buffer_3025 ( .C (clk), .D (new_AGEMA_signal_5800), .Q (new_AGEMA_signal_5801) ) ;
    buf_clk new_AGEMA_reg_buffer_3033 ( .C (clk), .D (new_AGEMA_signal_5808), .Q (new_AGEMA_signal_5809) ) ;
    buf_clk new_AGEMA_reg_buffer_3041 ( .C (clk), .D (new_AGEMA_signal_5816), .Q (new_AGEMA_signal_5817) ) ;
    buf_clk new_AGEMA_reg_buffer_3049 ( .C (clk), .D (new_AGEMA_signal_5824), .Q (new_AGEMA_signal_5825) ) ;
    buf_clk new_AGEMA_reg_buffer_3057 ( .C (clk), .D (new_AGEMA_signal_5832), .Q (new_AGEMA_signal_5833) ) ;
    buf_clk new_AGEMA_reg_buffer_3065 ( .C (clk), .D (new_AGEMA_signal_5840), .Q (new_AGEMA_signal_5841) ) ;
    buf_clk new_AGEMA_reg_buffer_3073 ( .C (clk), .D (new_AGEMA_signal_5848), .Q (new_AGEMA_signal_5849) ) ;
    buf_clk new_AGEMA_reg_buffer_3081 ( .C (clk), .D (new_AGEMA_signal_5856), .Q (new_AGEMA_signal_5857) ) ;
    buf_clk new_AGEMA_reg_buffer_3089 ( .C (clk), .D (new_AGEMA_signal_5864), .Q (new_AGEMA_signal_5865) ) ;
    buf_clk new_AGEMA_reg_buffer_3097 ( .C (clk), .D (new_AGEMA_signal_5872), .Q (new_AGEMA_signal_5873) ) ;
    buf_clk new_AGEMA_reg_buffer_3105 ( .C (clk), .D (new_AGEMA_signal_5880), .Q (new_AGEMA_signal_5881) ) ;
    buf_clk new_AGEMA_reg_buffer_3113 ( .C (clk), .D (new_AGEMA_signal_5888), .Q (new_AGEMA_signal_5889) ) ;
    buf_clk new_AGEMA_reg_buffer_3121 ( .C (clk), .D (new_AGEMA_signal_5896), .Q (new_AGEMA_signal_5897) ) ;
    buf_clk new_AGEMA_reg_buffer_3129 ( .C (clk), .D (new_AGEMA_signal_5904), .Q (new_AGEMA_signal_5905) ) ;
    buf_clk new_AGEMA_reg_buffer_3137 ( .C (clk), .D (new_AGEMA_signal_5912), .Q (new_AGEMA_signal_5913) ) ;
    buf_clk new_AGEMA_reg_buffer_3145 ( .C (clk), .D (new_AGEMA_signal_5920), .Q (new_AGEMA_signal_5921) ) ;
    buf_clk new_AGEMA_reg_buffer_3153 ( .C (clk), .D (new_AGEMA_signal_5928), .Q (new_AGEMA_signal_5929) ) ;
    buf_clk new_AGEMA_reg_buffer_3161 ( .C (clk), .D (new_AGEMA_signal_5936), .Q (new_AGEMA_signal_5937) ) ;
    buf_clk new_AGEMA_reg_buffer_3169 ( .C (clk), .D (new_AGEMA_signal_5944), .Q (new_AGEMA_signal_5945) ) ;
    buf_clk new_AGEMA_reg_buffer_3177 ( .C (clk), .D (new_AGEMA_signal_5952), .Q (new_AGEMA_signal_5953) ) ;
    buf_clk new_AGEMA_reg_buffer_3185 ( .C (clk), .D (new_AGEMA_signal_5960), .Q (new_AGEMA_signal_5961) ) ;
    buf_clk new_AGEMA_reg_buffer_3193 ( .C (clk), .D (new_AGEMA_signal_5968), .Q (new_AGEMA_signal_5969) ) ;
    buf_clk new_AGEMA_reg_buffer_3201 ( .C (clk), .D (new_AGEMA_signal_5976), .Q (new_AGEMA_signal_5977) ) ;
    buf_clk new_AGEMA_reg_buffer_3209 ( .C (clk), .D (new_AGEMA_signal_5984), .Q (new_AGEMA_signal_5985) ) ;
    buf_clk new_AGEMA_reg_buffer_3217 ( .C (clk), .D (new_AGEMA_signal_5992), .Q (new_AGEMA_signal_5993) ) ;
    buf_clk new_AGEMA_reg_buffer_3225 ( .C (clk), .D (new_AGEMA_signal_6000), .Q (new_AGEMA_signal_6001) ) ;
    buf_clk new_AGEMA_reg_buffer_3233 ( .C (clk), .D (new_AGEMA_signal_6008), .Q (new_AGEMA_signal_6009) ) ;
    buf_clk new_AGEMA_reg_buffer_3241 ( .C (clk), .D (new_AGEMA_signal_6016), .Q (new_AGEMA_signal_6017) ) ;
    buf_clk new_AGEMA_reg_buffer_3249 ( .C (clk), .D (new_AGEMA_signal_6024), .Q (new_AGEMA_signal_6025) ) ;
    buf_clk new_AGEMA_reg_buffer_3257 ( .C (clk), .D (new_AGEMA_signal_6032), .Q (new_AGEMA_signal_6033) ) ;
    buf_clk new_AGEMA_reg_buffer_3265 ( .C (clk), .D (new_AGEMA_signal_6040), .Q (new_AGEMA_signal_6041) ) ;
    buf_clk new_AGEMA_reg_buffer_3273 ( .C (clk), .D (new_AGEMA_signal_6048), .Q (new_AGEMA_signal_6049) ) ;
    buf_clk new_AGEMA_reg_buffer_3281 ( .C (clk), .D (new_AGEMA_signal_6056), .Q (new_AGEMA_signal_6057) ) ;
    buf_clk new_AGEMA_reg_buffer_3289 ( .C (clk), .D (new_AGEMA_signal_6064), .Q (new_AGEMA_signal_6065) ) ;
    buf_clk new_AGEMA_reg_buffer_3297 ( .C (clk), .D (new_AGEMA_signal_6072), .Q (new_AGEMA_signal_6073) ) ;
    buf_clk new_AGEMA_reg_buffer_3305 ( .C (clk), .D (new_AGEMA_signal_6080), .Q (new_AGEMA_signal_6081) ) ;
    buf_clk new_AGEMA_reg_buffer_3313 ( .C (clk), .D (new_AGEMA_signal_6088), .Q (new_AGEMA_signal_6089) ) ;
    buf_clk new_AGEMA_reg_buffer_3321 ( .C (clk), .D (new_AGEMA_signal_6096), .Q (new_AGEMA_signal_6097) ) ;
    buf_clk new_AGEMA_reg_buffer_3329 ( .C (clk), .D (new_AGEMA_signal_6104), .Q (new_AGEMA_signal_6105) ) ;
    buf_clk new_AGEMA_reg_buffer_3337 ( .C (clk), .D (new_AGEMA_signal_6112), .Q (new_AGEMA_signal_6113) ) ;
    buf_clk new_AGEMA_reg_buffer_3345 ( .C (clk), .D (new_AGEMA_signal_6120), .Q (new_AGEMA_signal_6121) ) ;
    buf_clk new_AGEMA_reg_buffer_3353 ( .C (clk), .D (new_AGEMA_signal_6128), .Q (new_AGEMA_signal_6129) ) ;
    buf_clk new_AGEMA_reg_buffer_3361 ( .C (clk), .D (new_AGEMA_signal_6136), .Q (new_AGEMA_signal_6137) ) ;
    buf_clk new_AGEMA_reg_buffer_3369 ( .C (clk), .D (new_AGEMA_signal_6144), .Q (new_AGEMA_signal_6145) ) ;
    buf_clk new_AGEMA_reg_buffer_3377 ( .C (clk), .D (new_AGEMA_signal_6152), .Q (new_AGEMA_signal_6153) ) ;
    buf_clk new_AGEMA_reg_buffer_3385 ( .C (clk), .D (new_AGEMA_signal_6160), .Q (new_AGEMA_signal_6161) ) ;
    buf_clk new_AGEMA_reg_buffer_3393 ( .C (clk), .D (new_AGEMA_signal_6168), .Q (new_AGEMA_signal_6169) ) ;
    buf_clk new_AGEMA_reg_buffer_3401 ( .C (clk), .D (new_AGEMA_signal_6176), .Q (new_AGEMA_signal_6177) ) ;
    buf_clk new_AGEMA_reg_buffer_3409 ( .C (clk), .D (new_AGEMA_signal_6184), .Q (new_AGEMA_signal_6185) ) ;
    buf_clk new_AGEMA_reg_buffer_3417 ( .C (clk), .D (new_AGEMA_signal_6192), .Q (new_AGEMA_signal_6193) ) ;
    buf_clk new_AGEMA_reg_buffer_3425 ( .C (clk), .D (new_AGEMA_signal_6200), .Q (new_AGEMA_signal_6201) ) ;
    buf_clk new_AGEMA_reg_buffer_3433 ( .C (clk), .D (new_AGEMA_signal_6208), .Q (new_AGEMA_signal_6209) ) ;
    buf_clk new_AGEMA_reg_buffer_3441 ( .C (clk), .D (new_AGEMA_signal_6216), .Q (new_AGEMA_signal_6217) ) ;
    buf_clk new_AGEMA_reg_buffer_3449 ( .C (clk), .D (new_AGEMA_signal_6224), .Q (new_AGEMA_signal_6225) ) ;
    buf_clk new_AGEMA_reg_buffer_3457 ( .C (clk), .D (new_AGEMA_signal_6232), .Q (new_AGEMA_signal_6233) ) ;
    buf_clk new_AGEMA_reg_buffer_3465 ( .C (clk), .D (new_AGEMA_signal_6240), .Q (new_AGEMA_signal_6241) ) ;
    buf_clk new_AGEMA_reg_buffer_3473 ( .C (clk), .D (new_AGEMA_signal_6248), .Q (new_AGEMA_signal_6249) ) ;
    buf_clk new_AGEMA_reg_buffer_3481 ( .C (clk), .D (new_AGEMA_signal_6256), .Q (new_AGEMA_signal_6257) ) ;
    buf_clk new_AGEMA_reg_buffer_3489 ( .C (clk), .D (new_AGEMA_signal_6264), .Q (new_AGEMA_signal_6265) ) ;
    buf_clk new_AGEMA_reg_buffer_3497 ( .C (clk), .D (new_AGEMA_signal_6272), .Q (new_AGEMA_signal_6273) ) ;
    buf_clk new_AGEMA_reg_buffer_3505 ( .C (clk), .D (new_AGEMA_signal_6280), .Q (new_AGEMA_signal_6281) ) ;
    buf_clk new_AGEMA_reg_buffer_3513 ( .C (clk), .D (new_AGEMA_signal_6288), .Q (new_AGEMA_signal_6289) ) ;
    buf_clk new_AGEMA_reg_buffer_3521 ( .C (clk), .D (new_AGEMA_signal_6296), .Q (new_AGEMA_signal_6297) ) ;
    buf_clk new_AGEMA_reg_buffer_3529 ( .C (clk), .D (new_AGEMA_signal_6304), .Q (new_AGEMA_signal_6305) ) ;
    buf_clk new_AGEMA_reg_buffer_3537 ( .C (clk), .D (new_AGEMA_signal_6312), .Q (new_AGEMA_signal_6313) ) ;
    buf_clk new_AGEMA_reg_buffer_3545 ( .C (clk), .D (new_AGEMA_signal_6320), .Q (new_AGEMA_signal_6321) ) ;
    buf_clk new_AGEMA_reg_buffer_3553 ( .C (clk), .D (new_AGEMA_signal_6328), .Q (new_AGEMA_signal_6329) ) ;
    buf_clk new_AGEMA_reg_buffer_3561 ( .C (clk), .D (new_AGEMA_signal_6336), .Q (new_AGEMA_signal_6337) ) ;
    buf_clk new_AGEMA_reg_buffer_3569 ( .C (clk), .D (new_AGEMA_signal_6344), .Q (new_AGEMA_signal_6345) ) ;
    buf_clk new_AGEMA_reg_buffer_3577 ( .C (clk), .D (new_AGEMA_signal_6352), .Q (new_AGEMA_signal_6353) ) ;
    buf_clk new_AGEMA_reg_buffer_3585 ( .C (clk), .D (new_AGEMA_signal_6360), .Q (new_AGEMA_signal_6361) ) ;
    buf_clk new_AGEMA_reg_buffer_3593 ( .C (clk), .D (new_AGEMA_signal_6368), .Q (new_AGEMA_signal_6369) ) ;
    buf_clk new_AGEMA_reg_buffer_3601 ( .C (clk), .D (new_AGEMA_signal_6376), .Q (new_AGEMA_signal_6377) ) ;
    buf_clk new_AGEMA_reg_buffer_3609 ( .C (clk), .D (new_AGEMA_signal_6384), .Q (new_AGEMA_signal_6385) ) ;
    buf_clk new_AGEMA_reg_buffer_3617 ( .C (clk), .D (new_AGEMA_signal_6392), .Q (new_AGEMA_signal_6393) ) ;
    buf_clk new_AGEMA_reg_buffer_3625 ( .C (clk), .D (new_AGEMA_signal_6400), .Q (new_AGEMA_signal_6401) ) ;
    buf_clk new_AGEMA_reg_buffer_3633 ( .C (clk), .D (new_AGEMA_signal_6408), .Q (new_AGEMA_signal_6409) ) ;
    buf_clk new_AGEMA_reg_buffer_3641 ( .C (clk), .D (new_AGEMA_signal_6416), .Q (new_AGEMA_signal_6417) ) ;
    buf_clk new_AGEMA_reg_buffer_3649 ( .C (clk), .D (new_AGEMA_signal_6424), .Q (new_AGEMA_signal_6425) ) ;
    buf_clk new_AGEMA_reg_buffer_3657 ( .C (clk), .D (new_AGEMA_signal_6432), .Q (new_AGEMA_signal_6433) ) ;
    buf_clk new_AGEMA_reg_buffer_3665 ( .C (clk), .D (new_AGEMA_signal_6440), .Q (new_AGEMA_signal_6441) ) ;
    buf_clk new_AGEMA_reg_buffer_3673 ( .C (clk), .D (new_AGEMA_signal_6448), .Q (new_AGEMA_signal_6449) ) ;
    buf_clk new_AGEMA_reg_buffer_3681 ( .C (clk), .D (new_AGEMA_signal_6456), .Q (new_AGEMA_signal_6457) ) ;
    buf_clk new_AGEMA_reg_buffer_3689 ( .C (clk), .D (new_AGEMA_signal_6464), .Q (new_AGEMA_signal_6465) ) ;
    buf_clk new_AGEMA_reg_buffer_3697 ( .C (clk), .D (new_AGEMA_signal_6472), .Q (new_AGEMA_signal_6473) ) ;
    buf_clk new_AGEMA_reg_buffer_3705 ( .C (clk), .D (new_AGEMA_signal_6480), .Q (new_AGEMA_signal_6481) ) ;
    buf_clk new_AGEMA_reg_buffer_3713 ( .C (clk), .D (new_AGEMA_signal_6488), .Q (new_AGEMA_signal_6489) ) ;
    buf_clk new_AGEMA_reg_buffer_3721 ( .C (clk), .D (new_AGEMA_signal_6496), .Q (new_AGEMA_signal_6497) ) ;
    buf_clk new_AGEMA_reg_buffer_3729 ( .C (clk), .D (new_AGEMA_signal_6504), .Q (new_AGEMA_signal_6505) ) ;
    buf_clk new_AGEMA_reg_buffer_3737 ( .C (clk), .D (new_AGEMA_signal_6512), .Q (new_AGEMA_signal_6513) ) ;
    buf_clk new_AGEMA_reg_buffer_3745 ( .C (clk), .D (new_AGEMA_signal_6520), .Q (new_AGEMA_signal_6521) ) ;
    buf_clk new_AGEMA_reg_buffer_3753 ( .C (clk), .D (new_AGEMA_signal_6528), .Q (new_AGEMA_signal_6529) ) ;
    buf_clk new_AGEMA_reg_buffer_3761 ( .C (clk), .D (new_AGEMA_signal_6536), .Q (new_AGEMA_signal_6537) ) ;
    buf_clk new_AGEMA_reg_buffer_3769 ( .C (clk), .D (new_AGEMA_signal_6544), .Q (new_AGEMA_signal_6545) ) ;
    buf_clk new_AGEMA_reg_buffer_3777 ( .C (clk), .D (new_AGEMA_signal_6552), .Q (new_AGEMA_signal_6553) ) ;
    buf_clk new_AGEMA_reg_buffer_3785 ( .C (clk), .D (new_AGEMA_signal_6560), .Q (new_AGEMA_signal_6561) ) ;
    buf_clk new_AGEMA_reg_buffer_3793 ( .C (clk), .D (new_AGEMA_signal_6568), .Q (new_AGEMA_signal_6569) ) ;
    buf_clk new_AGEMA_reg_buffer_3801 ( .C (clk), .D (new_AGEMA_signal_6576), .Q (new_AGEMA_signal_6577) ) ;
    buf_clk new_AGEMA_reg_buffer_3809 ( .C (clk), .D (new_AGEMA_signal_6584), .Q (new_AGEMA_signal_6585) ) ;
    buf_clk new_AGEMA_reg_buffer_3817 ( .C (clk), .D (new_AGEMA_signal_6592), .Q (new_AGEMA_signal_6593) ) ;
    buf_clk new_AGEMA_reg_buffer_3825 ( .C (clk), .D (new_AGEMA_signal_6600), .Q (new_AGEMA_signal_6601) ) ;
    buf_clk new_AGEMA_reg_buffer_3833 ( .C (clk), .D (new_AGEMA_signal_6608), .Q (new_AGEMA_signal_6609) ) ;
    buf_clk new_AGEMA_reg_buffer_3841 ( .C (clk), .D (new_AGEMA_signal_6616), .Q (new_AGEMA_signal_6617) ) ;
    buf_clk new_AGEMA_reg_buffer_3849 ( .C (clk), .D (new_AGEMA_signal_6624), .Q (new_AGEMA_signal_6625) ) ;
    buf_clk new_AGEMA_reg_buffer_3857 ( .C (clk), .D (new_AGEMA_signal_6632), .Q (new_AGEMA_signal_6633) ) ;
    buf_clk new_AGEMA_reg_buffer_3865 ( .C (clk), .D (new_AGEMA_signal_6640), .Q (new_AGEMA_signal_6641) ) ;
    buf_clk new_AGEMA_reg_buffer_3873 ( .C (clk), .D (new_AGEMA_signal_6648), .Q (new_AGEMA_signal_6649) ) ;
    buf_clk new_AGEMA_reg_buffer_3881 ( .C (clk), .D (new_AGEMA_signal_6656), .Q (new_AGEMA_signal_6657) ) ;
    buf_clk new_AGEMA_reg_buffer_3889 ( .C (clk), .D (new_AGEMA_signal_6664), .Q (new_AGEMA_signal_6665) ) ;
    buf_clk new_AGEMA_reg_buffer_3897 ( .C (clk), .D (new_AGEMA_signal_6672), .Q (new_AGEMA_signal_6673) ) ;
    buf_clk new_AGEMA_reg_buffer_3905 ( .C (clk), .D (new_AGEMA_signal_6680), .Q (new_AGEMA_signal_6681) ) ;
    buf_clk new_AGEMA_reg_buffer_3913 ( .C (clk), .D (new_AGEMA_signal_6688), .Q (new_AGEMA_signal_6689) ) ;
    buf_clk new_AGEMA_reg_buffer_3921 ( .C (clk), .D (new_AGEMA_signal_6696), .Q (new_AGEMA_signal_6697) ) ;
    buf_clk new_AGEMA_reg_buffer_3929 ( .C (clk), .D (new_AGEMA_signal_6704), .Q (new_AGEMA_signal_6705) ) ;
    buf_clk new_AGEMA_reg_buffer_3937 ( .C (clk), .D (new_AGEMA_signal_6712), .Q (new_AGEMA_signal_6713) ) ;
    buf_clk new_AGEMA_reg_buffer_3945 ( .C (clk), .D (new_AGEMA_signal_6720), .Q (new_AGEMA_signal_6721) ) ;
    buf_clk new_AGEMA_reg_buffer_3953 ( .C (clk), .D (new_AGEMA_signal_6728), .Q (new_AGEMA_signal_6729) ) ;
    buf_clk new_AGEMA_reg_buffer_3961 ( .C (clk), .D (new_AGEMA_signal_6736), .Q (new_AGEMA_signal_6737) ) ;
    buf_clk new_AGEMA_reg_buffer_3969 ( .C (clk), .D (new_AGEMA_signal_6744), .Q (new_AGEMA_signal_6745) ) ;
    buf_clk new_AGEMA_reg_buffer_3977 ( .C (clk), .D (new_AGEMA_signal_6752), .Q (new_AGEMA_signal_6753) ) ;
    buf_clk new_AGEMA_reg_buffer_3985 ( .C (clk), .D (new_AGEMA_signal_6760), .Q (new_AGEMA_signal_6761) ) ;
    buf_clk new_AGEMA_reg_buffer_3993 ( .C (clk), .D (new_AGEMA_signal_6768), .Q (new_AGEMA_signal_6769) ) ;
    buf_clk new_AGEMA_reg_buffer_4001 ( .C (clk), .D (new_AGEMA_signal_6776), .Q (new_AGEMA_signal_6777) ) ;
    buf_clk new_AGEMA_reg_buffer_4009 ( .C (clk), .D (new_AGEMA_signal_6784), .Q (new_AGEMA_signal_6785) ) ;
    buf_clk new_AGEMA_reg_buffer_4017 ( .C (clk), .D (new_AGEMA_signal_6792), .Q (new_AGEMA_signal_6793) ) ;
    buf_clk new_AGEMA_reg_buffer_4025 ( .C (clk), .D (new_AGEMA_signal_6800), .Q (new_AGEMA_signal_6801) ) ;
    buf_clk new_AGEMA_reg_buffer_4033 ( .C (clk), .D (new_AGEMA_signal_6808), .Q (new_AGEMA_signal_6809) ) ;
    buf_clk new_AGEMA_reg_buffer_4041 ( .C (clk), .D (new_AGEMA_signal_6816), .Q (new_AGEMA_signal_6817) ) ;
    buf_clk new_AGEMA_reg_buffer_4049 ( .C (clk), .D (new_AGEMA_signal_6824), .Q (new_AGEMA_signal_6825) ) ;
    buf_clk new_AGEMA_reg_buffer_4057 ( .C (clk), .D (new_AGEMA_signal_6832), .Q (new_AGEMA_signal_6833) ) ;
    buf_clk new_AGEMA_reg_buffer_4065 ( .C (clk), .D (new_AGEMA_signal_6840), .Q (new_AGEMA_signal_6841) ) ;
    buf_clk new_AGEMA_reg_buffer_4073 ( .C (clk), .D (new_AGEMA_signal_6848), .Q (new_AGEMA_signal_6849) ) ;
    buf_clk new_AGEMA_reg_buffer_4081 ( .C (clk), .D (new_AGEMA_signal_6856), .Q (new_AGEMA_signal_6857) ) ;
    buf_clk new_AGEMA_reg_buffer_4089 ( .C (clk), .D (new_AGEMA_signal_6864), .Q (new_AGEMA_signal_6865) ) ;
    buf_clk new_AGEMA_reg_buffer_4097 ( .C (clk), .D (new_AGEMA_signal_6872), .Q (new_AGEMA_signal_6873) ) ;
    buf_clk new_AGEMA_reg_buffer_4105 ( .C (clk), .D (new_AGEMA_signal_6880), .Q (new_AGEMA_signal_6881) ) ;
    buf_clk new_AGEMA_reg_buffer_4113 ( .C (clk), .D (new_AGEMA_signal_6888), .Q (new_AGEMA_signal_6889) ) ;
    buf_clk new_AGEMA_reg_buffer_4121 ( .C (clk), .D (new_AGEMA_signal_6896), .Q (new_AGEMA_signal_6897) ) ;
    buf_clk new_AGEMA_reg_buffer_4129 ( .C (clk), .D (new_AGEMA_signal_6904), .Q (new_AGEMA_signal_6905) ) ;
    buf_clk new_AGEMA_reg_buffer_4137 ( .C (clk), .D (new_AGEMA_signal_6912), .Q (new_AGEMA_signal_6913) ) ;
    buf_clk new_AGEMA_reg_buffer_4145 ( .C (clk), .D (new_AGEMA_signal_6920), .Q (new_AGEMA_signal_6921) ) ;
    buf_clk new_AGEMA_reg_buffer_4153 ( .C (clk), .D (new_AGEMA_signal_6928), .Q (new_AGEMA_signal_6929) ) ;
    buf_clk new_AGEMA_reg_buffer_4161 ( .C (clk), .D (new_AGEMA_signal_6936), .Q (new_AGEMA_signal_6937) ) ;
    buf_clk new_AGEMA_reg_buffer_4169 ( .C (clk), .D (new_AGEMA_signal_6944), .Q (new_AGEMA_signal_6945) ) ;
    buf_clk new_AGEMA_reg_buffer_4177 ( .C (clk), .D (new_AGEMA_signal_6952), .Q (new_AGEMA_signal_6953) ) ;
    buf_clk new_AGEMA_reg_buffer_4185 ( .C (clk), .D (new_AGEMA_signal_6960), .Q (new_AGEMA_signal_6961) ) ;
    buf_clk new_AGEMA_reg_buffer_4475 ( .C (clk), .D (AddRoundKeyOutput[63]), .Q (new_AGEMA_signal_7251) ) ;
    buf_clk new_AGEMA_reg_buffer_4477 ( .C (clk), .D (new_AGEMA_signal_2793), .Q (new_AGEMA_signal_7253) ) ;
    buf_clk new_AGEMA_reg_buffer_4479 ( .C (clk), .D (new_AGEMA_signal_2794), .Q (new_AGEMA_signal_7255) ) ;
    buf_clk new_AGEMA_reg_buffer_4481 ( .C (clk), .D (AddRoundKeyOutput[61]), .Q (new_AGEMA_signal_7257) ) ;
    buf_clk new_AGEMA_reg_buffer_4483 ( .C (clk), .D (new_AGEMA_signal_2789), .Q (new_AGEMA_signal_7259) ) ;
    buf_clk new_AGEMA_reg_buffer_4485 ( .C (clk), .D (new_AGEMA_signal_2790), .Q (new_AGEMA_signal_7261) ) ;
    buf_clk new_AGEMA_reg_buffer_4487 ( .C (clk), .D (AddRoundKeyOutput[59]), .Q (new_AGEMA_signal_7263) ) ;
    buf_clk new_AGEMA_reg_buffer_4489 ( .C (clk), .D (new_AGEMA_signal_2785), .Q (new_AGEMA_signal_7265) ) ;
    buf_clk new_AGEMA_reg_buffer_4491 ( .C (clk), .D (new_AGEMA_signal_2786), .Q (new_AGEMA_signal_7267) ) ;
    buf_clk new_AGEMA_reg_buffer_4493 ( .C (clk), .D (AddRoundKeyOutput[57]), .Q (new_AGEMA_signal_7269) ) ;
    buf_clk new_AGEMA_reg_buffer_4495 ( .C (clk), .D (new_AGEMA_signal_2781), .Q (new_AGEMA_signal_7271) ) ;
    buf_clk new_AGEMA_reg_buffer_4497 ( .C (clk), .D (new_AGEMA_signal_2782), .Q (new_AGEMA_signal_7273) ) ;
    buf_clk new_AGEMA_reg_buffer_4499 ( .C (clk), .D (AddRoundKeyOutput[55]), .Q (new_AGEMA_signal_7275) ) ;
    buf_clk new_AGEMA_reg_buffer_4501 ( .C (clk), .D (new_AGEMA_signal_2777), .Q (new_AGEMA_signal_7277) ) ;
    buf_clk new_AGEMA_reg_buffer_4503 ( .C (clk), .D (new_AGEMA_signal_2778), .Q (new_AGEMA_signal_7279) ) ;
    buf_clk new_AGEMA_reg_buffer_4505 ( .C (clk), .D (AddRoundKeyOutput[53]), .Q (new_AGEMA_signal_7281) ) ;
    buf_clk new_AGEMA_reg_buffer_4507 ( .C (clk), .D (new_AGEMA_signal_2773), .Q (new_AGEMA_signal_7283) ) ;
    buf_clk new_AGEMA_reg_buffer_4509 ( .C (clk), .D (new_AGEMA_signal_2774), .Q (new_AGEMA_signal_7285) ) ;
    buf_clk new_AGEMA_reg_buffer_4511 ( .C (clk), .D (AddRoundKeyOutput[51]), .Q (new_AGEMA_signal_7287) ) ;
    buf_clk new_AGEMA_reg_buffer_4513 ( .C (clk), .D (new_AGEMA_signal_2769), .Q (new_AGEMA_signal_7289) ) ;
    buf_clk new_AGEMA_reg_buffer_4515 ( .C (clk), .D (new_AGEMA_signal_2770), .Q (new_AGEMA_signal_7291) ) ;
    buf_clk new_AGEMA_reg_buffer_4517 ( .C (clk), .D (AddRoundKeyOutput[49]), .Q (new_AGEMA_signal_7293) ) ;
    buf_clk new_AGEMA_reg_buffer_4519 ( .C (clk), .D (new_AGEMA_signal_2765), .Q (new_AGEMA_signal_7295) ) ;
    buf_clk new_AGEMA_reg_buffer_4521 ( .C (clk), .D (new_AGEMA_signal_2766), .Q (new_AGEMA_signal_7297) ) ;
    buf_clk new_AGEMA_reg_buffer_4523 ( .C (clk), .D (AddRoundKeyOutput[47]), .Q (new_AGEMA_signal_7299) ) ;
    buf_clk new_AGEMA_reg_buffer_4525 ( .C (clk), .D (new_AGEMA_signal_2809), .Q (new_AGEMA_signal_7301) ) ;
    buf_clk new_AGEMA_reg_buffer_4527 ( .C (clk), .D (new_AGEMA_signal_2810), .Q (new_AGEMA_signal_7303) ) ;
    buf_clk new_AGEMA_reg_buffer_4529 ( .C (clk), .D (AddRoundKeyOutput[45]), .Q (new_AGEMA_signal_7305) ) ;
    buf_clk new_AGEMA_reg_buffer_4531 ( .C (clk), .D (new_AGEMA_signal_2805), .Q (new_AGEMA_signal_7307) ) ;
    buf_clk new_AGEMA_reg_buffer_4533 ( .C (clk), .D (new_AGEMA_signal_2806), .Q (new_AGEMA_signal_7309) ) ;
    buf_clk new_AGEMA_reg_buffer_4535 ( .C (clk), .D (AddRoundKeyOutput[43]), .Q (new_AGEMA_signal_7311) ) ;
    buf_clk new_AGEMA_reg_buffer_4537 ( .C (clk), .D (new_AGEMA_signal_2801), .Q (new_AGEMA_signal_7313) ) ;
    buf_clk new_AGEMA_reg_buffer_4539 ( .C (clk), .D (new_AGEMA_signal_2802), .Q (new_AGEMA_signal_7315) ) ;
    buf_clk new_AGEMA_reg_buffer_4541 ( .C (clk), .D (AddRoundKeyOutput[41]), .Q (new_AGEMA_signal_7317) ) ;
    buf_clk new_AGEMA_reg_buffer_4543 ( .C (clk), .D (new_AGEMA_signal_2797), .Q (new_AGEMA_signal_7319) ) ;
    buf_clk new_AGEMA_reg_buffer_4545 ( .C (clk), .D (new_AGEMA_signal_2798), .Q (new_AGEMA_signal_7321) ) ;
    buf_clk new_AGEMA_reg_buffer_4547 ( .C (clk), .D (AddRoundKeyOutput[39]), .Q (new_AGEMA_signal_7323) ) ;
    buf_clk new_AGEMA_reg_buffer_4549 ( .C (clk), .D (new_AGEMA_signal_2825), .Q (new_AGEMA_signal_7325) ) ;
    buf_clk new_AGEMA_reg_buffer_4551 ( .C (clk), .D (new_AGEMA_signal_2826), .Q (new_AGEMA_signal_7327) ) ;
    buf_clk new_AGEMA_reg_buffer_4553 ( .C (clk), .D (AddRoundKeyOutput[37]), .Q (new_AGEMA_signal_7329) ) ;
    buf_clk new_AGEMA_reg_buffer_4555 ( .C (clk), .D (new_AGEMA_signal_2821), .Q (new_AGEMA_signal_7331) ) ;
    buf_clk new_AGEMA_reg_buffer_4557 ( .C (clk), .D (new_AGEMA_signal_2822), .Q (new_AGEMA_signal_7333) ) ;
    buf_clk new_AGEMA_reg_buffer_4559 ( .C (clk), .D (AddRoundKeyOutput[35]), .Q (new_AGEMA_signal_7335) ) ;
    buf_clk new_AGEMA_reg_buffer_4561 ( .C (clk), .D (new_AGEMA_signal_2817), .Q (new_AGEMA_signal_7337) ) ;
    buf_clk new_AGEMA_reg_buffer_4563 ( .C (clk), .D (new_AGEMA_signal_2818), .Q (new_AGEMA_signal_7339) ) ;
    buf_clk new_AGEMA_reg_buffer_4565 ( .C (clk), .D (AddRoundKeyOutput[33]), .Q (new_AGEMA_signal_7341) ) ;
    buf_clk new_AGEMA_reg_buffer_4567 ( .C (clk), .D (new_AGEMA_signal_2813), .Q (new_AGEMA_signal_7343) ) ;
    buf_clk new_AGEMA_reg_buffer_4569 ( .C (clk), .D (new_AGEMA_signal_2814), .Q (new_AGEMA_signal_7345) ) ;
    buf_clk new_AGEMA_reg_buffer_4571 ( .C (clk), .D (AddRoundKeyOutput[31]), .Q (new_AGEMA_signal_7347) ) ;
    buf_clk new_AGEMA_reg_buffer_4573 ( .C (clk), .D (new_AGEMA_signal_2697), .Q (new_AGEMA_signal_7349) ) ;
    buf_clk new_AGEMA_reg_buffer_4575 ( .C (clk), .D (new_AGEMA_signal_2698), .Q (new_AGEMA_signal_7351) ) ;
    buf_clk new_AGEMA_reg_buffer_4577 ( .C (clk), .D (AddRoundKeyOutput[29]), .Q (new_AGEMA_signal_7353) ) ;
    buf_clk new_AGEMA_reg_buffer_4579 ( .C (clk), .D (new_AGEMA_signal_2693), .Q (new_AGEMA_signal_7355) ) ;
    buf_clk new_AGEMA_reg_buffer_4581 ( .C (clk), .D (new_AGEMA_signal_2694), .Q (new_AGEMA_signal_7357) ) ;
    buf_clk new_AGEMA_reg_buffer_4583 ( .C (clk), .D (AddRoundKeyOutput[27]), .Q (new_AGEMA_signal_7359) ) ;
    buf_clk new_AGEMA_reg_buffer_4585 ( .C (clk), .D (new_AGEMA_signal_2689), .Q (new_AGEMA_signal_7361) ) ;
    buf_clk new_AGEMA_reg_buffer_4587 ( .C (clk), .D (new_AGEMA_signal_2690), .Q (new_AGEMA_signal_7363) ) ;
    buf_clk new_AGEMA_reg_buffer_4589 ( .C (clk), .D (AddRoundKeyOutput[25]), .Q (new_AGEMA_signal_7365) ) ;
    buf_clk new_AGEMA_reg_buffer_4591 ( .C (clk), .D (new_AGEMA_signal_2685), .Q (new_AGEMA_signal_7367) ) ;
    buf_clk new_AGEMA_reg_buffer_4593 ( .C (clk), .D (new_AGEMA_signal_2686), .Q (new_AGEMA_signal_7369) ) ;
    buf_clk new_AGEMA_reg_buffer_4595 ( .C (clk), .D (AddRoundKeyOutput[23]), .Q (new_AGEMA_signal_7371) ) ;
    buf_clk new_AGEMA_reg_buffer_4597 ( .C (clk), .D (new_AGEMA_signal_2681), .Q (new_AGEMA_signal_7373) ) ;
    buf_clk new_AGEMA_reg_buffer_4599 ( .C (clk), .D (new_AGEMA_signal_2682), .Q (new_AGEMA_signal_7375) ) ;
    buf_clk new_AGEMA_reg_buffer_4601 ( .C (clk), .D (AddRoundKeyOutput[21]), .Q (new_AGEMA_signal_7377) ) ;
    buf_clk new_AGEMA_reg_buffer_4603 ( .C (clk), .D (new_AGEMA_signal_2677), .Q (new_AGEMA_signal_7379) ) ;
    buf_clk new_AGEMA_reg_buffer_4605 ( .C (clk), .D (new_AGEMA_signal_2678), .Q (new_AGEMA_signal_7381) ) ;
    buf_clk new_AGEMA_reg_buffer_4607 ( .C (clk), .D (AddRoundKeyOutput[19]), .Q (new_AGEMA_signal_7383) ) ;
    buf_clk new_AGEMA_reg_buffer_4609 ( .C (clk), .D (new_AGEMA_signal_2673), .Q (new_AGEMA_signal_7385) ) ;
    buf_clk new_AGEMA_reg_buffer_4611 ( .C (clk), .D (new_AGEMA_signal_2674), .Q (new_AGEMA_signal_7387) ) ;
    buf_clk new_AGEMA_reg_buffer_4613 ( .C (clk), .D (AddRoundKeyOutput[17]), .Q (new_AGEMA_signal_7389) ) ;
    buf_clk new_AGEMA_reg_buffer_4615 ( .C (clk), .D (new_AGEMA_signal_2669), .Q (new_AGEMA_signal_7391) ) ;
    buf_clk new_AGEMA_reg_buffer_4617 ( .C (clk), .D (new_AGEMA_signal_2670), .Q (new_AGEMA_signal_7393) ) ;
    buf_clk new_AGEMA_reg_buffer_4619 ( .C (clk), .D (AddRoundKeyOutput[15]), .Q (new_AGEMA_signal_7395) ) ;
    buf_clk new_AGEMA_reg_buffer_4621 ( .C (clk), .D (new_AGEMA_signal_2665), .Q (new_AGEMA_signal_7397) ) ;
    buf_clk new_AGEMA_reg_buffer_4623 ( .C (clk), .D (new_AGEMA_signal_2666), .Q (new_AGEMA_signal_7399) ) ;
    buf_clk new_AGEMA_reg_buffer_4625 ( .C (clk), .D (AddRoundKeyOutput[13]), .Q (new_AGEMA_signal_7401) ) ;
    buf_clk new_AGEMA_reg_buffer_4627 ( .C (clk), .D (new_AGEMA_signal_2661), .Q (new_AGEMA_signal_7403) ) ;
    buf_clk new_AGEMA_reg_buffer_4629 ( .C (clk), .D (new_AGEMA_signal_2662), .Q (new_AGEMA_signal_7405) ) ;
    buf_clk new_AGEMA_reg_buffer_4631 ( .C (clk), .D (AddRoundKeyOutput[11]), .Q (new_AGEMA_signal_7407) ) ;
    buf_clk new_AGEMA_reg_buffer_4633 ( .C (clk), .D (new_AGEMA_signal_2657), .Q (new_AGEMA_signal_7409) ) ;
    buf_clk new_AGEMA_reg_buffer_4635 ( .C (clk), .D (new_AGEMA_signal_2658), .Q (new_AGEMA_signal_7411) ) ;
    buf_clk new_AGEMA_reg_buffer_4637 ( .C (clk), .D (AddRoundKeyOutput[9]), .Q (new_AGEMA_signal_7413) ) ;
    buf_clk new_AGEMA_reg_buffer_4639 ( .C (clk), .D (new_AGEMA_signal_2653), .Q (new_AGEMA_signal_7415) ) ;
    buf_clk new_AGEMA_reg_buffer_4641 ( .C (clk), .D (new_AGEMA_signal_2654), .Q (new_AGEMA_signal_7417) ) ;
    buf_clk new_AGEMA_reg_buffer_4643 ( .C (clk), .D (AddRoundKeyOutput[7]), .Q (new_AGEMA_signal_7419) ) ;
    buf_clk new_AGEMA_reg_buffer_4645 ( .C (clk), .D (new_AGEMA_signal_2649), .Q (new_AGEMA_signal_7421) ) ;
    buf_clk new_AGEMA_reg_buffer_4647 ( .C (clk), .D (new_AGEMA_signal_2650), .Q (new_AGEMA_signal_7423) ) ;
    buf_clk new_AGEMA_reg_buffer_4649 ( .C (clk), .D (AddRoundKeyOutput[5]), .Q (new_AGEMA_signal_7425) ) ;
    buf_clk new_AGEMA_reg_buffer_4651 ( .C (clk), .D (new_AGEMA_signal_2645), .Q (new_AGEMA_signal_7427) ) ;
    buf_clk new_AGEMA_reg_buffer_4653 ( .C (clk), .D (new_AGEMA_signal_2646), .Q (new_AGEMA_signal_7429) ) ;
    buf_clk new_AGEMA_reg_buffer_4655 ( .C (clk), .D (AddRoundKeyOutput[3]), .Q (new_AGEMA_signal_7431) ) ;
    buf_clk new_AGEMA_reg_buffer_4657 ( .C (clk), .D (new_AGEMA_signal_2641), .Q (new_AGEMA_signal_7433) ) ;
    buf_clk new_AGEMA_reg_buffer_4659 ( .C (clk), .D (new_AGEMA_signal_2642), .Q (new_AGEMA_signal_7435) ) ;
    buf_clk new_AGEMA_reg_buffer_4661 ( .C (clk), .D (AddRoundKeyOutput[1]), .Q (new_AGEMA_signal_7437) ) ;
    buf_clk new_AGEMA_reg_buffer_4663 ( .C (clk), .D (new_AGEMA_signal_2637), .Q (new_AGEMA_signal_7439) ) ;
    buf_clk new_AGEMA_reg_buffer_4665 ( .C (clk), .D (new_AGEMA_signal_2638), .Q (new_AGEMA_signal_7441) ) ;
    buf_clk new_AGEMA_reg_buffer_4673 ( .C (clk), .D (new_AGEMA_signal_7448), .Q (new_AGEMA_signal_7449) ) ;
    buf_clk new_AGEMA_reg_buffer_4681 ( .C (clk), .D (new_AGEMA_signal_7456), .Q (new_AGEMA_signal_7457) ) ;
    buf_clk new_AGEMA_reg_buffer_4689 ( .C (clk), .D (new_AGEMA_signal_7464), .Q (new_AGEMA_signal_7465) ) ;
    buf_clk new_AGEMA_reg_buffer_4697 ( .C (clk), .D (new_AGEMA_signal_7472), .Q (new_AGEMA_signal_7473) ) ;
    buf_clk new_AGEMA_reg_buffer_4705 ( .C (clk), .D (new_AGEMA_signal_7480), .Q (new_AGEMA_signal_7481) ) ;
    buf_clk new_AGEMA_reg_buffer_4713 ( .C (clk), .D (new_AGEMA_signal_7488), .Q (new_AGEMA_signal_7489) ) ;
    buf_clk new_AGEMA_reg_buffer_4721 ( .C (clk), .D (new_AGEMA_signal_7496), .Q (new_AGEMA_signal_7497) ) ;
    buf_clk new_AGEMA_reg_buffer_4729 ( .C (clk), .D (new_AGEMA_signal_7504), .Q (new_AGEMA_signal_7505) ) ;
    buf_clk new_AGEMA_reg_buffer_4737 ( .C (clk), .D (new_AGEMA_signal_7512), .Q (new_AGEMA_signal_7513) ) ;
    buf_clk new_AGEMA_reg_buffer_4745 ( .C (clk), .D (new_AGEMA_signal_7520), .Q (new_AGEMA_signal_7521) ) ;

    /* cells in depth 8 */
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_0_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1730, new_AGEMA_signal_1729, Feedback[0]}), .a ({new_AGEMA_signal_5450, new_AGEMA_signal_5442, new_AGEMA_signal_5434}), .c ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, MCOutput[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_2_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1726, new_AGEMA_signal_1725, Feedback[2]}), .a ({new_AGEMA_signal_5474, new_AGEMA_signal_5466, new_AGEMA_signal_5458}), .c ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, MCOutput[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_4_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1738, new_AGEMA_signal_1737, Feedback[4]}), .a ({new_AGEMA_signal_5498, new_AGEMA_signal_5490, new_AGEMA_signal_5482}), .c ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, MCOutput[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_6_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1734, new_AGEMA_signal_1733, Feedback[6]}), .a ({new_AGEMA_signal_5522, new_AGEMA_signal_5514, new_AGEMA_signal_5506}), .c ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, MCOutput[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_8_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1746, new_AGEMA_signal_1745, Feedback[8]}), .a ({new_AGEMA_signal_5546, new_AGEMA_signal_5538, new_AGEMA_signal_5530}), .c ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, MCOutput[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_10_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1742, new_AGEMA_signal_1741, Feedback[10]}), .a ({new_AGEMA_signal_5570, new_AGEMA_signal_5562, new_AGEMA_signal_5554}), .c ({new_AGEMA_signal_2182, new_AGEMA_signal_2181, MCOutput[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_12_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1754, new_AGEMA_signal_1753, Feedback[12]}), .a ({new_AGEMA_signal_5594, new_AGEMA_signal_5586, new_AGEMA_signal_5578}), .c ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, MCOutput[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_14_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1750, new_AGEMA_signal_1749, Feedback[14]}), .a ({new_AGEMA_signal_5618, new_AGEMA_signal_5610, new_AGEMA_signal_5602}), .c ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, MCOutput[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_16_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1762, new_AGEMA_signal_1761, Feedback[16]}), .a ({new_AGEMA_signal_5642, new_AGEMA_signal_5634, new_AGEMA_signal_5626}), .c ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, MCOutput[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_18_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1758, new_AGEMA_signal_1757, Feedback[18]}), .a ({new_AGEMA_signal_5666, new_AGEMA_signal_5658, new_AGEMA_signal_5650}), .c ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, MCOutput[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_20_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, Feedback[20]}), .a ({new_AGEMA_signal_5690, new_AGEMA_signal_5682, new_AGEMA_signal_5674}), .c ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, MCOutput[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_22_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1766, new_AGEMA_signal_1765, Feedback[22]}), .a ({new_AGEMA_signal_5714, new_AGEMA_signal_5706, new_AGEMA_signal_5698}), .c ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, MCOutput[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_24_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1778, new_AGEMA_signal_1777, Feedback[24]}), .a ({new_AGEMA_signal_5738, new_AGEMA_signal_5730, new_AGEMA_signal_5722}), .c ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, MCOutput[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_26_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1774, new_AGEMA_signal_1773, Feedback[26]}), .a ({new_AGEMA_signal_5762, new_AGEMA_signal_5754, new_AGEMA_signal_5746}), .c ({new_AGEMA_signal_2246, new_AGEMA_signal_2245, MCOutput[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_28_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1786, new_AGEMA_signal_1785, Feedback[28]}), .a ({new_AGEMA_signal_5786, new_AGEMA_signal_5778, new_AGEMA_signal_5770}), .c ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, MCOutput[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_30_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1782, new_AGEMA_signal_1781, Feedback[30]}), .a ({new_AGEMA_signal_5810, new_AGEMA_signal_5802, new_AGEMA_signal_5794}), .c ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, MCOutput[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_32_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1794, new_AGEMA_signal_1793, Feedback[32]}), .a ({new_AGEMA_signal_5834, new_AGEMA_signal_5826, new_AGEMA_signal_5818}), .c ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, MCInput[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_34_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1790, new_AGEMA_signal_1789, Feedback[34]}), .a ({new_AGEMA_signal_5858, new_AGEMA_signal_5850, new_AGEMA_signal_5842}), .c ({new_AGEMA_signal_2278, new_AGEMA_signal_2277, MCInput[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_36_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, Feedback[36]}), .a ({new_AGEMA_signal_5882, new_AGEMA_signal_5874, new_AGEMA_signal_5866}), .c ({new_AGEMA_signal_2286, new_AGEMA_signal_2285, MCInput[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_38_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1798, new_AGEMA_signal_1797, Feedback[38]}), .a ({new_AGEMA_signal_5906, new_AGEMA_signal_5898, new_AGEMA_signal_5890}), .c ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, MCInput[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_40_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1810, new_AGEMA_signal_1809, Feedback[40]}), .a ({new_AGEMA_signal_5930, new_AGEMA_signal_5922, new_AGEMA_signal_5914}), .c ({new_AGEMA_signal_2302, new_AGEMA_signal_2301, MCInput[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_42_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1806, new_AGEMA_signal_1805, Feedback[42]}), .a ({new_AGEMA_signal_5954, new_AGEMA_signal_5946, new_AGEMA_signal_5938}), .c ({new_AGEMA_signal_2310, new_AGEMA_signal_2309, MCInput[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_44_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1818, new_AGEMA_signal_1817, Feedback[44]}), .a ({new_AGEMA_signal_5978, new_AGEMA_signal_5970, new_AGEMA_signal_5962}), .c ({new_AGEMA_signal_2318, new_AGEMA_signal_2317, MCInput[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_46_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1814, new_AGEMA_signal_1813, Feedback[46]}), .a ({new_AGEMA_signal_6002, new_AGEMA_signal_5994, new_AGEMA_signal_5986}), .c ({new_AGEMA_signal_2326, new_AGEMA_signal_2325, MCInput[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_48_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1826, new_AGEMA_signal_1825, Feedback[48]}), .a ({new_AGEMA_signal_6026, new_AGEMA_signal_6018, new_AGEMA_signal_6010}), .c ({new_AGEMA_signal_2334, new_AGEMA_signal_2333, MCInput[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_50_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1822, new_AGEMA_signal_1821, Feedback[50]}), .a ({new_AGEMA_signal_6050, new_AGEMA_signal_6042, new_AGEMA_signal_6034}), .c ({new_AGEMA_signal_2342, new_AGEMA_signal_2341, MCInput[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_52_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1834, new_AGEMA_signal_1833, Feedback[52]}), .a ({new_AGEMA_signal_6074, new_AGEMA_signal_6066, new_AGEMA_signal_6058}), .c ({new_AGEMA_signal_2350, new_AGEMA_signal_2349, MCInput[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_54_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1830, new_AGEMA_signal_1829, Feedback[54]}), .a ({new_AGEMA_signal_6098, new_AGEMA_signal_6090, new_AGEMA_signal_6082}), .c ({new_AGEMA_signal_2358, new_AGEMA_signal_2357, MCInput[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_56_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1842, new_AGEMA_signal_1841, Feedback[56]}), .a ({new_AGEMA_signal_6122, new_AGEMA_signal_6114, new_AGEMA_signal_6106}), .c ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, MCInput[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_58_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1838, new_AGEMA_signal_1837, Feedback[58]}), .a ({new_AGEMA_signal_6146, new_AGEMA_signal_6138, new_AGEMA_signal_6130}), .c ({new_AGEMA_signal_2374, new_AGEMA_signal_2373, MCInput[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_60_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, Feedback[60]}), .a ({new_AGEMA_signal_6170, new_AGEMA_signal_6162, new_AGEMA_signal_6154}), .c ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, MCInput[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) InputMUX_MUXInst_62_U1 ( .s (new_AGEMA_signal_5426), .b ({new_AGEMA_signal_1846, new_AGEMA_signal_1845, Feedback[62]}), .a ({new_AGEMA_signal_6194, new_AGEMA_signal_6186, new_AGEMA_signal_6178}), .c ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, MCInput[62]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_0_U3 ( .a ({new_AGEMA_signal_2414, new_AGEMA_signal_2413, MCInst_XOR_r0_Inst_0_n2}), .b ({new_AGEMA_signal_2412, new_AGEMA_signal_2411, MCInst_XOR_r0_Inst_0_n1}), .c ({new_AGEMA_signal_2572, new_AGEMA_signal_2571, MCOutput[48]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_0_U2 ( .a ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, MCOutput[16]}), .b ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, MCOutput[0]}), .c ({new_AGEMA_signal_2412, new_AGEMA_signal_2411, MCInst_XOR_r0_Inst_0_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2334, new_AGEMA_signal_2333, MCInput[48]}), .c ({new_AGEMA_signal_2414, new_AGEMA_signal_2413, MCInst_XOR_r0_Inst_0_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_0_U2 ( .a ({new_AGEMA_signal_2416, new_AGEMA_signal_2415, MCInst_XOR_r1_Inst_0_n1}), .b ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, MCOutput[0]}), .c ({new_AGEMA_signal_2574, new_AGEMA_signal_2573, MCOutput[32]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, MCInput[32]}), .c ({new_AGEMA_signal_2416, new_AGEMA_signal_2415, MCInst_XOR_r1_Inst_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_2_U3 ( .a ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, MCInst_XOR_r0_Inst_2_n2}), .b ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, MCInst_XOR_r0_Inst_2_n1}), .c ({new_AGEMA_signal_2580, new_AGEMA_signal_2579, MCOutput[50]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_2_U2 ( .a ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, MCOutput[18]}), .b ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, MCOutput[2]}), .c ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, MCInst_XOR_r0_Inst_2_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2342, new_AGEMA_signal_2341, MCInput[50]}), .c ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, MCInst_XOR_r0_Inst_2_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_2_U2 ( .a ({new_AGEMA_signal_2428, new_AGEMA_signal_2427, MCInst_XOR_r1_Inst_2_n1}), .b ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, MCOutput[2]}), .c ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, MCOutput[34]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2278, new_AGEMA_signal_2277, MCInput[34]}), .c ({new_AGEMA_signal_2428, new_AGEMA_signal_2427, MCInst_XOR_r1_Inst_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_4_U3 ( .a ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, MCInst_XOR_r0_Inst_4_n2}), .b ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, MCInst_XOR_r0_Inst_4_n1}), .c ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, MCOutput[52]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_4_U2 ( .a ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, MCOutput[20]}), .b ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, MCOutput[4]}), .c ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, MCInst_XOR_r0_Inst_4_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_4_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2350, new_AGEMA_signal_2349, MCInput[52]}), .c ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, MCInst_XOR_r0_Inst_4_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_4_U2 ( .a ({new_AGEMA_signal_2440, new_AGEMA_signal_2439, MCInst_XOR_r1_Inst_4_n1}), .b ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, MCOutput[4]}), .c ({new_AGEMA_signal_2590, new_AGEMA_signal_2589, MCOutput[36]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_4_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2286, new_AGEMA_signal_2285, MCInput[36]}), .c ({new_AGEMA_signal_2440, new_AGEMA_signal_2439, MCInst_XOR_r1_Inst_4_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_6_U3 ( .a ({new_AGEMA_signal_2450, new_AGEMA_signal_2449, MCInst_XOR_r0_Inst_6_n2}), .b ({new_AGEMA_signal_2448, new_AGEMA_signal_2447, MCInst_XOR_r0_Inst_6_n1}), .c ({new_AGEMA_signal_2596, new_AGEMA_signal_2595, MCOutput[54]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_6_U2 ( .a ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, MCOutput[22]}), .b ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, MCOutput[6]}), .c ({new_AGEMA_signal_2448, new_AGEMA_signal_2447, MCInst_XOR_r0_Inst_6_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_6_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2358, new_AGEMA_signal_2357, MCInput[54]}), .c ({new_AGEMA_signal_2450, new_AGEMA_signal_2449, MCInst_XOR_r0_Inst_6_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_6_U2 ( .a ({new_AGEMA_signal_2452, new_AGEMA_signal_2451, MCInst_XOR_r1_Inst_6_n1}), .b ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, MCOutput[6]}), .c ({new_AGEMA_signal_2598, new_AGEMA_signal_2597, MCOutput[38]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_6_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, MCInput[38]}), .c ({new_AGEMA_signal_2452, new_AGEMA_signal_2451, MCInst_XOR_r1_Inst_6_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_8_U3 ( .a ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, MCInst_XOR_r0_Inst_8_n2}), .b ({new_AGEMA_signal_2460, new_AGEMA_signal_2459, MCInst_XOR_r0_Inst_8_n1}), .c ({new_AGEMA_signal_2604, new_AGEMA_signal_2603, MCOutput[56]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_8_U2 ( .a ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, MCOutput[24]}), .b ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, MCOutput[8]}), .c ({new_AGEMA_signal_2460, new_AGEMA_signal_2459, MCInst_XOR_r0_Inst_8_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_8_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, MCInput[56]}), .c ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, MCInst_XOR_r0_Inst_8_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_8_U2 ( .a ({new_AGEMA_signal_2464, new_AGEMA_signal_2463, MCInst_XOR_r1_Inst_8_n1}), .b ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, MCOutput[8]}), .c ({new_AGEMA_signal_2606, new_AGEMA_signal_2605, MCOutput[40]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_8_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2302, new_AGEMA_signal_2301, MCInput[40]}), .c ({new_AGEMA_signal_2464, new_AGEMA_signal_2463, MCInst_XOR_r1_Inst_8_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_10_U3 ( .a ({new_AGEMA_signal_2474, new_AGEMA_signal_2473, MCInst_XOR_r0_Inst_10_n2}), .b ({new_AGEMA_signal_2472, new_AGEMA_signal_2471, MCInst_XOR_r0_Inst_10_n1}), .c ({new_AGEMA_signal_2612, new_AGEMA_signal_2611, MCOutput[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_10_U2 ( .a ({new_AGEMA_signal_2246, new_AGEMA_signal_2245, MCOutput[26]}), .b ({new_AGEMA_signal_2182, new_AGEMA_signal_2181, MCOutput[10]}), .c ({new_AGEMA_signal_2472, new_AGEMA_signal_2471, MCInst_XOR_r0_Inst_10_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_10_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2374, new_AGEMA_signal_2373, MCInput[58]}), .c ({new_AGEMA_signal_2474, new_AGEMA_signal_2473, MCInst_XOR_r0_Inst_10_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_10_U2 ( .a ({new_AGEMA_signal_2476, new_AGEMA_signal_2475, MCInst_XOR_r1_Inst_10_n1}), .b ({new_AGEMA_signal_2182, new_AGEMA_signal_2181, MCOutput[10]}), .c ({new_AGEMA_signal_2614, new_AGEMA_signal_2613, MCOutput[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_10_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2310, new_AGEMA_signal_2309, MCInput[42]}), .c ({new_AGEMA_signal_2476, new_AGEMA_signal_2475, MCInst_XOR_r1_Inst_10_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_12_U3 ( .a ({new_AGEMA_signal_2486, new_AGEMA_signal_2485, MCInst_XOR_r0_Inst_12_n2}), .b ({new_AGEMA_signal_2484, new_AGEMA_signal_2483, MCInst_XOR_r0_Inst_12_n1}), .c ({new_AGEMA_signal_2620, new_AGEMA_signal_2619, MCOutput[60]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_12_U2 ( .a ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, MCOutput[28]}), .b ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, MCOutput[12]}), .c ({new_AGEMA_signal_2484, new_AGEMA_signal_2483, MCInst_XOR_r0_Inst_12_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_12_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, MCInput[60]}), .c ({new_AGEMA_signal_2486, new_AGEMA_signal_2485, MCInst_XOR_r0_Inst_12_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_12_U2 ( .a ({new_AGEMA_signal_2488, new_AGEMA_signal_2487, MCInst_XOR_r1_Inst_12_n1}), .b ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, MCOutput[12]}), .c ({new_AGEMA_signal_2622, new_AGEMA_signal_2621, MCOutput[44]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_12_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2318, new_AGEMA_signal_2317, MCInput[44]}), .c ({new_AGEMA_signal_2488, new_AGEMA_signal_2487, MCInst_XOR_r1_Inst_12_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_14_U3 ( .a ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, MCInst_XOR_r0_Inst_14_n2}), .b ({new_AGEMA_signal_2496, new_AGEMA_signal_2495, MCInst_XOR_r0_Inst_14_n1}), .c ({new_AGEMA_signal_2628, new_AGEMA_signal_2627, MCOutput[62]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_14_U2 ( .a ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, MCOutput[30]}), .b ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, MCOutput[14]}), .c ({new_AGEMA_signal_2496, new_AGEMA_signal_2495, MCInst_XOR_r0_Inst_14_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r0_Inst_14_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, MCInput[62]}), .c ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, MCInst_XOR_r0_Inst_14_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_14_U2 ( .a ({new_AGEMA_signal_2500, new_AGEMA_signal_2499, MCInst_XOR_r1_Inst_14_n1}), .b ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, MCOutput[14]}), .c ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, MCOutput[46]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) MCInst_XOR_r1_Inst_14_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2326, new_AGEMA_signal_2325, MCInput[46]}), .c ({new_AGEMA_signal_2500, new_AGEMA_signal_2499, MCInst_XOR_r1_Inst_14_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2700, new_AGEMA_signal_2699, AddKeyXOR1_XORInst_0_0_n1}), .b ({new_AGEMA_signal_6218, new_AGEMA_signal_6210, new_AGEMA_signal_6202}), .c ({new_AGEMA_signal_2764, new_AGEMA_signal_2763, AddRoundKeyOutput[48]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2572, new_AGEMA_signal_2571, MCOutput[48]}), .c ({new_AGEMA_signal_2700, new_AGEMA_signal_2699, AddKeyXOR1_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, AddKeyXOR1_XORInst_0_2_n1}), .b ({new_AGEMA_signal_6242, new_AGEMA_signal_6234, new_AGEMA_signal_6226}), .c ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, AddRoundKeyOutput[50]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2580, new_AGEMA_signal_2579, MCOutput[50]}), .c ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, AddKeyXOR1_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2708, new_AGEMA_signal_2707, AddKeyXOR1_XORInst_1_0_n1}), .b ({new_AGEMA_signal_6266, new_AGEMA_signal_6258, new_AGEMA_signal_6250}), .c ({new_AGEMA_signal_2772, new_AGEMA_signal_2771, AddRoundKeyOutput[52]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, MCOutput[52]}), .c ({new_AGEMA_signal_2708, new_AGEMA_signal_2707, AddKeyXOR1_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2712, new_AGEMA_signal_2711, AddKeyXOR1_XORInst_1_2_n1}), .b ({new_AGEMA_signal_6290, new_AGEMA_signal_6282, new_AGEMA_signal_6274}), .c ({new_AGEMA_signal_2776, new_AGEMA_signal_2775, AddRoundKeyOutput[54]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2596, new_AGEMA_signal_2595, MCOutput[54]}), .c ({new_AGEMA_signal_2712, new_AGEMA_signal_2711, AddKeyXOR1_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_2716, new_AGEMA_signal_2715, AddKeyXOR1_XORInst_2_0_n1}), .b ({new_AGEMA_signal_6314, new_AGEMA_signal_6306, new_AGEMA_signal_6298}), .c ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, AddRoundKeyOutput[56]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2604, new_AGEMA_signal_2603, MCOutput[56]}), .c ({new_AGEMA_signal_2716, new_AGEMA_signal_2715, AddKeyXOR1_XORInst_2_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_2720, new_AGEMA_signal_2719, AddKeyXOR1_XORInst_2_2_n1}), .b ({new_AGEMA_signal_6338, new_AGEMA_signal_6330, new_AGEMA_signal_6322}), .c ({new_AGEMA_signal_2784, new_AGEMA_signal_2783, AddRoundKeyOutput[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2612, new_AGEMA_signal_2611, MCOutput[58]}), .c ({new_AGEMA_signal_2720, new_AGEMA_signal_2719, AddKeyXOR1_XORInst_2_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_2724, new_AGEMA_signal_2723, AddKeyXOR1_XORInst_3_0_n1}), .b ({new_AGEMA_signal_6362, new_AGEMA_signal_6354, new_AGEMA_signal_6346}), .c ({new_AGEMA_signal_2788, new_AGEMA_signal_2787, AddRoundKeyOutput[60]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2620, new_AGEMA_signal_2619, MCOutput[60]}), .c ({new_AGEMA_signal_2724, new_AGEMA_signal_2723, AddKeyXOR1_XORInst_3_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_2728, new_AGEMA_signal_2727, AddKeyXOR1_XORInst_3_2_n1}), .b ({new_AGEMA_signal_6386, new_AGEMA_signal_6378, new_AGEMA_signal_6370}), .c ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, AddRoundKeyOutput[62]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR1_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2628, new_AGEMA_signal_2627, MCOutput[62]}), .c ({new_AGEMA_signal_2728, new_AGEMA_signal_2727, AddKeyXOR1_XORInst_3_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_0_0_U3 ( .a ({new_AGEMA_signal_2732, new_AGEMA_signal_2731, AddKeyConstXOR_XORInst_0_0_n2}), .b ({new_AGEMA_signal_6410, new_AGEMA_signal_6402, new_AGEMA_signal_6394}), .c ({new_AGEMA_signal_2796, new_AGEMA_signal_2795, AddRoundKeyOutput[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2606, new_AGEMA_signal_2605, MCOutput[40]}), .c ({new_AGEMA_signal_2732, new_AGEMA_signal_2731, AddKeyConstXOR_XORInst_0_0_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_0_2_U3 ( .a ({new_AGEMA_signal_2736, new_AGEMA_signal_2735, AddKeyConstXOR_XORInst_0_2_n2}), .b ({new_AGEMA_signal_6434, new_AGEMA_signal_6426, new_AGEMA_signal_6418}), .c ({new_AGEMA_signal_2800, new_AGEMA_signal_2799, AddRoundKeyOutput[42]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2614, new_AGEMA_signal_2613, MCOutput[42]}), .c ({new_AGEMA_signal_2736, new_AGEMA_signal_2735, AddKeyConstXOR_XORInst_0_2_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_1_0_U3 ( .a ({new_AGEMA_signal_2740, new_AGEMA_signal_2739, AddKeyConstXOR_XORInst_1_0_n2}), .b ({new_AGEMA_signal_6458, new_AGEMA_signal_6450, new_AGEMA_signal_6442}), .c ({new_AGEMA_signal_2804, new_AGEMA_signal_2803, AddRoundKeyOutput[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2622, new_AGEMA_signal_2621, MCOutput[44]}), .c ({new_AGEMA_signal_2740, new_AGEMA_signal_2739, AddKeyConstXOR_XORInst_1_0_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_1_2_U3 ( .a ({new_AGEMA_signal_2744, new_AGEMA_signal_2743, AddKeyConstXOR_XORInst_1_2_n2}), .b ({new_AGEMA_signal_6482, new_AGEMA_signal_6474, new_AGEMA_signal_6466}), .c ({new_AGEMA_signal_2808, new_AGEMA_signal_2807, AddRoundKeyOutput[46]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyConstXOR_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, MCOutput[46]}), .c ({new_AGEMA_signal_2744, new_AGEMA_signal_2743, AddKeyConstXOR_XORInst_1_2_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2508, new_AGEMA_signal_2507, AddKeyXOR2_XORInst_0_0_n1}), .b ({new_AGEMA_signal_6506, new_AGEMA_signal_6498, new_AGEMA_signal_6490}), .c ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, AddRoundKeyOutput[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, MCOutput[0]}), .c ({new_AGEMA_signal_2508, new_AGEMA_signal_2507, AddKeyXOR2_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2512, new_AGEMA_signal_2511, AddKeyXOR2_XORInst_0_2_n1}), .b ({new_AGEMA_signal_6530, new_AGEMA_signal_6522, new_AGEMA_signal_6514}), .c ({new_AGEMA_signal_2640, new_AGEMA_signal_2639, AddRoundKeyOutput[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, MCOutput[2]}), .c ({new_AGEMA_signal_2512, new_AGEMA_signal_2511, AddKeyXOR2_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, AddKeyXOR2_XORInst_1_0_n1}), .b ({new_AGEMA_signal_6554, new_AGEMA_signal_6546, new_AGEMA_signal_6538}), .c ({new_AGEMA_signal_2644, new_AGEMA_signal_2643, AddRoundKeyOutput[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, MCOutput[4]}), .c ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, AddKeyXOR2_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2520, new_AGEMA_signal_2519, AddKeyXOR2_XORInst_1_2_n1}), .b ({new_AGEMA_signal_6578, new_AGEMA_signal_6570, new_AGEMA_signal_6562}), .c ({new_AGEMA_signal_2648, new_AGEMA_signal_2647, AddRoundKeyOutput[6]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, MCOutput[6]}), .c ({new_AGEMA_signal_2520, new_AGEMA_signal_2519, AddKeyXOR2_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_2524, new_AGEMA_signal_2523, AddKeyXOR2_XORInst_2_0_n1}), .b ({new_AGEMA_signal_6602, new_AGEMA_signal_6594, new_AGEMA_signal_6586}), .c ({new_AGEMA_signal_2652, new_AGEMA_signal_2651, AddRoundKeyOutput[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, MCOutput[8]}), .c ({new_AGEMA_signal_2524, new_AGEMA_signal_2523, AddKeyXOR2_XORInst_2_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_2528, new_AGEMA_signal_2527, AddKeyXOR2_XORInst_2_2_n1}), .b ({new_AGEMA_signal_6626, new_AGEMA_signal_6618, new_AGEMA_signal_6610}), .c ({new_AGEMA_signal_2656, new_AGEMA_signal_2655, AddRoundKeyOutput[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2182, new_AGEMA_signal_2181, MCOutput[10]}), .c ({new_AGEMA_signal_2528, new_AGEMA_signal_2527, AddKeyXOR2_XORInst_2_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_2532, new_AGEMA_signal_2531, AddKeyXOR2_XORInst_3_0_n1}), .b ({new_AGEMA_signal_6650, new_AGEMA_signal_6642, new_AGEMA_signal_6634}), .c ({new_AGEMA_signal_2660, new_AGEMA_signal_2659, AddRoundKeyOutput[12]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, MCOutput[12]}), .c ({new_AGEMA_signal_2532, new_AGEMA_signal_2531, AddKeyXOR2_XORInst_3_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_2536, new_AGEMA_signal_2535, AddKeyXOR2_XORInst_3_2_n1}), .b ({new_AGEMA_signal_6674, new_AGEMA_signal_6666, new_AGEMA_signal_6658}), .c ({new_AGEMA_signal_2664, new_AGEMA_signal_2663, AddRoundKeyOutput[14]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, MCOutput[14]}), .c ({new_AGEMA_signal_2536, new_AGEMA_signal_2535, AddKeyXOR2_XORInst_3_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_4_0_U2 ( .a ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, AddKeyXOR2_XORInst_4_0_n1}), .b ({new_AGEMA_signal_6698, new_AGEMA_signal_6690, new_AGEMA_signal_6682}), .c ({new_AGEMA_signal_2668, new_AGEMA_signal_2667, AddRoundKeyOutput[16]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_4_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, MCOutput[16]}), .c ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, AddKeyXOR2_XORInst_4_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_4_2_U2 ( .a ({new_AGEMA_signal_2544, new_AGEMA_signal_2543, AddKeyXOR2_XORInst_4_2_n1}), .b ({new_AGEMA_signal_6722, new_AGEMA_signal_6714, new_AGEMA_signal_6706}), .c ({new_AGEMA_signal_2672, new_AGEMA_signal_2671, AddRoundKeyOutput[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_4_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, MCOutput[18]}), .c ({new_AGEMA_signal_2544, new_AGEMA_signal_2543, AddKeyXOR2_XORInst_4_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_5_0_U2 ( .a ({new_AGEMA_signal_2548, new_AGEMA_signal_2547, AddKeyXOR2_XORInst_5_0_n1}), .b ({new_AGEMA_signal_6746, new_AGEMA_signal_6738, new_AGEMA_signal_6730}), .c ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, AddRoundKeyOutput[20]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_5_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, MCOutput[20]}), .c ({new_AGEMA_signal_2548, new_AGEMA_signal_2547, AddKeyXOR2_XORInst_5_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_5_2_U2 ( .a ({new_AGEMA_signal_2552, new_AGEMA_signal_2551, AddKeyXOR2_XORInst_5_2_n1}), .b ({new_AGEMA_signal_6770, new_AGEMA_signal_6762, new_AGEMA_signal_6754}), .c ({new_AGEMA_signal_2680, new_AGEMA_signal_2679, AddRoundKeyOutput[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_5_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, MCOutput[22]}), .c ({new_AGEMA_signal_2552, new_AGEMA_signal_2551, AddKeyXOR2_XORInst_5_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_6_0_U2 ( .a ({new_AGEMA_signal_2556, new_AGEMA_signal_2555, AddKeyXOR2_XORInst_6_0_n1}), .b ({new_AGEMA_signal_6794, new_AGEMA_signal_6786, new_AGEMA_signal_6778}), .c ({new_AGEMA_signal_2684, new_AGEMA_signal_2683, AddRoundKeyOutput[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_6_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, MCOutput[24]}), .c ({new_AGEMA_signal_2556, new_AGEMA_signal_2555, AddKeyXOR2_XORInst_6_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_6_2_U2 ( .a ({new_AGEMA_signal_2560, new_AGEMA_signal_2559, AddKeyXOR2_XORInst_6_2_n1}), .b ({new_AGEMA_signal_6818, new_AGEMA_signal_6810, new_AGEMA_signal_6802}), .c ({new_AGEMA_signal_2688, new_AGEMA_signal_2687, AddRoundKeyOutput[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_6_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2246, new_AGEMA_signal_2245, MCOutput[26]}), .c ({new_AGEMA_signal_2560, new_AGEMA_signal_2559, AddKeyXOR2_XORInst_6_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_7_0_U2 ( .a ({new_AGEMA_signal_2564, new_AGEMA_signal_2563, AddKeyXOR2_XORInst_7_0_n1}), .b ({new_AGEMA_signal_6842, new_AGEMA_signal_6834, new_AGEMA_signal_6826}), .c ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, AddRoundKeyOutput[28]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_7_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, MCOutput[28]}), .c ({new_AGEMA_signal_2564, new_AGEMA_signal_2563, AddKeyXOR2_XORInst_7_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_7_2_U2 ( .a ({new_AGEMA_signal_2568, new_AGEMA_signal_2567, AddKeyXOR2_XORInst_7_2_n1}), .b ({new_AGEMA_signal_6866, new_AGEMA_signal_6858, new_AGEMA_signal_6850}), .c ({new_AGEMA_signal_2696, new_AGEMA_signal_2695, AddRoundKeyOutput[30]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_7_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, MCOutput[30]}), .c ({new_AGEMA_signal_2568, new_AGEMA_signal_2567, AddKeyXOR2_XORInst_7_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_8_0_U2 ( .a ({new_AGEMA_signal_2748, new_AGEMA_signal_2747, AddKeyXOR2_XORInst_8_0_n1}), .b ({new_AGEMA_signal_6890, new_AGEMA_signal_6882, new_AGEMA_signal_6874}), .c ({new_AGEMA_signal_2812, new_AGEMA_signal_2811, AddRoundKeyOutput[32]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_8_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2574, new_AGEMA_signal_2573, MCOutput[32]}), .c ({new_AGEMA_signal_2748, new_AGEMA_signal_2747, AddKeyXOR2_XORInst_8_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_8_2_U2 ( .a ({new_AGEMA_signal_2752, new_AGEMA_signal_2751, AddKeyXOR2_XORInst_8_2_n1}), .b ({new_AGEMA_signal_6914, new_AGEMA_signal_6906, new_AGEMA_signal_6898}), .c ({new_AGEMA_signal_2816, new_AGEMA_signal_2815, AddRoundKeyOutput[34]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_8_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, MCOutput[34]}), .c ({new_AGEMA_signal_2752, new_AGEMA_signal_2751, AddKeyXOR2_XORInst_8_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_9_0_U2 ( .a ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, AddKeyXOR2_XORInst_9_0_n1}), .b ({new_AGEMA_signal_6938, new_AGEMA_signal_6930, new_AGEMA_signal_6922}), .c ({new_AGEMA_signal_2820, new_AGEMA_signal_2819, AddRoundKeyOutput[36]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_9_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2590, new_AGEMA_signal_2589, MCOutput[36]}), .c ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, AddKeyXOR2_XORInst_9_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_9_2_U2 ( .a ({new_AGEMA_signal_2760, new_AGEMA_signal_2759, AddKeyXOR2_XORInst_9_2_n1}), .b ({new_AGEMA_signal_6962, new_AGEMA_signal_6954, new_AGEMA_signal_6946}), .c ({new_AGEMA_signal_2824, new_AGEMA_signal_2823, AddRoundKeyOutput[38]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) AddKeyXOR2_XORInst_9_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2598, new_AGEMA_signal_2597, MCOutput[38]}), .c ({new_AGEMA_signal_2760, new_AGEMA_signal_2759, AddKeyXOR2_XORInst_9_2_n1}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U17 ( .a ({new_AGEMA_signal_6968, new_AGEMA_signal_6966, new_AGEMA_signal_6964}), .b ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, SubCellInst_SboxInst_0_n12}), .clk (clk), .r ({Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_1726, new_AGEMA_signal_1725, Feedback[2]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U8 ( .a ({new_AGEMA_signal_6980, new_AGEMA_signal_6976, new_AGEMA_signal_6972}), .b ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, SubCellInst_SboxInst_0_n3}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675]}), .c ({new_AGEMA_signal_1730, new_AGEMA_signal_1729, Feedback[0]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U17 ( .a ({new_AGEMA_signal_6986, new_AGEMA_signal_6984, new_AGEMA_signal_6982}), .b ({new_AGEMA_signal_1578, new_AGEMA_signal_1577, SubCellInst_SboxInst_1_n12}), .clk (clk), .r ({Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_1734, new_AGEMA_signal_1733, Feedback[6]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U8 ( .a ({new_AGEMA_signal_6998, new_AGEMA_signal_6994, new_AGEMA_signal_6990}), .b ({new_AGEMA_signal_1582, new_AGEMA_signal_1581, SubCellInst_SboxInst_1_n3}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681]}), .c ({new_AGEMA_signal_1738, new_AGEMA_signal_1737, Feedback[4]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U17 ( .a ({new_AGEMA_signal_7004, new_AGEMA_signal_7002, new_AGEMA_signal_7000}), .b ({new_AGEMA_signal_1588, new_AGEMA_signal_1587, SubCellInst_SboxInst_2_n12}), .clk (clk), .r ({Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_1742, new_AGEMA_signal_1741, Feedback[10]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U8 ( .a ({new_AGEMA_signal_7016, new_AGEMA_signal_7012, new_AGEMA_signal_7008}), .b ({new_AGEMA_signal_1592, new_AGEMA_signal_1591, SubCellInst_SboxInst_2_n3}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687]}), .c ({new_AGEMA_signal_1746, new_AGEMA_signal_1745, Feedback[8]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U17 ( .a ({new_AGEMA_signal_7022, new_AGEMA_signal_7020, new_AGEMA_signal_7018}), .b ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, SubCellInst_SboxInst_3_n12}), .clk (clk), .r ({Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_1750, new_AGEMA_signal_1749, Feedback[14]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U8 ( .a ({new_AGEMA_signal_7034, new_AGEMA_signal_7030, new_AGEMA_signal_7026}), .b ({new_AGEMA_signal_1602, new_AGEMA_signal_1601, SubCellInst_SboxInst_3_n3}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693]}), .c ({new_AGEMA_signal_1754, new_AGEMA_signal_1753, Feedback[12]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U17 ( .a ({new_AGEMA_signal_7040, new_AGEMA_signal_7038, new_AGEMA_signal_7036}), .b ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, SubCellInst_SboxInst_4_n12}), .clk (clk), .r ({Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_1758, new_AGEMA_signal_1757, Feedback[18]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U8 ( .a ({new_AGEMA_signal_7052, new_AGEMA_signal_7048, new_AGEMA_signal_7044}), .b ({new_AGEMA_signal_1612, new_AGEMA_signal_1611, SubCellInst_SboxInst_4_n3}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699]}), .c ({new_AGEMA_signal_1762, new_AGEMA_signal_1761, Feedback[16]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U17 ( .a ({new_AGEMA_signal_7058, new_AGEMA_signal_7056, new_AGEMA_signal_7054}), .b ({new_AGEMA_signal_1618, new_AGEMA_signal_1617, SubCellInst_SboxInst_5_n12}), .clk (clk), .r ({Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_1766, new_AGEMA_signal_1765, Feedback[22]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U8 ( .a ({new_AGEMA_signal_7070, new_AGEMA_signal_7066, new_AGEMA_signal_7062}), .b ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, SubCellInst_SboxInst_5_n3}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705]}), .c ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, Feedback[20]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U17 ( .a ({new_AGEMA_signal_7076, new_AGEMA_signal_7074, new_AGEMA_signal_7072}), .b ({new_AGEMA_signal_1628, new_AGEMA_signal_1627, SubCellInst_SboxInst_6_n12}), .clk (clk), .r ({Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_1774, new_AGEMA_signal_1773, Feedback[26]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U8 ( .a ({new_AGEMA_signal_7088, new_AGEMA_signal_7084, new_AGEMA_signal_7080}), .b ({new_AGEMA_signal_1632, new_AGEMA_signal_1631, SubCellInst_SboxInst_6_n3}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711]}), .c ({new_AGEMA_signal_1778, new_AGEMA_signal_1777, Feedback[24]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U17 ( .a ({new_AGEMA_signal_7094, new_AGEMA_signal_7092, new_AGEMA_signal_7090}), .b ({new_AGEMA_signal_1638, new_AGEMA_signal_1637, SubCellInst_SboxInst_7_n12}), .clk (clk), .r ({Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_1782, new_AGEMA_signal_1781, Feedback[30]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U8 ( .a ({new_AGEMA_signal_7106, new_AGEMA_signal_7102, new_AGEMA_signal_7098}), .b ({new_AGEMA_signal_1642, new_AGEMA_signal_1641, SubCellInst_SboxInst_7_n3}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717]}), .c ({new_AGEMA_signal_1786, new_AGEMA_signal_1785, Feedback[28]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U17 ( .a ({new_AGEMA_signal_7112, new_AGEMA_signal_7110, new_AGEMA_signal_7108}), .b ({new_AGEMA_signal_1648, new_AGEMA_signal_1647, SubCellInst_SboxInst_8_n12}), .clk (clk), .r ({Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_1790, new_AGEMA_signal_1789, Feedback[34]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U8 ( .a ({new_AGEMA_signal_7124, new_AGEMA_signal_7120, new_AGEMA_signal_7116}), .b ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, SubCellInst_SboxInst_8_n3}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723]}), .c ({new_AGEMA_signal_1794, new_AGEMA_signal_1793, Feedback[32]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U17 ( .a ({new_AGEMA_signal_7130, new_AGEMA_signal_7128, new_AGEMA_signal_7126}), .b ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, SubCellInst_SboxInst_9_n12}), .clk (clk), .r ({Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_1798, new_AGEMA_signal_1797, Feedback[38]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U8 ( .a ({new_AGEMA_signal_7142, new_AGEMA_signal_7138, new_AGEMA_signal_7134}), .b ({new_AGEMA_signal_1662, new_AGEMA_signal_1661, SubCellInst_SboxInst_9_n3}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729]}), .c ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, Feedback[36]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U17 ( .a ({new_AGEMA_signal_7148, new_AGEMA_signal_7146, new_AGEMA_signal_7144}), .b ({new_AGEMA_signal_1668, new_AGEMA_signal_1667, SubCellInst_SboxInst_10_n12}), .clk (clk), .r ({Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_1806, new_AGEMA_signal_1805, Feedback[42]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U8 ( .a ({new_AGEMA_signal_7160, new_AGEMA_signal_7156, new_AGEMA_signal_7152}), .b ({new_AGEMA_signal_1672, new_AGEMA_signal_1671, SubCellInst_SboxInst_10_n3}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735]}), .c ({new_AGEMA_signal_1810, new_AGEMA_signal_1809, Feedback[40]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U17 ( .a ({new_AGEMA_signal_7166, new_AGEMA_signal_7164, new_AGEMA_signal_7162}), .b ({new_AGEMA_signal_1678, new_AGEMA_signal_1677, SubCellInst_SboxInst_11_n12}), .clk (clk), .r ({Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_1814, new_AGEMA_signal_1813, Feedback[46]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U8 ( .a ({new_AGEMA_signal_7178, new_AGEMA_signal_7174, new_AGEMA_signal_7170}), .b ({new_AGEMA_signal_1682, new_AGEMA_signal_1681, SubCellInst_SboxInst_11_n3}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741]}), .c ({new_AGEMA_signal_1818, new_AGEMA_signal_1817, Feedback[44]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U17 ( .a ({new_AGEMA_signal_7184, new_AGEMA_signal_7182, new_AGEMA_signal_7180}), .b ({new_AGEMA_signal_1688, new_AGEMA_signal_1687, SubCellInst_SboxInst_12_n12}), .clk (clk), .r ({Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_1822, new_AGEMA_signal_1821, Feedback[50]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U8 ( .a ({new_AGEMA_signal_7196, new_AGEMA_signal_7192, new_AGEMA_signal_7188}), .b ({new_AGEMA_signal_1692, new_AGEMA_signal_1691, SubCellInst_SboxInst_12_n3}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747]}), .c ({new_AGEMA_signal_1826, new_AGEMA_signal_1825, Feedback[48]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U17 ( .a ({new_AGEMA_signal_7202, new_AGEMA_signal_7200, new_AGEMA_signal_7198}), .b ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, SubCellInst_SboxInst_13_n12}), .clk (clk), .r ({Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_1830, new_AGEMA_signal_1829, Feedback[54]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U8 ( .a ({new_AGEMA_signal_7214, new_AGEMA_signal_7210, new_AGEMA_signal_7206}), .b ({new_AGEMA_signal_1702, new_AGEMA_signal_1701, SubCellInst_SboxInst_13_n3}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753]}), .c ({new_AGEMA_signal_1834, new_AGEMA_signal_1833, Feedback[52]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U17 ( .a ({new_AGEMA_signal_7220, new_AGEMA_signal_7218, new_AGEMA_signal_7216}), .b ({new_AGEMA_signal_1708, new_AGEMA_signal_1707, SubCellInst_SboxInst_14_n12}), .clk (clk), .r ({Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_1838, new_AGEMA_signal_1837, Feedback[58]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U8 ( .a ({new_AGEMA_signal_7232, new_AGEMA_signal_7228, new_AGEMA_signal_7224}), .b ({new_AGEMA_signal_1712, new_AGEMA_signal_1711, SubCellInst_SboxInst_14_n3}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759]}), .c ({new_AGEMA_signal_1842, new_AGEMA_signal_1841, Feedback[56]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U17 ( .a ({new_AGEMA_signal_7238, new_AGEMA_signal_7236, new_AGEMA_signal_7234}), .b ({new_AGEMA_signal_1718, new_AGEMA_signal_1717, SubCellInst_SboxInst_15_n12}), .clk (clk), .r ({Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_1846, new_AGEMA_signal_1845, Feedback[62]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U8 ( .a ({new_AGEMA_signal_7250, new_AGEMA_signal_7246, new_AGEMA_signal_7242}), .b ({new_AGEMA_signal_1722, new_AGEMA_signal_1721, SubCellInst_SboxInst_15_n3}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765]}), .c ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, Feedback[60]}) ) ;
    buf_clk new_AGEMA_reg_buffer_2650 ( .C (clk), .D (new_AGEMA_signal_5425), .Q (new_AGEMA_signal_5426) ) ;
    buf_clk new_AGEMA_reg_buffer_2658 ( .C (clk), .D (new_AGEMA_signal_5433), .Q (new_AGEMA_signal_5434) ) ;
    buf_clk new_AGEMA_reg_buffer_2666 ( .C (clk), .D (new_AGEMA_signal_5441), .Q (new_AGEMA_signal_5442) ) ;
    buf_clk new_AGEMA_reg_buffer_2674 ( .C (clk), .D (new_AGEMA_signal_5449), .Q (new_AGEMA_signal_5450) ) ;
    buf_clk new_AGEMA_reg_buffer_2682 ( .C (clk), .D (new_AGEMA_signal_5457), .Q (new_AGEMA_signal_5458) ) ;
    buf_clk new_AGEMA_reg_buffer_2690 ( .C (clk), .D (new_AGEMA_signal_5465), .Q (new_AGEMA_signal_5466) ) ;
    buf_clk new_AGEMA_reg_buffer_2698 ( .C (clk), .D (new_AGEMA_signal_5473), .Q (new_AGEMA_signal_5474) ) ;
    buf_clk new_AGEMA_reg_buffer_2706 ( .C (clk), .D (new_AGEMA_signal_5481), .Q (new_AGEMA_signal_5482) ) ;
    buf_clk new_AGEMA_reg_buffer_2714 ( .C (clk), .D (new_AGEMA_signal_5489), .Q (new_AGEMA_signal_5490) ) ;
    buf_clk new_AGEMA_reg_buffer_2722 ( .C (clk), .D (new_AGEMA_signal_5497), .Q (new_AGEMA_signal_5498) ) ;
    buf_clk new_AGEMA_reg_buffer_2730 ( .C (clk), .D (new_AGEMA_signal_5505), .Q (new_AGEMA_signal_5506) ) ;
    buf_clk new_AGEMA_reg_buffer_2738 ( .C (clk), .D (new_AGEMA_signal_5513), .Q (new_AGEMA_signal_5514) ) ;
    buf_clk new_AGEMA_reg_buffer_2746 ( .C (clk), .D (new_AGEMA_signal_5521), .Q (new_AGEMA_signal_5522) ) ;
    buf_clk new_AGEMA_reg_buffer_2754 ( .C (clk), .D (new_AGEMA_signal_5529), .Q (new_AGEMA_signal_5530) ) ;
    buf_clk new_AGEMA_reg_buffer_2762 ( .C (clk), .D (new_AGEMA_signal_5537), .Q (new_AGEMA_signal_5538) ) ;
    buf_clk new_AGEMA_reg_buffer_2770 ( .C (clk), .D (new_AGEMA_signal_5545), .Q (new_AGEMA_signal_5546) ) ;
    buf_clk new_AGEMA_reg_buffer_2778 ( .C (clk), .D (new_AGEMA_signal_5553), .Q (new_AGEMA_signal_5554) ) ;
    buf_clk new_AGEMA_reg_buffer_2786 ( .C (clk), .D (new_AGEMA_signal_5561), .Q (new_AGEMA_signal_5562) ) ;
    buf_clk new_AGEMA_reg_buffer_2794 ( .C (clk), .D (new_AGEMA_signal_5569), .Q (new_AGEMA_signal_5570) ) ;
    buf_clk new_AGEMA_reg_buffer_2802 ( .C (clk), .D (new_AGEMA_signal_5577), .Q (new_AGEMA_signal_5578) ) ;
    buf_clk new_AGEMA_reg_buffer_2810 ( .C (clk), .D (new_AGEMA_signal_5585), .Q (new_AGEMA_signal_5586) ) ;
    buf_clk new_AGEMA_reg_buffer_2818 ( .C (clk), .D (new_AGEMA_signal_5593), .Q (new_AGEMA_signal_5594) ) ;
    buf_clk new_AGEMA_reg_buffer_2826 ( .C (clk), .D (new_AGEMA_signal_5601), .Q (new_AGEMA_signal_5602) ) ;
    buf_clk new_AGEMA_reg_buffer_2834 ( .C (clk), .D (new_AGEMA_signal_5609), .Q (new_AGEMA_signal_5610) ) ;
    buf_clk new_AGEMA_reg_buffer_2842 ( .C (clk), .D (new_AGEMA_signal_5617), .Q (new_AGEMA_signal_5618) ) ;
    buf_clk new_AGEMA_reg_buffer_2850 ( .C (clk), .D (new_AGEMA_signal_5625), .Q (new_AGEMA_signal_5626) ) ;
    buf_clk new_AGEMA_reg_buffer_2858 ( .C (clk), .D (new_AGEMA_signal_5633), .Q (new_AGEMA_signal_5634) ) ;
    buf_clk new_AGEMA_reg_buffer_2866 ( .C (clk), .D (new_AGEMA_signal_5641), .Q (new_AGEMA_signal_5642) ) ;
    buf_clk new_AGEMA_reg_buffer_2874 ( .C (clk), .D (new_AGEMA_signal_5649), .Q (new_AGEMA_signal_5650) ) ;
    buf_clk new_AGEMA_reg_buffer_2882 ( .C (clk), .D (new_AGEMA_signal_5657), .Q (new_AGEMA_signal_5658) ) ;
    buf_clk new_AGEMA_reg_buffer_2890 ( .C (clk), .D (new_AGEMA_signal_5665), .Q (new_AGEMA_signal_5666) ) ;
    buf_clk new_AGEMA_reg_buffer_2898 ( .C (clk), .D (new_AGEMA_signal_5673), .Q (new_AGEMA_signal_5674) ) ;
    buf_clk new_AGEMA_reg_buffer_2906 ( .C (clk), .D (new_AGEMA_signal_5681), .Q (new_AGEMA_signal_5682) ) ;
    buf_clk new_AGEMA_reg_buffer_2914 ( .C (clk), .D (new_AGEMA_signal_5689), .Q (new_AGEMA_signal_5690) ) ;
    buf_clk new_AGEMA_reg_buffer_2922 ( .C (clk), .D (new_AGEMA_signal_5697), .Q (new_AGEMA_signal_5698) ) ;
    buf_clk new_AGEMA_reg_buffer_2930 ( .C (clk), .D (new_AGEMA_signal_5705), .Q (new_AGEMA_signal_5706) ) ;
    buf_clk new_AGEMA_reg_buffer_2938 ( .C (clk), .D (new_AGEMA_signal_5713), .Q (new_AGEMA_signal_5714) ) ;
    buf_clk new_AGEMA_reg_buffer_2946 ( .C (clk), .D (new_AGEMA_signal_5721), .Q (new_AGEMA_signal_5722) ) ;
    buf_clk new_AGEMA_reg_buffer_2954 ( .C (clk), .D (new_AGEMA_signal_5729), .Q (new_AGEMA_signal_5730) ) ;
    buf_clk new_AGEMA_reg_buffer_2962 ( .C (clk), .D (new_AGEMA_signal_5737), .Q (new_AGEMA_signal_5738) ) ;
    buf_clk new_AGEMA_reg_buffer_2970 ( .C (clk), .D (new_AGEMA_signal_5745), .Q (new_AGEMA_signal_5746) ) ;
    buf_clk new_AGEMA_reg_buffer_2978 ( .C (clk), .D (new_AGEMA_signal_5753), .Q (new_AGEMA_signal_5754) ) ;
    buf_clk new_AGEMA_reg_buffer_2986 ( .C (clk), .D (new_AGEMA_signal_5761), .Q (new_AGEMA_signal_5762) ) ;
    buf_clk new_AGEMA_reg_buffer_2994 ( .C (clk), .D (new_AGEMA_signal_5769), .Q (new_AGEMA_signal_5770) ) ;
    buf_clk new_AGEMA_reg_buffer_3002 ( .C (clk), .D (new_AGEMA_signal_5777), .Q (new_AGEMA_signal_5778) ) ;
    buf_clk new_AGEMA_reg_buffer_3010 ( .C (clk), .D (new_AGEMA_signal_5785), .Q (new_AGEMA_signal_5786) ) ;
    buf_clk new_AGEMA_reg_buffer_3018 ( .C (clk), .D (new_AGEMA_signal_5793), .Q (new_AGEMA_signal_5794) ) ;
    buf_clk new_AGEMA_reg_buffer_3026 ( .C (clk), .D (new_AGEMA_signal_5801), .Q (new_AGEMA_signal_5802) ) ;
    buf_clk new_AGEMA_reg_buffer_3034 ( .C (clk), .D (new_AGEMA_signal_5809), .Q (new_AGEMA_signal_5810) ) ;
    buf_clk new_AGEMA_reg_buffer_3042 ( .C (clk), .D (new_AGEMA_signal_5817), .Q (new_AGEMA_signal_5818) ) ;
    buf_clk new_AGEMA_reg_buffer_3050 ( .C (clk), .D (new_AGEMA_signal_5825), .Q (new_AGEMA_signal_5826) ) ;
    buf_clk new_AGEMA_reg_buffer_3058 ( .C (clk), .D (new_AGEMA_signal_5833), .Q (new_AGEMA_signal_5834) ) ;
    buf_clk new_AGEMA_reg_buffer_3066 ( .C (clk), .D (new_AGEMA_signal_5841), .Q (new_AGEMA_signal_5842) ) ;
    buf_clk new_AGEMA_reg_buffer_3074 ( .C (clk), .D (new_AGEMA_signal_5849), .Q (new_AGEMA_signal_5850) ) ;
    buf_clk new_AGEMA_reg_buffer_3082 ( .C (clk), .D (new_AGEMA_signal_5857), .Q (new_AGEMA_signal_5858) ) ;
    buf_clk new_AGEMA_reg_buffer_3090 ( .C (clk), .D (new_AGEMA_signal_5865), .Q (new_AGEMA_signal_5866) ) ;
    buf_clk new_AGEMA_reg_buffer_3098 ( .C (clk), .D (new_AGEMA_signal_5873), .Q (new_AGEMA_signal_5874) ) ;
    buf_clk new_AGEMA_reg_buffer_3106 ( .C (clk), .D (new_AGEMA_signal_5881), .Q (new_AGEMA_signal_5882) ) ;
    buf_clk new_AGEMA_reg_buffer_3114 ( .C (clk), .D (new_AGEMA_signal_5889), .Q (new_AGEMA_signal_5890) ) ;
    buf_clk new_AGEMA_reg_buffer_3122 ( .C (clk), .D (new_AGEMA_signal_5897), .Q (new_AGEMA_signal_5898) ) ;
    buf_clk new_AGEMA_reg_buffer_3130 ( .C (clk), .D (new_AGEMA_signal_5905), .Q (new_AGEMA_signal_5906) ) ;
    buf_clk new_AGEMA_reg_buffer_3138 ( .C (clk), .D (new_AGEMA_signal_5913), .Q (new_AGEMA_signal_5914) ) ;
    buf_clk new_AGEMA_reg_buffer_3146 ( .C (clk), .D (new_AGEMA_signal_5921), .Q (new_AGEMA_signal_5922) ) ;
    buf_clk new_AGEMA_reg_buffer_3154 ( .C (clk), .D (new_AGEMA_signal_5929), .Q (new_AGEMA_signal_5930) ) ;
    buf_clk new_AGEMA_reg_buffer_3162 ( .C (clk), .D (new_AGEMA_signal_5937), .Q (new_AGEMA_signal_5938) ) ;
    buf_clk new_AGEMA_reg_buffer_3170 ( .C (clk), .D (new_AGEMA_signal_5945), .Q (new_AGEMA_signal_5946) ) ;
    buf_clk new_AGEMA_reg_buffer_3178 ( .C (clk), .D (new_AGEMA_signal_5953), .Q (new_AGEMA_signal_5954) ) ;
    buf_clk new_AGEMA_reg_buffer_3186 ( .C (clk), .D (new_AGEMA_signal_5961), .Q (new_AGEMA_signal_5962) ) ;
    buf_clk new_AGEMA_reg_buffer_3194 ( .C (clk), .D (new_AGEMA_signal_5969), .Q (new_AGEMA_signal_5970) ) ;
    buf_clk new_AGEMA_reg_buffer_3202 ( .C (clk), .D (new_AGEMA_signal_5977), .Q (new_AGEMA_signal_5978) ) ;
    buf_clk new_AGEMA_reg_buffer_3210 ( .C (clk), .D (new_AGEMA_signal_5985), .Q (new_AGEMA_signal_5986) ) ;
    buf_clk new_AGEMA_reg_buffer_3218 ( .C (clk), .D (new_AGEMA_signal_5993), .Q (new_AGEMA_signal_5994) ) ;
    buf_clk new_AGEMA_reg_buffer_3226 ( .C (clk), .D (new_AGEMA_signal_6001), .Q (new_AGEMA_signal_6002) ) ;
    buf_clk new_AGEMA_reg_buffer_3234 ( .C (clk), .D (new_AGEMA_signal_6009), .Q (new_AGEMA_signal_6010) ) ;
    buf_clk new_AGEMA_reg_buffer_3242 ( .C (clk), .D (new_AGEMA_signal_6017), .Q (new_AGEMA_signal_6018) ) ;
    buf_clk new_AGEMA_reg_buffer_3250 ( .C (clk), .D (new_AGEMA_signal_6025), .Q (new_AGEMA_signal_6026) ) ;
    buf_clk new_AGEMA_reg_buffer_3258 ( .C (clk), .D (new_AGEMA_signal_6033), .Q (new_AGEMA_signal_6034) ) ;
    buf_clk new_AGEMA_reg_buffer_3266 ( .C (clk), .D (new_AGEMA_signal_6041), .Q (new_AGEMA_signal_6042) ) ;
    buf_clk new_AGEMA_reg_buffer_3274 ( .C (clk), .D (new_AGEMA_signal_6049), .Q (new_AGEMA_signal_6050) ) ;
    buf_clk new_AGEMA_reg_buffer_3282 ( .C (clk), .D (new_AGEMA_signal_6057), .Q (new_AGEMA_signal_6058) ) ;
    buf_clk new_AGEMA_reg_buffer_3290 ( .C (clk), .D (new_AGEMA_signal_6065), .Q (new_AGEMA_signal_6066) ) ;
    buf_clk new_AGEMA_reg_buffer_3298 ( .C (clk), .D (new_AGEMA_signal_6073), .Q (new_AGEMA_signal_6074) ) ;
    buf_clk new_AGEMA_reg_buffer_3306 ( .C (clk), .D (new_AGEMA_signal_6081), .Q (new_AGEMA_signal_6082) ) ;
    buf_clk new_AGEMA_reg_buffer_3314 ( .C (clk), .D (new_AGEMA_signal_6089), .Q (new_AGEMA_signal_6090) ) ;
    buf_clk new_AGEMA_reg_buffer_3322 ( .C (clk), .D (new_AGEMA_signal_6097), .Q (new_AGEMA_signal_6098) ) ;
    buf_clk new_AGEMA_reg_buffer_3330 ( .C (clk), .D (new_AGEMA_signal_6105), .Q (new_AGEMA_signal_6106) ) ;
    buf_clk new_AGEMA_reg_buffer_3338 ( .C (clk), .D (new_AGEMA_signal_6113), .Q (new_AGEMA_signal_6114) ) ;
    buf_clk new_AGEMA_reg_buffer_3346 ( .C (clk), .D (new_AGEMA_signal_6121), .Q (new_AGEMA_signal_6122) ) ;
    buf_clk new_AGEMA_reg_buffer_3354 ( .C (clk), .D (new_AGEMA_signal_6129), .Q (new_AGEMA_signal_6130) ) ;
    buf_clk new_AGEMA_reg_buffer_3362 ( .C (clk), .D (new_AGEMA_signal_6137), .Q (new_AGEMA_signal_6138) ) ;
    buf_clk new_AGEMA_reg_buffer_3370 ( .C (clk), .D (new_AGEMA_signal_6145), .Q (new_AGEMA_signal_6146) ) ;
    buf_clk new_AGEMA_reg_buffer_3378 ( .C (clk), .D (new_AGEMA_signal_6153), .Q (new_AGEMA_signal_6154) ) ;
    buf_clk new_AGEMA_reg_buffer_3386 ( .C (clk), .D (new_AGEMA_signal_6161), .Q (new_AGEMA_signal_6162) ) ;
    buf_clk new_AGEMA_reg_buffer_3394 ( .C (clk), .D (new_AGEMA_signal_6169), .Q (new_AGEMA_signal_6170) ) ;
    buf_clk new_AGEMA_reg_buffer_3402 ( .C (clk), .D (new_AGEMA_signal_6177), .Q (new_AGEMA_signal_6178) ) ;
    buf_clk new_AGEMA_reg_buffer_3410 ( .C (clk), .D (new_AGEMA_signal_6185), .Q (new_AGEMA_signal_6186) ) ;
    buf_clk new_AGEMA_reg_buffer_3418 ( .C (clk), .D (new_AGEMA_signal_6193), .Q (new_AGEMA_signal_6194) ) ;
    buf_clk new_AGEMA_reg_buffer_3426 ( .C (clk), .D (new_AGEMA_signal_6201), .Q (new_AGEMA_signal_6202) ) ;
    buf_clk new_AGEMA_reg_buffer_3434 ( .C (clk), .D (new_AGEMA_signal_6209), .Q (new_AGEMA_signal_6210) ) ;
    buf_clk new_AGEMA_reg_buffer_3442 ( .C (clk), .D (new_AGEMA_signal_6217), .Q (new_AGEMA_signal_6218) ) ;
    buf_clk new_AGEMA_reg_buffer_3450 ( .C (clk), .D (new_AGEMA_signal_6225), .Q (new_AGEMA_signal_6226) ) ;
    buf_clk new_AGEMA_reg_buffer_3458 ( .C (clk), .D (new_AGEMA_signal_6233), .Q (new_AGEMA_signal_6234) ) ;
    buf_clk new_AGEMA_reg_buffer_3466 ( .C (clk), .D (new_AGEMA_signal_6241), .Q (new_AGEMA_signal_6242) ) ;
    buf_clk new_AGEMA_reg_buffer_3474 ( .C (clk), .D (new_AGEMA_signal_6249), .Q (new_AGEMA_signal_6250) ) ;
    buf_clk new_AGEMA_reg_buffer_3482 ( .C (clk), .D (new_AGEMA_signal_6257), .Q (new_AGEMA_signal_6258) ) ;
    buf_clk new_AGEMA_reg_buffer_3490 ( .C (clk), .D (new_AGEMA_signal_6265), .Q (new_AGEMA_signal_6266) ) ;
    buf_clk new_AGEMA_reg_buffer_3498 ( .C (clk), .D (new_AGEMA_signal_6273), .Q (new_AGEMA_signal_6274) ) ;
    buf_clk new_AGEMA_reg_buffer_3506 ( .C (clk), .D (new_AGEMA_signal_6281), .Q (new_AGEMA_signal_6282) ) ;
    buf_clk new_AGEMA_reg_buffer_3514 ( .C (clk), .D (new_AGEMA_signal_6289), .Q (new_AGEMA_signal_6290) ) ;
    buf_clk new_AGEMA_reg_buffer_3522 ( .C (clk), .D (new_AGEMA_signal_6297), .Q (new_AGEMA_signal_6298) ) ;
    buf_clk new_AGEMA_reg_buffer_3530 ( .C (clk), .D (new_AGEMA_signal_6305), .Q (new_AGEMA_signal_6306) ) ;
    buf_clk new_AGEMA_reg_buffer_3538 ( .C (clk), .D (new_AGEMA_signal_6313), .Q (new_AGEMA_signal_6314) ) ;
    buf_clk new_AGEMA_reg_buffer_3546 ( .C (clk), .D (new_AGEMA_signal_6321), .Q (new_AGEMA_signal_6322) ) ;
    buf_clk new_AGEMA_reg_buffer_3554 ( .C (clk), .D (new_AGEMA_signal_6329), .Q (new_AGEMA_signal_6330) ) ;
    buf_clk new_AGEMA_reg_buffer_3562 ( .C (clk), .D (new_AGEMA_signal_6337), .Q (new_AGEMA_signal_6338) ) ;
    buf_clk new_AGEMA_reg_buffer_3570 ( .C (clk), .D (new_AGEMA_signal_6345), .Q (new_AGEMA_signal_6346) ) ;
    buf_clk new_AGEMA_reg_buffer_3578 ( .C (clk), .D (new_AGEMA_signal_6353), .Q (new_AGEMA_signal_6354) ) ;
    buf_clk new_AGEMA_reg_buffer_3586 ( .C (clk), .D (new_AGEMA_signal_6361), .Q (new_AGEMA_signal_6362) ) ;
    buf_clk new_AGEMA_reg_buffer_3594 ( .C (clk), .D (new_AGEMA_signal_6369), .Q (new_AGEMA_signal_6370) ) ;
    buf_clk new_AGEMA_reg_buffer_3602 ( .C (clk), .D (new_AGEMA_signal_6377), .Q (new_AGEMA_signal_6378) ) ;
    buf_clk new_AGEMA_reg_buffer_3610 ( .C (clk), .D (new_AGEMA_signal_6385), .Q (new_AGEMA_signal_6386) ) ;
    buf_clk new_AGEMA_reg_buffer_3618 ( .C (clk), .D (new_AGEMA_signal_6393), .Q (new_AGEMA_signal_6394) ) ;
    buf_clk new_AGEMA_reg_buffer_3626 ( .C (clk), .D (new_AGEMA_signal_6401), .Q (new_AGEMA_signal_6402) ) ;
    buf_clk new_AGEMA_reg_buffer_3634 ( .C (clk), .D (new_AGEMA_signal_6409), .Q (new_AGEMA_signal_6410) ) ;
    buf_clk new_AGEMA_reg_buffer_3642 ( .C (clk), .D (new_AGEMA_signal_6417), .Q (new_AGEMA_signal_6418) ) ;
    buf_clk new_AGEMA_reg_buffer_3650 ( .C (clk), .D (new_AGEMA_signal_6425), .Q (new_AGEMA_signal_6426) ) ;
    buf_clk new_AGEMA_reg_buffer_3658 ( .C (clk), .D (new_AGEMA_signal_6433), .Q (new_AGEMA_signal_6434) ) ;
    buf_clk new_AGEMA_reg_buffer_3666 ( .C (clk), .D (new_AGEMA_signal_6441), .Q (new_AGEMA_signal_6442) ) ;
    buf_clk new_AGEMA_reg_buffer_3674 ( .C (clk), .D (new_AGEMA_signal_6449), .Q (new_AGEMA_signal_6450) ) ;
    buf_clk new_AGEMA_reg_buffer_3682 ( .C (clk), .D (new_AGEMA_signal_6457), .Q (new_AGEMA_signal_6458) ) ;
    buf_clk new_AGEMA_reg_buffer_3690 ( .C (clk), .D (new_AGEMA_signal_6465), .Q (new_AGEMA_signal_6466) ) ;
    buf_clk new_AGEMA_reg_buffer_3698 ( .C (clk), .D (new_AGEMA_signal_6473), .Q (new_AGEMA_signal_6474) ) ;
    buf_clk new_AGEMA_reg_buffer_3706 ( .C (clk), .D (new_AGEMA_signal_6481), .Q (new_AGEMA_signal_6482) ) ;
    buf_clk new_AGEMA_reg_buffer_3714 ( .C (clk), .D (new_AGEMA_signal_6489), .Q (new_AGEMA_signal_6490) ) ;
    buf_clk new_AGEMA_reg_buffer_3722 ( .C (clk), .D (new_AGEMA_signal_6497), .Q (new_AGEMA_signal_6498) ) ;
    buf_clk new_AGEMA_reg_buffer_3730 ( .C (clk), .D (new_AGEMA_signal_6505), .Q (new_AGEMA_signal_6506) ) ;
    buf_clk new_AGEMA_reg_buffer_3738 ( .C (clk), .D (new_AGEMA_signal_6513), .Q (new_AGEMA_signal_6514) ) ;
    buf_clk new_AGEMA_reg_buffer_3746 ( .C (clk), .D (new_AGEMA_signal_6521), .Q (new_AGEMA_signal_6522) ) ;
    buf_clk new_AGEMA_reg_buffer_3754 ( .C (clk), .D (new_AGEMA_signal_6529), .Q (new_AGEMA_signal_6530) ) ;
    buf_clk new_AGEMA_reg_buffer_3762 ( .C (clk), .D (new_AGEMA_signal_6537), .Q (new_AGEMA_signal_6538) ) ;
    buf_clk new_AGEMA_reg_buffer_3770 ( .C (clk), .D (new_AGEMA_signal_6545), .Q (new_AGEMA_signal_6546) ) ;
    buf_clk new_AGEMA_reg_buffer_3778 ( .C (clk), .D (new_AGEMA_signal_6553), .Q (new_AGEMA_signal_6554) ) ;
    buf_clk new_AGEMA_reg_buffer_3786 ( .C (clk), .D (new_AGEMA_signal_6561), .Q (new_AGEMA_signal_6562) ) ;
    buf_clk new_AGEMA_reg_buffer_3794 ( .C (clk), .D (new_AGEMA_signal_6569), .Q (new_AGEMA_signal_6570) ) ;
    buf_clk new_AGEMA_reg_buffer_3802 ( .C (clk), .D (new_AGEMA_signal_6577), .Q (new_AGEMA_signal_6578) ) ;
    buf_clk new_AGEMA_reg_buffer_3810 ( .C (clk), .D (new_AGEMA_signal_6585), .Q (new_AGEMA_signal_6586) ) ;
    buf_clk new_AGEMA_reg_buffer_3818 ( .C (clk), .D (new_AGEMA_signal_6593), .Q (new_AGEMA_signal_6594) ) ;
    buf_clk new_AGEMA_reg_buffer_3826 ( .C (clk), .D (new_AGEMA_signal_6601), .Q (new_AGEMA_signal_6602) ) ;
    buf_clk new_AGEMA_reg_buffer_3834 ( .C (clk), .D (new_AGEMA_signal_6609), .Q (new_AGEMA_signal_6610) ) ;
    buf_clk new_AGEMA_reg_buffer_3842 ( .C (clk), .D (new_AGEMA_signal_6617), .Q (new_AGEMA_signal_6618) ) ;
    buf_clk new_AGEMA_reg_buffer_3850 ( .C (clk), .D (new_AGEMA_signal_6625), .Q (new_AGEMA_signal_6626) ) ;
    buf_clk new_AGEMA_reg_buffer_3858 ( .C (clk), .D (new_AGEMA_signal_6633), .Q (new_AGEMA_signal_6634) ) ;
    buf_clk new_AGEMA_reg_buffer_3866 ( .C (clk), .D (new_AGEMA_signal_6641), .Q (new_AGEMA_signal_6642) ) ;
    buf_clk new_AGEMA_reg_buffer_3874 ( .C (clk), .D (new_AGEMA_signal_6649), .Q (new_AGEMA_signal_6650) ) ;
    buf_clk new_AGEMA_reg_buffer_3882 ( .C (clk), .D (new_AGEMA_signal_6657), .Q (new_AGEMA_signal_6658) ) ;
    buf_clk new_AGEMA_reg_buffer_3890 ( .C (clk), .D (new_AGEMA_signal_6665), .Q (new_AGEMA_signal_6666) ) ;
    buf_clk new_AGEMA_reg_buffer_3898 ( .C (clk), .D (new_AGEMA_signal_6673), .Q (new_AGEMA_signal_6674) ) ;
    buf_clk new_AGEMA_reg_buffer_3906 ( .C (clk), .D (new_AGEMA_signal_6681), .Q (new_AGEMA_signal_6682) ) ;
    buf_clk new_AGEMA_reg_buffer_3914 ( .C (clk), .D (new_AGEMA_signal_6689), .Q (new_AGEMA_signal_6690) ) ;
    buf_clk new_AGEMA_reg_buffer_3922 ( .C (clk), .D (new_AGEMA_signal_6697), .Q (new_AGEMA_signal_6698) ) ;
    buf_clk new_AGEMA_reg_buffer_3930 ( .C (clk), .D (new_AGEMA_signal_6705), .Q (new_AGEMA_signal_6706) ) ;
    buf_clk new_AGEMA_reg_buffer_3938 ( .C (clk), .D (new_AGEMA_signal_6713), .Q (new_AGEMA_signal_6714) ) ;
    buf_clk new_AGEMA_reg_buffer_3946 ( .C (clk), .D (new_AGEMA_signal_6721), .Q (new_AGEMA_signal_6722) ) ;
    buf_clk new_AGEMA_reg_buffer_3954 ( .C (clk), .D (new_AGEMA_signal_6729), .Q (new_AGEMA_signal_6730) ) ;
    buf_clk new_AGEMA_reg_buffer_3962 ( .C (clk), .D (new_AGEMA_signal_6737), .Q (new_AGEMA_signal_6738) ) ;
    buf_clk new_AGEMA_reg_buffer_3970 ( .C (clk), .D (new_AGEMA_signal_6745), .Q (new_AGEMA_signal_6746) ) ;
    buf_clk new_AGEMA_reg_buffer_3978 ( .C (clk), .D (new_AGEMA_signal_6753), .Q (new_AGEMA_signal_6754) ) ;
    buf_clk new_AGEMA_reg_buffer_3986 ( .C (clk), .D (new_AGEMA_signal_6761), .Q (new_AGEMA_signal_6762) ) ;
    buf_clk new_AGEMA_reg_buffer_3994 ( .C (clk), .D (new_AGEMA_signal_6769), .Q (new_AGEMA_signal_6770) ) ;
    buf_clk new_AGEMA_reg_buffer_4002 ( .C (clk), .D (new_AGEMA_signal_6777), .Q (new_AGEMA_signal_6778) ) ;
    buf_clk new_AGEMA_reg_buffer_4010 ( .C (clk), .D (new_AGEMA_signal_6785), .Q (new_AGEMA_signal_6786) ) ;
    buf_clk new_AGEMA_reg_buffer_4018 ( .C (clk), .D (new_AGEMA_signal_6793), .Q (new_AGEMA_signal_6794) ) ;
    buf_clk new_AGEMA_reg_buffer_4026 ( .C (clk), .D (new_AGEMA_signal_6801), .Q (new_AGEMA_signal_6802) ) ;
    buf_clk new_AGEMA_reg_buffer_4034 ( .C (clk), .D (new_AGEMA_signal_6809), .Q (new_AGEMA_signal_6810) ) ;
    buf_clk new_AGEMA_reg_buffer_4042 ( .C (clk), .D (new_AGEMA_signal_6817), .Q (new_AGEMA_signal_6818) ) ;
    buf_clk new_AGEMA_reg_buffer_4050 ( .C (clk), .D (new_AGEMA_signal_6825), .Q (new_AGEMA_signal_6826) ) ;
    buf_clk new_AGEMA_reg_buffer_4058 ( .C (clk), .D (new_AGEMA_signal_6833), .Q (new_AGEMA_signal_6834) ) ;
    buf_clk new_AGEMA_reg_buffer_4066 ( .C (clk), .D (new_AGEMA_signal_6841), .Q (new_AGEMA_signal_6842) ) ;
    buf_clk new_AGEMA_reg_buffer_4074 ( .C (clk), .D (new_AGEMA_signal_6849), .Q (new_AGEMA_signal_6850) ) ;
    buf_clk new_AGEMA_reg_buffer_4082 ( .C (clk), .D (new_AGEMA_signal_6857), .Q (new_AGEMA_signal_6858) ) ;
    buf_clk new_AGEMA_reg_buffer_4090 ( .C (clk), .D (new_AGEMA_signal_6865), .Q (new_AGEMA_signal_6866) ) ;
    buf_clk new_AGEMA_reg_buffer_4098 ( .C (clk), .D (new_AGEMA_signal_6873), .Q (new_AGEMA_signal_6874) ) ;
    buf_clk new_AGEMA_reg_buffer_4106 ( .C (clk), .D (new_AGEMA_signal_6881), .Q (new_AGEMA_signal_6882) ) ;
    buf_clk new_AGEMA_reg_buffer_4114 ( .C (clk), .D (new_AGEMA_signal_6889), .Q (new_AGEMA_signal_6890) ) ;
    buf_clk new_AGEMA_reg_buffer_4122 ( .C (clk), .D (new_AGEMA_signal_6897), .Q (new_AGEMA_signal_6898) ) ;
    buf_clk new_AGEMA_reg_buffer_4130 ( .C (clk), .D (new_AGEMA_signal_6905), .Q (new_AGEMA_signal_6906) ) ;
    buf_clk new_AGEMA_reg_buffer_4138 ( .C (clk), .D (new_AGEMA_signal_6913), .Q (new_AGEMA_signal_6914) ) ;
    buf_clk new_AGEMA_reg_buffer_4146 ( .C (clk), .D (new_AGEMA_signal_6921), .Q (new_AGEMA_signal_6922) ) ;
    buf_clk new_AGEMA_reg_buffer_4154 ( .C (clk), .D (new_AGEMA_signal_6929), .Q (new_AGEMA_signal_6930) ) ;
    buf_clk new_AGEMA_reg_buffer_4162 ( .C (clk), .D (new_AGEMA_signal_6937), .Q (new_AGEMA_signal_6938) ) ;
    buf_clk new_AGEMA_reg_buffer_4170 ( .C (clk), .D (new_AGEMA_signal_6945), .Q (new_AGEMA_signal_6946) ) ;
    buf_clk new_AGEMA_reg_buffer_4178 ( .C (clk), .D (new_AGEMA_signal_6953), .Q (new_AGEMA_signal_6954) ) ;
    buf_clk new_AGEMA_reg_buffer_4186 ( .C (clk), .D (new_AGEMA_signal_6961), .Q (new_AGEMA_signal_6962) ) ;
    buf_clk new_AGEMA_reg_buffer_4476 ( .C (clk), .D (new_AGEMA_signal_7251), .Q (new_AGEMA_signal_7252) ) ;
    buf_clk new_AGEMA_reg_buffer_4478 ( .C (clk), .D (new_AGEMA_signal_7253), .Q (new_AGEMA_signal_7254) ) ;
    buf_clk new_AGEMA_reg_buffer_4480 ( .C (clk), .D (new_AGEMA_signal_7255), .Q (new_AGEMA_signal_7256) ) ;
    buf_clk new_AGEMA_reg_buffer_4482 ( .C (clk), .D (new_AGEMA_signal_7257), .Q (new_AGEMA_signal_7258) ) ;
    buf_clk new_AGEMA_reg_buffer_4484 ( .C (clk), .D (new_AGEMA_signal_7259), .Q (new_AGEMA_signal_7260) ) ;
    buf_clk new_AGEMA_reg_buffer_4486 ( .C (clk), .D (new_AGEMA_signal_7261), .Q (new_AGEMA_signal_7262) ) ;
    buf_clk new_AGEMA_reg_buffer_4488 ( .C (clk), .D (new_AGEMA_signal_7263), .Q (new_AGEMA_signal_7264) ) ;
    buf_clk new_AGEMA_reg_buffer_4490 ( .C (clk), .D (new_AGEMA_signal_7265), .Q (new_AGEMA_signal_7266) ) ;
    buf_clk new_AGEMA_reg_buffer_4492 ( .C (clk), .D (new_AGEMA_signal_7267), .Q (new_AGEMA_signal_7268) ) ;
    buf_clk new_AGEMA_reg_buffer_4494 ( .C (clk), .D (new_AGEMA_signal_7269), .Q (new_AGEMA_signal_7270) ) ;
    buf_clk new_AGEMA_reg_buffer_4496 ( .C (clk), .D (new_AGEMA_signal_7271), .Q (new_AGEMA_signal_7272) ) ;
    buf_clk new_AGEMA_reg_buffer_4498 ( .C (clk), .D (new_AGEMA_signal_7273), .Q (new_AGEMA_signal_7274) ) ;
    buf_clk new_AGEMA_reg_buffer_4500 ( .C (clk), .D (new_AGEMA_signal_7275), .Q (new_AGEMA_signal_7276) ) ;
    buf_clk new_AGEMA_reg_buffer_4502 ( .C (clk), .D (new_AGEMA_signal_7277), .Q (new_AGEMA_signal_7278) ) ;
    buf_clk new_AGEMA_reg_buffer_4504 ( .C (clk), .D (new_AGEMA_signal_7279), .Q (new_AGEMA_signal_7280) ) ;
    buf_clk new_AGEMA_reg_buffer_4506 ( .C (clk), .D (new_AGEMA_signal_7281), .Q (new_AGEMA_signal_7282) ) ;
    buf_clk new_AGEMA_reg_buffer_4508 ( .C (clk), .D (new_AGEMA_signal_7283), .Q (new_AGEMA_signal_7284) ) ;
    buf_clk new_AGEMA_reg_buffer_4510 ( .C (clk), .D (new_AGEMA_signal_7285), .Q (new_AGEMA_signal_7286) ) ;
    buf_clk new_AGEMA_reg_buffer_4512 ( .C (clk), .D (new_AGEMA_signal_7287), .Q (new_AGEMA_signal_7288) ) ;
    buf_clk new_AGEMA_reg_buffer_4514 ( .C (clk), .D (new_AGEMA_signal_7289), .Q (new_AGEMA_signal_7290) ) ;
    buf_clk new_AGEMA_reg_buffer_4516 ( .C (clk), .D (new_AGEMA_signal_7291), .Q (new_AGEMA_signal_7292) ) ;
    buf_clk new_AGEMA_reg_buffer_4518 ( .C (clk), .D (new_AGEMA_signal_7293), .Q (new_AGEMA_signal_7294) ) ;
    buf_clk new_AGEMA_reg_buffer_4520 ( .C (clk), .D (new_AGEMA_signal_7295), .Q (new_AGEMA_signal_7296) ) ;
    buf_clk new_AGEMA_reg_buffer_4522 ( .C (clk), .D (new_AGEMA_signal_7297), .Q (new_AGEMA_signal_7298) ) ;
    buf_clk new_AGEMA_reg_buffer_4524 ( .C (clk), .D (new_AGEMA_signal_7299), .Q (new_AGEMA_signal_7300) ) ;
    buf_clk new_AGEMA_reg_buffer_4526 ( .C (clk), .D (new_AGEMA_signal_7301), .Q (new_AGEMA_signal_7302) ) ;
    buf_clk new_AGEMA_reg_buffer_4528 ( .C (clk), .D (new_AGEMA_signal_7303), .Q (new_AGEMA_signal_7304) ) ;
    buf_clk new_AGEMA_reg_buffer_4530 ( .C (clk), .D (new_AGEMA_signal_7305), .Q (new_AGEMA_signal_7306) ) ;
    buf_clk new_AGEMA_reg_buffer_4532 ( .C (clk), .D (new_AGEMA_signal_7307), .Q (new_AGEMA_signal_7308) ) ;
    buf_clk new_AGEMA_reg_buffer_4534 ( .C (clk), .D (new_AGEMA_signal_7309), .Q (new_AGEMA_signal_7310) ) ;
    buf_clk new_AGEMA_reg_buffer_4536 ( .C (clk), .D (new_AGEMA_signal_7311), .Q (new_AGEMA_signal_7312) ) ;
    buf_clk new_AGEMA_reg_buffer_4538 ( .C (clk), .D (new_AGEMA_signal_7313), .Q (new_AGEMA_signal_7314) ) ;
    buf_clk new_AGEMA_reg_buffer_4540 ( .C (clk), .D (new_AGEMA_signal_7315), .Q (new_AGEMA_signal_7316) ) ;
    buf_clk new_AGEMA_reg_buffer_4542 ( .C (clk), .D (new_AGEMA_signal_7317), .Q (new_AGEMA_signal_7318) ) ;
    buf_clk new_AGEMA_reg_buffer_4544 ( .C (clk), .D (new_AGEMA_signal_7319), .Q (new_AGEMA_signal_7320) ) ;
    buf_clk new_AGEMA_reg_buffer_4546 ( .C (clk), .D (new_AGEMA_signal_7321), .Q (new_AGEMA_signal_7322) ) ;
    buf_clk new_AGEMA_reg_buffer_4548 ( .C (clk), .D (new_AGEMA_signal_7323), .Q (new_AGEMA_signal_7324) ) ;
    buf_clk new_AGEMA_reg_buffer_4550 ( .C (clk), .D (new_AGEMA_signal_7325), .Q (new_AGEMA_signal_7326) ) ;
    buf_clk new_AGEMA_reg_buffer_4552 ( .C (clk), .D (new_AGEMA_signal_7327), .Q (new_AGEMA_signal_7328) ) ;
    buf_clk new_AGEMA_reg_buffer_4554 ( .C (clk), .D (new_AGEMA_signal_7329), .Q (new_AGEMA_signal_7330) ) ;
    buf_clk new_AGEMA_reg_buffer_4556 ( .C (clk), .D (new_AGEMA_signal_7331), .Q (new_AGEMA_signal_7332) ) ;
    buf_clk new_AGEMA_reg_buffer_4558 ( .C (clk), .D (new_AGEMA_signal_7333), .Q (new_AGEMA_signal_7334) ) ;
    buf_clk new_AGEMA_reg_buffer_4560 ( .C (clk), .D (new_AGEMA_signal_7335), .Q (new_AGEMA_signal_7336) ) ;
    buf_clk new_AGEMA_reg_buffer_4562 ( .C (clk), .D (new_AGEMA_signal_7337), .Q (new_AGEMA_signal_7338) ) ;
    buf_clk new_AGEMA_reg_buffer_4564 ( .C (clk), .D (new_AGEMA_signal_7339), .Q (new_AGEMA_signal_7340) ) ;
    buf_clk new_AGEMA_reg_buffer_4566 ( .C (clk), .D (new_AGEMA_signal_7341), .Q (new_AGEMA_signal_7342) ) ;
    buf_clk new_AGEMA_reg_buffer_4568 ( .C (clk), .D (new_AGEMA_signal_7343), .Q (new_AGEMA_signal_7344) ) ;
    buf_clk new_AGEMA_reg_buffer_4570 ( .C (clk), .D (new_AGEMA_signal_7345), .Q (new_AGEMA_signal_7346) ) ;
    buf_clk new_AGEMA_reg_buffer_4572 ( .C (clk), .D (new_AGEMA_signal_7347), .Q (new_AGEMA_signal_7348) ) ;
    buf_clk new_AGEMA_reg_buffer_4574 ( .C (clk), .D (new_AGEMA_signal_7349), .Q (new_AGEMA_signal_7350) ) ;
    buf_clk new_AGEMA_reg_buffer_4576 ( .C (clk), .D (new_AGEMA_signal_7351), .Q (new_AGEMA_signal_7352) ) ;
    buf_clk new_AGEMA_reg_buffer_4578 ( .C (clk), .D (new_AGEMA_signal_7353), .Q (new_AGEMA_signal_7354) ) ;
    buf_clk new_AGEMA_reg_buffer_4580 ( .C (clk), .D (new_AGEMA_signal_7355), .Q (new_AGEMA_signal_7356) ) ;
    buf_clk new_AGEMA_reg_buffer_4582 ( .C (clk), .D (new_AGEMA_signal_7357), .Q (new_AGEMA_signal_7358) ) ;
    buf_clk new_AGEMA_reg_buffer_4584 ( .C (clk), .D (new_AGEMA_signal_7359), .Q (new_AGEMA_signal_7360) ) ;
    buf_clk new_AGEMA_reg_buffer_4586 ( .C (clk), .D (new_AGEMA_signal_7361), .Q (new_AGEMA_signal_7362) ) ;
    buf_clk new_AGEMA_reg_buffer_4588 ( .C (clk), .D (new_AGEMA_signal_7363), .Q (new_AGEMA_signal_7364) ) ;
    buf_clk new_AGEMA_reg_buffer_4590 ( .C (clk), .D (new_AGEMA_signal_7365), .Q (new_AGEMA_signal_7366) ) ;
    buf_clk new_AGEMA_reg_buffer_4592 ( .C (clk), .D (new_AGEMA_signal_7367), .Q (new_AGEMA_signal_7368) ) ;
    buf_clk new_AGEMA_reg_buffer_4594 ( .C (clk), .D (new_AGEMA_signal_7369), .Q (new_AGEMA_signal_7370) ) ;
    buf_clk new_AGEMA_reg_buffer_4596 ( .C (clk), .D (new_AGEMA_signal_7371), .Q (new_AGEMA_signal_7372) ) ;
    buf_clk new_AGEMA_reg_buffer_4598 ( .C (clk), .D (new_AGEMA_signal_7373), .Q (new_AGEMA_signal_7374) ) ;
    buf_clk new_AGEMA_reg_buffer_4600 ( .C (clk), .D (new_AGEMA_signal_7375), .Q (new_AGEMA_signal_7376) ) ;
    buf_clk new_AGEMA_reg_buffer_4602 ( .C (clk), .D (new_AGEMA_signal_7377), .Q (new_AGEMA_signal_7378) ) ;
    buf_clk new_AGEMA_reg_buffer_4604 ( .C (clk), .D (new_AGEMA_signal_7379), .Q (new_AGEMA_signal_7380) ) ;
    buf_clk new_AGEMA_reg_buffer_4606 ( .C (clk), .D (new_AGEMA_signal_7381), .Q (new_AGEMA_signal_7382) ) ;
    buf_clk new_AGEMA_reg_buffer_4608 ( .C (clk), .D (new_AGEMA_signal_7383), .Q (new_AGEMA_signal_7384) ) ;
    buf_clk new_AGEMA_reg_buffer_4610 ( .C (clk), .D (new_AGEMA_signal_7385), .Q (new_AGEMA_signal_7386) ) ;
    buf_clk new_AGEMA_reg_buffer_4612 ( .C (clk), .D (new_AGEMA_signal_7387), .Q (new_AGEMA_signal_7388) ) ;
    buf_clk new_AGEMA_reg_buffer_4614 ( .C (clk), .D (new_AGEMA_signal_7389), .Q (new_AGEMA_signal_7390) ) ;
    buf_clk new_AGEMA_reg_buffer_4616 ( .C (clk), .D (new_AGEMA_signal_7391), .Q (new_AGEMA_signal_7392) ) ;
    buf_clk new_AGEMA_reg_buffer_4618 ( .C (clk), .D (new_AGEMA_signal_7393), .Q (new_AGEMA_signal_7394) ) ;
    buf_clk new_AGEMA_reg_buffer_4620 ( .C (clk), .D (new_AGEMA_signal_7395), .Q (new_AGEMA_signal_7396) ) ;
    buf_clk new_AGEMA_reg_buffer_4622 ( .C (clk), .D (new_AGEMA_signal_7397), .Q (new_AGEMA_signal_7398) ) ;
    buf_clk new_AGEMA_reg_buffer_4624 ( .C (clk), .D (new_AGEMA_signal_7399), .Q (new_AGEMA_signal_7400) ) ;
    buf_clk new_AGEMA_reg_buffer_4626 ( .C (clk), .D (new_AGEMA_signal_7401), .Q (new_AGEMA_signal_7402) ) ;
    buf_clk new_AGEMA_reg_buffer_4628 ( .C (clk), .D (new_AGEMA_signal_7403), .Q (new_AGEMA_signal_7404) ) ;
    buf_clk new_AGEMA_reg_buffer_4630 ( .C (clk), .D (new_AGEMA_signal_7405), .Q (new_AGEMA_signal_7406) ) ;
    buf_clk new_AGEMA_reg_buffer_4632 ( .C (clk), .D (new_AGEMA_signal_7407), .Q (new_AGEMA_signal_7408) ) ;
    buf_clk new_AGEMA_reg_buffer_4634 ( .C (clk), .D (new_AGEMA_signal_7409), .Q (new_AGEMA_signal_7410) ) ;
    buf_clk new_AGEMA_reg_buffer_4636 ( .C (clk), .D (new_AGEMA_signal_7411), .Q (new_AGEMA_signal_7412) ) ;
    buf_clk new_AGEMA_reg_buffer_4638 ( .C (clk), .D (new_AGEMA_signal_7413), .Q (new_AGEMA_signal_7414) ) ;
    buf_clk new_AGEMA_reg_buffer_4640 ( .C (clk), .D (new_AGEMA_signal_7415), .Q (new_AGEMA_signal_7416) ) ;
    buf_clk new_AGEMA_reg_buffer_4642 ( .C (clk), .D (new_AGEMA_signal_7417), .Q (new_AGEMA_signal_7418) ) ;
    buf_clk new_AGEMA_reg_buffer_4644 ( .C (clk), .D (new_AGEMA_signal_7419), .Q (new_AGEMA_signal_7420) ) ;
    buf_clk new_AGEMA_reg_buffer_4646 ( .C (clk), .D (new_AGEMA_signal_7421), .Q (new_AGEMA_signal_7422) ) ;
    buf_clk new_AGEMA_reg_buffer_4648 ( .C (clk), .D (new_AGEMA_signal_7423), .Q (new_AGEMA_signal_7424) ) ;
    buf_clk new_AGEMA_reg_buffer_4650 ( .C (clk), .D (new_AGEMA_signal_7425), .Q (new_AGEMA_signal_7426) ) ;
    buf_clk new_AGEMA_reg_buffer_4652 ( .C (clk), .D (new_AGEMA_signal_7427), .Q (new_AGEMA_signal_7428) ) ;
    buf_clk new_AGEMA_reg_buffer_4654 ( .C (clk), .D (new_AGEMA_signal_7429), .Q (new_AGEMA_signal_7430) ) ;
    buf_clk new_AGEMA_reg_buffer_4656 ( .C (clk), .D (new_AGEMA_signal_7431), .Q (new_AGEMA_signal_7432) ) ;
    buf_clk new_AGEMA_reg_buffer_4658 ( .C (clk), .D (new_AGEMA_signal_7433), .Q (new_AGEMA_signal_7434) ) ;
    buf_clk new_AGEMA_reg_buffer_4660 ( .C (clk), .D (new_AGEMA_signal_7435), .Q (new_AGEMA_signal_7436) ) ;
    buf_clk new_AGEMA_reg_buffer_4662 ( .C (clk), .D (new_AGEMA_signal_7437), .Q (new_AGEMA_signal_7438) ) ;
    buf_clk new_AGEMA_reg_buffer_4664 ( .C (clk), .D (new_AGEMA_signal_7439), .Q (new_AGEMA_signal_7440) ) ;
    buf_clk new_AGEMA_reg_buffer_4666 ( .C (clk), .D (new_AGEMA_signal_7441), .Q (new_AGEMA_signal_7442) ) ;
    buf_clk new_AGEMA_reg_buffer_4674 ( .C (clk), .D (new_AGEMA_signal_7449), .Q (new_AGEMA_signal_7450) ) ;
    buf_clk new_AGEMA_reg_buffer_4682 ( .C (clk), .D (new_AGEMA_signal_7457), .Q (new_AGEMA_signal_7458) ) ;
    buf_clk new_AGEMA_reg_buffer_4690 ( .C (clk), .D (new_AGEMA_signal_7465), .Q (new_AGEMA_signal_7466) ) ;
    buf_clk new_AGEMA_reg_buffer_4698 ( .C (clk), .D (new_AGEMA_signal_7473), .Q (new_AGEMA_signal_7474) ) ;
    buf_clk new_AGEMA_reg_buffer_4706 ( .C (clk), .D (new_AGEMA_signal_7481), .Q (new_AGEMA_signal_7482) ) ;
    buf_clk new_AGEMA_reg_buffer_4714 ( .C (clk), .D (new_AGEMA_signal_7489), .Q (new_AGEMA_signal_7490) ) ;
    buf_clk new_AGEMA_reg_buffer_4722 ( .C (clk), .D (new_AGEMA_signal_7497), .Q (new_AGEMA_signal_7498) ) ;
    buf_clk new_AGEMA_reg_buffer_4730 ( .C (clk), .D (new_AGEMA_signal_7505), .Q (new_AGEMA_signal_7506) ) ;
    buf_clk new_AGEMA_reg_buffer_4738 ( .C (clk), .D (new_AGEMA_signal_7513), .Q (new_AGEMA_signal_7514) ) ;
    buf_clk new_AGEMA_reg_buffer_4746 ( .C (clk), .D (new_AGEMA_signal_7521), .Q (new_AGEMA_signal_7522) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_63__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7256, new_AGEMA_signal_7254, new_AGEMA_signal_7252}), .Q ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_62__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, AddRoundKeyOutput[62]}), .Q ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_61__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7262, new_AGEMA_signal_7260, new_AGEMA_signal_7258}), .Q ({ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_60__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2788, new_AGEMA_signal_2787, AddRoundKeyOutput[60]}), .Q ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_59__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7268, new_AGEMA_signal_7266, new_AGEMA_signal_7264}), .Q ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_58__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2784, new_AGEMA_signal_2783, AddRoundKeyOutput[58]}), .Q ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_57__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7274, new_AGEMA_signal_7272, new_AGEMA_signal_7270}), .Q ({ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_56__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, AddRoundKeyOutput[56]}), .Q ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_55__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7280, new_AGEMA_signal_7278, new_AGEMA_signal_7276}), .Q ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_54__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2776, new_AGEMA_signal_2775, AddRoundKeyOutput[54]}), .Q ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_53__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7286, new_AGEMA_signal_7284, new_AGEMA_signal_7282}), .Q ({ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_52__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2772, new_AGEMA_signal_2771, AddRoundKeyOutput[52]}), .Q ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_51__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7292, new_AGEMA_signal_7290, new_AGEMA_signal_7288}), .Q ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_50__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, AddRoundKeyOutput[50]}), .Q ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_49__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7298, new_AGEMA_signal_7296, new_AGEMA_signal_7294}), .Q ({ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_48__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2764, new_AGEMA_signal_2763, AddRoundKeyOutput[48]}), .Q ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_47__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7304, new_AGEMA_signal_7302, new_AGEMA_signal_7300}), .Q ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_46__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2808, new_AGEMA_signal_2807, AddRoundKeyOutput[46]}), .Q ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_45__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7310, new_AGEMA_signal_7308, new_AGEMA_signal_7306}), .Q ({ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_44__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2804, new_AGEMA_signal_2803, AddRoundKeyOutput[44]}), .Q ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_43__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7316, new_AGEMA_signal_7314, new_AGEMA_signal_7312}), .Q ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_42__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2800, new_AGEMA_signal_2799, AddRoundKeyOutput[42]}), .Q ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_41__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7322, new_AGEMA_signal_7320, new_AGEMA_signal_7318}), .Q ({ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_40__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2796, new_AGEMA_signal_2795, AddRoundKeyOutput[40]}), .Q ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_39__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7328, new_AGEMA_signal_7326, new_AGEMA_signal_7324}), .Q ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_38__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2824, new_AGEMA_signal_2823, AddRoundKeyOutput[38]}), .Q ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_37__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7334, new_AGEMA_signal_7332, new_AGEMA_signal_7330}), .Q ({ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_36__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2820, new_AGEMA_signal_2819, AddRoundKeyOutput[36]}), .Q ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_35__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7340, new_AGEMA_signal_7338, new_AGEMA_signal_7336}), .Q ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_34__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2816, new_AGEMA_signal_2815, AddRoundKeyOutput[34]}), .Q ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_33__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7346, new_AGEMA_signal_7344, new_AGEMA_signal_7342}), .Q ({ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_32__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2812, new_AGEMA_signal_2811, AddRoundKeyOutput[32]}), .Q ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_31__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7352, new_AGEMA_signal_7350, new_AGEMA_signal_7348}), .Q ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_30__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2696, new_AGEMA_signal_2695, AddRoundKeyOutput[30]}), .Q ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_29__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7358, new_AGEMA_signal_7356, new_AGEMA_signal_7354}), .Q ({ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_28__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, AddRoundKeyOutput[28]}), .Q ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_27__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7364, new_AGEMA_signal_7362, new_AGEMA_signal_7360}), .Q ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_26__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2688, new_AGEMA_signal_2687, AddRoundKeyOutput[26]}), .Q ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_25__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7370, new_AGEMA_signal_7368, new_AGEMA_signal_7366}), .Q ({ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_24__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2684, new_AGEMA_signal_2683, AddRoundKeyOutput[24]}), .Q ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_23__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7376, new_AGEMA_signal_7374, new_AGEMA_signal_7372}), .Q ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_22__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2680, new_AGEMA_signal_2679, AddRoundKeyOutput[22]}), .Q ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_21__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7382, new_AGEMA_signal_7380, new_AGEMA_signal_7378}), .Q ({ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_20__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, AddRoundKeyOutput[20]}), .Q ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_19__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7388, new_AGEMA_signal_7386, new_AGEMA_signal_7384}), .Q ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_18__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2672, new_AGEMA_signal_2671, AddRoundKeyOutput[18]}), .Q ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_17__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7394, new_AGEMA_signal_7392, new_AGEMA_signal_7390}), .Q ({ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_16__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2668, new_AGEMA_signal_2667, AddRoundKeyOutput[16]}), .Q ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_15__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7400, new_AGEMA_signal_7398, new_AGEMA_signal_7396}), .Q ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_14__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2664, new_AGEMA_signal_2663, AddRoundKeyOutput[14]}), .Q ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_13__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7406, new_AGEMA_signal_7404, new_AGEMA_signal_7402}), .Q ({ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_12__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2660, new_AGEMA_signal_2659, AddRoundKeyOutput[12]}), .Q ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_11__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7412, new_AGEMA_signal_7410, new_AGEMA_signal_7408}), .Q ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_10__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2656, new_AGEMA_signal_2655, AddRoundKeyOutput[10]}), .Q ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_9__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7418, new_AGEMA_signal_7416, new_AGEMA_signal_7414}), .Q ({ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_8__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2652, new_AGEMA_signal_2651, AddRoundKeyOutput[8]}), .Q ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_7__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7424, new_AGEMA_signal_7422, new_AGEMA_signal_7420}), .Q ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_6__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2648, new_AGEMA_signal_2647, AddRoundKeyOutput[6]}), .Q ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_5__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7430, new_AGEMA_signal_7428, new_AGEMA_signal_7426}), .Q ({ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_4__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2644, new_AGEMA_signal_2643, AddRoundKeyOutput[4]}), .Q ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7436, new_AGEMA_signal_7434, new_AGEMA_signal_7432}), .Q ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2640, new_AGEMA_signal_2639, AddRoundKeyOutput[2]}), .Q ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7442, new_AGEMA_signal_7440, new_AGEMA_signal_7438}), .Q ({ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, AddRoundKeyOutput[0]}), .Q ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_6__FF_FF ( .CK (clk), .D (new_AGEMA_signal_7450), .Q (FSMReg[6]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_5__FF_FF ( .CK (clk), .D (new_AGEMA_signal_7458), .Q (FSMReg[5]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_4__FF_FF ( .CK (clk), .D (new_AGEMA_signal_7466), .Q (FSMReg[4]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_3__FF_FF ( .CK (clk), .D (new_AGEMA_signal_7474), .Q (FSMReg[3]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_2__FF_FF ( .CK (clk), .D (new_AGEMA_signal_7482), .Q (FSMReg[2]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_1__FF_FF ( .CK (clk), .D (new_AGEMA_signal_7490), .Q (FSMReg[1]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_0__FF_FF ( .CK (clk), .D (new_AGEMA_signal_7498), .Q (FSMReg[0]), .QN () ) ;
    DFF_X1 selectsRegInst_s_current_state_reg_1__FF_FF ( .CK (clk), .D (new_AGEMA_signal_7506), .Q (selectsReg[1]), .QN () ) ;
    DFF_X1 selectsRegInst_s_current_state_reg_0__FF_FF ( .CK (clk), .D (new_AGEMA_signal_7514), .Q (selectsReg[0]), .QN () ) ;
    DFF_X1 done_reg_FF_FF ( .CK (clk), .D (new_AGEMA_signal_7522), .Q (done), .QN () ) ;
endmodule
