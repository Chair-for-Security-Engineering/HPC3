////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module SkinnyTop in file /AGEMA/Designs/Skinny64_64_round-based/AGEMA/SkinnyTop.v */
/* clock gating is added to the circuit, the latency increased 4 time(s)  */

module SkinnyTop_HPC2_ClockGating_d1 (Plaintext_s0, Key_s0, clk, rst, Key_s1, Plaintext_s1, Fresh, Ciphertext_s0, done, Ciphertext_s1, Synch);
    input [63:0] Plaintext_s0 ;
    input [63:0] Key_s0 ;
    input clk ;
    input rst ;
    input [63:0] Key_s1 ;
    input [63:0] Plaintext_s1 ;
    input [63:0] Fresh ;
    output [63:0] Ciphertext_s0 ;
    output done ;
    output [63:0] Ciphertext_s1 ;
    output Synch ;
    wire SubCellInst_SboxInst_0_n3 ;
    wire SubCellInst_SboxInst_0_YY_0_ ;
    wire SubCellInst_SboxInst_0_YY_1_ ;
    wire SubCellInst_SboxInst_0_L3 ;
    wire SubCellInst_SboxInst_0_YY_3 ;
    wire SubCellInst_SboxInst_0_L2 ;
    wire SubCellInst_SboxInst_0_T3 ;
    wire SubCellInst_SboxInst_0_Q7 ;
    wire SubCellInst_SboxInst_0_L1 ;
    wire SubCellInst_SboxInst_0_Q6 ;
    wire SubCellInst_SboxInst_0_L0 ;
    wire SubCellInst_SboxInst_0_T2 ;
    wire SubCellInst_SboxInst_0_Q4 ;
    wire SubCellInst_SboxInst_0_T1 ;
    wire SubCellInst_SboxInst_0_Q2 ;
    wire SubCellInst_SboxInst_0_T0 ;
    wire SubCellInst_SboxInst_0_Q1 ;
    wire SubCellInst_SboxInst_0_Q0 ;
    wire SubCellInst_SboxInst_0_XX_1_ ;
    wire SubCellInst_SboxInst_0_XX_2_ ;
    wire SubCellInst_SboxInst_1_n3 ;
    wire SubCellInst_SboxInst_1_YY_0_ ;
    wire SubCellInst_SboxInst_1_YY_1_ ;
    wire SubCellInst_SboxInst_1_L3 ;
    wire SubCellInst_SboxInst_1_YY_3 ;
    wire SubCellInst_SboxInst_1_L2 ;
    wire SubCellInst_SboxInst_1_T3 ;
    wire SubCellInst_SboxInst_1_Q7 ;
    wire SubCellInst_SboxInst_1_L1 ;
    wire SubCellInst_SboxInst_1_Q6 ;
    wire SubCellInst_SboxInst_1_L0 ;
    wire SubCellInst_SboxInst_1_T2 ;
    wire SubCellInst_SboxInst_1_Q4 ;
    wire SubCellInst_SboxInst_1_T1 ;
    wire SubCellInst_SboxInst_1_Q2 ;
    wire SubCellInst_SboxInst_1_T0 ;
    wire SubCellInst_SboxInst_1_Q1 ;
    wire SubCellInst_SboxInst_1_Q0 ;
    wire SubCellInst_SboxInst_1_XX_1_ ;
    wire SubCellInst_SboxInst_1_XX_2_ ;
    wire SubCellInst_SboxInst_2_n3 ;
    wire SubCellInst_SboxInst_2_YY_0_ ;
    wire SubCellInst_SboxInst_2_YY_1_ ;
    wire SubCellInst_SboxInst_2_L3 ;
    wire SubCellInst_SboxInst_2_YY_3 ;
    wire SubCellInst_SboxInst_2_L2 ;
    wire SubCellInst_SboxInst_2_T3 ;
    wire SubCellInst_SboxInst_2_Q7 ;
    wire SubCellInst_SboxInst_2_L1 ;
    wire SubCellInst_SboxInst_2_Q6 ;
    wire SubCellInst_SboxInst_2_L0 ;
    wire SubCellInst_SboxInst_2_T2 ;
    wire SubCellInst_SboxInst_2_Q4 ;
    wire SubCellInst_SboxInst_2_T1 ;
    wire SubCellInst_SboxInst_2_Q2 ;
    wire SubCellInst_SboxInst_2_T0 ;
    wire SubCellInst_SboxInst_2_Q1 ;
    wire SubCellInst_SboxInst_2_Q0 ;
    wire SubCellInst_SboxInst_2_XX_1_ ;
    wire SubCellInst_SboxInst_2_XX_2_ ;
    wire SubCellInst_SboxInst_3_n3 ;
    wire SubCellInst_SboxInst_3_YY_0_ ;
    wire SubCellInst_SboxInst_3_YY_1_ ;
    wire SubCellInst_SboxInst_3_L3 ;
    wire SubCellInst_SboxInst_3_YY_3 ;
    wire SubCellInst_SboxInst_3_L2 ;
    wire SubCellInst_SboxInst_3_T3 ;
    wire SubCellInst_SboxInst_3_Q7 ;
    wire SubCellInst_SboxInst_3_L1 ;
    wire SubCellInst_SboxInst_3_Q6 ;
    wire SubCellInst_SboxInst_3_L0 ;
    wire SubCellInst_SboxInst_3_T2 ;
    wire SubCellInst_SboxInst_3_Q4 ;
    wire SubCellInst_SboxInst_3_T1 ;
    wire SubCellInst_SboxInst_3_Q2 ;
    wire SubCellInst_SboxInst_3_T0 ;
    wire SubCellInst_SboxInst_3_Q1 ;
    wire SubCellInst_SboxInst_3_Q0 ;
    wire SubCellInst_SboxInst_3_XX_1_ ;
    wire SubCellInst_SboxInst_3_XX_2_ ;
    wire SubCellInst_SboxInst_4_n3 ;
    wire SubCellInst_SboxInst_4_YY_0_ ;
    wire SubCellInst_SboxInst_4_YY_1_ ;
    wire SubCellInst_SboxInst_4_L3 ;
    wire SubCellInst_SboxInst_4_YY_3 ;
    wire SubCellInst_SboxInst_4_L2 ;
    wire SubCellInst_SboxInst_4_T3 ;
    wire SubCellInst_SboxInst_4_Q7 ;
    wire SubCellInst_SboxInst_4_L1 ;
    wire SubCellInst_SboxInst_4_Q6 ;
    wire SubCellInst_SboxInst_4_L0 ;
    wire SubCellInst_SboxInst_4_T2 ;
    wire SubCellInst_SboxInst_4_Q4 ;
    wire SubCellInst_SboxInst_4_T1 ;
    wire SubCellInst_SboxInst_4_Q2 ;
    wire SubCellInst_SboxInst_4_T0 ;
    wire SubCellInst_SboxInst_4_Q1 ;
    wire SubCellInst_SboxInst_4_Q0 ;
    wire SubCellInst_SboxInst_4_XX_1_ ;
    wire SubCellInst_SboxInst_4_XX_2_ ;
    wire SubCellInst_SboxInst_5_n3 ;
    wire SubCellInst_SboxInst_5_YY_0_ ;
    wire SubCellInst_SboxInst_5_YY_1_ ;
    wire SubCellInst_SboxInst_5_L3 ;
    wire SubCellInst_SboxInst_5_YY_3 ;
    wire SubCellInst_SboxInst_5_L2 ;
    wire SubCellInst_SboxInst_5_T3 ;
    wire SubCellInst_SboxInst_5_Q7 ;
    wire SubCellInst_SboxInst_5_L1 ;
    wire SubCellInst_SboxInst_5_Q6 ;
    wire SubCellInst_SboxInst_5_L0 ;
    wire SubCellInst_SboxInst_5_T2 ;
    wire SubCellInst_SboxInst_5_Q4 ;
    wire SubCellInst_SboxInst_5_T1 ;
    wire SubCellInst_SboxInst_5_Q2 ;
    wire SubCellInst_SboxInst_5_T0 ;
    wire SubCellInst_SboxInst_5_Q1 ;
    wire SubCellInst_SboxInst_5_Q0 ;
    wire SubCellInst_SboxInst_5_XX_1_ ;
    wire SubCellInst_SboxInst_5_XX_2_ ;
    wire SubCellInst_SboxInst_6_n3 ;
    wire SubCellInst_SboxInst_6_YY_0_ ;
    wire SubCellInst_SboxInst_6_YY_1_ ;
    wire SubCellInst_SboxInst_6_L3 ;
    wire SubCellInst_SboxInst_6_YY_3 ;
    wire SubCellInst_SboxInst_6_L2 ;
    wire SubCellInst_SboxInst_6_T3 ;
    wire SubCellInst_SboxInst_6_Q7 ;
    wire SubCellInst_SboxInst_6_L1 ;
    wire SubCellInst_SboxInst_6_Q6 ;
    wire SubCellInst_SboxInst_6_L0 ;
    wire SubCellInst_SboxInst_6_T2 ;
    wire SubCellInst_SboxInst_6_Q4 ;
    wire SubCellInst_SboxInst_6_T1 ;
    wire SubCellInst_SboxInst_6_Q2 ;
    wire SubCellInst_SboxInst_6_T0 ;
    wire SubCellInst_SboxInst_6_Q1 ;
    wire SubCellInst_SboxInst_6_Q0 ;
    wire SubCellInst_SboxInst_6_XX_1_ ;
    wire SubCellInst_SboxInst_6_XX_2_ ;
    wire SubCellInst_SboxInst_7_n3 ;
    wire SubCellInst_SboxInst_7_YY_0_ ;
    wire SubCellInst_SboxInst_7_YY_1_ ;
    wire SubCellInst_SboxInst_7_L3 ;
    wire SubCellInst_SboxInst_7_YY_3 ;
    wire SubCellInst_SboxInst_7_L2 ;
    wire SubCellInst_SboxInst_7_T3 ;
    wire SubCellInst_SboxInst_7_Q7 ;
    wire SubCellInst_SboxInst_7_L1 ;
    wire SubCellInst_SboxInst_7_Q6 ;
    wire SubCellInst_SboxInst_7_L0 ;
    wire SubCellInst_SboxInst_7_T2 ;
    wire SubCellInst_SboxInst_7_Q4 ;
    wire SubCellInst_SboxInst_7_T1 ;
    wire SubCellInst_SboxInst_7_Q2 ;
    wire SubCellInst_SboxInst_7_T0 ;
    wire SubCellInst_SboxInst_7_Q1 ;
    wire SubCellInst_SboxInst_7_Q0 ;
    wire SubCellInst_SboxInst_7_XX_1_ ;
    wire SubCellInst_SboxInst_7_XX_2_ ;
    wire SubCellInst_SboxInst_8_n3 ;
    wire SubCellInst_SboxInst_8_YY_0_ ;
    wire SubCellInst_SboxInst_8_YY_1_ ;
    wire SubCellInst_SboxInst_8_L3 ;
    wire SubCellInst_SboxInst_8_YY_3 ;
    wire SubCellInst_SboxInst_8_L2 ;
    wire SubCellInst_SboxInst_8_T3 ;
    wire SubCellInst_SboxInst_8_Q7 ;
    wire SubCellInst_SboxInst_8_L1 ;
    wire SubCellInst_SboxInst_8_Q6 ;
    wire SubCellInst_SboxInst_8_L0 ;
    wire SubCellInst_SboxInst_8_T2 ;
    wire SubCellInst_SboxInst_8_Q4 ;
    wire SubCellInst_SboxInst_8_T1 ;
    wire SubCellInst_SboxInst_8_Q2 ;
    wire SubCellInst_SboxInst_8_T0 ;
    wire SubCellInst_SboxInst_8_Q1 ;
    wire SubCellInst_SboxInst_8_Q0 ;
    wire SubCellInst_SboxInst_8_XX_1_ ;
    wire SubCellInst_SboxInst_8_XX_2_ ;
    wire SubCellInst_SboxInst_9_n3 ;
    wire SubCellInst_SboxInst_9_YY_0_ ;
    wire SubCellInst_SboxInst_9_YY_1_ ;
    wire SubCellInst_SboxInst_9_L3 ;
    wire SubCellInst_SboxInst_9_YY_3 ;
    wire SubCellInst_SboxInst_9_L2 ;
    wire SubCellInst_SboxInst_9_T3 ;
    wire SubCellInst_SboxInst_9_Q7 ;
    wire SubCellInst_SboxInst_9_L1 ;
    wire SubCellInst_SboxInst_9_Q6 ;
    wire SubCellInst_SboxInst_9_L0 ;
    wire SubCellInst_SboxInst_9_T2 ;
    wire SubCellInst_SboxInst_9_Q4 ;
    wire SubCellInst_SboxInst_9_T1 ;
    wire SubCellInst_SboxInst_9_Q2 ;
    wire SubCellInst_SboxInst_9_T0 ;
    wire SubCellInst_SboxInst_9_Q1 ;
    wire SubCellInst_SboxInst_9_Q0 ;
    wire SubCellInst_SboxInst_9_XX_1_ ;
    wire SubCellInst_SboxInst_9_XX_2_ ;
    wire SubCellInst_SboxInst_10_n3 ;
    wire SubCellInst_SboxInst_10_YY_0_ ;
    wire SubCellInst_SboxInst_10_YY_1_ ;
    wire SubCellInst_SboxInst_10_L3 ;
    wire SubCellInst_SboxInst_10_YY_3 ;
    wire SubCellInst_SboxInst_10_L2 ;
    wire SubCellInst_SboxInst_10_T3 ;
    wire SubCellInst_SboxInst_10_Q7 ;
    wire SubCellInst_SboxInst_10_L1 ;
    wire SubCellInst_SboxInst_10_Q6 ;
    wire SubCellInst_SboxInst_10_L0 ;
    wire SubCellInst_SboxInst_10_T2 ;
    wire SubCellInst_SboxInst_10_Q4 ;
    wire SubCellInst_SboxInst_10_T1 ;
    wire SubCellInst_SboxInst_10_Q2 ;
    wire SubCellInst_SboxInst_10_T0 ;
    wire SubCellInst_SboxInst_10_Q1 ;
    wire SubCellInst_SboxInst_10_Q0 ;
    wire SubCellInst_SboxInst_10_XX_1_ ;
    wire SubCellInst_SboxInst_10_XX_2_ ;
    wire SubCellInst_SboxInst_11_n3 ;
    wire SubCellInst_SboxInst_11_YY_0_ ;
    wire SubCellInst_SboxInst_11_YY_1_ ;
    wire SubCellInst_SboxInst_11_L3 ;
    wire SubCellInst_SboxInst_11_YY_3 ;
    wire SubCellInst_SboxInst_11_L2 ;
    wire SubCellInst_SboxInst_11_T3 ;
    wire SubCellInst_SboxInst_11_Q7 ;
    wire SubCellInst_SboxInst_11_L1 ;
    wire SubCellInst_SboxInst_11_Q6 ;
    wire SubCellInst_SboxInst_11_L0 ;
    wire SubCellInst_SboxInst_11_T2 ;
    wire SubCellInst_SboxInst_11_Q4 ;
    wire SubCellInst_SboxInst_11_T1 ;
    wire SubCellInst_SboxInst_11_Q2 ;
    wire SubCellInst_SboxInst_11_T0 ;
    wire SubCellInst_SboxInst_11_Q1 ;
    wire SubCellInst_SboxInst_11_Q0 ;
    wire SubCellInst_SboxInst_11_XX_1_ ;
    wire SubCellInst_SboxInst_11_XX_2_ ;
    wire SubCellInst_SboxInst_12_n3 ;
    wire SubCellInst_SboxInst_12_YY_0_ ;
    wire SubCellInst_SboxInst_12_YY_1_ ;
    wire SubCellInst_SboxInst_12_L3 ;
    wire SubCellInst_SboxInst_12_YY_3 ;
    wire SubCellInst_SboxInst_12_L2 ;
    wire SubCellInst_SboxInst_12_T3 ;
    wire SubCellInst_SboxInst_12_Q7 ;
    wire SubCellInst_SboxInst_12_L1 ;
    wire SubCellInst_SboxInst_12_Q6 ;
    wire SubCellInst_SboxInst_12_L0 ;
    wire SubCellInst_SboxInst_12_T2 ;
    wire SubCellInst_SboxInst_12_Q4 ;
    wire SubCellInst_SboxInst_12_T1 ;
    wire SubCellInst_SboxInst_12_Q2 ;
    wire SubCellInst_SboxInst_12_T0 ;
    wire SubCellInst_SboxInst_12_Q1 ;
    wire SubCellInst_SboxInst_12_Q0 ;
    wire SubCellInst_SboxInst_12_XX_1_ ;
    wire SubCellInst_SboxInst_12_XX_2_ ;
    wire SubCellInst_SboxInst_13_n3 ;
    wire SubCellInst_SboxInst_13_YY_0_ ;
    wire SubCellInst_SboxInst_13_YY_1_ ;
    wire SubCellInst_SboxInst_13_L3 ;
    wire SubCellInst_SboxInst_13_YY_3 ;
    wire SubCellInst_SboxInst_13_L2 ;
    wire SubCellInst_SboxInst_13_T3 ;
    wire SubCellInst_SboxInst_13_Q7 ;
    wire SubCellInst_SboxInst_13_L1 ;
    wire SubCellInst_SboxInst_13_Q6 ;
    wire SubCellInst_SboxInst_13_L0 ;
    wire SubCellInst_SboxInst_13_T2 ;
    wire SubCellInst_SboxInst_13_Q4 ;
    wire SubCellInst_SboxInst_13_T1 ;
    wire SubCellInst_SboxInst_13_Q2 ;
    wire SubCellInst_SboxInst_13_T0 ;
    wire SubCellInst_SboxInst_13_Q1 ;
    wire SubCellInst_SboxInst_13_Q0 ;
    wire SubCellInst_SboxInst_13_XX_1_ ;
    wire SubCellInst_SboxInst_13_XX_2_ ;
    wire SubCellInst_SboxInst_14_n3 ;
    wire SubCellInst_SboxInst_14_YY_0_ ;
    wire SubCellInst_SboxInst_14_YY_1_ ;
    wire SubCellInst_SboxInst_14_L3 ;
    wire SubCellInst_SboxInst_14_YY_3 ;
    wire SubCellInst_SboxInst_14_L2 ;
    wire SubCellInst_SboxInst_14_T3 ;
    wire SubCellInst_SboxInst_14_Q7 ;
    wire SubCellInst_SboxInst_14_L1 ;
    wire SubCellInst_SboxInst_14_Q6 ;
    wire SubCellInst_SboxInst_14_L0 ;
    wire SubCellInst_SboxInst_14_T2 ;
    wire SubCellInst_SboxInst_14_Q4 ;
    wire SubCellInst_SboxInst_14_T1 ;
    wire SubCellInst_SboxInst_14_Q2 ;
    wire SubCellInst_SboxInst_14_T0 ;
    wire SubCellInst_SboxInst_14_Q1 ;
    wire SubCellInst_SboxInst_14_Q0 ;
    wire SubCellInst_SboxInst_14_XX_1_ ;
    wire SubCellInst_SboxInst_14_XX_2_ ;
    wire SubCellInst_SboxInst_15_n3 ;
    wire SubCellInst_SboxInst_15_YY_0_ ;
    wire SubCellInst_SboxInst_15_YY_1_ ;
    wire SubCellInst_SboxInst_15_L3 ;
    wire SubCellInst_SboxInst_15_YY_3 ;
    wire SubCellInst_SboxInst_15_L2 ;
    wire SubCellInst_SboxInst_15_T3 ;
    wire SubCellInst_SboxInst_15_Q7 ;
    wire SubCellInst_SboxInst_15_L1 ;
    wire SubCellInst_SboxInst_15_Q6 ;
    wire SubCellInst_SboxInst_15_L0 ;
    wire SubCellInst_SboxInst_15_T2 ;
    wire SubCellInst_SboxInst_15_Q4 ;
    wire SubCellInst_SboxInst_15_T1 ;
    wire SubCellInst_SboxInst_15_Q2 ;
    wire SubCellInst_SboxInst_15_T0 ;
    wire SubCellInst_SboxInst_15_Q1 ;
    wire SubCellInst_SboxInst_15_Q0 ;
    wire SubCellInst_SboxInst_15_XX_1_ ;
    wire SubCellInst_SboxInst_15_XX_2_ ;
    wire AddConstXOR_AddConstXOR_XORInst_0_0_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_0_1_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_0_2_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_0_3_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_0_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_1_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_2_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_3_n1 ;
    wire MCInst_MCR0_XORInst_0_0_n2 ;
    wire MCInst_MCR0_XORInst_0_0_n1 ;
    wire MCInst_MCR0_XORInst_0_1_n2 ;
    wire MCInst_MCR0_XORInst_0_1_n1 ;
    wire MCInst_MCR0_XORInst_0_2_n2 ;
    wire MCInst_MCR0_XORInst_0_2_n1 ;
    wire MCInst_MCR0_XORInst_0_3_n2 ;
    wire MCInst_MCR0_XORInst_0_3_n1 ;
    wire MCInst_MCR0_XORInst_1_0_n2 ;
    wire MCInst_MCR0_XORInst_1_0_n1 ;
    wire MCInst_MCR0_XORInst_1_1_n2 ;
    wire MCInst_MCR0_XORInst_1_1_n1 ;
    wire MCInst_MCR0_XORInst_1_2_n2 ;
    wire MCInst_MCR0_XORInst_1_2_n1 ;
    wire MCInst_MCR0_XORInst_1_3_n2 ;
    wire MCInst_MCR0_XORInst_1_3_n1 ;
    wire MCInst_MCR0_XORInst_2_0_n2 ;
    wire MCInst_MCR0_XORInst_2_0_n1 ;
    wire MCInst_MCR0_XORInst_2_1_n2 ;
    wire MCInst_MCR0_XORInst_2_1_n1 ;
    wire MCInst_MCR0_XORInst_2_2_n2 ;
    wire MCInst_MCR0_XORInst_2_2_n1 ;
    wire MCInst_MCR0_XORInst_2_3_n2 ;
    wire MCInst_MCR0_XORInst_2_3_n1 ;
    wire MCInst_MCR0_XORInst_3_0_n2 ;
    wire MCInst_MCR0_XORInst_3_0_n1 ;
    wire MCInst_MCR0_XORInst_3_1_n2 ;
    wire MCInst_MCR0_XORInst_3_1_n1 ;
    wire MCInst_MCR0_XORInst_3_2_n2 ;
    wire MCInst_MCR0_XORInst_3_2_n1 ;
    wire MCInst_MCR0_XORInst_3_3_n2 ;
    wire MCInst_MCR0_XORInst_3_3_n1 ;
    wire MCInst_MCR2_XORInst_0_0_n1 ;
    wire MCInst_MCR2_XORInst_0_1_n1 ;
    wire MCInst_MCR2_XORInst_0_2_n1 ;
    wire MCInst_MCR2_XORInst_0_3_n1 ;
    wire MCInst_MCR2_XORInst_1_0_n1 ;
    wire MCInst_MCR2_XORInst_1_1_n1 ;
    wire MCInst_MCR2_XORInst_1_2_n1 ;
    wire MCInst_MCR2_XORInst_1_3_n1 ;
    wire MCInst_MCR2_XORInst_2_0_n1 ;
    wire MCInst_MCR2_XORInst_2_1_n1 ;
    wire MCInst_MCR2_XORInst_2_2_n1 ;
    wire MCInst_MCR2_XORInst_2_3_n1 ;
    wire MCInst_MCR2_XORInst_3_0_n1 ;
    wire MCInst_MCR2_XORInst_3_1_n1 ;
    wire MCInst_MCR2_XORInst_3_2_n1 ;
    wire MCInst_MCR2_XORInst_3_3_n1 ;
    wire MCInst_MCR3_XORInst_0_0_n1 ;
    wire MCInst_MCR3_XORInst_0_1_n1 ;
    wire MCInst_MCR3_XORInst_0_2_n1 ;
    wire MCInst_MCR3_XORInst_0_3_n1 ;
    wire MCInst_MCR3_XORInst_1_0_n1 ;
    wire MCInst_MCR3_XORInst_1_1_n1 ;
    wire MCInst_MCR3_XORInst_1_2_n1 ;
    wire MCInst_MCR3_XORInst_1_3_n1 ;
    wire MCInst_MCR3_XORInst_2_0_n1 ;
    wire MCInst_MCR3_XORInst_2_1_n1 ;
    wire MCInst_MCR3_XORInst_2_2_n1 ;
    wire MCInst_MCR3_XORInst_2_3_n1 ;
    wire MCInst_MCR3_XORInst_3_0_n1 ;
    wire MCInst_MCR3_XORInst_3_1_n1 ;
    wire MCInst_MCR3_XORInst_3_2_n1 ;
    wire MCInst_MCR3_XORInst_3_3_n1 ;
    wire FSMUpdateInst_StateUpdateInst_0_n4 ;
    wire FSMUpdateInst_StateUpdateInst_0_n3 ;
    wire FSMUpdateInst_StateUpdateInst_0_n2 ;
    wire FSMUpdateInst_StateUpdateInst_0_n1 ;
    wire FSMUpdateInst_StateUpdateInst_2_n4 ;
    wire FSMUpdateInst_StateUpdateInst_2_n3 ;
    wire FSMUpdateInst_StateUpdateInst_2_n2 ;
    wire FSMUpdateInst_StateUpdateInst_2_n1 ;
    wire FSMUpdateInst_StateUpdateInst_5_n4 ;
    wire FSMUpdateInst_StateUpdateInst_5_n3 ;
    wire FSMUpdateInst_StateUpdateInst_5_n2 ;
    wire FSMUpdateInst_StateUpdateInst_5_n1 ;
    wire FSMSignalsInst_doneInst_n5 ;
    wire FSMSignalsInst_doneInst_n4 ;
    wire FSMSignalsInst_doneInst_n3 ;
    wire FSMSignalsInst_doneInst_n2 ;
    wire FSMSignalsInst_doneInst_n1 ;
    wire [63:0] MCOutput ;
    wire [63:0] StateRegInput ;
    wire [63:29] SubCellOutput ;
    wire [5:1] FSM ;
    wire [63:32] AddRoundConstantOutput ;
    wire [47:0] ShiftRowsOutput ;
    wire [5:0] FSMUpdate ;
    wire [5:0] FSMSelected ;
    wire [63:0] TweakeyGeneration_StateRegInput ;
    wire [63:0] TweakeyGeneration_key_Feedback ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2124 ;
    wire clk_gated ;

    /* cells in depth 0 */
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_U1 ( .a ({Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({new_AGEMA_signal_1165, SubCellInst_SboxInst_0_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_XOR_i1_U1 ( .a ({Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({Ciphertext_s1[3], Ciphertext_s0[3]}), .c ({new_AGEMA_signal_1167, SubCellInst_SboxInst_0_XX_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_XOR_i2_U1 ( .a ({Ciphertext_s1[0], Ciphertext_s0[0]}), .b ({Ciphertext_s1[2], Ciphertext_s0[2]}), .c ({new_AGEMA_signal_1169, SubCellInst_SboxInst_0_XX_2_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_XOR0_U1 ( .a ({Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1169, SubCellInst_SboxInst_0_XX_2_}), .c ({new_AGEMA_signal_1453, SubCellInst_SboxInst_0_Q0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_XOR1_U1 ( .a ({Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1167, SubCellInst_SboxInst_0_XX_1_}), .c ({new_AGEMA_signal_1454, SubCellInst_SboxInst_0_Q1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_XOR3_U1 ( .a ({Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1165, SubCellInst_SboxInst_0_n3}), .c ({new_AGEMA_signal_1455, SubCellInst_SboxInst_0_Q4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_XOR5_U1 ( .a ({new_AGEMA_signal_1169, SubCellInst_SboxInst_0_XX_2_}), .b ({new_AGEMA_signal_1165, SubCellInst_SboxInst_0_n3}), .c ({new_AGEMA_signal_1456, SubCellInst_SboxInst_0_Q6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_XOR6_U1 ( .a ({new_AGEMA_signal_1454, SubCellInst_SboxInst_0_Q1}), .b ({new_AGEMA_signal_1456, SubCellInst_SboxInst_0_Q6}), .c ({new_AGEMA_signal_1550, SubCellInst_SboxInst_0_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_XOR8_U1 ( .a ({Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1165, SubCellInst_SboxInst_0_n3}), .c ({new_AGEMA_signal_1457, SubCellInst_SboxInst_0_L2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_U1 ( .a ({Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({new_AGEMA_signal_1171, SubCellInst_SboxInst_1_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_XOR_i1_U1 ( .a ({Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({Ciphertext_s1[7], Ciphertext_s0[7]}), .c ({new_AGEMA_signal_1173, SubCellInst_SboxInst_1_XX_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_XOR_i2_U1 ( .a ({Ciphertext_s1[4], Ciphertext_s0[4]}), .b ({Ciphertext_s1[6], Ciphertext_s0[6]}), .c ({new_AGEMA_signal_1175, SubCellInst_SboxInst_1_XX_2_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_XOR0_U1 ( .a ({Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1175, SubCellInst_SboxInst_1_XX_2_}), .c ({new_AGEMA_signal_1459, SubCellInst_SboxInst_1_Q0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_XOR1_U1 ( .a ({Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1173, SubCellInst_SboxInst_1_XX_1_}), .c ({new_AGEMA_signal_1460, SubCellInst_SboxInst_1_Q1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_XOR3_U1 ( .a ({Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1171, SubCellInst_SboxInst_1_n3}), .c ({new_AGEMA_signal_1461, SubCellInst_SboxInst_1_Q4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_XOR5_U1 ( .a ({new_AGEMA_signal_1175, SubCellInst_SboxInst_1_XX_2_}), .b ({new_AGEMA_signal_1171, SubCellInst_SboxInst_1_n3}), .c ({new_AGEMA_signal_1462, SubCellInst_SboxInst_1_Q6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_XOR6_U1 ( .a ({new_AGEMA_signal_1460, SubCellInst_SboxInst_1_Q1}), .b ({new_AGEMA_signal_1462, SubCellInst_SboxInst_1_Q6}), .c ({new_AGEMA_signal_1553, SubCellInst_SboxInst_1_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_XOR8_U1 ( .a ({Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1171, SubCellInst_SboxInst_1_n3}), .c ({new_AGEMA_signal_1463, SubCellInst_SboxInst_1_L2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_U1 ( .a ({Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({new_AGEMA_signal_1177, SubCellInst_SboxInst_2_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_XOR_i1_U1 ( .a ({Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({Ciphertext_s1[11], Ciphertext_s0[11]}), .c ({new_AGEMA_signal_1179, SubCellInst_SboxInst_2_XX_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_XOR_i2_U1 ( .a ({Ciphertext_s1[8], Ciphertext_s0[8]}), .b ({Ciphertext_s1[10], Ciphertext_s0[10]}), .c ({new_AGEMA_signal_1181, SubCellInst_SboxInst_2_XX_2_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_XOR0_U1 ( .a ({Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1181, SubCellInst_SboxInst_2_XX_2_}), .c ({new_AGEMA_signal_1465, SubCellInst_SboxInst_2_Q0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_XOR1_U1 ( .a ({Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1179, SubCellInst_SboxInst_2_XX_1_}), .c ({new_AGEMA_signal_1466, SubCellInst_SboxInst_2_Q1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_XOR3_U1 ( .a ({Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1177, SubCellInst_SboxInst_2_n3}), .c ({new_AGEMA_signal_1467, SubCellInst_SboxInst_2_Q4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_XOR5_U1 ( .a ({new_AGEMA_signal_1181, SubCellInst_SboxInst_2_XX_2_}), .b ({new_AGEMA_signal_1177, SubCellInst_SboxInst_2_n3}), .c ({new_AGEMA_signal_1468, SubCellInst_SboxInst_2_Q6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_XOR6_U1 ( .a ({new_AGEMA_signal_1466, SubCellInst_SboxInst_2_Q1}), .b ({new_AGEMA_signal_1468, SubCellInst_SboxInst_2_Q6}), .c ({new_AGEMA_signal_1556, SubCellInst_SboxInst_2_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_XOR8_U1 ( .a ({Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1177, SubCellInst_SboxInst_2_n3}), .c ({new_AGEMA_signal_1469, SubCellInst_SboxInst_2_L2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_U1 ( .a ({Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({new_AGEMA_signal_1183, SubCellInst_SboxInst_3_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_XOR_i1_U1 ( .a ({Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({Ciphertext_s1[15], Ciphertext_s0[15]}), .c ({new_AGEMA_signal_1185, SubCellInst_SboxInst_3_XX_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_XOR_i2_U1 ( .a ({Ciphertext_s1[12], Ciphertext_s0[12]}), .b ({Ciphertext_s1[14], Ciphertext_s0[14]}), .c ({new_AGEMA_signal_1187, SubCellInst_SboxInst_3_XX_2_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_XOR0_U1 ( .a ({Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1187, SubCellInst_SboxInst_3_XX_2_}), .c ({new_AGEMA_signal_1471, SubCellInst_SboxInst_3_Q0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_XOR1_U1 ( .a ({Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1185, SubCellInst_SboxInst_3_XX_1_}), .c ({new_AGEMA_signal_1472, SubCellInst_SboxInst_3_Q1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_XOR3_U1 ( .a ({Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1183, SubCellInst_SboxInst_3_n3}), .c ({new_AGEMA_signal_1473, SubCellInst_SboxInst_3_Q4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_XOR5_U1 ( .a ({new_AGEMA_signal_1187, SubCellInst_SboxInst_3_XX_2_}), .b ({new_AGEMA_signal_1183, SubCellInst_SboxInst_3_n3}), .c ({new_AGEMA_signal_1474, SubCellInst_SboxInst_3_Q6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_XOR6_U1 ( .a ({new_AGEMA_signal_1472, SubCellInst_SboxInst_3_Q1}), .b ({new_AGEMA_signal_1474, SubCellInst_SboxInst_3_Q6}), .c ({new_AGEMA_signal_1559, SubCellInst_SboxInst_3_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_XOR8_U1 ( .a ({Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1183, SubCellInst_SboxInst_3_n3}), .c ({new_AGEMA_signal_1475, SubCellInst_SboxInst_3_L2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_U1 ( .a ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({new_AGEMA_signal_1189, SubCellInst_SboxInst_4_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_XOR_i1_U1 ( .a ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({Ciphertext_s1[19], Ciphertext_s0[19]}), .c ({new_AGEMA_signal_1191, SubCellInst_SboxInst_4_XX_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_XOR_i2_U1 ( .a ({Ciphertext_s1[16], Ciphertext_s0[16]}), .b ({Ciphertext_s1[18], Ciphertext_s0[18]}), .c ({new_AGEMA_signal_1193, SubCellInst_SboxInst_4_XX_2_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_XOR0_U1 ( .a ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1193, SubCellInst_SboxInst_4_XX_2_}), .c ({new_AGEMA_signal_1477, SubCellInst_SboxInst_4_Q0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_XOR1_U1 ( .a ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1191, SubCellInst_SboxInst_4_XX_1_}), .c ({new_AGEMA_signal_1478, SubCellInst_SboxInst_4_Q1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_XOR3_U1 ( .a ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1189, SubCellInst_SboxInst_4_n3}), .c ({new_AGEMA_signal_1479, SubCellInst_SboxInst_4_Q4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_XOR5_U1 ( .a ({new_AGEMA_signal_1193, SubCellInst_SboxInst_4_XX_2_}), .b ({new_AGEMA_signal_1189, SubCellInst_SboxInst_4_n3}), .c ({new_AGEMA_signal_1480, SubCellInst_SboxInst_4_Q6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_XOR6_U1 ( .a ({new_AGEMA_signal_1478, SubCellInst_SboxInst_4_Q1}), .b ({new_AGEMA_signal_1480, SubCellInst_SboxInst_4_Q6}), .c ({new_AGEMA_signal_1562, SubCellInst_SboxInst_4_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_XOR8_U1 ( .a ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1189, SubCellInst_SboxInst_4_n3}), .c ({new_AGEMA_signal_1481, SubCellInst_SboxInst_4_L2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_U1 ( .a ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({new_AGEMA_signal_1195, SubCellInst_SboxInst_5_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_XOR_i1_U1 ( .a ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({Ciphertext_s1[23], Ciphertext_s0[23]}), .c ({new_AGEMA_signal_1197, SubCellInst_SboxInst_5_XX_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_XOR_i2_U1 ( .a ({Ciphertext_s1[20], Ciphertext_s0[20]}), .b ({Ciphertext_s1[22], Ciphertext_s0[22]}), .c ({new_AGEMA_signal_1199, SubCellInst_SboxInst_5_XX_2_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_XOR0_U1 ( .a ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1199, SubCellInst_SboxInst_5_XX_2_}), .c ({new_AGEMA_signal_1483, SubCellInst_SboxInst_5_Q0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_XOR1_U1 ( .a ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1197, SubCellInst_SboxInst_5_XX_1_}), .c ({new_AGEMA_signal_1484, SubCellInst_SboxInst_5_Q1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_XOR3_U1 ( .a ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1195, SubCellInst_SboxInst_5_n3}), .c ({new_AGEMA_signal_1485, SubCellInst_SboxInst_5_Q4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_XOR5_U1 ( .a ({new_AGEMA_signal_1199, SubCellInst_SboxInst_5_XX_2_}), .b ({new_AGEMA_signal_1195, SubCellInst_SboxInst_5_n3}), .c ({new_AGEMA_signal_1486, SubCellInst_SboxInst_5_Q6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_XOR6_U1 ( .a ({new_AGEMA_signal_1484, SubCellInst_SboxInst_5_Q1}), .b ({new_AGEMA_signal_1486, SubCellInst_SboxInst_5_Q6}), .c ({new_AGEMA_signal_1565, SubCellInst_SboxInst_5_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_XOR8_U1 ( .a ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1195, SubCellInst_SboxInst_5_n3}), .c ({new_AGEMA_signal_1487, SubCellInst_SboxInst_5_L2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_U1 ( .a ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({new_AGEMA_signal_1201, SubCellInst_SboxInst_6_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_XOR_i1_U1 ( .a ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({Ciphertext_s1[27], Ciphertext_s0[27]}), .c ({new_AGEMA_signal_1203, SubCellInst_SboxInst_6_XX_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_XOR_i2_U1 ( .a ({Ciphertext_s1[24], Ciphertext_s0[24]}), .b ({Ciphertext_s1[26], Ciphertext_s0[26]}), .c ({new_AGEMA_signal_1205, SubCellInst_SboxInst_6_XX_2_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_XOR0_U1 ( .a ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1205, SubCellInst_SboxInst_6_XX_2_}), .c ({new_AGEMA_signal_1489, SubCellInst_SboxInst_6_Q0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_XOR1_U1 ( .a ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1203, SubCellInst_SboxInst_6_XX_1_}), .c ({new_AGEMA_signal_1490, SubCellInst_SboxInst_6_Q1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_XOR3_U1 ( .a ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1201, SubCellInst_SboxInst_6_n3}), .c ({new_AGEMA_signal_1491, SubCellInst_SboxInst_6_Q4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_XOR5_U1 ( .a ({new_AGEMA_signal_1205, SubCellInst_SboxInst_6_XX_2_}), .b ({new_AGEMA_signal_1201, SubCellInst_SboxInst_6_n3}), .c ({new_AGEMA_signal_1492, SubCellInst_SboxInst_6_Q6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_XOR6_U1 ( .a ({new_AGEMA_signal_1490, SubCellInst_SboxInst_6_Q1}), .b ({new_AGEMA_signal_1492, SubCellInst_SboxInst_6_Q6}), .c ({new_AGEMA_signal_1568, SubCellInst_SboxInst_6_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_XOR8_U1 ( .a ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1201, SubCellInst_SboxInst_6_n3}), .c ({new_AGEMA_signal_1493, SubCellInst_SboxInst_6_L2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_U1 ( .a ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({new_AGEMA_signal_1207, SubCellInst_SboxInst_7_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_XOR_i1_U1 ( .a ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({Ciphertext_s1[31], Ciphertext_s0[31]}), .c ({new_AGEMA_signal_1209, SubCellInst_SboxInst_7_XX_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_XOR_i2_U1 ( .a ({Ciphertext_s1[28], Ciphertext_s0[28]}), .b ({Ciphertext_s1[30], Ciphertext_s0[30]}), .c ({new_AGEMA_signal_1211, SubCellInst_SboxInst_7_XX_2_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_XOR0_U1 ( .a ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1211, SubCellInst_SboxInst_7_XX_2_}), .c ({new_AGEMA_signal_1495, SubCellInst_SboxInst_7_Q0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_XOR1_U1 ( .a ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1209, SubCellInst_SboxInst_7_XX_1_}), .c ({new_AGEMA_signal_1496, SubCellInst_SboxInst_7_Q1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_XOR3_U1 ( .a ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1207, SubCellInst_SboxInst_7_n3}), .c ({new_AGEMA_signal_1497, SubCellInst_SboxInst_7_Q4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_XOR5_U1 ( .a ({new_AGEMA_signal_1211, SubCellInst_SboxInst_7_XX_2_}), .b ({new_AGEMA_signal_1207, SubCellInst_SboxInst_7_n3}), .c ({new_AGEMA_signal_1498, SubCellInst_SboxInst_7_Q6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_XOR6_U1 ( .a ({new_AGEMA_signal_1496, SubCellInst_SboxInst_7_Q1}), .b ({new_AGEMA_signal_1498, SubCellInst_SboxInst_7_Q6}), .c ({new_AGEMA_signal_1571, SubCellInst_SboxInst_7_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_XOR8_U1 ( .a ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1207, SubCellInst_SboxInst_7_n3}), .c ({new_AGEMA_signal_1499, SubCellInst_SboxInst_7_L2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_U1 ( .a ({Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({new_AGEMA_signal_1213, SubCellInst_SboxInst_8_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_XOR_i1_U1 ( .a ({Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({Ciphertext_s1[35], Ciphertext_s0[35]}), .c ({new_AGEMA_signal_1215, SubCellInst_SboxInst_8_XX_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_XOR_i2_U1 ( .a ({Ciphertext_s1[32], Ciphertext_s0[32]}), .b ({Ciphertext_s1[34], Ciphertext_s0[34]}), .c ({new_AGEMA_signal_1217, SubCellInst_SboxInst_8_XX_2_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_XOR0_U1 ( .a ({Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1217, SubCellInst_SboxInst_8_XX_2_}), .c ({new_AGEMA_signal_1501, SubCellInst_SboxInst_8_Q0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_XOR1_U1 ( .a ({Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1215, SubCellInst_SboxInst_8_XX_1_}), .c ({new_AGEMA_signal_1502, SubCellInst_SboxInst_8_Q1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_XOR3_U1 ( .a ({Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1213, SubCellInst_SboxInst_8_n3}), .c ({new_AGEMA_signal_1503, SubCellInst_SboxInst_8_Q4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_XOR5_U1 ( .a ({new_AGEMA_signal_1217, SubCellInst_SboxInst_8_XX_2_}), .b ({new_AGEMA_signal_1213, SubCellInst_SboxInst_8_n3}), .c ({new_AGEMA_signal_1504, SubCellInst_SboxInst_8_Q6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_XOR6_U1 ( .a ({new_AGEMA_signal_1502, SubCellInst_SboxInst_8_Q1}), .b ({new_AGEMA_signal_1504, SubCellInst_SboxInst_8_Q6}), .c ({new_AGEMA_signal_1574, SubCellInst_SboxInst_8_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_XOR8_U1 ( .a ({Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1213, SubCellInst_SboxInst_8_n3}), .c ({new_AGEMA_signal_1505, SubCellInst_SboxInst_8_L2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_U1 ( .a ({Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({new_AGEMA_signal_1219, SubCellInst_SboxInst_9_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_XOR_i1_U1 ( .a ({Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({Ciphertext_s1[39], Ciphertext_s0[39]}), .c ({new_AGEMA_signal_1221, SubCellInst_SboxInst_9_XX_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_XOR_i2_U1 ( .a ({Ciphertext_s1[36], Ciphertext_s0[36]}), .b ({Ciphertext_s1[38], Ciphertext_s0[38]}), .c ({new_AGEMA_signal_1223, SubCellInst_SboxInst_9_XX_2_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_XOR0_U1 ( .a ({Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1223, SubCellInst_SboxInst_9_XX_2_}), .c ({new_AGEMA_signal_1507, SubCellInst_SboxInst_9_Q0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_XOR1_U1 ( .a ({Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1221, SubCellInst_SboxInst_9_XX_1_}), .c ({new_AGEMA_signal_1508, SubCellInst_SboxInst_9_Q1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_XOR3_U1 ( .a ({Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1219, SubCellInst_SboxInst_9_n3}), .c ({new_AGEMA_signal_1509, SubCellInst_SboxInst_9_Q4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_XOR5_U1 ( .a ({new_AGEMA_signal_1223, SubCellInst_SboxInst_9_XX_2_}), .b ({new_AGEMA_signal_1219, SubCellInst_SboxInst_9_n3}), .c ({new_AGEMA_signal_1510, SubCellInst_SboxInst_9_Q6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_XOR6_U1 ( .a ({new_AGEMA_signal_1508, SubCellInst_SboxInst_9_Q1}), .b ({new_AGEMA_signal_1510, SubCellInst_SboxInst_9_Q6}), .c ({new_AGEMA_signal_1577, SubCellInst_SboxInst_9_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_XOR8_U1 ( .a ({Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1219, SubCellInst_SboxInst_9_n3}), .c ({new_AGEMA_signal_1511, SubCellInst_SboxInst_9_L2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_U1 ( .a ({Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({new_AGEMA_signal_1225, SubCellInst_SboxInst_10_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_XOR_i1_U1 ( .a ({Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({Ciphertext_s1[43], Ciphertext_s0[43]}), .c ({new_AGEMA_signal_1227, SubCellInst_SboxInst_10_XX_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_XOR_i2_U1 ( .a ({Ciphertext_s1[40], Ciphertext_s0[40]}), .b ({Ciphertext_s1[42], Ciphertext_s0[42]}), .c ({new_AGEMA_signal_1229, SubCellInst_SboxInst_10_XX_2_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_XOR0_U1 ( .a ({Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1229, SubCellInst_SboxInst_10_XX_2_}), .c ({new_AGEMA_signal_1513, SubCellInst_SboxInst_10_Q0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_XOR1_U1 ( .a ({Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1227, SubCellInst_SboxInst_10_XX_1_}), .c ({new_AGEMA_signal_1514, SubCellInst_SboxInst_10_Q1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_XOR3_U1 ( .a ({Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1225, SubCellInst_SboxInst_10_n3}), .c ({new_AGEMA_signal_1515, SubCellInst_SboxInst_10_Q4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_XOR5_U1 ( .a ({new_AGEMA_signal_1229, SubCellInst_SboxInst_10_XX_2_}), .b ({new_AGEMA_signal_1225, SubCellInst_SboxInst_10_n3}), .c ({new_AGEMA_signal_1516, SubCellInst_SboxInst_10_Q6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_XOR6_U1 ( .a ({new_AGEMA_signal_1514, SubCellInst_SboxInst_10_Q1}), .b ({new_AGEMA_signal_1516, SubCellInst_SboxInst_10_Q6}), .c ({new_AGEMA_signal_1580, SubCellInst_SboxInst_10_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_XOR8_U1 ( .a ({Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1225, SubCellInst_SboxInst_10_n3}), .c ({new_AGEMA_signal_1517, SubCellInst_SboxInst_10_L2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_U1 ( .a ({Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({new_AGEMA_signal_1231, SubCellInst_SboxInst_11_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_XOR_i1_U1 ( .a ({Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({Ciphertext_s1[47], Ciphertext_s0[47]}), .c ({new_AGEMA_signal_1233, SubCellInst_SboxInst_11_XX_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_XOR_i2_U1 ( .a ({Ciphertext_s1[44], Ciphertext_s0[44]}), .b ({Ciphertext_s1[46], Ciphertext_s0[46]}), .c ({new_AGEMA_signal_1235, SubCellInst_SboxInst_11_XX_2_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_XOR0_U1 ( .a ({Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1235, SubCellInst_SboxInst_11_XX_2_}), .c ({new_AGEMA_signal_1519, SubCellInst_SboxInst_11_Q0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_XOR1_U1 ( .a ({Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1233, SubCellInst_SboxInst_11_XX_1_}), .c ({new_AGEMA_signal_1520, SubCellInst_SboxInst_11_Q1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_XOR3_U1 ( .a ({Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1231, SubCellInst_SboxInst_11_n3}), .c ({new_AGEMA_signal_1521, SubCellInst_SboxInst_11_Q4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_XOR5_U1 ( .a ({new_AGEMA_signal_1235, SubCellInst_SboxInst_11_XX_2_}), .b ({new_AGEMA_signal_1231, SubCellInst_SboxInst_11_n3}), .c ({new_AGEMA_signal_1522, SubCellInst_SboxInst_11_Q6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_XOR6_U1 ( .a ({new_AGEMA_signal_1520, SubCellInst_SboxInst_11_Q1}), .b ({new_AGEMA_signal_1522, SubCellInst_SboxInst_11_Q6}), .c ({new_AGEMA_signal_1583, SubCellInst_SboxInst_11_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_XOR8_U1 ( .a ({Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1231, SubCellInst_SboxInst_11_n3}), .c ({new_AGEMA_signal_1523, SubCellInst_SboxInst_11_L2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_U1 ( .a ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({new_AGEMA_signal_1237, SubCellInst_SboxInst_12_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_XOR_i1_U1 ( .a ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({Ciphertext_s1[51], Ciphertext_s0[51]}), .c ({new_AGEMA_signal_1239, SubCellInst_SboxInst_12_XX_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_XOR_i2_U1 ( .a ({Ciphertext_s1[48], Ciphertext_s0[48]}), .b ({Ciphertext_s1[50], Ciphertext_s0[50]}), .c ({new_AGEMA_signal_1241, SubCellInst_SboxInst_12_XX_2_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_XOR0_U1 ( .a ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1241, SubCellInst_SboxInst_12_XX_2_}), .c ({new_AGEMA_signal_1525, SubCellInst_SboxInst_12_Q0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_XOR1_U1 ( .a ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1239, SubCellInst_SboxInst_12_XX_1_}), .c ({new_AGEMA_signal_1526, SubCellInst_SboxInst_12_Q1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_XOR3_U1 ( .a ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1237, SubCellInst_SboxInst_12_n3}), .c ({new_AGEMA_signal_1527, SubCellInst_SboxInst_12_Q4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_XOR5_U1 ( .a ({new_AGEMA_signal_1241, SubCellInst_SboxInst_12_XX_2_}), .b ({new_AGEMA_signal_1237, SubCellInst_SboxInst_12_n3}), .c ({new_AGEMA_signal_1528, SubCellInst_SboxInst_12_Q6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_XOR6_U1 ( .a ({new_AGEMA_signal_1526, SubCellInst_SboxInst_12_Q1}), .b ({new_AGEMA_signal_1528, SubCellInst_SboxInst_12_Q6}), .c ({new_AGEMA_signal_1586, SubCellInst_SboxInst_12_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_XOR8_U1 ( .a ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1237, SubCellInst_SboxInst_12_n3}), .c ({new_AGEMA_signal_1529, SubCellInst_SboxInst_12_L2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_U1 ( .a ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({new_AGEMA_signal_1243, SubCellInst_SboxInst_13_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_XOR_i1_U1 ( .a ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({Ciphertext_s1[55], Ciphertext_s0[55]}), .c ({new_AGEMA_signal_1245, SubCellInst_SboxInst_13_XX_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_XOR_i2_U1 ( .a ({Ciphertext_s1[52], Ciphertext_s0[52]}), .b ({Ciphertext_s1[54], Ciphertext_s0[54]}), .c ({new_AGEMA_signal_1247, SubCellInst_SboxInst_13_XX_2_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_XOR0_U1 ( .a ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1247, SubCellInst_SboxInst_13_XX_2_}), .c ({new_AGEMA_signal_1531, SubCellInst_SboxInst_13_Q0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_XOR1_U1 ( .a ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1245, SubCellInst_SboxInst_13_XX_1_}), .c ({new_AGEMA_signal_1532, SubCellInst_SboxInst_13_Q1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_XOR3_U1 ( .a ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1243, SubCellInst_SboxInst_13_n3}), .c ({new_AGEMA_signal_1533, SubCellInst_SboxInst_13_Q4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_XOR5_U1 ( .a ({new_AGEMA_signal_1247, SubCellInst_SboxInst_13_XX_2_}), .b ({new_AGEMA_signal_1243, SubCellInst_SboxInst_13_n3}), .c ({new_AGEMA_signal_1534, SubCellInst_SboxInst_13_Q6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_XOR6_U1 ( .a ({new_AGEMA_signal_1532, SubCellInst_SboxInst_13_Q1}), .b ({new_AGEMA_signal_1534, SubCellInst_SboxInst_13_Q6}), .c ({new_AGEMA_signal_1589, SubCellInst_SboxInst_13_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_XOR8_U1 ( .a ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1243, SubCellInst_SboxInst_13_n3}), .c ({new_AGEMA_signal_1535, SubCellInst_SboxInst_13_L2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_U1 ( .a ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({new_AGEMA_signal_1249, SubCellInst_SboxInst_14_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_XOR_i1_U1 ( .a ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({Ciphertext_s1[59], Ciphertext_s0[59]}), .c ({new_AGEMA_signal_1251, SubCellInst_SboxInst_14_XX_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_XOR_i2_U1 ( .a ({Ciphertext_s1[56], Ciphertext_s0[56]}), .b ({Ciphertext_s1[58], Ciphertext_s0[58]}), .c ({new_AGEMA_signal_1253, SubCellInst_SboxInst_14_XX_2_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_XOR0_U1 ( .a ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1253, SubCellInst_SboxInst_14_XX_2_}), .c ({new_AGEMA_signal_1537, SubCellInst_SboxInst_14_Q0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_XOR1_U1 ( .a ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1251, SubCellInst_SboxInst_14_XX_1_}), .c ({new_AGEMA_signal_1538, SubCellInst_SboxInst_14_Q1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_XOR3_U1 ( .a ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1249, SubCellInst_SboxInst_14_n3}), .c ({new_AGEMA_signal_1539, SubCellInst_SboxInst_14_Q4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_XOR5_U1 ( .a ({new_AGEMA_signal_1253, SubCellInst_SboxInst_14_XX_2_}), .b ({new_AGEMA_signal_1249, SubCellInst_SboxInst_14_n3}), .c ({new_AGEMA_signal_1540, SubCellInst_SboxInst_14_Q6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_XOR6_U1 ( .a ({new_AGEMA_signal_1538, SubCellInst_SboxInst_14_Q1}), .b ({new_AGEMA_signal_1540, SubCellInst_SboxInst_14_Q6}), .c ({new_AGEMA_signal_1592, SubCellInst_SboxInst_14_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_XOR8_U1 ( .a ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1249, SubCellInst_SboxInst_14_n3}), .c ({new_AGEMA_signal_1541, SubCellInst_SboxInst_14_L2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_U1 ( .a ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({new_AGEMA_signal_1255, SubCellInst_SboxInst_15_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_XOR_i1_U1 ( .a ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({Ciphertext_s1[63], Ciphertext_s0[63]}), .c ({new_AGEMA_signal_1257, SubCellInst_SboxInst_15_XX_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_XOR_i2_U1 ( .a ({Ciphertext_s1[60], Ciphertext_s0[60]}), .b ({Ciphertext_s1[62], Ciphertext_s0[62]}), .c ({new_AGEMA_signal_1259, SubCellInst_SboxInst_15_XX_2_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_XOR0_U1 ( .a ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1259, SubCellInst_SboxInst_15_XX_2_}), .c ({new_AGEMA_signal_1543, SubCellInst_SboxInst_15_Q0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_XOR1_U1 ( .a ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1257, SubCellInst_SboxInst_15_XX_1_}), .c ({new_AGEMA_signal_1544, SubCellInst_SboxInst_15_Q1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_XOR3_U1 ( .a ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1255, SubCellInst_SboxInst_15_n3}), .c ({new_AGEMA_signal_1545, SubCellInst_SboxInst_15_Q4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_XOR5_U1 ( .a ({new_AGEMA_signal_1259, SubCellInst_SboxInst_15_XX_2_}), .b ({new_AGEMA_signal_1255, SubCellInst_SboxInst_15_n3}), .c ({new_AGEMA_signal_1546, SubCellInst_SboxInst_15_Q6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_XOR6_U1 ( .a ({new_AGEMA_signal_1544, SubCellInst_SboxInst_15_Q1}), .b ({new_AGEMA_signal_1546, SubCellInst_SboxInst_15_Q6}), .c ({new_AGEMA_signal_1595, SubCellInst_SboxInst_15_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_XOR8_U1 ( .a ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1255, SubCellInst_SboxInst_15_n3}), .c ({new_AGEMA_signal_1547, SubCellInst_SboxInst_15_L2}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_0_U1 ( .s (rst), .b ({new_AGEMA_signal_1260, TweakeyGeneration_key_Feedback[0]}), .a ({Key_s1[0], Key_s0[0]}), .c ({new_AGEMA_signal_1262, TweakeyGeneration_StateRegInput[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_1_U1 ( .s (rst), .b ({new_AGEMA_signal_1263, TweakeyGeneration_key_Feedback[1]}), .a ({Key_s1[1], Key_s0[1]}), .c ({new_AGEMA_signal_1265, TweakeyGeneration_StateRegInput[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_2_U1 ( .s (rst), .b ({new_AGEMA_signal_1266, TweakeyGeneration_key_Feedback[2]}), .a ({Key_s1[2], Key_s0[2]}), .c ({new_AGEMA_signal_1268, TweakeyGeneration_StateRegInput[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_3_U1 ( .s (rst), .b ({new_AGEMA_signal_1269, TweakeyGeneration_key_Feedback[3]}), .a ({Key_s1[3], Key_s0[3]}), .c ({new_AGEMA_signal_1271, TweakeyGeneration_StateRegInput[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_4_U1 ( .s (rst), .b ({new_AGEMA_signal_1272, TweakeyGeneration_key_Feedback[4]}), .a ({Key_s1[4], Key_s0[4]}), .c ({new_AGEMA_signal_1274, TweakeyGeneration_StateRegInput[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_5_U1 ( .s (rst), .b ({new_AGEMA_signal_1275, TweakeyGeneration_key_Feedback[5]}), .a ({Key_s1[5], Key_s0[5]}), .c ({new_AGEMA_signal_1277, TweakeyGeneration_StateRegInput[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_6_U1 ( .s (rst), .b ({new_AGEMA_signal_1278, TweakeyGeneration_key_Feedback[6]}), .a ({Key_s1[6], Key_s0[6]}), .c ({new_AGEMA_signal_1280, TweakeyGeneration_StateRegInput[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_7_U1 ( .s (rst), .b ({new_AGEMA_signal_1281, TweakeyGeneration_key_Feedback[7]}), .a ({Key_s1[7], Key_s0[7]}), .c ({new_AGEMA_signal_1283, TweakeyGeneration_StateRegInput[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_8_U1 ( .s (rst), .b ({new_AGEMA_signal_1284, TweakeyGeneration_key_Feedback[8]}), .a ({Key_s1[8], Key_s0[8]}), .c ({new_AGEMA_signal_1286, TweakeyGeneration_StateRegInput[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_9_U1 ( .s (rst), .b ({new_AGEMA_signal_1287, TweakeyGeneration_key_Feedback[9]}), .a ({Key_s1[9], Key_s0[9]}), .c ({new_AGEMA_signal_1289, TweakeyGeneration_StateRegInput[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_10_U1 ( .s (rst), .b ({new_AGEMA_signal_1290, TweakeyGeneration_key_Feedback[10]}), .a ({Key_s1[10], Key_s0[10]}), .c ({new_AGEMA_signal_1292, TweakeyGeneration_StateRegInput[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_11_U1 ( .s (rst), .b ({new_AGEMA_signal_1293, TweakeyGeneration_key_Feedback[11]}), .a ({Key_s1[11], Key_s0[11]}), .c ({new_AGEMA_signal_1295, TweakeyGeneration_StateRegInput[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_12_U1 ( .s (rst), .b ({new_AGEMA_signal_1296, TweakeyGeneration_key_Feedback[12]}), .a ({Key_s1[12], Key_s0[12]}), .c ({new_AGEMA_signal_1298, TweakeyGeneration_StateRegInput[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_13_U1 ( .s (rst), .b ({new_AGEMA_signal_1299, TweakeyGeneration_key_Feedback[13]}), .a ({Key_s1[13], Key_s0[13]}), .c ({new_AGEMA_signal_1301, TweakeyGeneration_StateRegInput[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_14_U1 ( .s (rst), .b ({new_AGEMA_signal_1302, TweakeyGeneration_key_Feedback[14]}), .a ({Key_s1[14], Key_s0[14]}), .c ({new_AGEMA_signal_1304, TweakeyGeneration_StateRegInput[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_15_U1 ( .s (rst), .b ({new_AGEMA_signal_1305, TweakeyGeneration_key_Feedback[15]}), .a ({Key_s1[15], Key_s0[15]}), .c ({new_AGEMA_signal_1307, TweakeyGeneration_StateRegInput[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_16_U1 ( .s (rst), .b ({new_AGEMA_signal_1308, TweakeyGeneration_key_Feedback[16]}), .a ({Key_s1[16], Key_s0[16]}), .c ({new_AGEMA_signal_1310, TweakeyGeneration_StateRegInput[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_17_U1 ( .s (rst), .b ({new_AGEMA_signal_1311, TweakeyGeneration_key_Feedback[17]}), .a ({Key_s1[17], Key_s0[17]}), .c ({new_AGEMA_signal_1313, TweakeyGeneration_StateRegInput[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_18_U1 ( .s (rst), .b ({new_AGEMA_signal_1314, TweakeyGeneration_key_Feedback[18]}), .a ({Key_s1[18], Key_s0[18]}), .c ({new_AGEMA_signal_1316, TweakeyGeneration_StateRegInput[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_19_U1 ( .s (rst), .b ({new_AGEMA_signal_1317, TweakeyGeneration_key_Feedback[19]}), .a ({Key_s1[19], Key_s0[19]}), .c ({new_AGEMA_signal_1319, TweakeyGeneration_StateRegInput[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_20_U1 ( .s (rst), .b ({new_AGEMA_signal_1320, TweakeyGeneration_key_Feedback[20]}), .a ({Key_s1[20], Key_s0[20]}), .c ({new_AGEMA_signal_1322, TweakeyGeneration_StateRegInput[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_21_U1 ( .s (rst), .b ({new_AGEMA_signal_1323, TweakeyGeneration_key_Feedback[21]}), .a ({Key_s1[21], Key_s0[21]}), .c ({new_AGEMA_signal_1325, TweakeyGeneration_StateRegInput[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_22_U1 ( .s (rst), .b ({new_AGEMA_signal_1326, TweakeyGeneration_key_Feedback[22]}), .a ({Key_s1[22], Key_s0[22]}), .c ({new_AGEMA_signal_1328, TweakeyGeneration_StateRegInput[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_23_U1 ( .s (rst), .b ({new_AGEMA_signal_1329, TweakeyGeneration_key_Feedback[23]}), .a ({Key_s1[23], Key_s0[23]}), .c ({new_AGEMA_signal_1331, TweakeyGeneration_StateRegInput[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_24_U1 ( .s (rst), .b ({new_AGEMA_signal_1332, TweakeyGeneration_key_Feedback[24]}), .a ({Key_s1[24], Key_s0[24]}), .c ({new_AGEMA_signal_1334, TweakeyGeneration_StateRegInput[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_25_U1 ( .s (rst), .b ({new_AGEMA_signal_1335, TweakeyGeneration_key_Feedback[25]}), .a ({Key_s1[25], Key_s0[25]}), .c ({new_AGEMA_signal_1337, TweakeyGeneration_StateRegInput[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_26_U1 ( .s (rst), .b ({new_AGEMA_signal_1338, TweakeyGeneration_key_Feedback[26]}), .a ({Key_s1[26], Key_s0[26]}), .c ({new_AGEMA_signal_1340, TweakeyGeneration_StateRegInput[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_27_U1 ( .s (rst), .b ({new_AGEMA_signal_1341, TweakeyGeneration_key_Feedback[27]}), .a ({Key_s1[27], Key_s0[27]}), .c ({new_AGEMA_signal_1343, TweakeyGeneration_StateRegInput[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_28_U1 ( .s (rst), .b ({new_AGEMA_signal_1344, TweakeyGeneration_key_Feedback[28]}), .a ({Key_s1[28], Key_s0[28]}), .c ({new_AGEMA_signal_1346, TweakeyGeneration_StateRegInput[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_29_U1 ( .s (rst), .b ({new_AGEMA_signal_1347, TweakeyGeneration_key_Feedback[29]}), .a ({Key_s1[29], Key_s0[29]}), .c ({new_AGEMA_signal_1349, TweakeyGeneration_StateRegInput[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_30_U1 ( .s (rst), .b ({new_AGEMA_signal_1350, TweakeyGeneration_key_Feedback[30]}), .a ({Key_s1[30], Key_s0[30]}), .c ({new_AGEMA_signal_1352, TweakeyGeneration_StateRegInput[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_31_U1 ( .s (rst), .b ({new_AGEMA_signal_1353, TweakeyGeneration_key_Feedback[31]}), .a ({Key_s1[31], Key_s0[31]}), .c ({new_AGEMA_signal_1355, TweakeyGeneration_StateRegInput[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_32_U1 ( .s (rst), .b ({new_AGEMA_signal_1356, TweakeyGeneration_key_Feedback[32]}), .a ({Key_s1[32], Key_s0[32]}), .c ({new_AGEMA_signal_1358, TweakeyGeneration_StateRegInput[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_33_U1 ( .s (rst), .b ({new_AGEMA_signal_1359, TweakeyGeneration_key_Feedback[33]}), .a ({Key_s1[33], Key_s0[33]}), .c ({new_AGEMA_signal_1361, TweakeyGeneration_StateRegInput[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_34_U1 ( .s (rst), .b ({new_AGEMA_signal_1362, TweakeyGeneration_key_Feedback[34]}), .a ({Key_s1[34], Key_s0[34]}), .c ({new_AGEMA_signal_1364, TweakeyGeneration_StateRegInput[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_35_U1 ( .s (rst), .b ({new_AGEMA_signal_1365, TweakeyGeneration_key_Feedback[35]}), .a ({Key_s1[35], Key_s0[35]}), .c ({new_AGEMA_signal_1367, TweakeyGeneration_StateRegInput[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_36_U1 ( .s (rst), .b ({new_AGEMA_signal_1368, TweakeyGeneration_key_Feedback[36]}), .a ({Key_s1[36], Key_s0[36]}), .c ({new_AGEMA_signal_1370, TweakeyGeneration_StateRegInput[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_37_U1 ( .s (rst), .b ({new_AGEMA_signal_1371, TweakeyGeneration_key_Feedback[37]}), .a ({Key_s1[37], Key_s0[37]}), .c ({new_AGEMA_signal_1373, TweakeyGeneration_StateRegInput[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_38_U1 ( .s (rst), .b ({new_AGEMA_signal_1374, TweakeyGeneration_key_Feedback[38]}), .a ({Key_s1[38], Key_s0[38]}), .c ({new_AGEMA_signal_1376, TweakeyGeneration_StateRegInput[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_39_U1 ( .s (rst), .b ({new_AGEMA_signal_1377, TweakeyGeneration_key_Feedback[39]}), .a ({Key_s1[39], Key_s0[39]}), .c ({new_AGEMA_signal_1379, TweakeyGeneration_StateRegInput[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_40_U1 ( .s (rst), .b ({new_AGEMA_signal_1380, TweakeyGeneration_key_Feedback[40]}), .a ({Key_s1[40], Key_s0[40]}), .c ({new_AGEMA_signal_1382, TweakeyGeneration_StateRegInput[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_41_U1 ( .s (rst), .b ({new_AGEMA_signal_1383, TweakeyGeneration_key_Feedback[41]}), .a ({Key_s1[41], Key_s0[41]}), .c ({new_AGEMA_signal_1385, TweakeyGeneration_StateRegInput[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_42_U1 ( .s (rst), .b ({new_AGEMA_signal_1386, TweakeyGeneration_key_Feedback[42]}), .a ({Key_s1[42], Key_s0[42]}), .c ({new_AGEMA_signal_1388, TweakeyGeneration_StateRegInput[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_43_U1 ( .s (rst), .b ({new_AGEMA_signal_1389, TweakeyGeneration_key_Feedback[43]}), .a ({Key_s1[43], Key_s0[43]}), .c ({new_AGEMA_signal_1391, TweakeyGeneration_StateRegInput[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_44_U1 ( .s (rst), .b ({new_AGEMA_signal_1392, TweakeyGeneration_key_Feedback[44]}), .a ({Key_s1[44], Key_s0[44]}), .c ({new_AGEMA_signal_1394, TweakeyGeneration_StateRegInput[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_45_U1 ( .s (rst), .b ({new_AGEMA_signal_1395, TweakeyGeneration_key_Feedback[45]}), .a ({Key_s1[45], Key_s0[45]}), .c ({new_AGEMA_signal_1397, TweakeyGeneration_StateRegInput[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_46_U1 ( .s (rst), .b ({new_AGEMA_signal_1398, TweakeyGeneration_key_Feedback[46]}), .a ({Key_s1[46], Key_s0[46]}), .c ({new_AGEMA_signal_1400, TweakeyGeneration_StateRegInput[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_47_U1 ( .s (rst), .b ({new_AGEMA_signal_1401, TweakeyGeneration_key_Feedback[47]}), .a ({Key_s1[47], Key_s0[47]}), .c ({new_AGEMA_signal_1403, TweakeyGeneration_StateRegInput[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_48_U1 ( .s (rst), .b ({new_AGEMA_signal_1404, TweakeyGeneration_key_Feedback[48]}), .a ({Key_s1[48], Key_s0[48]}), .c ({new_AGEMA_signal_1406, TweakeyGeneration_StateRegInput[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_49_U1 ( .s (rst), .b ({new_AGEMA_signal_1407, TweakeyGeneration_key_Feedback[49]}), .a ({Key_s1[49], Key_s0[49]}), .c ({new_AGEMA_signal_1409, TweakeyGeneration_StateRegInput[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_50_U1 ( .s (rst), .b ({new_AGEMA_signal_1410, TweakeyGeneration_key_Feedback[50]}), .a ({Key_s1[50], Key_s0[50]}), .c ({new_AGEMA_signal_1412, TweakeyGeneration_StateRegInput[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_51_U1 ( .s (rst), .b ({new_AGEMA_signal_1413, TweakeyGeneration_key_Feedback[51]}), .a ({Key_s1[51], Key_s0[51]}), .c ({new_AGEMA_signal_1415, TweakeyGeneration_StateRegInput[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_52_U1 ( .s (rst), .b ({new_AGEMA_signal_1416, TweakeyGeneration_key_Feedback[52]}), .a ({Key_s1[52], Key_s0[52]}), .c ({new_AGEMA_signal_1418, TweakeyGeneration_StateRegInput[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_53_U1 ( .s (rst), .b ({new_AGEMA_signal_1419, TweakeyGeneration_key_Feedback[53]}), .a ({Key_s1[53], Key_s0[53]}), .c ({new_AGEMA_signal_1421, TweakeyGeneration_StateRegInput[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_54_U1 ( .s (rst), .b ({new_AGEMA_signal_1422, TweakeyGeneration_key_Feedback[54]}), .a ({Key_s1[54], Key_s0[54]}), .c ({new_AGEMA_signal_1424, TweakeyGeneration_StateRegInput[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_55_U1 ( .s (rst), .b ({new_AGEMA_signal_1425, TweakeyGeneration_key_Feedback[55]}), .a ({Key_s1[55], Key_s0[55]}), .c ({new_AGEMA_signal_1427, TweakeyGeneration_StateRegInput[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_56_U1 ( .s (rst), .b ({new_AGEMA_signal_1428, TweakeyGeneration_key_Feedback[56]}), .a ({Key_s1[56], Key_s0[56]}), .c ({new_AGEMA_signal_1430, TweakeyGeneration_StateRegInput[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_57_U1 ( .s (rst), .b ({new_AGEMA_signal_1431, TweakeyGeneration_key_Feedback[57]}), .a ({Key_s1[57], Key_s0[57]}), .c ({new_AGEMA_signal_1433, TweakeyGeneration_StateRegInput[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_58_U1 ( .s (rst), .b ({new_AGEMA_signal_1434, TweakeyGeneration_key_Feedback[58]}), .a ({Key_s1[58], Key_s0[58]}), .c ({new_AGEMA_signal_1436, TweakeyGeneration_StateRegInput[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_59_U1 ( .s (rst), .b ({new_AGEMA_signal_1437, TweakeyGeneration_key_Feedback[59]}), .a ({Key_s1[59], Key_s0[59]}), .c ({new_AGEMA_signal_1439, TweakeyGeneration_StateRegInput[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_60_U1 ( .s (rst), .b ({new_AGEMA_signal_1440, TweakeyGeneration_key_Feedback[60]}), .a ({Key_s1[60], Key_s0[60]}), .c ({new_AGEMA_signal_1442, TweakeyGeneration_StateRegInput[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_61_U1 ( .s (rst), .b ({new_AGEMA_signal_1443, TweakeyGeneration_key_Feedback[61]}), .a ({Key_s1[61], Key_s0[61]}), .c ({new_AGEMA_signal_1445, TweakeyGeneration_StateRegInput[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_62_U1 ( .s (rst), .b ({new_AGEMA_signal_1446, TweakeyGeneration_key_Feedback[62]}), .a ({Key_s1[62], Key_s0[62]}), .c ({new_AGEMA_signal_1448, TweakeyGeneration_StateRegInput[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_63_U1 ( .s (rst), .b ({new_AGEMA_signal_1449, TweakeyGeneration_key_Feedback[63]}), .a ({Key_s1[63], Key_s0[63]}), .c ({new_AGEMA_signal_1451, TweakeyGeneration_StateRegInput[63]}) ) ;
    MUX2_X1 FSMMUX_MUXInst_0_U1 ( .S (rst), .A (FSMUpdate[0]), .B (1'b1), .Z (FSMSelected[0]) ) ;
    MUX2_X1 FSMMUX_MUXInst_1_U1 ( .S (rst), .A (FSMUpdate[1]), .B (1'b0), .Z (FSMSelected[1]) ) ;
    MUX2_X1 FSMMUX_MUXInst_2_U1 ( .S (rst), .A (FSMUpdate[2]), .B (1'b0), .Z (FSMSelected[2]) ) ;
    MUX2_X1 FSMMUX_MUXInst_3_U1 ( .S (rst), .A (FSMUpdate[3]), .B (1'b0), .Z (FSMSelected[3]) ) ;
    MUX2_X1 FSMMUX_MUXInst_4_U1 ( .S (rst), .A (FSMUpdate[4]), .B (1'b0), .Z (FSMSelected[4]) ) ;
    MUX2_X1 FSMMUX_MUXInst_5_U1 ( .S (rst), .A (FSMUpdate[5]), .B (1'b0), .Z (FSMSelected[5]) ) ;
    MUX2_X1 FSMUpdateInst_StateUpdateInst_0_U5 ( .S (FSM[4]), .A (FSMUpdateInst_StateUpdateInst_0_n4), .B (FSM[5]), .Z (FSMUpdate[0]) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_0_U4 ( .A1 (FSM[5]), .A2 (FSMUpdateInst_StateUpdateInst_0_n3), .ZN (FSMUpdateInst_StateUpdateInst_0_n4) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_0_U3 ( .A1 (FSMUpdateInst_StateUpdateInst_0_n2), .A2 (FSMUpdateInst_StateUpdateInst_0_n1), .ZN (FSMUpdateInst_StateUpdateInst_0_n3) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_0_U2 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdate[4]), .ZN (FSMUpdateInst_StateUpdateInst_0_n1) ) ;
    AND2_X1 FSMUpdateInst_StateUpdateInst_0_U1 ( .A1 (FSMUpdate[1]), .A2 (FSM[1]), .ZN (FSMUpdateInst_StateUpdateInst_0_n2) ) ;
    AND2_X1 FSMUpdateInst_StateUpdateInst_2_U5 ( .A1 (FSMUpdateInst_StateUpdateInst_2_n4), .A2 (FSM[1]), .ZN (FSMUpdate[2]) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_2_U4 ( .A1 (FSMUpdateInst_StateUpdateInst_2_n3), .A2 (FSM[5]), .ZN (FSMUpdateInst_StateUpdateInst_2_n4) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_2_U3 ( .A1 (FSM[4]), .A2 (FSMUpdateInst_StateUpdateInst_2_n2), .ZN (FSMUpdateInst_StateUpdateInst_2_n3) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_2_U2 ( .A1 (FSMUpdate[1]), .A2 (FSMUpdateInst_StateUpdateInst_2_n1), .ZN (FSMUpdateInst_StateUpdateInst_2_n2) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_2_U1 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdate[4]), .ZN (FSMUpdateInst_StateUpdateInst_2_n1) ) ;
    OR2_X1 FSMUpdateInst_StateUpdateInst_5_U5 ( .A1 (FSM[4]), .A2 (FSMUpdateInst_StateUpdateInst_5_n4), .ZN (FSMUpdate[5]) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_5_U4 ( .A1 (FSMUpdate[4]), .A2 (FSMUpdateInst_StateUpdateInst_5_n3), .ZN (FSMUpdateInst_StateUpdateInst_5_n4) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_5_U3 ( .A1 (FSM[5]), .A2 (FSMUpdateInst_StateUpdateInst_5_n2), .ZN (FSMUpdateInst_StateUpdateInst_5_n3) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_5_U2 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdateInst_StateUpdateInst_5_n1), .ZN (FSMUpdateInst_StateUpdateInst_5_n2) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_5_U1 ( .A1 (FSMUpdate[1]), .A2 (FSM[1]), .ZN (FSMUpdateInst_StateUpdateInst_5_n1) ) ;
    NOR2_X1 FSMSignalsInst_doneInst_U6 ( .A1 (FSMSignalsInst_doneInst_n5), .A2 (FSMSignalsInst_doneInst_n4), .ZN (done) ) ;
    NAND2_X1 FSMSignalsInst_doneInst_U5 ( .A1 (FSM[4]), .A2 (FSM[5]), .ZN (FSMSignalsInst_doneInst_n4) ) ;
    NAND2_X1 FSMSignalsInst_doneInst_U4 ( .A1 (FSMSignalsInst_doneInst_n3), .A2 (FSMSignalsInst_doneInst_n2), .ZN (FSMSignalsInst_doneInst_n5) ) ;
    NOR2_X1 FSMSignalsInst_doneInst_U3 ( .A1 (FSMUpdate[4]), .A2 (FSMSignalsInst_doneInst_n1), .ZN (FSMSignalsInst_doneInst_n2) ) ;
    INV_X1 FSMSignalsInst_doneInst_U2 ( .A (FSMUpdate[1]), .ZN (FSMSignalsInst_doneInst_n1) ) ;
    NOR2_X1 FSMSignalsInst_doneInst_U1 ( .A1 (FSM[1]), .A2 (FSMUpdate[3]), .ZN (FSMSignalsInst_doneInst_n3) ) ;
    ClockGatingController #(5) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_2_U1 ( .s (rst), .b ({new_AGEMA_signal_1915, MCOutput[2]}), .a ({Plaintext_s1[2], Plaintext_s0[2]}), .c ({new_AGEMA_signal_1922, StateRegInput[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_3_U1 ( .s (rst), .b ({new_AGEMA_signal_1975, MCOutput[3]}), .a ({Plaintext_s1[3], Plaintext_s0[3]}), .c ({new_AGEMA_signal_1982, StateRegInput[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_6_U1 ( .s (rst), .b ({new_AGEMA_signal_1917, MCOutput[6]}), .a ({Plaintext_s1[6], Plaintext_s0[6]}), .c ({new_AGEMA_signal_1924, StateRegInput[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_7_U1 ( .s (rst), .b ({new_AGEMA_signal_1977, MCOutput[7]}), .a ({Plaintext_s1[7], Plaintext_s0[7]}), .c ({new_AGEMA_signal_1984, StateRegInput[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_10_U1 ( .s (rst), .b ({new_AGEMA_signal_1919, MCOutput[10]}), .a ({Plaintext_s1[10], Plaintext_s0[10]}), .c ({new_AGEMA_signal_1926, StateRegInput[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_11_U1 ( .s (rst), .b ({new_AGEMA_signal_1979, MCOutput[11]}), .a ({Plaintext_s1[11], Plaintext_s0[11]}), .c ({new_AGEMA_signal_1986, StateRegInput[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_14_U1 ( .s (rst), .b ({new_AGEMA_signal_2033, MCOutput[14]}), .a ({Plaintext_s1[14], Plaintext_s0[14]}), .c ({new_AGEMA_signal_2042, StateRegInput[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_15_U1 ( .s (rst), .b ({new_AGEMA_signal_2077, MCOutput[15]}), .a ({Plaintext_s1[15], Plaintext_s0[15]}), .c ({new_AGEMA_signal_2085, StateRegInput[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_18_U1 ( .s (rst), .b ({new_AGEMA_signal_1909, MCOutput[18]}), .a ({Plaintext_s1[18], Plaintext_s0[18]}), .c ({new_AGEMA_signal_1928, StateRegInput[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_19_U1 ( .s (rst), .b ({new_AGEMA_signal_1968, MCOutput[19]}), .a ({Plaintext_s1[19], Plaintext_s0[19]}), .c ({new_AGEMA_signal_1988, StateRegInput[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_22_U1 ( .s (rst), .b ({new_AGEMA_signal_1911, MCOutput[22]}), .a ({Plaintext_s1[22], Plaintext_s0[22]}), .c ({new_AGEMA_signal_1930, StateRegInput[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_23_U1 ( .s (rst), .b ({new_AGEMA_signal_1970, MCOutput[23]}), .a ({Plaintext_s1[23], Plaintext_s0[23]}), .c ({new_AGEMA_signal_1990, StateRegInput[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_26_U1 ( .s (rst), .b ({new_AGEMA_signal_2023, MCOutput[26]}), .a ({Plaintext_s1[26], Plaintext_s0[26]}), .c ({new_AGEMA_signal_2048, StateRegInput[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_27_U1 ( .s (rst), .b ({new_AGEMA_signal_2071, MCOutput[27]}), .a ({Plaintext_s1[27], Plaintext_s0[27]}), .c ({new_AGEMA_signal_2091, StateRegInput[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_30_U1 ( .s (rst), .b ({new_AGEMA_signal_1913, MCOutput[30]}), .a ({Plaintext_s1[30], Plaintext_s0[30]}), .c ({new_AGEMA_signal_1932, StateRegInput[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_31_U1 ( .s (rst), .b ({new_AGEMA_signal_1973, MCOutput[31]}), .a ({Plaintext_s1[31], Plaintext_s0[31]}), .c ({new_AGEMA_signal_1992, StateRegInput[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_34_U1 ( .s (rst), .b ({new_AGEMA_signal_1810, MCOutput[34]}), .a ({Plaintext_s1[34], Plaintext_s0[34]}), .c ({new_AGEMA_signal_1821, StateRegInput[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_35_U1 ( .s (rst), .b ({new_AGEMA_signal_1854, MCOutput[35]}), .a ({Plaintext_s1[35], Plaintext_s0[35]}), .c ({new_AGEMA_signal_1874, StateRegInput[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_38_U1 ( .s (rst), .b ({new_AGEMA_signal_1812, MCOutput[38]}), .a ({Plaintext_s1[38], Plaintext_s0[38]}), .c ({new_AGEMA_signal_1823, StateRegInput[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_39_U1 ( .s (rst), .b ({new_AGEMA_signal_1856, MCOutput[39]}), .a ({Plaintext_s1[39], Plaintext_s0[39]}), .c ({new_AGEMA_signal_1876, StateRegInput[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_42_U1 ( .s (rst), .b ({new_AGEMA_signal_1814, MCOutput[42]}), .a ({Plaintext_s1[42], Plaintext_s0[42]}), .c ({new_AGEMA_signal_1825, StateRegInput[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_43_U1 ( .s (rst), .b ({new_AGEMA_signal_1858, MCOutput[43]}), .a ({Plaintext_s1[43], Plaintext_s0[43]}), .c ({new_AGEMA_signal_1878, StateRegInput[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_46_U1 ( .s (rst), .b ({new_AGEMA_signal_1898, MCOutput[46]}), .a ({Plaintext_s1[46], Plaintext_s0[46]}), .c ({new_AGEMA_signal_1940, StateRegInput[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_47_U1 ( .s (rst), .b ({new_AGEMA_signal_1958, MCOutput[47]}), .a ({Plaintext_s1[47], Plaintext_s0[47]}), .c ({new_AGEMA_signal_2000, StateRegInput[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_50_U1 ( .s (rst), .b ({new_AGEMA_signal_1901, MCOutput[50]}), .a ({Plaintext_s1[50], Plaintext_s0[50]}), .c ({new_AGEMA_signal_1942, StateRegInput[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_51_U1 ( .s (rst), .b ({new_AGEMA_signal_1960, MCOutput[51]}), .a ({Plaintext_s1[51], Plaintext_s0[51]}), .c ({new_AGEMA_signal_2002, StateRegInput[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_54_U1 ( .s (rst), .b ({new_AGEMA_signal_1903, MCOutput[54]}), .a ({Plaintext_s1[54], Plaintext_s0[54]}), .c ({new_AGEMA_signal_1944, StateRegInput[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_55_U1 ( .s (rst), .b ({new_AGEMA_signal_1963, MCOutput[55]}), .a ({Plaintext_s1[55], Plaintext_s0[55]}), .c ({new_AGEMA_signal_2004, StateRegInput[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_58_U1 ( .s (rst), .b ({new_AGEMA_signal_1906, MCOutput[58]}), .a ({Plaintext_s1[58], Plaintext_s0[58]}), .c ({new_AGEMA_signal_1946, StateRegInput[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_59_U1 ( .s (rst), .b ({new_AGEMA_signal_1965, MCOutput[59]}), .a ({Plaintext_s1[59], Plaintext_s0[59]}), .c ({new_AGEMA_signal_2006, StateRegInput[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_62_U1 ( .s (rst), .b ({new_AGEMA_signal_2017, MCOutput[62]}), .a ({Plaintext_s1[62], Plaintext_s0[62]}), .c ({new_AGEMA_signal_2060, StateRegInput[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_63_U1 ( .s (rst), .b ({new_AGEMA_signal_2067, MCOutput[63]}), .a ({Plaintext_s1[63], Plaintext_s0[63]}), .c ({new_AGEMA_signal_2103, StateRegInput[63]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_U3 ( .a ({new_AGEMA_signal_1663, SubCellInst_SboxInst_0_YY_1_}), .b ({new_AGEMA_signal_1724, ShiftRowsOutput[7]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_U2 ( .a ({new_AGEMA_signal_1599, SubCellInst_SboxInst_0_YY_0_}), .b ({new_AGEMA_signal_1660, ShiftRowsOutput[6]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_AND1_U1 ( .a ({new_AGEMA_signal_1165, SubCellInst_SboxInst_0_n3}), .b ({new_AGEMA_signal_1454, SubCellInst_SboxInst_0_Q1}), .clk (clk), .r (Fresh[0]), .c ({new_AGEMA_signal_1548, SubCellInst_SboxInst_0_T0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_XOR2_U1 ( .a ({new_AGEMA_signal_1453, SubCellInst_SboxInst_0_Q0}), .b ({new_AGEMA_signal_1548, SubCellInst_SboxInst_0_T0}), .c ({new_AGEMA_signal_1596, SubCellInst_SboxInst_0_Q2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_AND3_U1 ( .a ({new_AGEMA_signal_1165, SubCellInst_SboxInst_0_n3}), .b ({new_AGEMA_signal_1455, SubCellInst_SboxInst_0_Q4}), .clk (clk), .r (Fresh[1]), .c ({new_AGEMA_signal_1549, SubCellInst_SboxInst_0_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_XOR7_U1 ( .a ({new_AGEMA_signal_1550, SubCellInst_SboxInst_0_L1}), .b ({new_AGEMA_signal_1549, SubCellInst_SboxInst_0_T2}), .c ({new_AGEMA_signal_1597, SubCellInst_SboxInst_0_Q7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_XOR11_U1 ( .a ({new_AGEMA_signal_1169, SubCellInst_SboxInst_0_XX_2_}), .b ({new_AGEMA_signal_1548, SubCellInst_SboxInst_0_T0}), .c ({new_AGEMA_signal_1598, SubCellInst_SboxInst_0_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_XOR12_U1 ( .a ({new_AGEMA_signal_1598, SubCellInst_SboxInst_0_L3}), .b ({new_AGEMA_signal_1549, SubCellInst_SboxInst_0_T2}), .c ({new_AGEMA_signal_1663, SubCellInst_SboxInst_0_YY_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_XOR13_U1 ( .a ({new_AGEMA_signal_1167, SubCellInst_SboxInst_0_XX_1_}), .b ({new_AGEMA_signal_1549, SubCellInst_SboxInst_0_T2}), .c ({new_AGEMA_signal_1599, SubCellInst_SboxInst_0_YY_0_}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_U3 ( .a ({new_AGEMA_signal_1667, SubCellInst_SboxInst_1_YY_1_}), .b ({new_AGEMA_signal_1726, ShiftRowsOutput[11]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_U2 ( .a ({new_AGEMA_signal_1603, SubCellInst_SboxInst_1_YY_0_}), .b ({new_AGEMA_signal_1664, ShiftRowsOutput[10]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_AND1_U1 ( .a ({new_AGEMA_signal_1171, SubCellInst_SboxInst_1_n3}), .b ({new_AGEMA_signal_1460, SubCellInst_SboxInst_1_Q1}), .clk (clk), .r (Fresh[2]), .c ({new_AGEMA_signal_1551, SubCellInst_SboxInst_1_T0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_XOR2_U1 ( .a ({new_AGEMA_signal_1459, SubCellInst_SboxInst_1_Q0}), .b ({new_AGEMA_signal_1551, SubCellInst_SboxInst_1_T0}), .c ({new_AGEMA_signal_1600, SubCellInst_SboxInst_1_Q2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_AND3_U1 ( .a ({new_AGEMA_signal_1171, SubCellInst_SboxInst_1_n3}), .b ({new_AGEMA_signal_1461, SubCellInst_SboxInst_1_Q4}), .clk (clk), .r (Fresh[3]), .c ({new_AGEMA_signal_1552, SubCellInst_SboxInst_1_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_XOR7_U1 ( .a ({new_AGEMA_signal_1553, SubCellInst_SboxInst_1_L1}), .b ({new_AGEMA_signal_1552, SubCellInst_SboxInst_1_T2}), .c ({new_AGEMA_signal_1601, SubCellInst_SboxInst_1_Q7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_XOR11_U1 ( .a ({new_AGEMA_signal_1175, SubCellInst_SboxInst_1_XX_2_}), .b ({new_AGEMA_signal_1551, SubCellInst_SboxInst_1_T0}), .c ({new_AGEMA_signal_1602, SubCellInst_SboxInst_1_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_XOR12_U1 ( .a ({new_AGEMA_signal_1602, SubCellInst_SboxInst_1_L3}), .b ({new_AGEMA_signal_1552, SubCellInst_SboxInst_1_T2}), .c ({new_AGEMA_signal_1667, SubCellInst_SboxInst_1_YY_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_XOR13_U1 ( .a ({new_AGEMA_signal_1173, SubCellInst_SboxInst_1_XX_1_}), .b ({new_AGEMA_signal_1552, SubCellInst_SboxInst_1_T2}), .c ({new_AGEMA_signal_1603, SubCellInst_SboxInst_1_YY_0_}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_U3 ( .a ({new_AGEMA_signal_1671, SubCellInst_SboxInst_2_YY_1_}), .b ({new_AGEMA_signal_1728, ShiftRowsOutput[15]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_U2 ( .a ({new_AGEMA_signal_1607, SubCellInst_SboxInst_2_YY_0_}), .b ({new_AGEMA_signal_1668, ShiftRowsOutput[14]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_AND1_U1 ( .a ({new_AGEMA_signal_1177, SubCellInst_SboxInst_2_n3}), .b ({new_AGEMA_signal_1466, SubCellInst_SboxInst_2_Q1}), .clk (clk), .r (Fresh[4]), .c ({new_AGEMA_signal_1554, SubCellInst_SboxInst_2_T0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_XOR2_U1 ( .a ({new_AGEMA_signal_1465, SubCellInst_SboxInst_2_Q0}), .b ({new_AGEMA_signal_1554, SubCellInst_SboxInst_2_T0}), .c ({new_AGEMA_signal_1604, SubCellInst_SboxInst_2_Q2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_AND3_U1 ( .a ({new_AGEMA_signal_1177, SubCellInst_SboxInst_2_n3}), .b ({new_AGEMA_signal_1467, SubCellInst_SboxInst_2_Q4}), .clk (clk), .r (Fresh[5]), .c ({new_AGEMA_signal_1555, SubCellInst_SboxInst_2_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_XOR7_U1 ( .a ({new_AGEMA_signal_1556, SubCellInst_SboxInst_2_L1}), .b ({new_AGEMA_signal_1555, SubCellInst_SboxInst_2_T2}), .c ({new_AGEMA_signal_1605, SubCellInst_SboxInst_2_Q7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_XOR11_U1 ( .a ({new_AGEMA_signal_1181, SubCellInst_SboxInst_2_XX_2_}), .b ({new_AGEMA_signal_1554, SubCellInst_SboxInst_2_T0}), .c ({new_AGEMA_signal_1606, SubCellInst_SboxInst_2_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_XOR12_U1 ( .a ({new_AGEMA_signal_1606, SubCellInst_SboxInst_2_L3}), .b ({new_AGEMA_signal_1555, SubCellInst_SboxInst_2_T2}), .c ({new_AGEMA_signal_1671, SubCellInst_SboxInst_2_YY_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_XOR13_U1 ( .a ({new_AGEMA_signal_1179, SubCellInst_SboxInst_2_XX_1_}), .b ({new_AGEMA_signal_1555, SubCellInst_SboxInst_2_T2}), .c ({new_AGEMA_signal_1607, SubCellInst_SboxInst_2_YY_0_}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_U3 ( .a ({new_AGEMA_signal_1675, SubCellInst_SboxInst_3_YY_1_}), .b ({new_AGEMA_signal_1730, ShiftRowsOutput[3]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_U2 ( .a ({new_AGEMA_signal_1611, SubCellInst_SboxInst_3_YY_0_}), .b ({new_AGEMA_signal_1672, ShiftRowsOutput[2]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_AND1_U1 ( .a ({new_AGEMA_signal_1183, SubCellInst_SboxInst_3_n3}), .b ({new_AGEMA_signal_1472, SubCellInst_SboxInst_3_Q1}), .clk (clk), .r (Fresh[6]), .c ({new_AGEMA_signal_1557, SubCellInst_SboxInst_3_T0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_XOR2_U1 ( .a ({new_AGEMA_signal_1471, SubCellInst_SboxInst_3_Q0}), .b ({new_AGEMA_signal_1557, SubCellInst_SboxInst_3_T0}), .c ({new_AGEMA_signal_1608, SubCellInst_SboxInst_3_Q2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_AND3_U1 ( .a ({new_AGEMA_signal_1183, SubCellInst_SboxInst_3_n3}), .b ({new_AGEMA_signal_1473, SubCellInst_SboxInst_3_Q4}), .clk (clk), .r (Fresh[7]), .c ({new_AGEMA_signal_1558, SubCellInst_SboxInst_3_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_XOR7_U1 ( .a ({new_AGEMA_signal_1559, SubCellInst_SboxInst_3_L1}), .b ({new_AGEMA_signal_1558, SubCellInst_SboxInst_3_T2}), .c ({new_AGEMA_signal_1609, SubCellInst_SboxInst_3_Q7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_XOR11_U1 ( .a ({new_AGEMA_signal_1187, SubCellInst_SboxInst_3_XX_2_}), .b ({new_AGEMA_signal_1557, SubCellInst_SboxInst_3_T0}), .c ({new_AGEMA_signal_1610, SubCellInst_SboxInst_3_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_XOR12_U1 ( .a ({new_AGEMA_signal_1610, SubCellInst_SboxInst_3_L3}), .b ({new_AGEMA_signal_1558, SubCellInst_SboxInst_3_T2}), .c ({new_AGEMA_signal_1675, SubCellInst_SboxInst_3_YY_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_XOR13_U1 ( .a ({new_AGEMA_signal_1185, SubCellInst_SboxInst_3_XX_1_}), .b ({new_AGEMA_signal_1558, SubCellInst_SboxInst_3_T2}), .c ({new_AGEMA_signal_1611, SubCellInst_SboxInst_3_YY_0_}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_U3 ( .a ({new_AGEMA_signal_1679, SubCellInst_SboxInst_4_YY_1_}), .b ({new_AGEMA_signal_1732, ShiftRowsOutput[27]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_U2 ( .a ({new_AGEMA_signal_1615, SubCellInst_SboxInst_4_YY_0_}), .b ({new_AGEMA_signal_1676, ShiftRowsOutput[26]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_AND1_U1 ( .a ({new_AGEMA_signal_1189, SubCellInst_SboxInst_4_n3}), .b ({new_AGEMA_signal_1478, SubCellInst_SboxInst_4_Q1}), .clk (clk), .r (Fresh[8]), .c ({new_AGEMA_signal_1560, SubCellInst_SboxInst_4_T0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_XOR2_U1 ( .a ({new_AGEMA_signal_1477, SubCellInst_SboxInst_4_Q0}), .b ({new_AGEMA_signal_1560, SubCellInst_SboxInst_4_T0}), .c ({new_AGEMA_signal_1612, SubCellInst_SboxInst_4_Q2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_AND3_U1 ( .a ({new_AGEMA_signal_1189, SubCellInst_SboxInst_4_n3}), .b ({new_AGEMA_signal_1479, SubCellInst_SboxInst_4_Q4}), .clk (clk), .r (Fresh[9]), .c ({new_AGEMA_signal_1561, SubCellInst_SboxInst_4_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_XOR7_U1 ( .a ({new_AGEMA_signal_1562, SubCellInst_SboxInst_4_L1}), .b ({new_AGEMA_signal_1561, SubCellInst_SboxInst_4_T2}), .c ({new_AGEMA_signal_1613, SubCellInst_SboxInst_4_Q7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_XOR11_U1 ( .a ({new_AGEMA_signal_1193, SubCellInst_SboxInst_4_XX_2_}), .b ({new_AGEMA_signal_1560, SubCellInst_SboxInst_4_T0}), .c ({new_AGEMA_signal_1614, SubCellInst_SboxInst_4_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_XOR12_U1 ( .a ({new_AGEMA_signal_1614, SubCellInst_SboxInst_4_L3}), .b ({new_AGEMA_signal_1561, SubCellInst_SboxInst_4_T2}), .c ({new_AGEMA_signal_1679, SubCellInst_SboxInst_4_YY_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_XOR13_U1 ( .a ({new_AGEMA_signal_1191, SubCellInst_SboxInst_4_XX_1_}), .b ({new_AGEMA_signal_1561, SubCellInst_SboxInst_4_T2}), .c ({new_AGEMA_signal_1615, SubCellInst_SboxInst_4_YY_0_}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_U3 ( .a ({new_AGEMA_signal_1683, SubCellInst_SboxInst_5_YY_1_}), .b ({new_AGEMA_signal_1734, ShiftRowsOutput[31]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_U2 ( .a ({new_AGEMA_signal_1619, SubCellInst_SboxInst_5_YY_0_}), .b ({new_AGEMA_signal_1680, ShiftRowsOutput[30]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_AND1_U1 ( .a ({new_AGEMA_signal_1195, SubCellInst_SboxInst_5_n3}), .b ({new_AGEMA_signal_1484, SubCellInst_SboxInst_5_Q1}), .clk (clk), .r (Fresh[10]), .c ({new_AGEMA_signal_1563, SubCellInst_SboxInst_5_T0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_XOR2_U1 ( .a ({new_AGEMA_signal_1483, SubCellInst_SboxInst_5_Q0}), .b ({new_AGEMA_signal_1563, SubCellInst_SboxInst_5_T0}), .c ({new_AGEMA_signal_1616, SubCellInst_SboxInst_5_Q2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_AND3_U1 ( .a ({new_AGEMA_signal_1195, SubCellInst_SboxInst_5_n3}), .b ({new_AGEMA_signal_1485, SubCellInst_SboxInst_5_Q4}), .clk (clk), .r (Fresh[11]), .c ({new_AGEMA_signal_1564, SubCellInst_SboxInst_5_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_XOR7_U1 ( .a ({new_AGEMA_signal_1565, SubCellInst_SboxInst_5_L1}), .b ({new_AGEMA_signal_1564, SubCellInst_SboxInst_5_T2}), .c ({new_AGEMA_signal_1617, SubCellInst_SboxInst_5_Q7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_XOR11_U1 ( .a ({new_AGEMA_signal_1199, SubCellInst_SboxInst_5_XX_2_}), .b ({new_AGEMA_signal_1563, SubCellInst_SboxInst_5_T0}), .c ({new_AGEMA_signal_1618, SubCellInst_SboxInst_5_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_XOR12_U1 ( .a ({new_AGEMA_signal_1618, SubCellInst_SboxInst_5_L3}), .b ({new_AGEMA_signal_1564, SubCellInst_SboxInst_5_T2}), .c ({new_AGEMA_signal_1683, SubCellInst_SboxInst_5_YY_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_XOR13_U1 ( .a ({new_AGEMA_signal_1197, SubCellInst_SboxInst_5_XX_1_}), .b ({new_AGEMA_signal_1564, SubCellInst_SboxInst_5_T2}), .c ({new_AGEMA_signal_1619, SubCellInst_SboxInst_5_YY_0_}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_U3 ( .a ({new_AGEMA_signal_1687, SubCellInst_SboxInst_6_YY_1_}), .b ({new_AGEMA_signal_1736, ShiftRowsOutput[19]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_U2 ( .a ({new_AGEMA_signal_1623, SubCellInst_SboxInst_6_YY_0_}), .b ({new_AGEMA_signal_1684, ShiftRowsOutput[18]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_AND1_U1 ( .a ({new_AGEMA_signal_1201, SubCellInst_SboxInst_6_n3}), .b ({new_AGEMA_signal_1490, SubCellInst_SboxInst_6_Q1}), .clk (clk), .r (Fresh[12]), .c ({new_AGEMA_signal_1566, SubCellInst_SboxInst_6_T0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_XOR2_U1 ( .a ({new_AGEMA_signal_1489, SubCellInst_SboxInst_6_Q0}), .b ({new_AGEMA_signal_1566, SubCellInst_SboxInst_6_T0}), .c ({new_AGEMA_signal_1620, SubCellInst_SboxInst_6_Q2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_AND3_U1 ( .a ({new_AGEMA_signal_1201, SubCellInst_SboxInst_6_n3}), .b ({new_AGEMA_signal_1491, SubCellInst_SboxInst_6_Q4}), .clk (clk), .r (Fresh[13]), .c ({new_AGEMA_signal_1567, SubCellInst_SboxInst_6_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_XOR7_U1 ( .a ({new_AGEMA_signal_1568, SubCellInst_SboxInst_6_L1}), .b ({new_AGEMA_signal_1567, SubCellInst_SboxInst_6_T2}), .c ({new_AGEMA_signal_1621, SubCellInst_SboxInst_6_Q7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_XOR11_U1 ( .a ({new_AGEMA_signal_1205, SubCellInst_SboxInst_6_XX_2_}), .b ({new_AGEMA_signal_1566, SubCellInst_SboxInst_6_T0}), .c ({new_AGEMA_signal_1622, SubCellInst_SboxInst_6_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_XOR12_U1 ( .a ({new_AGEMA_signal_1622, SubCellInst_SboxInst_6_L3}), .b ({new_AGEMA_signal_1567, SubCellInst_SboxInst_6_T2}), .c ({new_AGEMA_signal_1687, SubCellInst_SboxInst_6_YY_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_XOR13_U1 ( .a ({new_AGEMA_signal_1203, SubCellInst_SboxInst_6_XX_1_}), .b ({new_AGEMA_signal_1567, SubCellInst_SboxInst_6_T2}), .c ({new_AGEMA_signal_1623, SubCellInst_SboxInst_6_YY_0_}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_U3 ( .a ({new_AGEMA_signal_1691, SubCellInst_SboxInst_7_YY_1_}), .b ({new_AGEMA_signal_1738, ShiftRowsOutput[23]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_U2 ( .a ({new_AGEMA_signal_1627, SubCellInst_SboxInst_7_YY_0_}), .b ({new_AGEMA_signal_1688, ShiftRowsOutput[22]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_AND1_U1 ( .a ({new_AGEMA_signal_1207, SubCellInst_SboxInst_7_n3}), .b ({new_AGEMA_signal_1496, SubCellInst_SboxInst_7_Q1}), .clk (clk), .r (Fresh[14]), .c ({new_AGEMA_signal_1569, SubCellInst_SboxInst_7_T0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_XOR2_U1 ( .a ({new_AGEMA_signal_1495, SubCellInst_SboxInst_7_Q0}), .b ({new_AGEMA_signal_1569, SubCellInst_SboxInst_7_T0}), .c ({new_AGEMA_signal_1624, SubCellInst_SboxInst_7_Q2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_AND3_U1 ( .a ({new_AGEMA_signal_1207, SubCellInst_SboxInst_7_n3}), .b ({new_AGEMA_signal_1497, SubCellInst_SboxInst_7_Q4}), .clk (clk), .r (Fresh[15]), .c ({new_AGEMA_signal_1570, SubCellInst_SboxInst_7_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_XOR7_U1 ( .a ({new_AGEMA_signal_1571, SubCellInst_SboxInst_7_L1}), .b ({new_AGEMA_signal_1570, SubCellInst_SboxInst_7_T2}), .c ({new_AGEMA_signal_1625, SubCellInst_SboxInst_7_Q7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_XOR11_U1 ( .a ({new_AGEMA_signal_1211, SubCellInst_SboxInst_7_XX_2_}), .b ({new_AGEMA_signal_1569, SubCellInst_SboxInst_7_T0}), .c ({new_AGEMA_signal_1626, SubCellInst_SboxInst_7_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_XOR12_U1 ( .a ({new_AGEMA_signal_1626, SubCellInst_SboxInst_7_L3}), .b ({new_AGEMA_signal_1570, SubCellInst_SboxInst_7_T2}), .c ({new_AGEMA_signal_1691, SubCellInst_SboxInst_7_YY_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_XOR13_U1 ( .a ({new_AGEMA_signal_1209, SubCellInst_SboxInst_7_XX_1_}), .b ({new_AGEMA_signal_1570, SubCellInst_SboxInst_7_T2}), .c ({new_AGEMA_signal_1627, SubCellInst_SboxInst_7_YY_0_}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_U3 ( .a ({new_AGEMA_signal_1695, SubCellInst_SboxInst_8_YY_1_}), .b ({new_AGEMA_signal_1740, AddRoundConstantOutput[35]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_U2 ( .a ({new_AGEMA_signal_1631, SubCellInst_SboxInst_8_YY_0_}), .b ({new_AGEMA_signal_1692, AddRoundConstantOutput[34]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_AND1_U1 ( .a ({new_AGEMA_signal_1213, SubCellInst_SboxInst_8_n3}), .b ({new_AGEMA_signal_1502, SubCellInst_SboxInst_8_Q1}), .clk (clk), .r (Fresh[16]), .c ({new_AGEMA_signal_1572, SubCellInst_SboxInst_8_T0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_XOR2_U1 ( .a ({new_AGEMA_signal_1501, SubCellInst_SboxInst_8_Q0}), .b ({new_AGEMA_signal_1572, SubCellInst_SboxInst_8_T0}), .c ({new_AGEMA_signal_1628, SubCellInst_SboxInst_8_Q2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_AND3_U1 ( .a ({new_AGEMA_signal_1213, SubCellInst_SboxInst_8_n3}), .b ({new_AGEMA_signal_1503, SubCellInst_SboxInst_8_Q4}), .clk (clk), .r (Fresh[17]), .c ({new_AGEMA_signal_1573, SubCellInst_SboxInst_8_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_XOR7_U1 ( .a ({new_AGEMA_signal_1574, SubCellInst_SboxInst_8_L1}), .b ({new_AGEMA_signal_1573, SubCellInst_SboxInst_8_T2}), .c ({new_AGEMA_signal_1629, SubCellInst_SboxInst_8_Q7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_XOR11_U1 ( .a ({new_AGEMA_signal_1217, SubCellInst_SboxInst_8_XX_2_}), .b ({new_AGEMA_signal_1572, SubCellInst_SboxInst_8_T0}), .c ({new_AGEMA_signal_1630, SubCellInst_SboxInst_8_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_XOR12_U1 ( .a ({new_AGEMA_signal_1630, SubCellInst_SboxInst_8_L3}), .b ({new_AGEMA_signal_1573, SubCellInst_SboxInst_8_T2}), .c ({new_AGEMA_signal_1695, SubCellInst_SboxInst_8_YY_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_XOR13_U1 ( .a ({new_AGEMA_signal_1215, SubCellInst_SboxInst_8_XX_1_}), .b ({new_AGEMA_signal_1573, SubCellInst_SboxInst_8_T2}), .c ({new_AGEMA_signal_1631, SubCellInst_SboxInst_8_YY_0_}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_U3 ( .a ({new_AGEMA_signal_1699, SubCellInst_SboxInst_9_YY_1_}), .b ({new_AGEMA_signal_1742, AddRoundConstantOutput[39]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_U2 ( .a ({new_AGEMA_signal_1635, SubCellInst_SboxInst_9_YY_0_}), .b ({new_AGEMA_signal_1696, AddRoundConstantOutput[38]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_AND1_U1 ( .a ({new_AGEMA_signal_1219, SubCellInst_SboxInst_9_n3}), .b ({new_AGEMA_signal_1508, SubCellInst_SboxInst_9_Q1}), .clk (clk), .r (Fresh[18]), .c ({new_AGEMA_signal_1575, SubCellInst_SboxInst_9_T0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_XOR2_U1 ( .a ({new_AGEMA_signal_1507, SubCellInst_SboxInst_9_Q0}), .b ({new_AGEMA_signal_1575, SubCellInst_SboxInst_9_T0}), .c ({new_AGEMA_signal_1632, SubCellInst_SboxInst_9_Q2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_AND3_U1 ( .a ({new_AGEMA_signal_1219, SubCellInst_SboxInst_9_n3}), .b ({new_AGEMA_signal_1509, SubCellInst_SboxInst_9_Q4}), .clk (clk), .r (Fresh[19]), .c ({new_AGEMA_signal_1576, SubCellInst_SboxInst_9_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_XOR7_U1 ( .a ({new_AGEMA_signal_1577, SubCellInst_SboxInst_9_L1}), .b ({new_AGEMA_signal_1576, SubCellInst_SboxInst_9_T2}), .c ({new_AGEMA_signal_1633, SubCellInst_SboxInst_9_Q7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_XOR11_U1 ( .a ({new_AGEMA_signal_1223, SubCellInst_SboxInst_9_XX_2_}), .b ({new_AGEMA_signal_1575, SubCellInst_SboxInst_9_T0}), .c ({new_AGEMA_signal_1634, SubCellInst_SboxInst_9_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_XOR12_U1 ( .a ({new_AGEMA_signal_1634, SubCellInst_SboxInst_9_L3}), .b ({new_AGEMA_signal_1576, SubCellInst_SboxInst_9_T2}), .c ({new_AGEMA_signal_1699, SubCellInst_SboxInst_9_YY_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_XOR13_U1 ( .a ({new_AGEMA_signal_1221, SubCellInst_SboxInst_9_XX_1_}), .b ({new_AGEMA_signal_1576, SubCellInst_SboxInst_9_T2}), .c ({new_AGEMA_signal_1635, SubCellInst_SboxInst_9_YY_0_}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_U3 ( .a ({new_AGEMA_signal_1703, SubCellInst_SboxInst_10_YY_1_}), .b ({new_AGEMA_signal_1744, AddRoundConstantOutput[43]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_U2 ( .a ({new_AGEMA_signal_1639, SubCellInst_SboxInst_10_YY_0_}), .b ({new_AGEMA_signal_1700, AddRoundConstantOutput[42]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_AND1_U1 ( .a ({new_AGEMA_signal_1225, SubCellInst_SboxInst_10_n3}), .b ({new_AGEMA_signal_1514, SubCellInst_SboxInst_10_Q1}), .clk (clk), .r (Fresh[20]), .c ({new_AGEMA_signal_1578, SubCellInst_SboxInst_10_T0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_XOR2_U1 ( .a ({new_AGEMA_signal_1513, SubCellInst_SboxInst_10_Q0}), .b ({new_AGEMA_signal_1578, SubCellInst_SboxInst_10_T0}), .c ({new_AGEMA_signal_1636, SubCellInst_SboxInst_10_Q2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_AND3_U1 ( .a ({new_AGEMA_signal_1225, SubCellInst_SboxInst_10_n3}), .b ({new_AGEMA_signal_1515, SubCellInst_SboxInst_10_Q4}), .clk (clk), .r (Fresh[21]), .c ({new_AGEMA_signal_1579, SubCellInst_SboxInst_10_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_XOR7_U1 ( .a ({new_AGEMA_signal_1580, SubCellInst_SboxInst_10_L1}), .b ({new_AGEMA_signal_1579, SubCellInst_SboxInst_10_T2}), .c ({new_AGEMA_signal_1637, SubCellInst_SboxInst_10_Q7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_XOR11_U1 ( .a ({new_AGEMA_signal_1229, SubCellInst_SboxInst_10_XX_2_}), .b ({new_AGEMA_signal_1578, SubCellInst_SboxInst_10_T0}), .c ({new_AGEMA_signal_1638, SubCellInst_SboxInst_10_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_XOR12_U1 ( .a ({new_AGEMA_signal_1638, SubCellInst_SboxInst_10_L3}), .b ({new_AGEMA_signal_1579, SubCellInst_SboxInst_10_T2}), .c ({new_AGEMA_signal_1703, SubCellInst_SboxInst_10_YY_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_XOR13_U1 ( .a ({new_AGEMA_signal_1227, SubCellInst_SboxInst_10_XX_1_}), .b ({new_AGEMA_signal_1579, SubCellInst_SboxInst_10_T2}), .c ({new_AGEMA_signal_1639, SubCellInst_SboxInst_10_YY_0_}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_U3 ( .a ({new_AGEMA_signal_1707, SubCellInst_SboxInst_11_YY_1_}), .b ({new_AGEMA_signal_1746, SubCellOutput[47]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_U2 ( .a ({new_AGEMA_signal_1643, SubCellInst_SboxInst_11_YY_0_}), .b ({new_AGEMA_signal_1704, SubCellOutput[46]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_AND1_U1 ( .a ({new_AGEMA_signal_1231, SubCellInst_SboxInst_11_n3}), .b ({new_AGEMA_signal_1520, SubCellInst_SboxInst_11_Q1}), .clk (clk), .r (Fresh[22]), .c ({new_AGEMA_signal_1581, SubCellInst_SboxInst_11_T0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_XOR2_U1 ( .a ({new_AGEMA_signal_1519, SubCellInst_SboxInst_11_Q0}), .b ({new_AGEMA_signal_1581, SubCellInst_SboxInst_11_T0}), .c ({new_AGEMA_signal_1640, SubCellInst_SboxInst_11_Q2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_AND3_U1 ( .a ({new_AGEMA_signal_1231, SubCellInst_SboxInst_11_n3}), .b ({new_AGEMA_signal_1521, SubCellInst_SboxInst_11_Q4}), .clk (clk), .r (Fresh[23]), .c ({new_AGEMA_signal_1582, SubCellInst_SboxInst_11_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_XOR7_U1 ( .a ({new_AGEMA_signal_1583, SubCellInst_SboxInst_11_L1}), .b ({new_AGEMA_signal_1582, SubCellInst_SboxInst_11_T2}), .c ({new_AGEMA_signal_1641, SubCellInst_SboxInst_11_Q7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_XOR11_U1 ( .a ({new_AGEMA_signal_1235, SubCellInst_SboxInst_11_XX_2_}), .b ({new_AGEMA_signal_1581, SubCellInst_SboxInst_11_T0}), .c ({new_AGEMA_signal_1642, SubCellInst_SboxInst_11_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_XOR12_U1 ( .a ({new_AGEMA_signal_1642, SubCellInst_SboxInst_11_L3}), .b ({new_AGEMA_signal_1582, SubCellInst_SboxInst_11_T2}), .c ({new_AGEMA_signal_1707, SubCellInst_SboxInst_11_YY_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_XOR13_U1 ( .a ({new_AGEMA_signal_1233, SubCellInst_SboxInst_11_XX_1_}), .b ({new_AGEMA_signal_1582, SubCellInst_SboxInst_11_T2}), .c ({new_AGEMA_signal_1643, SubCellInst_SboxInst_11_YY_0_}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_U3 ( .a ({new_AGEMA_signal_1711, SubCellInst_SboxInst_12_YY_1_}), .b ({new_AGEMA_signal_1748, AddRoundConstantOutput[51]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_U2 ( .a ({new_AGEMA_signal_1647, SubCellInst_SboxInst_12_YY_0_}), .b ({new_AGEMA_signal_1708, AddRoundConstantOutput[50]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_AND1_U1 ( .a ({new_AGEMA_signal_1237, SubCellInst_SboxInst_12_n3}), .b ({new_AGEMA_signal_1526, SubCellInst_SboxInst_12_Q1}), .clk (clk), .r (Fresh[24]), .c ({new_AGEMA_signal_1584, SubCellInst_SboxInst_12_T0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_XOR2_U1 ( .a ({new_AGEMA_signal_1525, SubCellInst_SboxInst_12_Q0}), .b ({new_AGEMA_signal_1584, SubCellInst_SboxInst_12_T0}), .c ({new_AGEMA_signal_1644, SubCellInst_SboxInst_12_Q2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_AND3_U1 ( .a ({new_AGEMA_signal_1237, SubCellInst_SboxInst_12_n3}), .b ({new_AGEMA_signal_1527, SubCellInst_SboxInst_12_Q4}), .clk (clk), .r (Fresh[25]), .c ({new_AGEMA_signal_1585, SubCellInst_SboxInst_12_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_XOR7_U1 ( .a ({new_AGEMA_signal_1586, SubCellInst_SboxInst_12_L1}), .b ({new_AGEMA_signal_1585, SubCellInst_SboxInst_12_T2}), .c ({new_AGEMA_signal_1645, SubCellInst_SboxInst_12_Q7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_XOR11_U1 ( .a ({new_AGEMA_signal_1241, SubCellInst_SboxInst_12_XX_2_}), .b ({new_AGEMA_signal_1584, SubCellInst_SboxInst_12_T0}), .c ({new_AGEMA_signal_1646, SubCellInst_SboxInst_12_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_XOR12_U1 ( .a ({new_AGEMA_signal_1646, SubCellInst_SboxInst_12_L3}), .b ({new_AGEMA_signal_1585, SubCellInst_SboxInst_12_T2}), .c ({new_AGEMA_signal_1711, SubCellInst_SboxInst_12_YY_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_XOR13_U1 ( .a ({new_AGEMA_signal_1239, SubCellInst_SboxInst_12_XX_1_}), .b ({new_AGEMA_signal_1585, SubCellInst_SboxInst_12_T2}), .c ({new_AGEMA_signal_1647, SubCellInst_SboxInst_12_YY_0_}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_U3 ( .a ({new_AGEMA_signal_1715, SubCellInst_SboxInst_13_YY_1_}), .b ({new_AGEMA_signal_1750, AddRoundConstantOutput[55]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_U2 ( .a ({new_AGEMA_signal_1651, SubCellInst_SboxInst_13_YY_0_}), .b ({new_AGEMA_signal_1712, AddRoundConstantOutput[54]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_AND1_U1 ( .a ({new_AGEMA_signal_1243, SubCellInst_SboxInst_13_n3}), .b ({new_AGEMA_signal_1532, SubCellInst_SboxInst_13_Q1}), .clk (clk), .r (Fresh[26]), .c ({new_AGEMA_signal_1587, SubCellInst_SboxInst_13_T0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_XOR2_U1 ( .a ({new_AGEMA_signal_1531, SubCellInst_SboxInst_13_Q0}), .b ({new_AGEMA_signal_1587, SubCellInst_SboxInst_13_T0}), .c ({new_AGEMA_signal_1648, SubCellInst_SboxInst_13_Q2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_AND3_U1 ( .a ({new_AGEMA_signal_1243, SubCellInst_SboxInst_13_n3}), .b ({new_AGEMA_signal_1533, SubCellInst_SboxInst_13_Q4}), .clk (clk), .r (Fresh[27]), .c ({new_AGEMA_signal_1588, SubCellInst_SboxInst_13_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_XOR7_U1 ( .a ({new_AGEMA_signal_1589, SubCellInst_SboxInst_13_L1}), .b ({new_AGEMA_signal_1588, SubCellInst_SboxInst_13_T2}), .c ({new_AGEMA_signal_1649, SubCellInst_SboxInst_13_Q7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_XOR11_U1 ( .a ({new_AGEMA_signal_1247, SubCellInst_SboxInst_13_XX_2_}), .b ({new_AGEMA_signal_1587, SubCellInst_SboxInst_13_T0}), .c ({new_AGEMA_signal_1650, SubCellInst_SboxInst_13_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_XOR12_U1 ( .a ({new_AGEMA_signal_1650, SubCellInst_SboxInst_13_L3}), .b ({new_AGEMA_signal_1588, SubCellInst_SboxInst_13_T2}), .c ({new_AGEMA_signal_1715, SubCellInst_SboxInst_13_YY_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_XOR13_U1 ( .a ({new_AGEMA_signal_1245, SubCellInst_SboxInst_13_XX_1_}), .b ({new_AGEMA_signal_1588, SubCellInst_SboxInst_13_T2}), .c ({new_AGEMA_signal_1651, SubCellInst_SboxInst_13_YY_0_}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_U3 ( .a ({new_AGEMA_signal_1719, SubCellInst_SboxInst_14_YY_1_}), .b ({new_AGEMA_signal_1752, AddRoundConstantOutput[59]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_U2 ( .a ({new_AGEMA_signal_1655, SubCellInst_SboxInst_14_YY_0_}), .b ({new_AGEMA_signal_1716, AddRoundConstantOutput[58]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_AND1_U1 ( .a ({new_AGEMA_signal_1249, SubCellInst_SboxInst_14_n3}), .b ({new_AGEMA_signal_1538, SubCellInst_SboxInst_14_Q1}), .clk (clk), .r (Fresh[28]), .c ({new_AGEMA_signal_1590, SubCellInst_SboxInst_14_T0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_XOR2_U1 ( .a ({new_AGEMA_signal_1537, SubCellInst_SboxInst_14_Q0}), .b ({new_AGEMA_signal_1590, SubCellInst_SboxInst_14_T0}), .c ({new_AGEMA_signal_1652, SubCellInst_SboxInst_14_Q2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_AND3_U1 ( .a ({new_AGEMA_signal_1249, SubCellInst_SboxInst_14_n3}), .b ({new_AGEMA_signal_1539, SubCellInst_SboxInst_14_Q4}), .clk (clk), .r (Fresh[29]), .c ({new_AGEMA_signal_1591, SubCellInst_SboxInst_14_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_XOR7_U1 ( .a ({new_AGEMA_signal_1592, SubCellInst_SboxInst_14_L1}), .b ({new_AGEMA_signal_1591, SubCellInst_SboxInst_14_T2}), .c ({new_AGEMA_signal_1653, SubCellInst_SboxInst_14_Q7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_XOR11_U1 ( .a ({new_AGEMA_signal_1253, SubCellInst_SboxInst_14_XX_2_}), .b ({new_AGEMA_signal_1590, SubCellInst_SboxInst_14_T0}), .c ({new_AGEMA_signal_1654, SubCellInst_SboxInst_14_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_XOR12_U1 ( .a ({new_AGEMA_signal_1654, SubCellInst_SboxInst_14_L3}), .b ({new_AGEMA_signal_1591, SubCellInst_SboxInst_14_T2}), .c ({new_AGEMA_signal_1719, SubCellInst_SboxInst_14_YY_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_XOR13_U1 ( .a ({new_AGEMA_signal_1251, SubCellInst_SboxInst_14_XX_1_}), .b ({new_AGEMA_signal_1591, SubCellInst_SboxInst_14_T2}), .c ({new_AGEMA_signal_1655, SubCellInst_SboxInst_14_YY_0_}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_U3 ( .a ({new_AGEMA_signal_1723, SubCellInst_SboxInst_15_YY_1_}), .b ({new_AGEMA_signal_1754, SubCellOutput[63]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_U2 ( .a ({new_AGEMA_signal_1659, SubCellInst_SboxInst_15_YY_0_}), .b ({new_AGEMA_signal_1720, SubCellOutput[62]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_AND1_U1 ( .a ({new_AGEMA_signal_1255, SubCellInst_SboxInst_15_n3}), .b ({new_AGEMA_signal_1544, SubCellInst_SboxInst_15_Q1}), .clk (clk), .r (Fresh[30]), .c ({new_AGEMA_signal_1593, SubCellInst_SboxInst_15_T0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_XOR2_U1 ( .a ({new_AGEMA_signal_1543, SubCellInst_SboxInst_15_Q0}), .b ({new_AGEMA_signal_1593, SubCellInst_SboxInst_15_T0}), .c ({new_AGEMA_signal_1656, SubCellInst_SboxInst_15_Q2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_AND3_U1 ( .a ({new_AGEMA_signal_1255, SubCellInst_SboxInst_15_n3}), .b ({new_AGEMA_signal_1545, SubCellInst_SboxInst_15_Q4}), .clk (clk), .r (Fresh[31]), .c ({new_AGEMA_signal_1594, SubCellInst_SboxInst_15_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_XOR7_U1 ( .a ({new_AGEMA_signal_1595, SubCellInst_SboxInst_15_L1}), .b ({new_AGEMA_signal_1594, SubCellInst_SboxInst_15_T2}), .c ({new_AGEMA_signal_1657, SubCellInst_SboxInst_15_Q7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_XOR11_U1 ( .a ({new_AGEMA_signal_1259, SubCellInst_SboxInst_15_XX_2_}), .b ({new_AGEMA_signal_1593, SubCellInst_SboxInst_15_T0}), .c ({new_AGEMA_signal_1658, SubCellInst_SboxInst_15_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_XOR12_U1 ( .a ({new_AGEMA_signal_1658, SubCellInst_SboxInst_15_L3}), .b ({new_AGEMA_signal_1594, SubCellInst_SboxInst_15_T2}), .c ({new_AGEMA_signal_1723, SubCellInst_SboxInst_15_YY_1_}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_XOR13_U1 ( .a ({new_AGEMA_signal_1257, SubCellInst_SboxInst_15_XX_1_}), .b ({new_AGEMA_signal_1594, SubCellInst_SboxInst_15_T2}), .c ({new_AGEMA_signal_1659, SubCellInst_SboxInst_15_YY_0_}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_1756, AddConstXOR_AddConstXOR_XORInst_0_2_n1}), .b ({1'b0, FSMUpdate[3]}), .c ({new_AGEMA_signal_1800, AddRoundConstantOutput[62]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1720, SubCellOutput[62]}), .c ({new_AGEMA_signal_1756, AddConstXOR_AddConstXOR_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_1801, AddConstXOR_AddConstXOR_XORInst_0_3_n1}), .b ({1'b0, FSMUpdate[4]}), .c ({new_AGEMA_signal_1843, AddRoundConstantOutput[63]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1754, SubCellOutput[63]}), .c ({new_AGEMA_signal_1801, AddConstXOR_AddConstXOR_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_1757, AddConstXOR_AddConstXOR_XORInst_1_2_n1}), .b ({1'b0, 1'b0}), .c ({new_AGEMA_signal_1802, AddRoundConstantOutput[46]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1704, SubCellOutput[46]}), .c ({new_AGEMA_signal_1757, AddConstXOR_AddConstXOR_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_1803, AddConstXOR_AddConstXOR_XORInst_1_3_n1}), .b ({1'b0, 1'b0}), .c ({new_AGEMA_signal_1845, AddRoundConstantOutput[47]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1746, SubCellOutput[47]}), .c ({new_AGEMA_signal_1803, AddConstXOR_AddConstXOR_XORInst_1_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_1758, AddRoundTweakeyXOR_XORInst_0_2_n1}), .b ({new_AGEMA_signal_1266, TweakeyGeneration_key_Feedback[2]}), .c ({new_AGEMA_signal_1804, ShiftRowsOutput[46]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1692, AddRoundConstantOutput[34]}), .c ({new_AGEMA_signal_1758, AddRoundTweakeyXOR_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_1805, AddRoundTweakeyXOR_XORInst_0_3_n1}), .b ({new_AGEMA_signal_1269, TweakeyGeneration_key_Feedback[3]}), .c ({new_AGEMA_signal_1847, ShiftRowsOutput[47]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1740, AddRoundConstantOutput[35]}), .c ({new_AGEMA_signal_1805, AddRoundTweakeyXOR_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_1759, AddRoundTweakeyXOR_XORInst_1_2_n1}), .b ({new_AGEMA_signal_1278, TweakeyGeneration_key_Feedback[6]}), .c ({new_AGEMA_signal_1806, ShiftRowsOutput[34]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1696, AddRoundConstantOutput[38]}), .c ({new_AGEMA_signal_1759, AddRoundTweakeyXOR_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_1807, AddRoundTweakeyXOR_XORInst_1_3_n1}), .b ({new_AGEMA_signal_1281, TweakeyGeneration_key_Feedback[7]}), .c ({new_AGEMA_signal_1849, ShiftRowsOutput[35]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1742, AddRoundConstantOutput[39]}), .c ({new_AGEMA_signal_1807, AddRoundTweakeyXOR_XORInst_1_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_1760, AddRoundTweakeyXOR_XORInst_2_2_n1}), .b ({new_AGEMA_signal_1290, TweakeyGeneration_key_Feedback[10]}), .c ({new_AGEMA_signal_1808, ShiftRowsOutput[38]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1700, AddRoundConstantOutput[42]}), .c ({new_AGEMA_signal_1760, AddRoundTweakeyXOR_XORInst_2_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_1809, AddRoundTweakeyXOR_XORInst_2_3_n1}), .b ({new_AGEMA_signal_1293, TweakeyGeneration_key_Feedback[11]}), .c ({new_AGEMA_signal_1851, ShiftRowsOutput[39]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1744, AddRoundConstantOutput[43]}), .c ({new_AGEMA_signal_1809, AddRoundTweakeyXOR_XORInst_2_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_1852, AddRoundTweakeyXOR_XORInst_3_2_n1}), .b ({new_AGEMA_signal_1302, TweakeyGeneration_key_Feedback[14]}), .c ({new_AGEMA_signal_1890, ShiftRowsOutput[42]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1802, AddRoundConstantOutput[46]}), .c ({new_AGEMA_signal_1852, AddRoundTweakeyXOR_XORInst_3_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_1891, AddRoundTweakeyXOR_XORInst_3_3_n1}), .b ({new_AGEMA_signal_1305, TweakeyGeneration_key_Feedback[15]}), .c ({new_AGEMA_signal_1953, ShiftRowsOutput[43]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1845, AddRoundConstantOutput[47]}), .c ({new_AGEMA_signal_1891, AddRoundTweakeyXOR_XORInst_3_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_2_U2 ( .a ({new_AGEMA_signal_1761, AddRoundTweakeyXOR_XORInst_4_2_n1}), .b ({new_AGEMA_signal_1314, TweakeyGeneration_key_Feedback[18]}), .c ({new_AGEMA_signal_1810, MCOutput[34]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1708, AddRoundConstantOutput[50]}), .c ({new_AGEMA_signal_1761, AddRoundTweakeyXOR_XORInst_4_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_3_U2 ( .a ({new_AGEMA_signal_1811, AddRoundTweakeyXOR_XORInst_4_3_n1}), .b ({new_AGEMA_signal_1317, TweakeyGeneration_key_Feedback[19]}), .c ({new_AGEMA_signal_1854, MCOutput[35]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1748, AddRoundConstantOutput[51]}), .c ({new_AGEMA_signal_1811, AddRoundTweakeyXOR_XORInst_4_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_2_U2 ( .a ({new_AGEMA_signal_1762, AddRoundTweakeyXOR_XORInst_5_2_n1}), .b ({new_AGEMA_signal_1326, TweakeyGeneration_key_Feedback[22]}), .c ({new_AGEMA_signal_1812, MCOutput[38]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1712, AddRoundConstantOutput[54]}), .c ({new_AGEMA_signal_1762, AddRoundTweakeyXOR_XORInst_5_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_3_U2 ( .a ({new_AGEMA_signal_1813, AddRoundTweakeyXOR_XORInst_5_3_n1}), .b ({new_AGEMA_signal_1329, TweakeyGeneration_key_Feedback[23]}), .c ({new_AGEMA_signal_1856, MCOutput[39]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1750, AddRoundConstantOutput[55]}), .c ({new_AGEMA_signal_1813, AddRoundTweakeyXOR_XORInst_5_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_2_U2 ( .a ({new_AGEMA_signal_1763, AddRoundTweakeyXOR_XORInst_6_2_n1}), .b ({new_AGEMA_signal_1338, TweakeyGeneration_key_Feedback[26]}), .c ({new_AGEMA_signal_1814, MCOutput[42]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1716, AddRoundConstantOutput[58]}), .c ({new_AGEMA_signal_1763, AddRoundTweakeyXOR_XORInst_6_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_3_U2 ( .a ({new_AGEMA_signal_1815, AddRoundTweakeyXOR_XORInst_6_3_n1}), .b ({new_AGEMA_signal_1341, TweakeyGeneration_key_Feedback[27]}), .c ({new_AGEMA_signal_1858, MCOutput[43]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1752, AddRoundConstantOutput[59]}), .c ({new_AGEMA_signal_1815, AddRoundTweakeyXOR_XORInst_6_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_2_U2 ( .a ({new_AGEMA_signal_1859, AddRoundTweakeyXOR_XORInst_7_2_n1}), .b ({new_AGEMA_signal_1350, TweakeyGeneration_key_Feedback[30]}), .c ({new_AGEMA_signal_1898, MCOutput[46]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1800, AddRoundConstantOutput[62]}), .c ({new_AGEMA_signal_1859, AddRoundTweakeyXOR_XORInst_7_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_3_U2 ( .a ({new_AGEMA_signal_1899, AddRoundTweakeyXOR_XORInst_7_3_n1}), .b ({new_AGEMA_signal_1353, TweakeyGeneration_key_Feedback[31]}), .c ({new_AGEMA_signal_1958, MCOutput[47]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1843, AddRoundConstantOutput[63]}), .c ({new_AGEMA_signal_1899, AddRoundTweakeyXOR_XORInst_7_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_0_2_U3 ( .a ({new_AGEMA_signal_1861, MCInst_MCR0_XORInst_0_2_n2}), .b ({new_AGEMA_signal_1764, MCInst_MCR0_XORInst_0_2_n1}), .c ({new_AGEMA_signal_1901, MCOutput[50]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_1684, ShiftRowsOutput[18]}), .b ({new_AGEMA_signal_1672, ShiftRowsOutput[2]}), .c ({new_AGEMA_signal_1764, MCInst_MCR0_XORInst_0_2_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_0_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1810, MCOutput[34]}), .c ({new_AGEMA_signal_1861, MCInst_MCR0_XORInst_0_2_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_0_3_U3 ( .a ({new_AGEMA_signal_1902, MCInst_MCR0_XORInst_0_3_n2}), .b ({new_AGEMA_signal_1816, MCInst_MCR0_XORInst_0_3_n1}), .c ({new_AGEMA_signal_1960, MCOutput[51]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_1736, ShiftRowsOutput[19]}), .b ({new_AGEMA_signal_1730, ShiftRowsOutput[3]}), .c ({new_AGEMA_signal_1816, MCInst_MCR0_XORInst_0_3_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_0_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1854, MCOutput[35]}), .c ({new_AGEMA_signal_1902, MCInst_MCR0_XORInst_0_3_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_1_2_U3 ( .a ({new_AGEMA_signal_1863, MCInst_MCR0_XORInst_1_2_n2}), .b ({new_AGEMA_signal_1765, MCInst_MCR0_XORInst_1_2_n1}), .c ({new_AGEMA_signal_1903, MCOutput[54]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_1688, ShiftRowsOutput[22]}), .b ({new_AGEMA_signal_1660, ShiftRowsOutput[6]}), .c ({new_AGEMA_signal_1765, MCInst_MCR0_XORInst_1_2_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_1_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1812, MCOutput[38]}), .c ({new_AGEMA_signal_1863, MCInst_MCR0_XORInst_1_2_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_1_3_U3 ( .a ({new_AGEMA_signal_1904, MCInst_MCR0_XORInst_1_3_n2}), .b ({new_AGEMA_signal_1817, MCInst_MCR0_XORInst_1_3_n1}), .c ({new_AGEMA_signal_1963, MCOutput[55]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_1738, ShiftRowsOutput[23]}), .b ({new_AGEMA_signal_1724, ShiftRowsOutput[7]}), .c ({new_AGEMA_signal_1817, MCInst_MCR0_XORInst_1_3_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_1_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1856, MCOutput[39]}), .c ({new_AGEMA_signal_1904, MCInst_MCR0_XORInst_1_3_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_2_2_U3 ( .a ({new_AGEMA_signal_1865, MCInst_MCR0_XORInst_2_2_n2}), .b ({new_AGEMA_signal_1766, MCInst_MCR0_XORInst_2_2_n1}), .c ({new_AGEMA_signal_1906, MCOutput[58]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_1676, ShiftRowsOutput[26]}), .b ({new_AGEMA_signal_1664, ShiftRowsOutput[10]}), .c ({new_AGEMA_signal_1766, MCInst_MCR0_XORInst_2_2_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_2_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1814, MCOutput[42]}), .c ({new_AGEMA_signal_1865, MCInst_MCR0_XORInst_2_2_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_2_3_U3 ( .a ({new_AGEMA_signal_1907, MCInst_MCR0_XORInst_2_3_n2}), .b ({new_AGEMA_signal_1818, MCInst_MCR0_XORInst_2_3_n1}), .c ({new_AGEMA_signal_1965, MCOutput[59]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_1732, ShiftRowsOutput[27]}), .b ({new_AGEMA_signal_1726, ShiftRowsOutput[11]}), .c ({new_AGEMA_signal_1818, MCInst_MCR0_XORInst_2_3_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_2_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1858, MCOutput[43]}), .c ({new_AGEMA_signal_1907, MCInst_MCR0_XORInst_2_3_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_3_2_U3 ( .a ({new_AGEMA_signal_1966, MCInst_MCR0_XORInst_3_2_n2}), .b ({new_AGEMA_signal_1767, MCInst_MCR0_XORInst_3_2_n1}), .c ({new_AGEMA_signal_2017, MCOutput[62]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_1680, ShiftRowsOutput[30]}), .b ({new_AGEMA_signal_1668, ShiftRowsOutput[14]}), .c ({new_AGEMA_signal_1767, MCInst_MCR0_XORInst_3_2_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_3_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1898, MCOutput[46]}), .c ({new_AGEMA_signal_1966, MCInst_MCR0_XORInst_3_2_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_3_3_U3 ( .a ({new_AGEMA_signal_2018, MCInst_MCR0_XORInst_3_3_n2}), .b ({new_AGEMA_signal_1819, MCInst_MCR0_XORInst_3_3_n1}), .c ({new_AGEMA_signal_2067, MCOutput[63]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_1734, ShiftRowsOutput[31]}), .b ({new_AGEMA_signal_1728, ShiftRowsOutput[15]}), .c ({new_AGEMA_signal_1819, MCInst_MCR0_XORInst_3_3_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_3_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1958, MCOutput[47]}), .c ({new_AGEMA_signal_2018, MCInst_MCR0_XORInst_3_3_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_1867, MCInst_MCR2_XORInst_0_2_n1}), .b ({new_AGEMA_signal_1684, ShiftRowsOutput[18]}), .c ({new_AGEMA_signal_1909, MCOutput[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_0_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1806, ShiftRowsOutput[34]}), .c ({new_AGEMA_signal_1867, MCInst_MCR2_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_1910, MCInst_MCR2_XORInst_0_3_n1}), .b ({new_AGEMA_signal_1736, ShiftRowsOutput[19]}), .c ({new_AGEMA_signal_1968, MCOutput[19]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_0_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1849, ShiftRowsOutput[35]}), .c ({new_AGEMA_signal_1910, MCInst_MCR2_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_1868, MCInst_MCR2_XORInst_1_2_n1}), .b ({new_AGEMA_signal_1688, ShiftRowsOutput[22]}), .c ({new_AGEMA_signal_1911, MCOutput[22]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_1_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1808, ShiftRowsOutput[38]}), .c ({new_AGEMA_signal_1868, MCInst_MCR2_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_1912, MCInst_MCR2_XORInst_1_3_n1}), .b ({new_AGEMA_signal_1738, ShiftRowsOutput[23]}), .c ({new_AGEMA_signal_1970, MCOutput[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_1_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1851, ShiftRowsOutput[39]}), .c ({new_AGEMA_signal_1912, MCInst_MCR2_XORInst_1_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_1971, MCInst_MCR2_XORInst_2_2_n1}), .b ({new_AGEMA_signal_1676, ShiftRowsOutput[26]}), .c ({new_AGEMA_signal_2023, MCOutput[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_2_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1890, ShiftRowsOutput[42]}), .c ({new_AGEMA_signal_1971, MCInst_MCR2_XORInst_2_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_2024, MCInst_MCR2_XORInst_2_3_n1}), .b ({new_AGEMA_signal_1732, ShiftRowsOutput[27]}), .c ({new_AGEMA_signal_2071, MCOutput[27]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_2_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1953, ShiftRowsOutput[43]}), .c ({new_AGEMA_signal_2024, MCInst_MCR2_XORInst_2_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_1869, MCInst_MCR2_XORInst_3_2_n1}), .b ({new_AGEMA_signal_1680, ShiftRowsOutput[30]}), .c ({new_AGEMA_signal_1913, MCOutput[30]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_3_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1804, ShiftRowsOutput[46]}), .c ({new_AGEMA_signal_1869, MCInst_MCR2_XORInst_3_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_1914, MCInst_MCR2_XORInst_3_3_n1}), .b ({new_AGEMA_signal_1734, ShiftRowsOutput[31]}), .c ({new_AGEMA_signal_1973, MCOutput[31]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_3_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1847, ShiftRowsOutput[47]}), .c ({new_AGEMA_signal_1914, MCInst_MCR2_XORInst_3_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_1870, MCInst_MCR3_XORInst_0_2_n1}), .b ({new_AGEMA_signal_1684, ShiftRowsOutput[18]}), .c ({new_AGEMA_signal_1915, MCOutput[2]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_0_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1810, MCOutput[34]}), .c ({new_AGEMA_signal_1870, MCInst_MCR3_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_1916, MCInst_MCR3_XORInst_0_3_n1}), .b ({new_AGEMA_signal_1736, ShiftRowsOutput[19]}), .c ({new_AGEMA_signal_1975, MCOutput[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_0_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1854, MCOutput[35]}), .c ({new_AGEMA_signal_1916, MCInst_MCR3_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_1871, MCInst_MCR3_XORInst_1_2_n1}), .b ({new_AGEMA_signal_1688, ShiftRowsOutput[22]}), .c ({new_AGEMA_signal_1917, MCOutput[6]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_1_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1812, MCOutput[38]}), .c ({new_AGEMA_signal_1871, MCInst_MCR3_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_1918, MCInst_MCR3_XORInst_1_3_n1}), .b ({new_AGEMA_signal_1738, ShiftRowsOutput[23]}), .c ({new_AGEMA_signal_1977, MCOutput[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_1_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1856, MCOutput[39]}), .c ({new_AGEMA_signal_1918, MCInst_MCR3_XORInst_1_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_1872, MCInst_MCR3_XORInst_2_2_n1}), .b ({new_AGEMA_signal_1676, ShiftRowsOutput[26]}), .c ({new_AGEMA_signal_1919, MCOutput[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_2_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1814, MCOutput[42]}), .c ({new_AGEMA_signal_1872, MCInst_MCR3_XORInst_2_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_1920, MCInst_MCR3_XORInst_2_3_n1}), .b ({new_AGEMA_signal_1732, ShiftRowsOutput[27]}), .c ({new_AGEMA_signal_1979, MCOutput[11]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_2_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1858, MCOutput[43]}), .c ({new_AGEMA_signal_1920, MCInst_MCR3_XORInst_2_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_1980, MCInst_MCR3_XORInst_3_2_n1}), .b ({new_AGEMA_signal_1680, ShiftRowsOutput[30]}), .c ({new_AGEMA_signal_2033, MCOutput[14]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_3_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1898, MCOutput[46]}), .c ({new_AGEMA_signal_1980, MCInst_MCR3_XORInst_3_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_2034, MCInst_MCR3_XORInst_3_3_n1}), .b ({new_AGEMA_signal_1734, ShiftRowsOutput[31]}), .c ({new_AGEMA_signal_2077, MCOutput[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_3_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1958, MCOutput[47]}), .c ({new_AGEMA_signal_2034, MCInst_MCR3_XORInst_3_3_n1}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_0_U1 ( .s (rst), .b ({new_AGEMA_signal_2027, MCOutput[0]}), .a ({Plaintext_s1[0], Plaintext_s0[0]}), .c ({new_AGEMA_signal_2036, StateRegInput[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_1_U1 ( .s (rst), .b ({new_AGEMA_signal_2073, MCOutput[1]}), .a ({Plaintext_s1[1], Plaintext_s0[1]}), .c ({new_AGEMA_signal_2079, StateRegInput[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_4_U1 ( .s (rst), .b ({new_AGEMA_signal_2029, MCOutput[4]}), .a ({Plaintext_s1[4], Plaintext_s0[4]}), .c ({new_AGEMA_signal_2038, StateRegInput[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_5_U1 ( .s (rst), .b ({new_AGEMA_signal_2074, MCOutput[5]}), .a ({Plaintext_s1[5], Plaintext_s0[5]}), .c ({new_AGEMA_signal_2081, StateRegInput[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_8_U1 ( .s (rst), .b ({new_AGEMA_signal_2031, MCOutput[8]}), .a ({Plaintext_s1[8], Plaintext_s0[8]}), .c ({new_AGEMA_signal_2040, StateRegInput[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_9_U1 ( .s (rst), .b ({new_AGEMA_signal_2075, MCOutput[9]}), .a ({Plaintext_s1[9], Plaintext_s0[9]}), .c ({new_AGEMA_signal_2083, StateRegInput[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_12_U1 ( .s (rst), .b ({new_AGEMA_signal_2108, MCOutput[12]}), .a ({Plaintext_s1[12], Plaintext_s0[12]}), .c ({new_AGEMA_signal_2111, StateRegInput[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_13_U1 ( .s (rst), .b ({new_AGEMA_signal_2118, MCOutput[13]}), .a ({Plaintext_s1[13], Plaintext_s0[13]}), .c ({new_AGEMA_signal_2120, StateRegInput[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_16_U1 ( .s (rst), .b ({new_AGEMA_signal_2019, MCOutput[16]}), .a ({Plaintext_s1[16], Plaintext_s0[16]}), .c ({new_AGEMA_signal_2044, StateRegInput[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_17_U1 ( .s (rst), .b ({new_AGEMA_signal_2068, MCOutput[17]}), .a ({Plaintext_s1[17], Plaintext_s0[17]}), .c ({new_AGEMA_signal_2087, StateRegInput[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_20_U1 ( .s (rst), .b ({new_AGEMA_signal_2021, MCOutput[20]}), .a ({Plaintext_s1[20], Plaintext_s0[20]}), .c ({new_AGEMA_signal_2046, StateRegInput[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_21_U1 ( .s (rst), .b ({new_AGEMA_signal_2069, MCOutput[21]}), .a ({Plaintext_s1[21], Plaintext_s0[21]}), .c ({new_AGEMA_signal_2089, StateRegInput[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_24_U1 ( .s (rst), .b ({new_AGEMA_signal_2106, MCOutput[24]}), .a ({Plaintext_s1[24], Plaintext_s0[24]}), .c ({new_AGEMA_signal_2113, StateRegInput[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_25_U1 ( .s (rst), .b ({new_AGEMA_signal_2117, MCOutput[25]}), .a ({Plaintext_s1[25], Plaintext_s0[25]}), .c ({new_AGEMA_signal_2122, StateRegInput[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_28_U1 ( .s (rst), .b ({new_AGEMA_signal_2025, MCOutput[28]}), .a ({Plaintext_s1[28], Plaintext_s0[28]}), .c ({new_AGEMA_signal_2050, StateRegInput[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_29_U1 ( .s (rst), .b ({new_AGEMA_signal_2072, MCOutput[29]}), .a ({Plaintext_s1[29], Plaintext_s0[29]}), .c ({new_AGEMA_signal_2093, StateRegInput[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_32_U1 ( .s (rst), .b ({new_AGEMA_signal_1892, MCOutput[32]}), .a ({Plaintext_s1[32], Plaintext_s0[32]}), .c ({new_AGEMA_signal_1934, StateRegInput[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_33_U1 ( .s (rst), .b ({new_AGEMA_signal_1954, MCOutput[33]}), .a ({Plaintext_s1[33], Plaintext_s0[33]}), .c ({new_AGEMA_signal_1994, StateRegInput[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_36_U1 ( .s (rst), .b ({new_AGEMA_signal_1894, MCOutput[36]}), .a ({Plaintext_s1[36], Plaintext_s0[36]}), .c ({new_AGEMA_signal_1936, StateRegInput[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_37_U1 ( .s (rst), .b ({new_AGEMA_signal_1955, MCOutput[37]}), .a ({Plaintext_s1[37], Plaintext_s0[37]}), .c ({new_AGEMA_signal_1996, StateRegInput[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_40_U1 ( .s (rst), .b ({new_AGEMA_signal_1896, MCOutput[40]}), .a ({Plaintext_s1[40], Plaintext_s0[40]}), .c ({new_AGEMA_signal_1938, StateRegInput[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_41_U1 ( .s (rst), .b ({new_AGEMA_signal_1956, MCOutput[41]}), .a ({Plaintext_s1[41], Plaintext_s0[41]}), .c ({new_AGEMA_signal_1998, StateRegInput[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_44_U1 ( .s (rst), .b ({new_AGEMA_signal_2009, MCOutput[44]}), .a ({Plaintext_s1[44], Plaintext_s0[44]}), .c ({new_AGEMA_signal_2052, StateRegInput[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_45_U1 ( .s (rst), .b ({new_AGEMA_signal_2062, MCOutput[45]}), .a ({Plaintext_s1[45], Plaintext_s0[45]}), .c ({new_AGEMA_signal_2095, StateRegInput[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_48_U1 ( .s (rst), .b ({new_AGEMA_signal_2011, MCOutput[48]}), .a ({Plaintext_s1[48], Plaintext_s0[48]}), .c ({new_AGEMA_signal_2054, StateRegInput[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_49_U1 ( .s (rst), .b ({new_AGEMA_signal_2063, MCOutput[49]}), .a ({Plaintext_s1[49], Plaintext_s0[49]}), .c ({new_AGEMA_signal_2097, StateRegInput[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_52_U1 ( .s (rst), .b ({new_AGEMA_signal_2013, MCOutput[52]}), .a ({Plaintext_s1[52], Plaintext_s0[52]}), .c ({new_AGEMA_signal_2056, StateRegInput[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_53_U1 ( .s (rst), .b ({new_AGEMA_signal_2064, MCOutput[53]}), .a ({Plaintext_s1[53], Plaintext_s0[53]}), .c ({new_AGEMA_signal_2099, StateRegInput[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_56_U1 ( .s (rst), .b ({new_AGEMA_signal_2015, MCOutput[56]}), .a ({Plaintext_s1[56], Plaintext_s0[56]}), .c ({new_AGEMA_signal_2058, StateRegInput[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_57_U1 ( .s (rst), .b ({new_AGEMA_signal_2065, MCOutput[57]}), .a ({Plaintext_s1[57], Plaintext_s0[57]}), .c ({new_AGEMA_signal_2101, StateRegInput[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_60_U1 ( .s (rst), .b ({new_AGEMA_signal_2104, MCOutput[60]}), .a ({Plaintext_s1[60], Plaintext_s0[60]}), .c ({new_AGEMA_signal_2115, StateRegInput[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) PlaintextMUX_MUXInst_61_U1 ( .s (rst), .b ({new_AGEMA_signal_2116, MCOutput[61]}), .a ({Plaintext_s1[61], Plaintext_s0[61]}), .c ({new_AGEMA_signal_2124, StateRegInput[61]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_AND2_U1 ( .a ({Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1596, SubCellInst_SboxInst_0_Q2}), .clk (clk), .r (Fresh[32]), .c ({new_AGEMA_signal_1661, SubCellInst_SboxInst_0_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_XOR4_U1 ( .a ({new_AGEMA_signal_1661, SubCellInst_SboxInst_0_T1}), .b ({new_AGEMA_signal_1549, SubCellInst_SboxInst_0_T2}), .c ({new_AGEMA_signal_1725, SubCellInst_SboxInst_0_L0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_AND4_U1 ( .a ({new_AGEMA_signal_1456, SubCellInst_SboxInst_0_Q6}), .b ({new_AGEMA_signal_1597, SubCellInst_SboxInst_0_Q7}), .clk (clk), .r (Fresh[33]), .c ({new_AGEMA_signal_1662, SubCellInst_SboxInst_0_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_XOR9_U1 ( .a ({new_AGEMA_signal_1725, SubCellInst_SboxInst_0_L0}), .b ({new_AGEMA_signal_1457, SubCellInst_SboxInst_0_L2}), .c ({new_AGEMA_signal_1768, SubCellInst_SboxInst_0_YY_3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_XOR10_U1 ( .a ({new_AGEMA_signal_1725, SubCellInst_SboxInst_0_L0}), .b ({new_AGEMA_signal_1662, SubCellInst_SboxInst_0_T3}), .c ({new_AGEMA_signal_1769, ShiftRowsOutput[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_0_XOR_o1_U1 ( .a ({new_AGEMA_signal_1663, SubCellInst_SboxInst_0_YY_1_}), .b ({new_AGEMA_signal_1768, SubCellInst_SboxInst_0_YY_3}), .c ({new_AGEMA_signal_1826, ShiftRowsOutput[5]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_AND2_U1 ( .a ({Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1600, SubCellInst_SboxInst_1_Q2}), .clk (clk), .r (Fresh[34]), .c ({new_AGEMA_signal_1665, SubCellInst_SboxInst_1_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_XOR4_U1 ( .a ({new_AGEMA_signal_1665, SubCellInst_SboxInst_1_T1}), .b ({new_AGEMA_signal_1552, SubCellInst_SboxInst_1_T2}), .c ({new_AGEMA_signal_1727, SubCellInst_SboxInst_1_L0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_AND4_U1 ( .a ({new_AGEMA_signal_1462, SubCellInst_SboxInst_1_Q6}), .b ({new_AGEMA_signal_1601, SubCellInst_SboxInst_1_Q7}), .clk (clk), .r (Fresh[35]), .c ({new_AGEMA_signal_1666, SubCellInst_SboxInst_1_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_XOR9_U1 ( .a ({new_AGEMA_signal_1727, SubCellInst_SboxInst_1_L0}), .b ({new_AGEMA_signal_1463, SubCellInst_SboxInst_1_L2}), .c ({new_AGEMA_signal_1770, SubCellInst_SboxInst_1_YY_3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_XOR10_U1 ( .a ({new_AGEMA_signal_1727, SubCellInst_SboxInst_1_L0}), .b ({new_AGEMA_signal_1666, SubCellInst_SboxInst_1_T3}), .c ({new_AGEMA_signal_1771, ShiftRowsOutput[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_1_XOR_o1_U1 ( .a ({new_AGEMA_signal_1667, SubCellInst_SboxInst_1_YY_1_}), .b ({new_AGEMA_signal_1770, SubCellInst_SboxInst_1_YY_3}), .c ({new_AGEMA_signal_1827, ShiftRowsOutput[9]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_AND2_U1 ( .a ({Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1604, SubCellInst_SboxInst_2_Q2}), .clk (clk), .r (Fresh[36]), .c ({new_AGEMA_signal_1669, SubCellInst_SboxInst_2_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_XOR4_U1 ( .a ({new_AGEMA_signal_1669, SubCellInst_SboxInst_2_T1}), .b ({new_AGEMA_signal_1555, SubCellInst_SboxInst_2_T2}), .c ({new_AGEMA_signal_1729, SubCellInst_SboxInst_2_L0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_AND4_U1 ( .a ({new_AGEMA_signal_1468, SubCellInst_SboxInst_2_Q6}), .b ({new_AGEMA_signal_1605, SubCellInst_SboxInst_2_Q7}), .clk (clk), .r (Fresh[37]), .c ({new_AGEMA_signal_1670, SubCellInst_SboxInst_2_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_XOR9_U1 ( .a ({new_AGEMA_signal_1729, SubCellInst_SboxInst_2_L0}), .b ({new_AGEMA_signal_1469, SubCellInst_SboxInst_2_L2}), .c ({new_AGEMA_signal_1772, SubCellInst_SboxInst_2_YY_3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_XOR10_U1 ( .a ({new_AGEMA_signal_1729, SubCellInst_SboxInst_2_L0}), .b ({new_AGEMA_signal_1670, SubCellInst_SboxInst_2_T3}), .c ({new_AGEMA_signal_1773, ShiftRowsOutput[12]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_2_XOR_o1_U1 ( .a ({new_AGEMA_signal_1671, SubCellInst_SboxInst_2_YY_1_}), .b ({new_AGEMA_signal_1772, SubCellInst_SboxInst_2_YY_3}), .c ({new_AGEMA_signal_1828, ShiftRowsOutput[13]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_AND2_U1 ( .a ({Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1608, SubCellInst_SboxInst_3_Q2}), .clk (clk), .r (Fresh[38]), .c ({new_AGEMA_signal_1673, SubCellInst_SboxInst_3_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_XOR4_U1 ( .a ({new_AGEMA_signal_1673, SubCellInst_SboxInst_3_T1}), .b ({new_AGEMA_signal_1558, SubCellInst_SboxInst_3_T2}), .c ({new_AGEMA_signal_1731, SubCellInst_SboxInst_3_L0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_AND4_U1 ( .a ({new_AGEMA_signal_1474, SubCellInst_SboxInst_3_Q6}), .b ({new_AGEMA_signal_1609, SubCellInst_SboxInst_3_Q7}), .clk (clk), .r (Fresh[39]), .c ({new_AGEMA_signal_1674, SubCellInst_SboxInst_3_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_XOR9_U1 ( .a ({new_AGEMA_signal_1731, SubCellInst_SboxInst_3_L0}), .b ({new_AGEMA_signal_1475, SubCellInst_SboxInst_3_L2}), .c ({new_AGEMA_signal_1774, SubCellInst_SboxInst_3_YY_3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_XOR10_U1 ( .a ({new_AGEMA_signal_1731, SubCellInst_SboxInst_3_L0}), .b ({new_AGEMA_signal_1674, SubCellInst_SboxInst_3_T3}), .c ({new_AGEMA_signal_1775, ShiftRowsOutput[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_3_XOR_o1_U1 ( .a ({new_AGEMA_signal_1675, SubCellInst_SboxInst_3_YY_1_}), .b ({new_AGEMA_signal_1774, SubCellInst_SboxInst_3_YY_3}), .c ({new_AGEMA_signal_1829, ShiftRowsOutput[1]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_AND2_U1 ( .a ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1612, SubCellInst_SboxInst_4_Q2}), .clk (clk), .r (Fresh[40]), .c ({new_AGEMA_signal_1677, SubCellInst_SboxInst_4_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_XOR4_U1 ( .a ({new_AGEMA_signal_1677, SubCellInst_SboxInst_4_T1}), .b ({new_AGEMA_signal_1561, SubCellInst_SboxInst_4_T2}), .c ({new_AGEMA_signal_1733, SubCellInst_SboxInst_4_L0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_AND4_U1 ( .a ({new_AGEMA_signal_1480, SubCellInst_SboxInst_4_Q6}), .b ({new_AGEMA_signal_1613, SubCellInst_SboxInst_4_Q7}), .clk (clk), .r (Fresh[41]), .c ({new_AGEMA_signal_1678, SubCellInst_SboxInst_4_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_XOR9_U1 ( .a ({new_AGEMA_signal_1733, SubCellInst_SboxInst_4_L0}), .b ({new_AGEMA_signal_1481, SubCellInst_SboxInst_4_L2}), .c ({new_AGEMA_signal_1776, SubCellInst_SboxInst_4_YY_3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_XOR10_U1 ( .a ({new_AGEMA_signal_1733, SubCellInst_SboxInst_4_L0}), .b ({new_AGEMA_signal_1678, SubCellInst_SboxInst_4_T3}), .c ({new_AGEMA_signal_1777, ShiftRowsOutput[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_4_XOR_o1_U1 ( .a ({new_AGEMA_signal_1679, SubCellInst_SboxInst_4_YY_1_}), .b ({new_AGEMA_signal_1776, SubCellInst_SboxInst_4_YY_3}), .c ({new_AGEMA_signal_1830, ShiftRowsOutput[25]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_AND2_U1 ( .a ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1616, SubCellInst_SboxInst_5_Q2}), .clk (clk), .r (Fresh[42]), .c ({new_AGEMA_signal_1681, SubCellInst_SboxInst_5_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_XOR4_U1 ( .a ({new_AGEMA_signal_1681, SubCellInst_SboxInst_5_T1}), .b ({new_AGEMA_signal_1564, SubCellInst_SboxInst_5_T2}), .c ({new_AGEMA_signal_1735, SubCellInst_SboxInst_5_L0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_AND4_U1 ( .a ({new_AGEMA_signal_1486, SubCellInst_SboxInst_5_Q6}), .b ({new_AGEMA_signal_1617, SubCellInst_SboxInst_5_Q7}), .clk (clk), .r (Fresh[43]), .c ({new_AGEMA_signal_1682, SubCellInst_SboxInst_5_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_XOR9_U1 ( .a ({new_AGEMA_signal_1735, SubCellInst_SboxInst_5_L0}), .b ({new_AGEMA_signal_1487, SubCellInst_SboxInst_5_L2}), .c ({new_AGEMA_signal_1778, SubCellInst_SboxInst_5_YY_3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_XOR10_U1 ( .a ({new_AGEMA_signal_1735, SubCellInst_SboxInst_5_L0}), .b ({new_AGEMA_signal_1682, SubCellInst_SboxInst_5_T3}), .c ({new_AGEMA_signal_1779, ShiftRowsOutput[28]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_5_XOR_o1_U1 ( .a ({new_AGEMA_signal_1683, SubCellInst_SboxInst_5_YY_1_}), .b ({new_AGEMA_signal_1778, SubCellInst_SboxInst_5_YY_3}), .c ({new_AGEMA_signal_1831, ShiftRowsOutput[29]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_AND2_U1 ( .a ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1620, SubCellInst_SboxInst_6_Q2}), .clk (clk), .r (Fresh[44]), .c ({new_AGEMA_signal_1685, SubCellInst_SboxInst_6_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_XOR4_U1 ( .a ({new_AGEMA_signal_1685, SubCellInst_SboxInst_6_T1}), .b ({new_AGEMA_signal_1567, SubCellInst_SboxInst_6_T2}), .c ({new_AGEMA_signal_1737, SubCellInst_SboxInst_6_L0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_AND4_U1 ( .a ({new_AGEMA_signal_1492, SubCellInst_SboxInst_6_Q6}), .b ({new_AGEMA_signal_1621, SubCellInst_SboxInst_6_Q7}), .clk (clk), .r (Fresh[45]), .c ({new_AGEMA_signal_1686, SubCellInst_SboxInst_6_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_XOR9_U1 ( .a ({new_AGEMA_signal_1737, SubCellInst_SboxInst_6_L0}), .b ({new_AGEMA_signal_1493, SubCellInst_SboxInst_6_L2}), .c ({new_AGEMA_signal_1780, SubCellInst_SboxInst_6_YY_3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_XOR10_U1 ( .a ({new_AGEMA_signal_1737, SubCellInst_SboxInst_6_L0}), .b ({new_AGEMA_signal_1686, SubCellInst_SboxInst_6_T3}), .c ({new_AGEMA_signal_1781, ShiftRowsOutput[16]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_6_XOR_o1_U1 ( .a ({new_AGEMA_signal_1687, SubCellInst_SboxInst_6_YY_1_}), .b ({new_AGEMA_signal_1780, SubCellInst_SboxInst_6_YY_3}), .c ({new_AGEMA_signal_1832, ShiftRowsOutput[17]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_AND2_U1 ( .a ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1624, SubCellInst_SboxInst_7_Q2}), .clk (clk), .r (Fresh[46]), .c ({new_AGEMA_signal_1689, SubCellInst_SboxInst_7_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_XOR4_U1 ( .a ({new_AGEMA_signal_1689, SubCellInst_SboxInst_7_T1}), .b ({new_AGEMA_signal_1570, SubCellInst_SboxInst_7_T2}), .c ({new_AGEMA_signal_1739, SubCellInst_SboxInst_7_L0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_AND4_U1 ( .a ({new_AGEMA_signal_1498, SubCellInst_SboxInst_7_Q6}), .b ({new_AGEMA_signal_1625, SubCellInst_SboxInst_7_Q7}), .clk (clk), .r (Fresh[47]), .c ({new_AGEMA_signal_1690, SubCellInst_SboxInst_7_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_XOR9_U1 ( .a ({new_AGEMA_signal_1739, SubCellInst_SboxInst_7_L0}), .b ({new_AGEMA_signal_1499, SubCellInst_SboxInst_7_L2}), .c ({new_AGEMA_signal_1782, SubCellInst_SboxInst_7_YY_3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_XOR10_U1 ( .a ({new_AGEMA_signal_1739, SubCellInst_SboxInst_7_L0}), .b ({new_AGEMA_signal_1690, SubCellInst_SboxInst_7_T3}), .c ({new_AGEMA_signal_1783, ShiftRowsOutput[20]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_7_XOR_o1_U1 ( .a ({new_AGEMA_signal_1691, SubCellInst_SboxInst_7_YY_1_}), .b ({new_AGEMA_signal_1782, SubCellInst_SboxInst_7_YY_3}), .c ({new_AGEMA_signal_1833, SubCellOutput[29]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_AND2_U1 ( .a ({Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1628, SubCellInst_SboxInst_8_Q2}), .clk (clk), .r (Fresh[48]), .c ({new_AGEMA_signal_1693, SubCellInst_SboxInst_8_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_XOR4_U1 ( .a ({new_AGEMA_signal_1693, SubCellInst_SboxInst_8_T1}), .b ({new_AGEMA_signal_1573, SubCellInst_SboxInst_8_T2}), .c ({new_AGEMA_signal_1741, SubCellInst_SboxInst_8_L0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_AND4_U1 ( .a ({new_AGEMA_signal_1504, SubCellInst_SboxInst_8_Q6}), .b ({new_AGEMA_signal_1629, SubCellInst_SboxInst_8_Q7}), .clk (clk), .r (Fresh[49]), .c ({new_AGEMA_signal_1694, SubCellInst_SboxInst_8_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_XOR9_U1 ( .a ({new_AGEMA_signal_1741, SubCellInst_SboxInst_8_L0}), .b ({new_AGEMA_signal_1505, SubCellInst_SboxInst_8_L2}), .c ({new_AGEMA_signal_1784, SubCellInst_SboxInst_8_YY_3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_XOR10_U1 ( .a ({new_AGEMA_signal_1741, SubCellInst_SboxInst_8_L0}), .b ({new_AGEMA_signal_1694, SubCellInst_SboxInst_8_T3}), .c ({new_AGEMA_signal_1785, AddRoundConstantOutput[32]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_8_XOR_o1_U1 ( .a ({new_AGEMA_signal_1695, SubCellInst_SboxInst_8_YY_1_}), .b ({new_AGEMA_signal_1784, SubCellInst_SboxInst_8_YY_3}), .c ({new_AGEMA_signal_1834, AddRoundConstantOutput[33]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_AND2_U1 ( .a ({Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1632, SubCellInst_SboxInst_9_Q2}), .clk (clk), .r (Fresh[50]), .c ({new_AGEMA_signal_1697, SubCellInst_SboxInst_9_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_XOR4_U1 ( .a ({new_AGEMA_signal_1697, SubCellInst_SboxInst_9_T1}), .b ({new_AGEMA_signal_1576, SubCellInst_SboxInst_9_T2}), .c ({new_AGEMA_signal_1743, SubCellInst_SboxInst_9_L0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_AND4_U1 ( .a ({new_AGEMA_signal_1510, SubCellInst_SboxInst_9_Q6}), .b ({new_AGEMA_signal_1633, SubCellInst_SboxInst_9_Q7}), .clk (clk), .r (Fresh[51]), .c ({new_AGEMA_signal_1698, SubCellInst_SboxInst_9_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_XOR9_U1 ( .a ({new_AGEMA_signal_1743, SubCellInst_SboxInst_9_L0}), .b ({new_AGEMA_signal_1511, SubCellInst_SboxInst_9_L2}), .c ({new_AGEMA_signal_1786, SubCellInst_SboxInst_9_YY_3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_XOR10_U1 ( .a ({new_AGEMA_signal_1743, SubCellInst_SboxInst_9_L0}), .b ({new_AGEMA_signal_1698, SubCellInst_SboxInst_9_T3}), .c ({new_AGEMA_signal_1787, AddRoundConstantOutput[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_9_XOR_o1_U1 ( .a ({new_AGEMA_signal_1699, SubCellInst_SboxInst_9_YY_1_}), .b ({new_AGEMA_signal_1786, SubCellInst_SboxInst_9_YY_3}), .c ({new_AGEMA_signal_1835, AddRoundConstantOutput[37]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_AND2_U1 ( .a ({Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1636, SubCellInst_SboxInst_10_Q2}), .clk (clk), .r (Fresh[52]), .c ({new_AGEMA_signal_1701, SubCellInst_SboxInst_10_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_XOR4_U1 ( .a ({new_AGEMA_signal_1701, SubCellInst_SboxInst_10_T1}), .b ({new_AGEMA_signal_1579, SubCellInst_SboxInst_10_T2}), .c ({new_AGEMA_signal_1745, SubCellInst_SboxInst_10_L0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_AND4_U1 ( .a ({new_AGEMA_signal_1516, SubCellInst_SboxInst_10_Q6}), .b ({new_AGEMA_signal_1637, SubCellInst_SboxInst_10_Q7}), .clk (clk), .r (Fresh[53]), .c ({new_AGEMA_signal_1702, SubCellInst_SboxInst_10_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_XOR9_U1 ( .a ({new_AGEMA_signal_1745, SubCellInst_SboxInst_10_L0}), .b ({new_AGEMA_signal_1517, SubCellInst_SboxInst_10_L2}), .c ({new_AGEMA_signal_1788, SubCellInst_SboxInst_10_YY_3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_XOR10_U1 ( .a ({new_AGEMA_signal_1745, SubCellInst_SboxInst_10_L0}), .b ({new_AGEMA_signal_1702, SubCellInst_SboxInst_10_T3}), .c ({new_AGEMA_signal_1789, AddRoundConstantOutput[40]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_10_XOR_o1_U1 ( .a ({new_AGEMA_signal_1703, SubCellInst_SboxInst_10_YY_1_}), .b ({new_AGEMA_signal_1788, SubCellInst_SboxInst_10_YY_3}), .c ({new_AGEMA_signal_1836, AddRoundConstantOutput[41]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_AND2_U1 ( .a ({Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1640, SubCellInst_SboxInst_11_Q2}), .clk (clk), .r (Fresh[54]), .c ({new_AGEMA_signal_1705, SubCellInst_SboxInst_11_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_XOR4_U1 ( .a ({new_AGEMA_signal_1705, SubCellInst_SboxInst_11_T1}), .b ({new_AGEMA_signal_1582, SubCellInst_SboxInst_11_T2}), .c ({new_AGEMA_signal_1747, SubCellInst_SboxInst_11_L0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_AND4_U1 ( .a ({new_AGEMA_signal_1522, SubCellInst_SboxInst_11_Q6}), .b ({new_AGEMA_signal_1641, SubCellInst_SboxInst_11_Q7}), .clk (clk), .r (Fresh[55]), .c ({new_AGEMA_signal_1706, SubCellInst_SboxInst_11_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_XOR9_U1 ( .a ({new_AGEMA_signal_1747, SubCellInst_SboxInst_11_L0}), .b ({new_AGEMA_signal_1523, SubCellInst_SboxInst_11_L2}), .c ({new_AGEMA_signal_1790, SubCellInst_SboxInst_11_YY_3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_XOR10_U1 ( .a ({new_AGEMA_signal_1747, SubCellInst_SboxInst_11_L0}), .b ({new_AGEMA_signal_1706, SubCellInst_SboxInst_11_T3}), .c ({new_AGEMA_signal_1791, SubCellOutput[44]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_11_XOR_o1_U1 ( .a ({new_AGEMA_signal_1707, SubCellInst_SboxInst_11_YY_1_}), .b ({new_AGEMA_signal_1790, SubCellInst_SboxInst_11_YY_3}), .c ({new_AGEMA_signal_1837, SubCellOutput[45]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_AND2_U1 ( .a ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1644, SubCellInst_SboxInst_12_Q2}), .clk (clk), .r (Fresh[56]), .c ({new_AGEMA_signal_1709, SubCellInst_SboxInst_12_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_XOR4_U1 ( .a ({new_AGEMA_signal_1709, SubCellInst_SboxInst_12_T1}), .b ({new_AGEMA_signal_1585, SubCellInst_SboxInst_12_T2}), .c ({new_AGEMA_signal_1749, SubCellInst_SboxInst_12_L0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_AND4_U1 ( .a ({new_AGEMA_signal_1528, SubCellInst_SboxInst_12_Q6}), .b ({new_AGEMA_signal_1645, SubCellInst_SboxInst_12_Q7}), .clk (clk), .r (Fresh[57]), .c ({new_AGEMA_signal_1710, SubCellInst_SboxInst_12_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_XOR9_U1 ( .a ({new_AGEMA_signal_1749, SubCellInst_SboxInst_12_L0}), .b ({new_AGEMA_signal_1529, SubCellInst_SboxInst_12_L2}), .c ({new_AGEMA_signal_1792, SubCellInst_SboxInst_12_YY_3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_XOR10_U1 ( .a ({new_AGEMA_signal_1749, SubCellInst_SboxInst_12_L0}), .b ({new_AGEMA_signal_1710, SubCellInst_SboxInst_12_T3}), .c ({new_AGEMA_signal_1793, AddRoundConstantOutput[48]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_12_XOR_o1_U1 ( .a ({new_AGEMA_signal_1711, SubCellInst_SboxInst_12_YY_1_}), .b ({new_AGEMA_signal_1792, SubCellInst_SboxInst_12_YY_3}), .c ({new_AGEMA_signal_1838, AddRoundConstantOutput[49]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_AND2_U1 ( .a ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1648, SubCellInst_SboxInst_13_Q2}), .clk (clk), .r (Fresh[58]), .c ({new_AGEMA_signal_1713, SubCellInst_SboxInst_13_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_XOR4_U1 ( .a ({new_AGEMA_signal_1713, SubCellInst_SboxInst_13_T1}), .b ({new_AGEMA_signal_1588, SubCellInst_SboxInst_13_T2}), .c ({new_AGEMA_signal_1751, SubCellInst_SboxInst_13_L0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_AND4_U1 ( .a ({new_AGEMA_signal_1534, SubCellInst_SboxInst_13_Q6}), .b ({new_AGEMA_signal_1649, SubCellInst_SboxInst_13_Q7}), .clk (clk), .r (Fresh[59]), .c ({new_AGEMA_signal_1714, SubCellInst_SboxInst_13_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_XOR9_U1 ( .a ({new_AGEMA_signal_1751, SubCellInst_SboxInst_13_L0}), .b ({new_AGEMA_signal_1535, SubCellInst_SboxInst_13_L2}), .c ({new_AGEMA_signal_1794, SubCellInst_SboxInst_13_YY_3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_XOR10_U1 ( .a ({new_AGEMA_signal_1751, SubCellInst_SboxInst_13_L0}), .b ({new_AGEMA_signal_1714, SubCellInst_SboxInst_13_T3}), .c ({new_AGEMA_signal_1795, AddRoundConstantOutput[52]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_13_XOR_o1_U1 ( .a ({new_AGEMA_signal_1715, SubCellInst_SboxInst_13_YY_1_}), .b ({new_AGEMA_signal_1794, SubCellInst_SboxInst_13_YY_3}), .c ({new_AGEMA_signal_1839, AddRoundConstantOutput[53]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_AND2_U1 ( .a ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1652, SubCellInst_SboxInst_14_Q2}), .clk (clk), .r (Fresh[60]), .c ({new_AGEMA_signal_1717, SubCellInst_SboxInst_14_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_XOR4_U1 ( .a ({new_AGEMA_signal_1717, SubCellInst_SboxInst_14_T1}), .b ({new_AGEMA_signal_1591, SubCellInst_SboxInst_14_T2}), .c ({new_AGEMA_signal_1753, SubCellInst_SboxInst_14_L0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_AND4_U1 ( .a ({new_AGEMA_signal_1540, SubCellInst_SboxInst_14_Q6}), .b ({new_AGEMA_signal_1653, SubCellInst_SboxInst_14_Q7}), .clk (clk), .r (Fresh[61]), .c ({new_AGEMA_signal_1718, SubCellInst_SboxInst_14_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_XOR9_U1 ( .a ({new_AGEMA_signal_1753, SubCellInst_SboxInst_14_L0}), .b ({new_AGEMA_signal_1541, SubCellInst_SboxInst_14_L2}), .c ({new_AGEMA_signal_1796, SubCellInst_SboxInst_14_YY_3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_XOR10_U1 ( .a ({new_AGEMA_signal_1753, SubCellInst_SboxInst_14_L0}), .b ({new_AGEMA_signal_1718, SubCellInst_SboxInst_14_T3}), .c ({new_AGEMA_signal_1797, AddRoundConstantOutput[56]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_14_XOR_o1_U1 ( .a ({new_AGEMA_signal_1719, SubCellInst_SboxInst_14_YY_1_}), .b ({new_AGEMA_signal_1796, SubCellInst_SboxInst_14_YY_3}), .c ({new_AGEMA_signal_1840, AddRoundConstantOutput[57]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_AND2_U1 ( .a ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1656, SubCellInst_SboxInst_15_Q2}), .clk (clk), .r (Fresh[62]), .c ({new_AGEMA_signal_1721, SubCellInst_SboxInst_15_T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_XOR4_U1 ( .a ({new_AGEMA_signal_1721, SubCellInst_SboxInst_15_T1}), .b ({new_AGEMA_signal_1594, SubCellInst_SboxInst_15_T2}), .c ({new_AGEMA_signal_1755, SubCellInst_SboxInst_15_L0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_AND4_U1 ( .a ({new_AGEMA_signal_1546, SubCellInst_SboxInst_15_Q6}), .b ({new_AGEMA_signal_1657, SubCellInst_SboxInst_15_Q7}), .clk (clk), .r (Fresh[63]), .c ({new_AGEMA_signal_1722, SubCellInst_SboxInst_15_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_XOR9_U1 ( .a ({new_AGEMA_signal_1755, SubCellInst_SboxInst_15_L0}), .b ({new_AGEMA_signal_1547, SubCellInst_SboxInst_15_L2}), .c ({new_AGEMA_signal_1798, SubCellInst_SboxInst_15_YY_3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_XOR10_U1 ( .a ({new_AGEMA_signal_1755, SubCellInst_SboxInst_15_L0}), .b ({new_AGEMA_signal_1722, SubCellInst_SboxInst_15_T3}), .c ({new_AGEMA_signal_1799, SubCellOutput[60]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SubCellInst_SboxInst_15_XOR_o1_U1 ( .a ({new_AGEMA_signal_1723, SubCellInst_SboxInst_15_YY_1_}), .b ({new_AGEMA_signal_1798, SubCellInst_SboxInst_15_YY_3}), .c ({new_AGEMA_signal_1841, SubCellOutput[61]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) AddConstXOR_U2 ( .a ({new_AGEMA_signal_1833, SubCellOutput[29]}), .b ({new_AGEMA_signal_1879, ShiftRowsOutput[21]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_1842, AddConstXOR_AddConstXOR_XORInst_0_0_n1}), .b ({1'b0, FSMUpdate[1]}), .c ({new_AGEMA_signal_1880, AddRoundConstantOutput[60]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1799, SubCellOutput[60]}), .c ({new_AGEMA_signal_1842, AddConstXOR_AddConstXOR_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_1881, AddConstXOR_AddConstXOR_XORInst_0_1_n1}), .b ({1'b0, FSM[1]}), .c ({new_AGEMA_signal_1947, AddRoundConstantOutput[61]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1841, SubCellOutput[61]}), .c ({new_AGEMA_signal_1881, AddConstXOR_AddConstXOR_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_1844, AddConstXOR_AddConstXOR_XORInst_1_0_n1}), .b ({1'b0, FSM[4]}), .c ({new_AGEMA_signal_1882, AddRoundConstantOutput[44]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1791, SubCellOutput[44]}), .c ({new_AGEMA_signal_1844, AddConstXOR_AddConstXOR_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_1883, AddConstXOR_AddConstXOR_XORInst_1_1_n1}), .b ({1'b0, FSM[5]}), .c ({new_AGEMA_signal_1948, AddRoundConstantOutput[45]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1837, SubCellOutput[45]}), .c ({new_AGEMA_signal_1883, AddConstXOR_AddConstXOR_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_1846, AddRoundTweakeyXOR_XORInst_0_0_n1}), .b ({new_AGEMA_signal_1260, TweakeyGeneration_key_Feedback[0]}), .c ({new_AGEMA_signal_1884, ShiftRowsOutput[44]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1785, AddRoundConstantOutput[32]}), .c ({new_AGEMA_signal_1846, AddRoundTweakeyXOR_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_1885, AddRoundTweakeyXOR_XORInst_0_1_n1}), .b ({new_AGEMA_signal_1263, TweakeyGeneration_key_Feedback[1]}), .c ({new_AGEMA_signal_1949, ShiftRowsOutput[45]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1834, AddRoundConstantOutput[33]}), .c ({new_AGEMA_signal_1885, AddRoundTweakeyXOR_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_1848, AddRoundTweakeyXOR_XORInst_1_0_n1}), .b ({new_AGEMA_signal_1272, TweakeyGeneration_key_Feedback[4]}), .c ({new_AGEMA_signal_1886, ShiftRowsOutput[32]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1787, AddRoundConstantOutput[36]}), .c ({new_AGEMA_signal_1848, AddRoundTweakeyXOR_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_1887, AddRoundTweakeyXOR_XORInst_1_1_n1}), .b ({new_AGEMA_signal_1275, TweakeyGeneration_key_Feedback[5]}), .c ({new_AGEMA_signal_1950, ShiftRowsOutput[33]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1835, AddRoundConstantOutput[37]}), .c ({new_AGEMA_signal_1887, AddRoundTweakeyXOR_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_1850, AddRoundTweakeyXOR_XORInst_2_0_n1}), .b ({new_AGEMA_signal_1284, TweakeyGeneration_key_Feedback[8]}), .c ({new_AGEMA_signal_1888, ShiftRowsOutput[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1789, AddRoundConstantOutput[40]}), .c ({new_AGEMA_signal_1850, AddRoundTweakeyXOR_XORInst_2_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_1889, AddRoundTweakeyXOR_XORInst_2_1_n1}), .b ({new_AGEMA_signal_1287, TweakeyGeneration_key_Feedback[9]}), .c ({new_AGEMA_signal_1951, ShiftRowsOutput[37]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1836, AddRoundConstantOutput[41]}), .c ({new_AGEMA_signal_1889, AddRoundTweakeyXOR_XORInst_2_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_1952, AddRoundTweakeyXOR_XORInst_3_0_n1}), .b ({new_AGEMA_signal_1296, TweakeyGeneration_key_Feedback[12]}), .c ({new_AGEMA_signal_2007, ShiftRowsOutput[40]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1882, AddRoundConstantOutput[44]}), .c ({new_AGEMA_signal_1952, AddRoundTweakeyXOR_XORInst_3_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_2008, AddRoundTweakeyXOR_XORInst_3_1_n1}), .b ({new_AGEMA_signal_1299, TweakeyGeneration_key_Feedback[13]}), .c ({new_AGEMA_signal_2061, ShiftRowsOutput[41]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1948, AddRoundConstantOutput[45]}), .c ({new_AGEMA_signal_2008, AddRoundTweakeyXOR_XORInst_3_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_0_U2 ( .a ({new_AGEMA_signal_1853, AddRoundTweakeyXOR_XORInst_4_0_n1}), .b ({new_AGEMA_signal_1308, TweakeyGeneration_key_Feedback[16]}), .c ({new_AGEMA_signal_1892, MCOutput[32]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1793, AddRoundConstantOutput[48]}), .c ({new_AGEMA_signal_1853, AddRoundTweakeyXOR_XORInst_4_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_1_U2 ( .a ({new_AGEMA_signal_1893, AddRoundTweakeyXOR_XORInst_4_1_n1}), .b ({new_AGEMA_signal_1311, TweakeyGeneration_key_Feedback[17]}), .c ({new_AGEMA_signal_1954, MCOutput[33]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1838, AddRoundConstantOutput[49]}), .c ({new_AGEMA_signal_1893, AddRoundTweakeyXOR_XORInst_4_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_0_U2 ( .a ({new_AGEMA_signal_1855, AddRoundTweakeyXOR_XORInst_5_0_n1}), .b ({new_AGEMA_signal_1320, TweakeyGeneration_key_Feedback[20]}), .c ({new_AGEMA_signal_1894, MCOutput[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1795, AddRoundConstantOutput[52]}), .c ({new_AGEMA_signal_1855, AddRoundTweakeyXOR_XORInst_5_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_1_U2 ( .a ({new_AGEMA_signal_1895, AddRoundTweakeyXOR_XORInst_5_1_n1}), .b ({new_AGEMA_signal_1323, TweakeyGeneration_key_Feedback[21]}), .c ({new_AGEMA_signal_1955, MCOutput[37]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1839, AddRoundConstantOutput[53]}), .c ({new_AGEMA_signal_1895, AddRoundTweakeyXOR_XORInst_5_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_0_U2 ( .a ({new_AGEMA_signal_1857, AddRoundTweakeyXOR_XORInst_6_0_n1}), .b ({new_AGEMA_signal_1332, TweakeyGeneration_key_Feedback[24]}), .c ({new_AGEMA_signal_1896, MCOutput[40]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1797, AddRoundConstantOutput[56]}), .c ({new_AGEMA_signal_1857, AddRoundTweakeyXOR_XORInst_6_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_1_U2 ( .a ({new_AGEMA_signal_1897, AddRoundTweakeyXOR_XORInst_6_1_n1}), .b ({new_AGEMA_signal_1335, TweakeyGeneration_key_Feedback[25]}), .c ({new_AGEMA_signal_1956, MCOutput[41]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1840, AddRoundConstantOutput[57]}), .c ({new_AGEMA_signal_1897, AddRoundTweakeyXOR_XORInst_6_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_0_U2 ( .a ({new_AGEMA_signal_1957, AddRoundTweakeyXOR_XORInst_7_0_n1}), .b ({new_AGEMA_signal_1344, TweakeyGeneration_key_Feedback[28]}), .c ({new_AGEMA_signal_2009, MCOutput[44]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1880, AddRoundConstantOutput[60]}), .c ({new_AGEMA_signal_1957, AddRoundTweakeyXOR_XORInst_7_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_1_U2 ( .a ({new_AGEMA_signal_2010, AddRoundTweakeyXOR_XORInst_7_1_n1}), .b ({new_AGEMA_signal_1347, TweakeyGeneration_key_Feedback[29]}), .c ({new_AGEMA_signal_2062, MCOutput[45]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1947, AddRoundConstantOutput[61]}), .c ({new_AGEMA_signal_2010, AddRoundTweakeyXOR_XORInst_7_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_0_0_U3 ( .a ({new_AGEMA_signal_1959, MCInst_MCR0_XORInst_0_0_n2}), .b ({new_AGEMA_signal_1860, MCInst_MCR0_XORInst_0_0_n1}), .c ({new_AGEMA_signal_2011, MCOutput[48]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_1781, ShiftRowsOutput[16]}), .b ({new_AGEMA_signal_1775, ShiftRowsOutput[0]}), .c ({new_AGEMA_signal_1860, MCInst_MCR0_XORInst_0_0_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_0_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1892, MCOutput[32]}), .c ({new_AGEMA_signal_1959, MCInst_MCR0_XORInst_0_0_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_0_1_U3 ( .a ({new_AGEMA_signal_2012, MCInst_MCR0_XORInst_0_1_n2}), .b ({new_AGEMA_signal_1900, MCInst_MCR0_XORInst_0_1_n1}), .c ({new_AGEMA_signal_2063, MCOutput[49]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_1832, ShiftRowsOutput[17]}), .b ({new_AGEMA_signal_1829, ShiftRowsOutput[1]}), .c ({new_AGEMA_signal_1900, MCInst_MCR0_XORInst_0_1_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_0_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1954, MCOutput[33]}), .c ({new_AGEMA_signal_2012, MCInst_MCR0_XORInst_0_1_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_1_0_U3 ( .a ({new_AGEMA_signal_1961, MCInst_MCR0_XORInst_1_0_n2}), .b ({new_AGEMA_signal_1862, MCInst_MCR0_XORInst_1_0_n1}), .c ({new_AGEMA_signal_2013, MCOutput[52]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_1783, ShiftRowsOutput[20]}), .b ({new_AGEMA_signal_1769, ShiftRowsOutput[4]}), .c ({new_AGEMA_signal_1862, MCInst_MCR0_XORInst_1_0_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_1_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1894, MCOutput[36]}), .c ({new_AGEMA_signal_1961, MCInst_MCR0_XORInst_1_0_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_1_1_U3 ( .a ({new_AGEMA_signal_2014, MCInst_MCR0_XORInst_1_1_n2}), .b ({new_AGEMA_signal_1962, MCInst_MCR0_XORInst_1_1_n1}), .c ({new_AGEMA_signal_2064, MCOutput[53]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_1879, ShiftRowsOutput[21]}), .b ({new_AGEMA_signal_1826, ShiftRowsOutput[5]}), .c ({new_AGEMA_signal_1962, MCInst_MCR0_XORInst_1_1_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_1_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1955, MCOutput[37]}), .c ({new_AGEMA_signal_2014, MCInst_MCR0_XORInst_1_1_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_2_0_U3 ( .a ({new_AGEMA_signal_1964, MCInst_MCR0_XORInst_2_0_n2}), .b ({new_AGEMA_signal_1864, MCInst_MCR0_XORInst_2_0_n1}), .c ({new_AGEMA_signal_2015, MCOutput[56]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_1777, ShiftRowsOutput[24]}), .b ({new_AGEMA_signal_1771, ShiftRowsOutput[8]}), .c ({new_AGEMA_signal_1864, MCInst_MCR0_XORInst_2_0_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_2_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1896, MCOutput[40]}), .c ({new_AGEMA_signal_1964, MCInst_MCR0_XORInst_2_0_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_2_1_U3 ( .a ({new_AGEMA_signal_2016, MCInst_MCR0_XORInst_2_1_n2}), .b ({new_AGEMA_signal_1905, MCInst_MCR0_XORInst_2_1_n1}), .c ({new_AGEMA_signal_2065, MCOutput[57]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_1830, ShiftRowsOutput[25]}), .b ({new_AGEMA_signal_1827, ShiftRowsOutput[9]}), .c ({new_AGEMA_signal_1905, MCInst_MCR0_XORInst_2_1_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_2_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1956, MCOutput[41]}), .c ({new_AGEMA_signal_2016, MCInst_MCR0_XORInst_2_1_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_3_0_U3 ( .a ({new_AGEMA_signal_2066, MCInst_MCR0_XORInst_3_0_n2}), .b ({new_AGEMA_signal_1866, MCInst_MCR0_XORInst_3_0_n1}), .c ({new_AGEMA_signal_2104, MCOutput[60]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_1779, ShiftRowsOutput[28]}), .b ({new_AGEMA_signal_1773, ShiftRowsOutput[12]}), .c ({new_AGEMA_signal_1866, MCInst_MCR0_XORInst_3_0_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_3_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_2009, MCOutput[44]}), .c ({new_AGEMA_signal_2066, MCInst_MCR0_XORInst_3_0_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_3_1_U3 ( .a ({new_AGEMA_signal_2105, MCInst_MCR0_XORInst_3_1_n2}), .b ({new_AGEMA_signal_1908, MCInst_MCR0_XORInst_3_1_n1}), .c ({new_AGEMA_signal_2116, MCOutput[61]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_1831, ShiftRowsOutput[29]}), .b ({new_AGEMA_signal_1828, ShiftRowsOutput[13]}), .c ({new_AGEMA_signal_1908, MCInst_MCR0_XORInst_3_1_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR0_XORInst_3_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_2062, MCOutput[45]}), .c ({new_AGEMA_signal_2105, MCInst_MCR0_XORInst_3_1_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_1967, MCInst_MCR2_XORInst_0_0_n1}), .b ({new_AGEMA_signal_1781, ShiftRowsOutput[16]}), .c ({new_AGEMA_signal_2019, MCOutput[16]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_0_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1886, ShiftRowsOutput[32]}), .c ({new_AGEMA_signal_1967, MCInst_MCR2_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2020, MCInst_MCR2_XORInst_0_1_n1}), .b ({new_AGEMA_signal_1832, ShiftRowsOutput[17]}), .c ({new_AGEMA_signal_2068, MCOutput[17]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_0_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1950, ShiftRowsOutput[33]}), .c ({new_AGEMA_signal_2020, MCInst_MCR2_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_1969, MCInst_MCR2_XORInst_1_0_n1}), .b ({new_AGEMA_signal_1783, ShiftRowsOutput[20]}), .c ({new_AGEMA_signal_2021, MCOutput[20]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_1_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1888, ShiftRowsOutput[36]}), .c ({new_AGEMA_signal_1969, MCInst_MCR2_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2022, MCInst_MCR2_XORInst_1_1_n1}), .b ({new_AGEMA_signal_1879, ShiftRowsOutput[21]}), .c ({new_AGEMA_signal_2069, MCOutput[21]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_1_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1951, ShiftRowsOutput[37]}), .c ({new_AGEMA_signal_2022, MCInst_MCR2_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_2070, MCInst_MCR2_XORInst_2_0_n1}), .b ({new_AGEMA_signal_1777, ShiftRowsOutput[24]}), .c ({new_AGEMA_signal_2106, MCOutput[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_2_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_2007, ShiftRowsOutput[40]}), .c ({new_AGEMA_signal_2070, MCInst_MCR2_XORInst_2_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_2107, MCInst_MCR2_XORInst_2_1_n1}), .b ({new_AGEMA_signal_1830, ShiftRowsOutput[25]}), .c ({new_AGEMA_signal_2117, MCOutput[25]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_2_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_2061, ShiftRowsOutput[41]}), .c ({new_AGEMA_signal_2107, MCInst_MCR2_XORInst_2_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_1972, MCInst_MCR2_XORInst_3_0_n1}), .b ({new_AGEMA_signal_1779, ShiftRowsOutput[28]}), .c ({new_AGEMA_signal_2025, MCOutput[28]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_3_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1884, ShiftRowsOutput[44]}), .c ({new_AGEMA_signal_1972, MCInst_MCR2_XORInst_3_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_2026, MCInst_MCR2_XORInst_3_1_n1}), .b ({new_AGEMA_signal_1831, ShiftRowsOutput[29]}), .c ({new_AGEMA_signal_2072, MCOutput[29]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR2_XORInst_3_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1949, ShiftRowsOutput[45]}), .c ({new_AGEMA_signal_2026, MCInst_MCR2_XORInst_3_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_1974, MCInst_MCR3_XORInst_0_0_n1}), .b ({new_AGEMA_signal_1781, ShiftRowsOutput[16]}), .c ({new_AGEMA_signal_2027, MCOutput[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_0_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1892, MCOutput[32]}), .c ({new_AGEMA_signal_1974, MCInst_MCR3_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2028, MCInst_MCR3_XORInst_0_1_n1}), .b ({new_AGEMA_signal_1832, ShiftRowsOutput[17]}), .c ({new_AGEMA_signal_2073, MCOutput[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_0_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1954, MCOutput[33]}), .c ({new_AGEMA_signal_2028, MCInst_MCR3_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_1976, MCInst_MCR3_XORInst_1_0_n1}), .b ({new_AGEMA_signal_1783, ShiftRowsOutput[20]}), .c ({new_AGEMA_signal_2029, MCOutput[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_1_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1894, MCOutput[36]}), .c ({new_AGEMA_signal_1976, MCInst_MCR3_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2030, MCInst_MCR3_XORInst_1_1_n1}), .b ({new_AGEMA_signal_1879, ShiftRowsOutput[21]}), .c ({new_AGEMA_signal_2074, MCOutput[5]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_1_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1955, MCOutput[37]}), .c ({new_AGEMA_signal_2030, MCInst_MCR3_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_1978, MCInst_MCR3_XORInst_2_0_n1}), .b ({new_AGEMA_signal_1777, ShiftRowsOutput[24]}), .c ({new_AGEMA_signal_2031, MCOutput[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_2_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1896, MCOutput[40]}), .c ({new_AGEMA_signal_1978, MCInst_MCR3_XORInst_2_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_2032, MCInst_MCR3_XORInst_2_1_n1}), .b ({new_AGEMA_signal_1830, ShiftRowsOutput[25]}), .c ({new_AGEMA_signal_2075, MCOutput[9]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_2_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1956, MCOutput[41]}), .c ({new_AGEMA_signal_2032, MCInst_MCR3_XORInst_2_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_2076, MCInst_MCR3_XORInst_3_0_n1}), .b ({new_AGEMA_signal_1779, ShiftRowsOutput[28]}), .c ({new_AGEMA_signal_2108, MCOutput[12]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_3_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_2009, MCOutput[44]}), .c ({new_AGEMA_signal_2076, MCInst_MCR3_XORInst_3_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_2109, MCInst_MCR3_XORInst_3_1_n1}), .b ({new_AGEMA_signal_1831, ShiftRowsOutput[29]}), .c ({new_AGEMA_signal_2118, MCOutput[13]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) MCInst_MCR3_XORInst_3_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_2062, MCOutput[45]}), .c ({new_AGEMA_signal_2109, MCInst_MCR3_XORInst_3_1_n1}) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_63__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2103, StateRegInput[63]}), .Q ({Ciphertext_s1[63], Ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_62__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2060, StateRegInput[62]}), .Q ({Ciphertext_s1[62], Ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_61__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2124, StateRegInput[61]}), .Q ({Ciphertext_s1[61], Ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_60__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2115, StateRegInput[60]}), .Q ({Ciphertext_s1[60], Ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_59__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2006, StateRegInput[59]}), .Q ({Ciphertext_s1[59], Ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_58__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1946, StateRegInput[58]}), .Q ({Ciphertext_s1[58], Ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_57__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2101, StateRegInput[57]}), .Q ({Ciphertext_s1[57], Ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_56__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2058, StateRegInput[56]}), .Q ({Ciphertext_s1[56], Ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_55__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2004, StateRegInput[55]}), .Q ({Ciphertext_s1[55], Ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_54__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1944, StateRegInput[54]}), .Q ({Ciphertext_s1[54], Ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_53__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2099, StateRegInput[53]}), .Q ({Ciphertext_s1[53], Ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_52__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2056, StateRegInput[52]}), .Q ({Ciphertext_s1[52], Ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_51__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2002, StateRegInput[51]}), .Q ({Ciphertext_s1[51], Ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_50__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1942, StateRegInput[50]}), .Q ({Ciphertext_s1[50], Ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_49__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2097, StateRegInput[49]}), .Q ({Ciphertext_s1[49], Ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_48__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2054, StateRegInput[48]}), .Q ({Ciphertext_s1[48], Ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_47__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2000, StateRegInput[47]}), .Q ({Ciphertext_s1[47], Ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_46__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1940, StateRegInput[46]}), .Q ({Ciphertext_s1[46], Ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_45__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2095, StateRegInput[45]}), .Q ({Ciphertext_s1[45], Ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_44__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2052, StateRegInput[44]}), .Q ({Ciphertext_s1[44], Ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_43__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1878, StateRegInput[43]}), .Q ({Ciphertext_s1[43], Ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_42__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1825, StateRegInput[42]}), .Q ({Ciphertext_s1[42], Ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_41__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1998, StateRegInput[41]}), .Q ({Ciphertext_s1[41], Ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_40__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1938, StateRegInput[40]}), .Q ({Ciphertext_s1[40], Ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_39__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1876, StateRegInput[39]}), .Q ({Ciphertext_s1[39], Ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_38__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1823, StateRegInput[38]}), .Q ({Ciphertext_s1[38], Ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_37__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1996, StateRegInput[37]}), .Q ({Ciphertext_s1[37], Ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_36__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1936, StateRegInput[36]}), .Q ({Ciphertext_s1[36], Ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_35__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1874, StateRegInput[35]}), .Q ({Ciphertext_s1[35], Ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_34__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1821, StateRegInput[34]}), .Q ({Ciphertext_s1[34], Ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_33__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1994, StateRegInput[33]}), .Q ({Ciphertext_s1[33], Ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_32__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1934, StateRegInput[32]}), .Q ({Ciphertext_s1[32], Ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_31__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1992, StateRegInput[31]}), .Q ({Ciphertext_s1[31], Ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_30__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1932, StateRegInput[30]}), .Q ({Ciphertext_s1[30], Ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_29__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2093, StateRegInput[29]}), .Q ({Ciphertext_s1[29], Ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_28__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2050, StateRegInput[28]}), .Q ({Ciphertext_s1[28], Ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_27__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2091, StateRegInput[27]}), .Q ({Ciphertext_s1[27], Ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_26__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2048, StateRegInput[26]}), .Q ({Ciphertext_s1[26], Ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_25__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2122, StateRegInput[25]}), .Q ({Ciphertext_s1[25], Ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_24__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2113, StateRegInput[24]}), .Q ({Ciphertext_s1[24], Ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_23__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1990, StateRegInput[23]}), .Q ({Ciphertext_s1[23], Ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_22__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1930, StateRegInput[22]}), .Q ({Ciphertext_s1[22], Ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_21__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2089, StateRegInput[21]}), .Q ({Ciphertext_s1[21], Ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_20__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2046, StateRegInput[20]}), .Q ({Ciphertext_s1[20], Ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_19__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1988, StateRegInput[19]}), .Q ({Ciphertext_s1[19], Ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_18__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1928, StateRegInput[18]}), .Q ({Ciphertext_s1[18], Ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_17__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2087, StateRegInput[17]}), .Q ({Ciphertext_s1[17], Ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_16__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2044, StateRegInput[16]}), .Q ({Ciphertext_s1[16], Ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_15__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2085, StateRegInput[15]}), .Q ({Ciphertext_s1[15], Ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_14__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2042, StateRegInput[14]}), .Q ({Ciphertext_s1[14], Ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_13__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2120, StateRegInput[13]}), .Q ({Ciphertext_s1[13], Ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_12__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2111, StateRegInput[12]}), .Q ({Ciphertext_s1[12], Ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_11__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1986, StateRegInput[11]}), .Q ({Ciphertext_s1[11], Ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_10__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1926, StateRegInput[10]}), .Q ({Ciphertext_s1[10], Ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_9__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2083, StateRegInput[9]}), .Q ({Ciphertext_s1[9], Ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_8__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2040, StateRegInput[8]}), .Q ({Ciphertext_s1[8], Ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_7__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1984, StateRegInput[7]}), .Q ({Ciphertext_s1[7], Ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_6__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1924, StateRegInput[6]}), .Q ({Ciphertext_s1[6], Ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_5__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2081, StateRegInput[5]}), .Q ({Ciphertext_s1[5], Ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_4__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2038, StateRegInput[4]}), .Q ({Ciphertext_s1[4], Ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1982, StateRegInput[3]}), .Q ({Ciphertext_s1[3], Ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1922, StateRegInput[2]}), .Q ({Ciphertext_s1[2], Ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2079, StateRegInput[1]}), .Q ({Ciphertext_s1[1], Ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) StateReg_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2036, StateRegInput[0]}), .Q ({Ciphertext_s1[0], Ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1451, TweakeyGeneration_StateRegInput[63]}), .Q ({new_AGEMA_signal_1353, TweakeyGeneration_key_Feedback[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1448, TweakeyGeneration_StateRegInput[62]}), .Q ({new_AGEMA_signal_1350, TweakeyGeneration_key_Feedback[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1445, TweakeyGeneration_StateRegInput[61]}), .Q ({new_AGEMA_signal_1347, TweakeyGeneration_key_Feedback[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1442, TweakeyGeneration_StateRegInput[60]}), .Q ({new_AGEMA_signal_1344, TweakeyGeneration_key_Feedback[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1439, TweakeyGeneration_StateRegInput[59]}), .Q ({new_AGEMA_signal_1341, TweakeyGeneration_key_Feedback[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1436, TweakeyGeneration_StateRegInput[58]}), .Q ({new_AGEMA_signal_1338, TweakeyGeneration_key_Feedback[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1433, TweakeyGeneration_StateRegInput[57]}), .Q ({new_AGEMA_signal_1335, TweakeyGeneration_key_Feedback[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1430, TweakeyGeneration_StateRegInput[56]}), .Q ({new_AGEMA_signal_1332, TweakeyGeneration_key_Feedback[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1427, TweakeyGeneration_StateRegInput[55]}), .Q ({new_AGEMA_signal_1329, TweakeyGeneration_key_Feedback[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1424, TweakeyGeneration_StateRegInput[54]}), .Q ({new_AGEMA_signal_1326, TweakeyGeneration_key_Feedback[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1421, TweakeyGeneration_StateRegInput[53]}), .Q ({new_AGEMA_signal_1323, TweakeyGeneration_key_Feedback[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1418, TweakeyGeneration_StateRegInput[52]}), .Q ({new_AGEMA_signal_1320, TweakeyGeneration_key_Feedback[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1415, TweakeyGeneration_StateRegInput[51]}), .Q ({new_AGEMA_signal_1317, TweakeyGeneration_key_Feedback[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1412, TweakeyGeneration_StateRegInput[50]}), .Q ({new_AGEMA_signal_1314, TweakeyGeneration_key_Feedback[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1409, TweakeyGeneration_StateRegInput[49]}), .Q ({new_AGEMA_signal_1311, TweakeyGeneration_key_Feedback[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1406, TweakeyGeneration_StateRegInput[48]}), .Q ({new_AGEMA_signal_1308, TweakeyGeneration_key_Feedback[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1403, TweakeyGeneration_StateRegInput[47]}), .Q ({new_AGEMA_signal_1305, TweakeyGeneration_key_Feedback[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1400, TweakeyGeneration_StateRegInput[46]}), .Q ({new_AGEMA_signal_1302, TweakeyGeneration_key_Feedback[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1397, TweakeyGeneration_StateRegInput[45]}), .Q ({new_AGEMA_signal_1299, TweakeyGeneration_key_Feedback[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1394, TweakeyGeneration_StateRegInput[44]}), .Q ({new_AGEMA_signal_1296, TweakeyGeneration_key_Feedback[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1391, TweakeyGeneration_StateRegInput[43]}), .Q ({new_AGEMA_signal_1293, TweakeyGeneration_key_Feedback[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1388, TweakeyGeneration_StateRegInput[42]}), .Q ({new_AGEMA_signal_1290, TweakeyGeneration_key_Feedback[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1385, TweakeyGeneration_StateRegInput[41]}), .Q ({new_AGEMA_signal_1287, TweakeyGeneration_key_Feedback[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1382, TweakeyGeneration_StateRegInput[40]}), .Q ({new_AGEMA_signal_1284, TweakeyGeneration_key_Feedback[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1379, TweakeyGeneration_StateRegInput[39]}), .Q ({new_AGEMA_signal_1281, TweakeyGeneration_key_Feedback[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1376, TweakeyGeneration_StateRegInput[38]}), .Q ({new_AGEMA_signal_1278, TweakeyGeneration_key_Feedback[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1373, TweakeyGeneration_StateRegInput[37]}), .Q ({new_AGEMA_signal_1275, TweakeyGeneration_key_Feedback[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1370, TweakeyGeneration_StateRegInput[36]}), .Q ({new_AGEMA_signal_1272, TweakeyGeneration_key_Feedback[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1367, TweakeyGeneration_StateRegInput[35]}), .Q ({new_AGEMA_signal_1269, TweakeyGeneration_key_Feedback[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1364, TweakeyGeneration_StateRegInput[34]}), .Q ({new_AGEMA_signal_1266, TweakeyGeneration_key_Feedback[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1361, TweakeyGeneration_StateRegInput[33]}), .Q ({new_AGEMA_signal_1263, TweakeyGeneration_key_Feedback[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1358, TweakeyGeneration_StateRegInput[32]}), .Q ({new_AGEMA_signal_1260, TweakeyGeneration_key_Feedback[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1355, TweakeyGeneration_StateRegInput[31]}), .Q ({new_AGEMA_signal_1425, TweakeyGeneration_key_Feedback[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1352, TweakeyGeneration_StateRegInput[30]}), .Q ({new_AGEMA_signal_1422, TweakeyGeneration_key_Feedback[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1349, TweakeyGeneration_StateRegInput[29]}), .Q ({new_AGEMA_signal_1419, TweakeyGeneration_key_Feedback[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1346, TweakeyGeneration_StateRegInput[28]}), .Q ({new_AGEMA_signal_1416, TweakeyGeneration_key_Feedback[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1343, TweakeyGeneration_StateRegInput[27]}), .Q ({new_AGEMA_signal_1449, TweakeyGeneration_key_Feedback[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1340, TweakeyGeneration_StateRegInput[26]}), .Q ({new_AGEMA_signal_1446, TweakeyGeneration_key_Feedback[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1337, TweakeyGeneration_StateRegInput[25]}), .Q ({new_AGEMA_signal_1443, TweakeyGeneration_key_Feedback[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1334, TweakeyGeneration_StateRegInput[24]}), .Q ({new_AGEMA_signal_1440, TweakeyGeneration_key_Feedback[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1331, TweakeyGeneration_StateRegInput[23]}), .Q ({new_AGEMA_signal_1401, TweakeyGeneration_key_Feedback[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1328, TweakeyGeneration_StateRegInput[22]}), .Q ({new_AGEMA_signal_1398, TweakeyGeneration_key_Feedback[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1325, TweakeyGeneration_StateRegInput[21]}), .Q ({new_AGEMA_signal_1395, TweakeyGeneration_key_Feedback[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1322, TweakeyGeneration_StateRegInput[20]}), .Q ({new_AGEMA_signal_1392, TweakeyGeneration_key_Feedback[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1319, TweakeyGeneration_StateRegInput[19]}), .Q ({new_AGEMA_signal_1365, TweakeyGeneration_key_Feedback[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1316, TweakeyGeneration_StateRegInput[18]}), .Q ({new_AGEMA_signal_1362, TweakeyGeneration_key_Feedback[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1313, TweakeyGeneration_StateRegInput[17]}), .Q ({new_AGEMA_signal_1359, TweakeyGeneration_key_Feedback[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1310, TweakeyGeneration_StateRegInput[16]}), .Q ({new_AGEMA_signal_1356, TweakeyGeneration_key_Feedback[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1307, TweakeyGeneration_StateRegInput[15]}), .Q ({new_AGEMA_signal_1377, TweakeyGeneration_key_Feedback[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1304, TweakeyGeneration_StateRegInput[14]}), .Q ({new_AGEMA_signal_1374, TweakeyGeneration_key_Feedback[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1301, TweakeyGeneration_StateRegInput[13]}), .Q ({new_AGEMA_signal_1371, TweakeyGeneration_key_Feedback[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1298, TweakeyGeneration_StateRegInput[12]}), .Q ({new_AGEMA_signal_1368, TweakeyGeneration_key_Feedback[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1295, TweakeyGeneration_StateRegInput[11]}), .Q ({new_AGEMA_signal_1413, TweakeyGeneration_key_Feedback[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1292, TweakeyGeneration_StateRegInput[10]}), .Q ({new_AGEMA_signal_1410, TweakeyGeneration_key_Feedback[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1289, TweakeyGeneration_StateRegInput[9]}), .Q ({new_AGEMA_signal_1407, TweakeyGeneration_key_Feedback[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1286, TweakeyGeneration_StateRegInput[8]}), .Q ({new_AGEMA_signal_1404, TweakeyGeneration_key_Feedback[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1283, TweakeyGeneration_StateRegInput[7]}), .Q ({new_AGEMA_signal_1389, TweakeyGeneration_key_Feedback[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1280, TweakeyGeneration_StateRegInput[6]}), .Q ({new_AGEMA_signal_1386, TweakeyGeneration_key_Feedback[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1277, TweakeyGeneration_StateRegInput[5]}), .Q ({new_AGEMA_signal_1383, TweakeyGeneration_key_Feedback[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1274, TweakeyGeneration_StateRegInput[4]}), .Q ({new_AGEMA_signal_1380, TweakeyGeneration_key_Feedback[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1271, TweakeyGeneration_StateRegInput[3]}), .Q ({new_AGEMA_signal_1437, TweakeyGeneration_key_Feedback[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1268, TweakeyGeneration_StateRegInput[2]}), .Q ({new_AGEMA_signal_1434, TweakeyGeneration_key_Feedback[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1265, TweakeyGeneration_StateRegInput[1]}), .Q ({new_AGEMA_signal_1431, TweakeyGeneration_key_Feedback[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1262, TweakeyGeneration_StateRegInput[0]}), .Q ({new_AGEMA_signal_1428, TweakeyGeneration_key_Feedback[56]}) ) ;
    DFF_X1 FSMReg_s_current_state_reg_5__FF_FF ( .CK (clk_gated), .D (FSMSelected[5]), .Q (FSM[5]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_4__FF_FF ( .CK (clk_gated), .D (FSMSelected[4]), .Q (FSM[4]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_3__FF_FF ( .CK (clk_gated), .D (FSMSelected[3]), .Q (FSMUpdate[4]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_2__FF_FF ( .CK (clk_gated), .D (FSMSelected[2]), .Q (FSMUpdate[3]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_1__FF_FF ( .CK (clk_gated), .D (FSMSelected[1]), .Q (FSM[1]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_0__FF_FF ( .CK (clk_gated), .D (FSMSelected[0]), .Q (FSMUpdate[1]), .QN () ) ;
endmodule
