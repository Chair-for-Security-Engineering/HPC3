////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module Midori64 in file /AGEMA/Designs/Midori_round_based/AGEMA/Midori64.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module Midori64_HPC2_Pipeline_d2 (DataIn_s0, key_s0, clk, reset, enc_dec, key_s1, key_s2, DataIn_s1, DataIn_s2, Fresh, DataOut_s0, done, DataOut_s1, DataOut_s2);
    input [63:0] DataIn_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input enc_dec ;
    input [127:0] key_s1 ;
    input [127:0] key_s2 ;
    input [63:0] DataIn_s1 ;
    input [63:0] DataIn_s2 ;
    input [767:0] Fresh ;
    output [63:0] DataOut_s0 ;
    output done ;
    output [63:0] DataOut_s1 ;
    output [63:0] DataOut_s2 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4784 ;
    wire controller_n2 ;
    wire controller_n1 ;
    wire controller_roundCounter_n13 ;
    wire controller_roundCounter_n12 ;
    wire controller_roundCounter_n11 ;
    wire controller_roundCounter_n10 ;
    wire controller_roundCounter_n9 ;
    wire controller_roundCounter_n8 ;
    wire controller_roundCounter_n7 ;
    wire controller_roundCounter_n5 ;
    wire controller_roundCounter_n4 ;
    wire controller_roundCounter_n3 ;
    wire controller_roundCounter_n2 ;
    wire controller_roundCounter_n1 ;
    wire controller_roundCounter_N10 ;
    wire controller_roundCounter_n6 ;
    wire controller_roundCounter_N8 ;
    wire controller_roundCounter_N7 ;
    wire Midori_rounds_n16 ;
    wire Midori_rounds_n15 ;
    wire Midori_rounds_n14 ;
    wire Midori_rounds_n13 ;
    wire Midori_rounds_n12 ;
    wire Midori_rounds_n11 ;
    wire Midori_rounds_n10 ;
    wire Midori_rounds_n9 ;
    wire Midori_rounds_n8 ;
    wire Midori_rounds_n7 ;
    wire Midori_rounds_n6 ;
    wire Midori_rounds_n5 ;
    wire Midori_rounds_n4 ;
    wire Midori_rounds_n3 ;
    wire Midori_rounds_n2 ;
    wire Midori_rounds_n1 ;
    wire Midori_rounds_SelectedKey_0_ ;
    wire Midori_rounds_SelectedKey_1_ ;
    wire Midori_rounds_SelectedKey_2_ ;
    wire Midori_rounds_SelectedKey_3_ ;
    wire Midori_rounds_SelectedKey_4_ ;
    wire Midori_rounds_SelectedKey_5_ ;
    wire Midori_rounds_SelectedKey_6_ ;
    wire Midori_rounds_SelectedKey_7_ ;
    wire Midori_rounds_SelectedKey_8_ ;
    wire Midori_rounds_SelectedKey_9_ ;
    wire Midori_rounds_SelectedKey_10_ ;
    wire Midori_rounds_SelectedKey_11_ ;
    wire Midori_rounds_SelectedKey_12_ ;
    wire Midori_rounds_SelectedKey_13_ ;
    wire Midori_rounds_SelectedKey_14_ ;
    wire Midori_rounds_SelectedKey_15_ ;
    wire Midori_rounds_SelectedKey_16_ ;
    wire Midori_rounds_SelectedKey_17_ ;
    wire Midori_rounds_SelectedKey_18_ ;
    wire Midori_rounds_SelectedKey_19_ ;
    wire Midori_rounds_SelectedKey_20_ ;
    wire Midori_rounds_SelectedKey_21_ ;
    wire Midori_rounds_SelectedKey_22_ ;
    wire Midori_rounds_SelectedKey_23_ ;
    wire Midori_rounds_SelectedKey_24_ ;
    wire Midori_rounds_SelectedKey_25_ ;
    wire Midori_rounds_SelectedKey_26_ ;
    wire Midori_rounds_SelectedKey_27_ ;
    wire Midori_rounds_SelectedKey_28_ ;
    wire Midori_rounds_SelectedKey_29_ ;
    wire Midori_rounds_SelectedKey_30_ ;
    wire Midori_rounds_SelectedKey_31_ ;
    wire Midori_rounds_SelectedKey_32_ ;
    wire Midori_rounds_SelectedKey_33_ ;
    wire Midori_rounds_SelectedKey_34_ ;
    wire Midori_rounds_SelectedKey_35_ ;
    wire Midori_rounds_SelectedKey_36_ ;
    wire Midori_rounds_SelectedKey_37_ ;
    wire Midori_rounds_SelectedKey_38_ ;
    wire Midori_rounds_SelectedKey_39_ ;
    wire Midori_rounds_SelectedKey_40_ ;
    wire Midori_rounds_SelectedKey_41_ ;
    wire Midori_rounds_SelectedKey_42_ ;
    wire Midori_rounds_SelectedKey_43_ ;
    wire Midori_rounds_SelectedKey_44_ ;
    wire Midori_rounds_SelectedKey_45_ ;
    wire Midori_rounds_SelectedKey_46_ ;
    wire Midori_rounds_SelectedKey_47_ ;
    wire Midori_rounds_SelectedKey_48_ ;
    wire Midori_rounds_SelectedKey_49_ ;
    wire Midori_rounds_SelectedKey_50_ ;
    wire Midori_rounds_SelectedKey_51_ ;
    wire Midori_rounds_SelectedKey_52_ ;
    wire Midori_rounds_SelectedKey_53_ ;
    wire Midori_rounds_SelectedKey_54_ ;
    wire Midori_rounds_SelectedKey_55_ ;
    wire Midori_rounds_SelectedKey_56_ ;
    wire Midori_rounds_SelectedKey_57_ ;
    wire Midori_rounds_SelectedKey_58_ ;
    wire Midori_rounds_SelectedKey_59_ ;
    wire Midori_rounds_SelectedKey_60_ ;
    wire Midori_rounds_SelectedKey_61_ ;
    wire Midori_rounds_SelectedKey_62_ ;
    wire Midori_rounds_SelectedKey_63_ ;
    wire Midori_rounds_constant_MUX_n217 ;
    wire Midori_rounds_constant_MUX_n216 ;
    wire Midori_rounds_constant_MUX_n215 ;
    wire Midori_rounds_constant_MUX_n214 ;
    wire Midori_rounds_constant_MUX_n213 ;
    wire Midori_rounds_constant_MUX_n212 ;
    wire Midori_rounds_constant_MUX_n211 ;
    wire Midori_rounds_constant_MUX_n210 ;
    wire Midori_rounds_constant_MUX_n209 ;
    wire Midori_rounds_constant_MUX_n208 ;
    wire Midori_rounds_constant_MUX_n207 ;
    wire Midori_rounds_constant_MUX_n206 ;
    wire Midori_rounds_constant_MUX_n205 ;
    wire Midori_rounds_constant_MUX_n204 ;
    wire Midori_rounds_constant_MUX_n203 ;
    wire Midori_rounds_constant_MUX_n202 ;
    wire Midori_rounds_constant_MUX_n201 ;
    wire Midori_rounds_constant_MUX_n200 ;
    wire Midori_rounds_constant_MUX_n199 ;
    wire Midori_rounds_constant_MUX_n198 ;
    wire Midori_rounds_constant_MUX_n197 ;
    wire Midori_rounds_constant_MUX_n196 ;
    wire Midori_rounds_constant_MUX_n195 ;
    wire Midori_rounds_constant_MUX_n194 ;
    wire Midori_rounds_constant_MUX_n193 ;
    wire Midori_rounds_constant_MUX_n192 ;
    wire Midori_rounds_constant_MUX_n191 ;
    wire Midori_rounds_constant_MUX_n190 ;
    wire Midori_rounds_constant_MUX_n189 ;
    wire Midori_rounds_constant_MUX_n188 ;
    wire Midori_rounds_constant_MUX_n187 ;
    wire Midori_rounds_constant_MUX_n186 ;
    wire Midori_rounds_constant_MUX_n185 ;
    wire Midori_rounds_constant_MUX_n184 ;
    wire Midori_rounds_constant_MUX_n183 ;
    wire Midori_rounds_constant_MUX_n182 ;
    wire Midori_rounds_constant_MUX_n181 ;
    wire Midori_rounds_constant_MUX_n180 ;
    wire Midori_rounds_constant_MUX_n179 ;
    wire Midori_rounds_constant_MUX_n178 ;
    wire Midori_rounds_constant_MUX_n177 ;
    wire Midori_rounds_constant_MUX_n176 ;
    wire Midori_rounds_constant_MUX_n175 ;
    wire Midori_rounds_constant_MUX_n174 ;
    wire Midori_rounds_constant_MUX_n173 ;
    wire Midori_rounds_constant_MUX_n172 ;
    wire Midori_rounds_constant_MUX_n171 ;
    wire Midori_rounds_constant_MUX_n170 ;
    wire Midori_rounds_constant_MUX_n169 ;
    wire Midori_rounds_constant_MUX_n168 ;
    wire Midori_rounds_constant_MUX_n167 ;
    wire Midori_rounds_constant_MUX_n166 ;
    wire Midori_rounds_constant_MUX_n165 ;
    wire Midori_rounds_constant_MUX_n164 ;
    wire Midori_rounds_constant_MUX_n163 ;
    wire Midori_rounds_constant_MUX_n162 ;
    wire Midori_rounds_constant_MUX_n161 ;
    wire Midori_rounds_constant_MUX_n160 ;
    wire Midori_rounds_constant_MUX_n159 ;
    wire Midori_rounds_constant_MUX_n158 ;
    wire Midori_rounds_constant_MUX_n157 ;
    wire Midori_rounds_constant_MUX_n156 ;
    wire Midori_rounds_constant_MUX_n155 ;
    wire Midori_rounds_constant_MUX_n154 ;
    wire Midori_rounds_constant_MUX_n153 ;
    wire Midori_rounds_constant_MUX_n152 ;
    wire Midori_rounds_constant_MUX_n151 ;
    wire Midori_rounds_constant_MUX_n150 ;
    wire Midori_rounds_constant_MUX_n149 ;
    wire Midori_rounds_constant_MUX_n148 ;
    wire Midori_rounds_constant_MUX_n147 ;
    wire Midori_rounds_constant_MUX_n146 ;
    wire Midori_rounds_constant_MUX_n145 ;
    wire Midori_rounds_constant_MUX_n144 ;
    wire Midori_rounds_constant_MUX_n143 ;
    wire Midori_rounds_constant_MUX_n142 ;
    wire Midori_rounds_constant_MUX_n141 ;
    wire Midori_rounds_constant_MUX_n140 ;
    wire Midori_rounds_constant_MUX_n139 ;
    wire Midori_rounds_constant_MUX_n138 ;
    wire Midori_rounds_constant_MUX_n137 ;
    wire Midori_rounds_constant_MUX_n136 ;
    wire Midori_rounds_constant_MUX_n135 ;
    wire Midori_rounds_constant_MUX_n134 ;
    wire Midori_rounds_constant_MUX_n133 ;
    wire Midori_rounds_constant_MUX_n132 ;
    wire Midori_rounds_constant_MUX_n131 ;
    wire Midori_rounds_constant_MUX_n130 ;
    wire Midori_rounds_constant_MUX_n129 ;
    wire Midori_rounds_constant_MUX_n128 ;
    wire Midori_rounds_MUXInst_n11 ;
    wire Midori_rounds_MUXInst_n10 ;
    wire Midori_rounds_MUXInst_n9 ;
    wire Midori_rounds_MUXInst_n8 ;
    wire Midori_rounds_roundResult_Reg_SFF_0_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_1_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_2_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_3_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_4_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_5_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_6_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_7_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_8_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_9_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_10_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_11_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_12_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_13_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_14_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_15_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_16_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_17_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_18_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_19_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_20_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_21_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_22_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_23_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_24_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_25_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_26_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_27_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_28_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_29_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_30_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_31_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_32_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_33_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_34_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_35_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_36_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_37_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_38_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_39_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_40_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_41_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_42_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_43_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_44_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_45_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_46_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_47_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_48_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_49_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_50_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_51_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_52_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_53_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_54_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_55_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_56_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_57_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_58_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_59_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_60_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_61_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_62_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_63_DQ ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n1 ;
    wire Midori_rounds_mul_MC1_n8 ;
    wire Midori_rounds_mul_MC1_n7 ;
    wire Midori_rounds_mul_MC1_n6 ;
    wire Midori_rounds_mul_MC1_n5 ;
    wire Midori_rounds_mul_MC1_n4 ;
    wire Midori_rounds_mul_MC1_n3 ;
    wire Midori_rounds_mul_MC1_n2 ;
    wire Midori_rounds_mul_MC1_n1 ;
    wire Midori_rounds_mul_MC2_n8 ;
    wire Midori_rounds_mul_MC2_n7 ;
    wire Midori_rounds_mul_MC2_n6 ;
    wire Midori_rounds_mul_MC2_n5 ;
    wire Midori_rounds_mul_MC2_n4 ;
    wire Midori_rounds_mul_MC2_n3 ;
    wire Midori_rounds_mul_MC2_n2 ;
    wire Midori_rounds_mul_MC2_n1 ;
    wire Midori_rounds_mul_MC3_n8 ;
    wire Midori_rounds_mul_MC3_n7 ;
    wire Midori_rounds_mul_MC3_n6 ;
    wire Midori_rounds_mul_MC3_n5 ;
    wire Midori_rounds_mul_MC3_n4 ;
    wire Midori_rounds_mul_MC3_n3 ;
    wire Midori_rounds_mul_MC3_n2 ;
    wire Midori_rounds_mul_MC3_n1 ;
    wire Midori_rounds_mul_MC4_n8 ;
    wire Midori_rounds_mul_MC4_n7 ;
    wire Midori_rounds_mul_MC4_n6 ;
    wire Midori_rounds_mul_MC4_n5 ;
    wire Midori_rounds_mul_MC4_n4 ;
    wire Midori_rounds_mul_MC4_n3 ;
    wire Midori_rounds_mul_MC4_n2 ;
    wire Midori_rounds_mul_MC4_n1 ;
    wire [63:0] wk ;
    wire [3:0] round_Signal ;
    wire [63:0] Midori_add_Result_Start ;
    wire [63:0] Midori_rounds_mul_ResultXORkey ;
    wire [63:0] Midori_rounds_SR_Inv_Result ;
    wire [63:0] Midori_rounds_mul_input ;
    wire [63:0] Midori_rounds_sub_ResultXORkey ;
    wire [63:0] Midori_rounds_SR_Result ;
    wire [63:0] Midori_rounds_roundReg_out ;
    wire [63:0] Midori_rounds_round_Result ;
    wire [15:0] Midori_rounds_round_Constant ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5195 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5202 ;
    wire new_AGEMA_signal_5203 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5207 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5213 ;
    wire new_AGEMA_signal_5214 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5219 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5226 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5231 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5238 ;
    wire new_AGEMA_signal_5239 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5249 ;
    wire new_AGEMA_signal_5250 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5255 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5262 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5273 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5291 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5303 ;
    wire new_AGEMA_signal_5304 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5309 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6654 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;
    wire new_AGEMA_signal_6672 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6677 ;
    wire new_AGEMA_signal_6678 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6682 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6688 ;
    wire new_AGEMA_signal_6689 ;
    wire new_AGEMA_signal_6690 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6695 ;
    wire new_AGEMA_signal_6696 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6700 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6706 ;
    wire new_AGEMA_signal_6707 ;
    wire new_AGEMA_signal_6708 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6713 ;
    wire new_AGEMA_signal_6714 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6718 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6724 ;
    wire new_AGEMA_signal_6725 ;
    wire new_AGEMA_signal_6726 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7036 ;
    wire new_AGEMA_signal_7037 ;
    wire new_AGEMA_signal_7038 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7042 ;
    wire new_AGEMA_signal_7043 ;
    wire new_AGEMA_signal_7044 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7048 ;
    wire new_AGEMA_signal_7049 ;
    wire new_AGEMA_signal_7050 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7054 ;
    wire new_AGEMA_signal_7055 ;
    wire new_AGEMA_signal_7056 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7060 ;
    wire new_AGEMA_signal_7061 ;
    wire new_AGEMA_signal_7062 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7066 ;
    wire new_AGEMA_signal_7067 ;
    wire new_AGEMA_signal_7068 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7072 ;
    wire new_AGEMA_signal_7073 ;
    wire new_AGEMA_signal_7074 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7078 ;
    wire new_AGEMA_signal_7079 ;
    wire new_AGEMA_signal_7080 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7084 ;
    wire new_AGEMA_signal_7085 ;
    wire new_AGEMA_signal_7086 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7090 ;
    wire new_AGEMA_signal_7091 ;
    wire new_AGEMA_signal_7092 ;
    wire new_AGEMA_signal_7093 ;
    wire new_AGEMA_signal_7094 ;
    wire new_AGEMA_signal_7095 ;
    wire new_AGEMA_signal_7096 ;
    wire new_AGEMA_signal_7097 ;
    wire new_AGEMA_signal_7098 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7102 ;
    wire new_AGEMA_signal_7103 ;
    wire new_AGEMA_signal_7104 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7108 ;
    wire new_AGEMA_signal_7109 ;
    wire new_AGEMA_signal_7110 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7114 ;
    wire new_AGEMA_signal_7115 ;
    wire new_AGEMA_signal_7116 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7120 ;
    wire new_AGEMA_signal_7121 ;
    wire new_AGEMA_signal_7122 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7126 ;
    wire new_AGEMA_signal_7127 ;
    wire new_AGEMA_signal_7128 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7132 ;
    wire new_AGEMA_signal_7133 ;
    wire new_AGEMA_signal_7134 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7138 ;
    wire new_AGEMA_signal_7139 ;
    wire new_AGEMA_signal_7140 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7144 ;
    wire new_AGEMA_signal_7145 ;
    wire new_AGEMA_signal_7146 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7150 ;
    wire new_AGEMA_signal_7151 ;
    wire new_AGEMA_signal_7152 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7156 ;
    wire new_AGEMA_signal_7157 ;
    wire new_AGEMA_signal_7158 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7162 ;
    wire new_AGEMA_signal_7163 ;
    wire new_AGEMA_signal_7164 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7168 ;
    wire new_AGEMA_signal_7169 ;
    wire new_AGEMA_signal_7170 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7174 ;
    wire new_AGEMA_signal_7175 ;
    wire new_AGEMA_signal_7176 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7180 ;
    wire new_AGEMA_signal_7181 ;
    wire new_AGEMA_signal_7182 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7186 ;
    wire new_AGEMA_signal_7187 ;
    wire new_AGEMA_signal_7188 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7192 ;
    wire new_AGEMA_signal_7193 ;
    wire new_AGEMA_signal_7194 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7198 ;
    wire new_AGEMA_signal_7199 ;
    wire new_AGEMA_signal_7200 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7204 ;
    wire new_AGEMA_signal_7205 ;
    wire new_AGEMA_signal_7206 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7489 ;
    wire new_AGEMA_signal_7490 ;
    wire new_AGEMA_signal_7491 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7495 ;
    wire new_AGEMA_signal_7496 ;
    wire new_AGEMA_signal_7497 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7499 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7501 ;
    wire new_AGEMA_signal_7502 ;
    wire new_AGEMA_signal_7503 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7507 ;
    wire new_AGEMA_signal_7508 ;
    wire new_AGEMA_signal_7509 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7513 ;
    wire new_AGEMA_signal_7514 ;
    wire new_AGEMA_signal_7515 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7519 ;
    wire new_AGEMA_signal_7520 ;
    wire new_AGEMA_signal_7521 ;
    wire new_AGEMA_signal_7522 ;
    wire new_AGEMA_signal_7523 ;
    wire new_AGEMA_signal_7524 ;
    wire new_AGEMA_signal_7525 ;
    wire new_AGEMA_signal_7526 ;
    wire new_AGEMA_signal_7527 ;
    wire new_AGEMA_signal_7528 ;
    wire new_AGEMA_signal_7529 ;
    wire new_AGEMA_signal_7530 ;
    wire new_AGEMA_signal_7531 ;
    wire new_AGEMA_signal_7532 ;
    wire new_AGEMA_signal_7533 ;
    wire new_AGEMA_signal_7534 ;
    wire new_AGEMA_signal_7535 ;
    wire new_AGEMA_signal_7536 ;
    wire new_AGEMA_signal_7537 ;
    wire new_AGEMA_signal_7538 ;
    wire new_AGEMA_signal_7539 ;
    wire new_AGEMA_signal_7540 ;
    wire new_AGEMA_signal_7541 ;
    wire new_AGEMA_signal_7542 ;
    wire new_AGEMA_signal_7543 ;
    wire new_AGEMA_signal_7544 ;
    wire new_AGEMA_signal_7545 ;
    wire new_AGEMA_signal_7546 ;
    wire new_AGEMA_signal_7547 ;
    wire new_AGEMA_signal_7548 ;
    wire new_AGEMA_signal_7549 ;
    wire new_AGEMA_signal_7550 ;
    wire new_AGEMA_signal_7551 ;
    wire new_AGEMA_signal_7552 ;
    wire new_AGEMA_signal_7553 ;
    wire new_AGEMA_signal_7554 ;
    wire new_AGEMA_signal_7555 ;
    wire new_AGEMA_signal_7556 ;
    wire new_AGEMA_signal_7557 ;
    wire new_AGEMA_signal_7558 ;
    wire new_AGEMA_signal_7559 ;
    wire new_AGEMA_signal_7560 ;
    wire new_AGEMA_signal_7561 ;
    wire new_AGEMA_signal_7562 ;
    wire new_AGEMA_signal_7563 ;
    wire new_AGEMA_signal_7564 ;
    wire new_AGEMA_signal_7565 ;
    wire new_AGEMA_signal_7566 ;
    wire new_AGEMA_signal_7567 ;
    wire new_AGEMA_signal_7568 ;
    wire new_AGEMA_signal_7569 ;
    wire new_AGEMA_signal_7570 ;
    wire new_AGEMA_signal_7571 ;
    wire new_AGEMA_signal_7572 ;
    wire new_AGEMA_signal_7573 ;
    wire new_AGEMA_signal_7574 ;
    wire new_AGEMA_signal_7575 ;
    wire new_AGEMA_signal_7576 ;
    wire new_AGEMA_signal_7577 ;
    wire new_AGEMA_signal_7578 ;
    wire new_AGEMA_signal_7579 ;
    wire new_AGEMA_signal_7580 ;
    wire new_AGEMA_signal_7581 ;
    wire new_AGEMA_signal_7582 ;
    wire new_AGEMA_signal_7583 ;
    wire new_AGEMA_signal_7584 ;
    wire new_AGEMA_signal_7585 ;
    wire new_AGEMA_signal_7586 ;
    wire new_AGEMA_signal_7587 ;
    wire new_AGEMA_signal_7588 ;
    wire new_AGEMA_signal_7589 ;
    wire new_AGEMA_signal_7590 ;
    wire new_AGEMA_signal_7591 ;
    wire new_AGEMA_signal_7592 ;
    wire new_AGEMA_signal_7593 ;
    wire new_AGEMA_signal_7594 ;
    wire new_AGEMA_signal_7595 ;
    wire new_AGEMA_signal_7596 ;
    wire new_AGEMA_signal_7597 ;
    wire new_AGEMA_signal_7598 ;
    wire new_AGEMA_signal_7599 ;
    wire new_AGEMA_signal_7600 ;
    wire new_AGEMA_signal_7601 ;
    wire new_AGEMA_signal_7602 ;
    wire new_AGEMA_signal_7603 ;
    wire new_AGEMA_signal_7604 ;
    wire new_AGEMA_signal_7605 ;
    wire new_AGEMA_signal_7606 ;
    wire new_AGEMA_signal_7607 ;
    wire new_AGEMA_signal_7608 ;
    wire new_AGEMA_signal_7609 ;
    wire new_AGEMA_signal_7610 ;
    wire new_AGEMA_signal_7611 ;
    wire new_AGEMA_signal_7612 ;
    wire new_AGEMA_signal_7613 ;
    wire new_AGEMA_signal_7614 ;
    wire new_AGEMA_signal_7615 ;
    wire new_AGEMA_signal_7616 ;
    wire new_AGEMA_signal_7617 ;
    wire new_AGEMA_signal_7618 ;
    wire new_AGEMA_signal_7619 ;
    wire new_AGEMA_signal_7620 ;
    wire new_AGEMA_signal_7621 ;
    wire new_AGEMA_signal_7622 ;
    wire new_AGEMA_signal_7623 ;
    wire new_AGEMA_signal_7624 ;
    wire new_AGEMA_signal_7625 ;
    wire new_AGEMA_signal_7626 ;
    wire new_AGEMA_signal_7627 ;
    wire new_AGEMA_signal_7628 ;
    wire new_AGEMA_signal_7629 ;
    wire new_AGEMA_signal_7630 ;
    wire new_AGEMA_signal_7631 ;
    wire new_AGEMA_signal_7632 ;
    wire new_AGEMA_signal_7633 ;
    wire new_AGEMA_signal_7634 ;
    wire new_AGEMA_signal_7635 ;
    wire new_AGEMA_signal_7636 ;
    wire new_AGEMA_signal_7637 ;
    wire new_AGEMA_signal_7638 ;
    wire new_AGEMA_signal_7639 ;
    wire new_AGEMA_signal_7640 ;
    wire new_AGEMA_signal_7641 ;
    wire new_AGEMA_signal_7642 ;
    wire new_AGEMA_signal_7643 ;
    wire new_AGEMA_signal_7644 ;
    wire new_AGEMA_signal_7645 ;
    wire new_AGEMA_signal_7646 ;
    wire new_AGEMA_signal_7647 ;
    wire new_AGEMA_signal_7648 ;
    wire new_AGEMA_signal_7649 ;
    wire new_AGEMA_signal_7650 ;
    wire new_AGEMA_signal_7651 ;
    wire new_AGEMA_signal_7652 ;
    wire new_AGEMA_signal_7653 ;
    wire new_AGEMA_signal_7654 ;
    wire new_AGEMA_signal_7655 ;
    wire new_AGEMA_signal_7656 ;
    wire new_AGEMA_signal_7657 ;
    wire new_AGEMA_signal_7658 ;
    wire new_AGEMA_signal_7659 ;
    wire new_AGEMA_signal_7660 ;
    wire new_AGEMA_signal_7661 ;
    wire new_AGEMA_signal_7662 ;
    wire new_AGEMA_signal_7663 ;
    wire new_AGEMA_signal_7664 ;
    wire new_AGEMA_signal_7665 ;
    wire new_AGEMA_signal_7666 ;
    wire new_AGEMA_signal_7667 ;
    wire new_AGEMA_signal_7668 ;
    wire new_AGEMA_signal_7669 ;
    wire new_AGEMA_signal_7670 ;
    wire new_AGEMA_signal_7671 ;
    wire new_AGEMA_signal_7672 ;
    wire new_AGEMA_signal_7673 ;
    wire new_AGEMA_signal_7674 ;
    wire new_AGEMA_signal_7675 ;
    wire new_AGEMA_signal_7676 ;
    wire new_AGEMA_signal_7677 ;
    wire new_AGEMA_signal_7678 ;
    wire new_AGEMA_signal_7679 ;
    wire new_AGEMA_signal_7680 ;
    wire new_AGEMA_signal_7681 ;
    wire new_AGEMA_signal_7682 ;
    wire new_AGEMA_signal_7683 ;
    wire new_AGEMA_signal_7684 ;
    wire new_AGEMA_signal_7685 ;
    wire new_AGEMA_signal_7686 ;
    wire new_AGEMA_signal_7687 ;
    wire new_AGEMA_signal_7688 ;
    wire new_AGEMA_signal_7689 ;
    wire new_AGEMA_signal_7690 ;
    wire new_AGEMA_signal_7691 ;
    wire new_AGEMA_signal_7692 ;
    wire new_AGEMA_signal_7693 ;
    wire new_AGEMA_signal_7694 ;
    wire new_AGEMA_signal_7695 ;
    wire new_AGEMA_signal_7696 ;
    wire new_AGEMA_signal_7697 ;
    wire new_AGEMA_signal_7698 ;
    wire new_AGEMA_signal_7699 ;
    wire new_AGEMA_signal_7700 ;
    wire new_AGEMA_signal_7701 ;
    wire new_AGEMA_signal_7702 ;
    wire new_AGEMA_signal_7703 ;
    wire new_AGEMA_signal_7704 ;
    wire new_AGEMA_signal_7705 ;
    wire new_AGEMA_signal_7706 ;
    wire new_AGEMA_signal_7707 ;
    wire new_AGEMA_signal_7708 ;
    wire new_AGEMA_signal_7709 ;
    wire new_AGEMA_signal_7710 ;
    wire new_AGEMA_signal_7711 ;
    wire new_AGEMA_signal_7712 ;
    wire new_AGEMA_signal_7713 ;
    wire new_AGEMA_signal_7714 ;
    wire new_AGEMA_signal_7715 ;
    wire new_AGEMA_signal_7716 ;
    wire new_AGEMA_signal_7717 ;
    wire new_AGEMA_signal_7718 ;
    wire new_AGEMA_signal_7719 ;
    wire new_AGEMA_signal_7720 ;
    wire new_AGEMA_signal_7721 ;
    wire new_AGEMA_signal_7722 ;
    wire new_AGEMA_signal_7723 ;
    wire new_AGEMA_signal_7724 ;
    wire new_AGEMA_signal_7725 ;
    wire new_AGEMA_signal_7726 ;
    wire new_AGEMA_signal_7727 ;
    wire new_AGEMA_signal_7728 ;
    wire new_AGEMA_signal_7729 ;
    wire new_AGEMA_signal_7730 ;
    wire new_AGEMA_signal_7731 ;
    wire new_AGEMA_signal_7732 ;
    wire new_AGEMA_signal_7733 ;
    wire new_AGEMA_signal_7734 ;
    wire new_AGEMA_signal_7735 ;
    wire new_AGEMA_signal_7736 ;
    wire new_AGEMA_signal_7737 ;
    wire new_AGEMA_signal_7738 ;
    wire new_AGEMA_signal_7739 ;
    wire new_AGEMA_signal_7740 ;
    wire new_AGEMA_signal_7741 ;
    wire new_AGEMA_signal_7742 ;
    wire new_AGEMA_signal_7743 ;
    wire new_AGEMA_signal_7744 ;
    wire new_AGEMA_signal_7745 ;
    wire new_AGEMA_signal_7746 ;
    wire new_AGEMA_signal_7747 ;
    wire new_AGEMA_signal_7748 ;
    wire new_AGEMA_signal_7749 ;
    wire new_AGEMA_signal_7750 ;
    wire new_AGEMA_signal_7751 ;
    wire new_AGEMA_signal_7752 ;
    wire new_AGEMA_signal_7753 ;
    wire new_AGEMA_signal_7754 ;
    wire new_AGEMA_signal_7755 ;
    wire new_AGEMA_signal_7756 ;
    wire new_AGEMA_signal_7757 ;
    wire new_AGEMA_signal_7758 ;
    wire new_AGEMA_signal_7759 ;
    wire new_AGEMA_signal_7760 ;
    wire new_AGEMA_signal_7761 ;
    wire new_AGEMA_signal_7762 ;
    wire new_AGEMA_signal_7763 ;
    wire new_AGEMA_signal_7764 ;
    wire new_AGEMA_signal_7765 ;
    wire new_AGEMA_signal_7766 ;
    wire new_AGEMA_signal_7767 ;
    wire new_AGEMA_signal_7768 ;
    wire new_AGEMA_signal_7769 ;
    wire new_AGEMA_signal_7770 ;
    wire new_AGEMA_signal_7771 ;
    wire new_AGEMA_signal_7772 ;
    wire new_AGEMA_signal_7773 ;
    wire new_AGEMA_signal_7774 ;
    wire new_AGEMA_signal_7775 ;
    wire new_AGEMA_signal_7776 ;
    wire new_AGEMA_signal_7777 ;
    wire new_AGEMA_signal_7778 ;
    wire new_AGEMA_signal_7779 ;
    wire new_AGEMA_signal_7780 ;
    wire new_AGEMA_signal_7781 ;
    wire new_AGEMA_signal_7782 ;
    wire new_AGEMA_signal_7783 ;
    wire new_AGEMA_signal_7784 ;
    wire new_AGEMA_signal_7785 ;
    wire new_AGEMA_signal_7786 ;
    wire new_AGEMA_signal_7787 ;
    wire new_AGEMA_signal_7788 ;
    wire new_AGEMA_signal_7789 ;
    wire new_AGEMA_signal_7790 ;
    wire new_AGEMA_signal_7791 ;
    wire new_AGEMA_signal_7792 ;
    wire new_AGEMA_signal_7793 ;
    wire new_AGEMA_signal_7794 ;
    wire new_AGEMA_signal_7795 ;
    wire new_AGEMA_signal_7796 ;
    wire new_AGEMA_signal_7797 ;
    wire new_AGEMA_signal_7798 ;
    wire new_AGEMA_signal_7799 ;
    wire new_AGEMA_signal_7800 ;
    wire new_AGEMA_signal_7801 ;
    wire new_AGEMA_signal_7802 ;
    wire new_AGEMA_signal_7803 ;
    wire new_AGEMA_signal_7804 ;
    wire new_AGEMA_signal_7805 ;
    wire new_AGEMA_signal_7806 ;
    wire new_AGEMA_signal_7807 ;
    wire new_AGEMA_signal_7808 ;
    wire new_AGEMA_signal_7809 ;
    wire new_AGEMA_signal_7810 ;
    wire new_AGEMA_signal_7811 ;
    wire new_AGEMA_signal_7812 ;
    wire new_AGEMA_signal_7813 ;
    wire new_AGEMA_signal_7814 ;
    wire new_AGEMA_signal_7815 ;
    wire new_AGEMA_signal_7816 ;
    wire new_AGEMA_signal_7817 ;
    wire new_AGEMA_signal_7818 ;
    wire new_AGEMA_signal_7819 ;
    wire new_AGEMA_signal_7820 ;
    wire new_AGEMA_signal_7821 ;
    wire new_AGEMA_signal_7822 ;
    wire new_AGEMA_signal_7823 ;
    wire new_AGEMA_signal_7824 ;
    wire new_AGEMA_signal_7825 ;
    wire new_AGEMA_signal_7826 ;
    wire new_AGEMA_signal_7827 ;
    wire new_AGEMA_signal_7828 ;
    wire new_AGEMA_signal_7829 ;
    wire new_AGEMA_signal_7830 ;
    wire new_AGEMA_signal_7831 ;
    wire new_AGEMA_signal_7832 ;
    wire new_AGEMA_signal_7833 ;
    wire new_AGEMA_signal_7834 ;
    wire new_AGEMA_signal_7835 ;
    wire new_AGEMA_signal_7836 ;
    wire new_AGEMA_signal_7837 ;
    wire new_AGEMA_signal_7838 ;
    wire new_AGEMA_signal_7839 ;
    wire new_AGEMA_signal_7840 ;
    wire new_AGEMA_signal_7841 ;
    wire new_AGEMA_signal_7842 ;
    wire new_AGEMA_signal_7843 ;
    wire new_AGEMA_signal_7844 ;
    wire new_AGEMA_signal_7845 ;
    wire new_AGEMA_signal_7846 ;
    wire new_AGEMA_signal_7847 ;
    wire new_AGEMA_signal_7848 ;
    wire new_AGEMA_signal_7849 ;
    wire new_AGEMA_signal_7850 ;
    wire new_AGEMA_signal_7851 ;
    wire new_AGEMA_signal_7852 ;
    wire new_AGEMA_signal_7853 ;
    wire new_AGEMA_signal_7854 ;
    wire new_AGEMA_signal_7855 ;
    wire new_AGEMA_signal_7856 ;
    wire new_AGEMA_signal_7857 ;
    wire new_AGEMA_signal_7858 ;
    wire new_AGEMA_signal_7859 ;
    wire new_AGEMA_signal_7860 ;
    wire new_AGEMA_signal_7861 ;
    wire new_AGEMA_signal_7862 ;
    wire new_AGEMA_signal_7863 ;
    wire new_AGEMA_signal_7864 ;
    wire new_AGEMA_signal_7865 ;
    wire new_AGEMA_signal_7866 ;
    wire new_AGEMA_signal_7867 ;
    wire new_AGEMA_signal_7868 ;
    wire new_AGEMA_signal_7869 ;
    wire new_AGEMA_signal_7870 ;
    wire new_AGEMA_signal_7871 ;
    wire new_AGEMA_signal_7872 ;
    wire new_AGEMA_signal_7873 ;
    wire new_AGEMA_signal_7874 ;
    wire new_AGEMA_signal_7875 ;
    wire new_AGEMA_signal_7876 ;
    wire new_AGEMA_signal_7877 ;
    wire new_AGEMA_signal_7878 ;
    wire new_AGEMA_signal_7879 ;
    wire new_AGEMA_signal_7880 ;
    wire new_AGEMA_signal_7881 ;
    wire new_AGEMA_signal_7882 ;
    wire new_AGEMA_signal_7883 ;
    wire new_AGEMA_signal_7884 ;
    wire new_AGEMA_signal_7885 ;
    wire new_AGEMA_signal_7886 ;
    wire new_AGEMA_signal_7887 ;
    wire new_AGEMA_signal_7888 ;
    wire new_AGEMA_signal_7889 ;
    wire new_AGEMA_signal_7890 ;
    wire new_AGEMA_signal_7891 ;
    wire new_AGEMA_signal_7892 ;
    wire new_AGEMA_signal_7893 ;
    wire new_AGEMA_signal_7894 ;
    wire new_AGEMA_signal_7895 ;
    wire new_AGEMA_signal_7896 ;
    wire new_AGEMA_signal_7897 ;
    wire new_AGEMA_signal_7898 ;
    wire new_AGEMA_signal_7899 ;
    wire new_AGEMA_signal_7900 ;
    wire new_AGEMA_signal_7901 ;
    wire new_AGEMA_signal_7902 ;
    wire new_AGEMA_signal_7903 ;
    wire new_AGEMA_signal_7904 ;
    wire new_AGEMA_signal_7905 ;
    wire new_AGEMA_signal_7906 ;
    wire new_AGEMA_signal_7907 ;
    wire new_AGEMA_signal_7908 ;
    wire new_AGEMA_signal_7909 ;
    wire new_AGEMA_signal_7910 ;
    wire new_AGEMA_signal_7911 ;
    wire new_AGEMA_signal_7912 ;
    wire new_AGEMA_signal_7913 ;
    wire new_AGEMA_signal_7914 ;
    wire new_AGEMA_signal_7915 ;
    wire new_AGEMA_signal_7916 ;
    wire new_AGEMA_signal_7917 ;
    wire new_AGEMA_signal_7918 ;
    wire new_AGEMA_signal_7919 ;
    wire new_AGEMA_signal_7920 ;
    wire new_AGEMA_signal_7921 ;
    wire new_AGEMA_signal_7922 ;
    wire new_AGEMA_signal_7923 ;
    wire new_AGEMA_signal_7924 ;
    wire new_AGEMA_signal_7925 ;
    wire new_AGEMA_signal_7926 ;
    wire new_AGEMA_signal_7927 ;
    wire new_AGEMA_signal_7928 ;
    wire new_AGEMA_signal_7929 ;
    wire new_AGEMA_signal_7930 ;
    wire new_AGEMA_signal_7931 ;
    wire new_AGEMA_signal_7932 ;
    wire new_AGEMA_signal_7933 ;
    wire new_AGEMA_signal_7934 ;
    wire new_AGEMA_signal_7935 ;
    wire new_AGEMA_signal_7936 ;
    wire new_AGEMA_signal_7937 ;
    wire new_AGEMA_signal_7938 ;
    wire new_AGEMA_signal_7939 ;
    wire new_AGEMA_signal_7940 ;
    wire new_AGEMA_signal_7941 ;
    wire new_AGEMA_signal_7942 ;
    wire new_AGEMA_signal_7943 ;
    wire new_AGEMA_signal_7944 ;
    wire new_AGEMA_signal_7945 ;
    wire new_AGEMA_signal_7946 ;
    wire new_AGEMA_signal_7947 ;
    wire new_AGEMA_signal_7948 ;
    wire new_AGEMA_signal_7949 ;
    wire new_AGEMA_signal_7950 ;
    wire new_AGEMA_signal_7951 ;
    wire new_AGEMA_signal_7952 ;
    wire new_AGEMA_signal_7953 ;
    wire new_AGEMA_signal_7954 ;
    wire new_AGEMA_signal_7955 ;
    wire new_AGEMA_signal_7956 ;
    wire new_AGEMA_signal_7957 ;
    wire new_AGEMA_signal_7958 ;
    wire new_AGEMA_signal_7959 ;
    wire new_AGEMA_signal_7960 ;
    wire new_AGEMA_signal_7961 ;
    wire new_AGEMA_signal_7962 ;
    wire new_AGEMA_signal_7963 ;
    wire new_AGEMA_signal_7964 ;
    wire new_AGEMA_signal_7965 ;
    wire new_AGEMA_signal_7966 ;
    wire new_AGEMA_signal_7967 ;
    wire new_AGEMA_signal_7968 ;
    wire new_AGEMA_signal_7969 ;
    wire new_AGEMA_signal_7970 ;
    wire new_AGEMA_signal_7971 ;
    wire new_AGEMA_signal_7972 ;
    wire new_AGEMA_signal_7973 ;
    wire new_AGEMA_signal_7974 ;
    wire new_AGEMA_signal_7975 ;
    wire new_AGEMA_signal_7976 ;
    wire new_AGEMA_signal_7977 ;
    wire new_AGEMA_signal_7978 ;
    wire new_AGEMA_signal_7979 ;
    wire new_AGEMA_signal_7980 ;
    wire new_AGEMA_signal_7981 ;
    wire new_AGEMA_signal_7982 ;
    wire new_AGEMA_signal_7983 ;
    wire new_AGEMA_signal_7984 ;
    wire new_AGEMA_signal_7985 ;
    wire new_AGEMA_signal_7986 ;
    wire new_AGEMA_signal_7987 ;
    wire new_AGEMA_signal_7988 ;
    wire new_AGEMA_signal_7989 ;
    wire new_AGEMA_signal_7990 ;
    wire new_AGEMA_signal_7991 ;
    wire new_AGEMA_signal_7992 ;
    wire new_AGEMA_signal_7993 ;
    wire new_AGEMA_signal_7994 ;
    wire new_AGEMA_signal_7995 ;
    wire new_AGEMA_signal_7996 ;
    wire new_AGEMA_signal_7997 ;
    wire new_AGEMA_signal_7998 ;
    wire new_AGEMA_signal_7999 ;
    wire new_AGEMA_signal_8000 ;
    wire new_AGEMA_signal_8001 ;
    wire new_AGEMA_signal_8002 ;
    wire new_AGEMA_signal_8003 ;
    wire new_AGEMA_signal_8004 ;
    wire new_AGEMA_signal_8005 ;
    wire new_AGEMA_signal_8006 ;
    wire new_AGEMA_signal_8007 ;
    wire new_AGEMA_signal_8008 ;
    wire new_AGEMA_signal_8009 ;
    wire new_AGEMA_signal_8010 ;
    wire new_AGEMA_signal_8011 ;
    wire new_AGEMA_signal_8012 ;
    wire new_AGEMA_signal_8013 ;
    wire new_AGEMA_signal_8014 ;
    wire new_AGEMA_signal_8015 ;
    wire new_AGEMA_signal_8016 ;
    wire new_AGEMA_signal_8017 ;
    wire new_AGEMA_signal_8018 ;
    wire new_AGEMA_signal_8019 ;
    wire new_AGEMA_signal_8020 ;
    wire new_AGEMA_signal_8021 ;
    wire new_AGEMA_signal_8022 ;
    wire new_AGEMA_signal_8023 ;
    wire new_AGEMA_signal_8024 ;
    wire new_AGEMA_signal_8025 ;
    wire new_AGEMA_signal_8026 ;
    wire new_AGEMA_signal_8027 ;
    wire new_AGEMA_signal_8028 ;
    wire new_AGEMA_signal_8029 ;
    wire new_AGEMA_signal_8030 ;
    wire new_AGEMA_signal_8031 ;
    wire new_AGEMA_signal_8032 ;
    wire new_AGEMA_signal_8033 ;
    wire new_AGEMA_signal_8034 ;
    wire new_AGEMA_signal_8035 ;
    wire new_AGEMA_signal_8036 ;
    wire new_AGEMA_signal_8037 ;
    wire new_AGEMA_signal_8038 ;
    wire new_AGEMA_signal_8039 ;
    wire new_AGEMA_signal_8040 ;
    wire new_AGEMA_signal_8041 ;
    wire new_AGEMA_signal_8042 ;
    wire new_AGEMA_signal_8043 ;
    wire new_AGEMA_signal_8044 ;
    wire new_AGEMA_signal_8045 ;
    wire new_AGEMA_signal_8046 ;
    wire new_AGEMA_signal_8047 ;
    wire new_AGEMA_signal_8048 ;
    wire new_AGEMA_signal_8049 ;
    wire new_AGEMA_signal_8050 ;
    wire new_AGEMA_signal_8051 ;
    wire new_AGEMA_signal_8052 ;
    wire new_AGEMA_signal_8053 ;
    wire new_AGEMA_signal_8054 ;
    wire new_AGEMA_signal_8055 ;
    wire new_AGEMA_signal_8056 ;
    wire new_AGEMA_signal_8057 ;
    wire new_AGEMA_signal_8058 ;
    wire new_AGEMA_signal_8059 ;
    wire new_AGEMA_signal_8060 ;
    wire new_AGEMA_signal_8061 ;
    wire new_AGEMA_signal_8062 ;
    wire new_AGEMA_signal_8063 ;
    wire new_AGEMA_signal_8064 ;
    wire new_AGEMA_signal_8065 ;
    wire new_AGEMA_signal_8066 ;
    wire new_AGEMA_signal_8067 ;
    wire new_AGEMA_signal_8068 ;
    wire new_AGEMA_signal_8069 ;
    wire new_AGEMA_signal_8070 ;
    wire new_AGEMA_signal_8071 ;
    wire new_AGEMA_signal_8072 ;
    wire new_AGEMA_signal_8073 ;
    wire new_AGEMA_signal_8074 ;
    wire new_AGEMA_signal_8075 ;
    wire new_AGEMA_signal_8076 ;
    wire new_AGEMA_signal_8077 ;
    wire new_AGEMA_signal_8078 ;
    wire new_AGEMA_signal_8079 ;
    wire new_AGEMA_signal_8080 ;
    wire new_AGEMA_signal_8081 ;
    wire new_AGEMA_signal_8082 ;
    wire new_AGEMA_signal_8083 ;
    wire new_AGEMA_signal_8084 ;
    wire new_AGEMA_signal_8085 ;
    wire new_AGEMA_signal_8086 ;
    wire new_AGEMA_signal_8087 ;
    wire new_AGEMA_signal_8088 ;
    wire new_AGEMA_signal_8089 ;
    wire new_AGEMA_signal_8090 ;
    wire new_AGEMA_signal_8091 ;
    wire new_AGEMA_signal_8092 ;
    wire new_AGEMA_signal_8093 ;
    wire new_AGEMA_signal_8094 ;
    wire new_AGEMA_signal_8095 ;
    wire new_AGEMA_signal_8096 ;
    wire new_AGEMA_signal_8097 ;
    wire new_AGEMA_signal_8098 ;
    wire new_AGEMA_signal_8099 ;
    wire new_AGEMA_signal_8100 ;
    wire new_AGEMA_signal_8101 ;
    wire new_AGEMA_signal_8102 ;
    wire new_AGEMA_signal_8103 ;
    wire new_AGEMA_signal_8104 ;
    wire new_AGEMA_signal_8105 ;
    wire new_AGEMA_signal_8106 ;
    wire new_AGEMA_signal_8107 ;
    wire new_AGEMA_signal_8108 ;
    wire new_AGEMA_signal_8109 ;
    wire new_AGEMA_signal_8110 ;
    wire new_AGEMA_signal_8111 ;
    wire new_AGEMA_signal_8112 ;
    wire new_AGEMA_signal_8113 ;
    wire new_AGEMA_signal_8114 ;
    wire new_AGEMA_signal_8115 ;
    wire new_AGEMA_signal_8116 ;
    wire new_AGEMA_signal_8117 ;
    wire new_AGEMA_signal_8118 ;
    wire new_AGEMA_signal_8119 ;
    wire new_AGEMA_signal_8120 ;
    wire new_AGEMA_signal_8121 ;
    wire new_AGEMA_signal_8122 ;
    wire new_AGEMA_signal_8123 ;
    wire new_AGEMA_signal_8124 ;
    wire new_AGEMA_signal_8125 ;
    wire new_AGEMA_signal_8126 ;
    wire new_AGEMA_signal_8127 ;
    wire new_AGEMA_signal_8128 ;
    wire new_AGEMA_signal_8129 ;
    wire new_AGEMA_signal_8130 ;
    wire new_AGEMA_signal_8131 ;
    wire new_AGEMA_signal_8132 ;
    wire new_AGEMA_signal_8133 ;
    wire new_AGEMA_signal_8134 ;
    wire new_AGEMA_signal_8135 ;
    wire new_AGEMA_signal_8136 ;
    wire new_AGEMA_signal_8137 ;
    wire new_AGEMA_signal_8138 ;
    wire new_AGEMA_signal_8139 ;
    wire new_AGEMA_signal_8140 ;
    wire new_AGEMA_signal_8141 ;
    wire new_AGEMA_signal_8142 ;
    wire new_AGEMA_signal_8143 ;
    wire new_AGEMA_signal_8144 ;
    wire new_AGEMA_signal_8145 ;
    wire new_AGEMA_signal_8146 ;
    wire new_AGEMA_signal_8147 ;
    wire new_AGEMA_signal_8148 ;
    wire new_AGEMA_signal_8149 ;
    wire new_AGEMA_signal_8150 ;
    wire new_AGEMA_signal_8151 ;
    wire new_AGEMA_signal_8152 ;
    wire new_AGEMA_signal_8153 ;
    wire new_AGEMA_signal_8154 ;
    wire new_AGEMA_signal_8155 ;
    wire new_AGEMA_signal_8156 ;
    wire new_AGEMA_signal_8157 ;
    wire new_AGEMA_signal_8158 ;
    wire new_AGEMA_signal_8159 ;
    wire new_AGEMA_signal_8160 ;
    wire new_AGEMA_signal_8161 ;
    wire new_AGEMA_signal_8162 ;
    wire new_AGEMA_signal_8163 ;
    wire new_AGEMA_signal_8164 ;
    wire new_AGEMA_signal_8165 ;
    wire new_AGEMA_signal_8166 ;
    wire new_AGEMA_signal_8167 ;
    wire new_AGEMA_signal_8168 ;
    wire new_AGEMA_signal_8169 ;
    wire new_AGEMA_signal_8170 ;
    wire new_AGEMA_signal_8171 ;
    wire new_AGEMA_signal_8172 ;
    wire new_AGEMA_signal_8173 ;
    wire new_AGEMA_signal_8174 ;
    wire new_AGEMA_signal_8175 ;
    wire new_AGEMA_signal_8176 ;
    wire new_AGEMA_signal_8177 ;
    wire new_AGEMA_signal_8178 ;
    wire new_AGEMA_signal_8179 ;
    wire new_AGEMA_signal_8180 ;
    wire new_AGEMA_signal_8181 ;
    wire new_AGEMA_signal_8182 ;
    wire new_AGEMA_signal_8183 ;
    wire new_AGEMA_signal_8184 ;
    wire new_AGEMA_signal_8185 ;
    wire new_AGEMA_signal_8186 ;
    wire new_AGEMA_signal_8187 ;
    wire new_AGEMA_signal_8188 ;
    wire new_AGEMA_signal_8189 ;
    wire new_AGEMA_signal_8190 ;
    wire new_AGEMA_signal_8191 ;
    wire new_AGEMA_signal_8192 ;
    wire new_AGEMA_signal_8193 ;
    wire new_AGEMA_signal_8194 ;
    wire new_AGEMA_signal_8195 ;
    wire new_AGEMA_signal_8196 ;
    wire new_AGEMA_signal_8197 ;
    wire new_AGEMA_signal_8198 ;
    wire new_AGEMA_signal_8199 ;
    wire new_AGEMA_signal_8200 ;
    wire new_AGEMA_signal_8201 ;
    wire new_AGEMA_signal_8202 ;
    wire new_AGEMA_signal_8203 ;
    wire new_AGEMA_signal_8204 ;
    wire new_AGEMA_signal_8205 ;
    wire new_AGEMA_signal_8206 ;
    wire new_AGEMA_signal_8207 ;
    wire new_AGEMA_signal_8208 ;
    wire new_AGEMA_signal_8209 ;
    wire new_AGEMA_signal_8210 ;
    wire new_AGEMA_signal_8211 ;
    wire new_AGEMA_signal_8212 ;
    wire new_AGEMA_signal_8213 ;
    wire new_AGEMA_signal_8214 ;
    wire new_AGEMA_signal_8215 ;
    wire new_AGEMA_signal_8216 ;
    wire new_AGEMA_signal_8217 ;
    wire new_AGEMA_signal_8218 ;
    wire new_AGEMA_signal_8219 ;
    wire new_AGEMA_signal_8220 ;
    wire new_AGEMA_signal_8221 ;
    wire new_AGEMA_signal_8222 ;
    wire new_AGEMA_signal_8223 ;
    wire new_AGEMA_signal_8224 ;
    wire new_AGEMA_signal_8225 ;
    wire new_AGEMA_signal_8226 ;
    wire new_AGEMA_signal_8227 ;
    wire new_AGEMA_signal_8228 ;
    wire new_AGEMA_signal_8229 ;
    wire new_AGEMA_signal_8230 ;
    wire new_AGEMA_signal_8231 ;
    wire new_AGEMA_signal_8232 ;
    wire new_AGEMA_signal_8233 ;
    wire new_AGEMA_signal_8234 ;
    wire new_AGEMA_signal_8235 ;
    wire new_AGEMA_signal_8236 ;
    wire new_AGEMA_signal_8237 ;
    wire new_AGEMA_signal_8238 ;
    wire new_AGEMA_signal_8239 ;
    wire new_AGEMA_signal_8240 ;
    wire new_AGEMA_signal_8241 ;
    wire new_AGEMA_signal_8242 ;
    wire new_AGEMA_signal_8243 ;
    wire new_AGEMA_signal_8244 ;
    wire new_AGEMA_signal_8245 ;
    wire new_AGEMA_signal_8246 ;
    wire new_AGEMA_signal_8247 ;
    wire new_AGEMA_signal_8248 ;
    wire new_AGEMA_signal_8249 ;
    wire new_AGEMA_signal_8250 ;
    wire new_AGEMA_signal_8251 ;
    wire new_AGEMA_signal_8252 ;
    wire new_AGEMA_signal_8253 ;
    wire new_AGEMA_signal_8254 ;
    wire new_AGEMA_signal_8255 ;
    wire new_AGEMA_signal_8256 ;
    wire new_AGEMA_signal_8257 ;
    wire new_AGEMA_signal_8258 ;
    wire new_AGEMA_signal_8259 ;
    wire new_AGEMA_signal_8260 ;
    wire new_AGEMA_signal_8261 ;
    wire new_AGEMA_signal_8262 ;
    wire new_AGEMA_signal_8263 ;
    wire new_AGEMA_signal_8264 ;
    wire new_AGEMA_signal_8265 ;
    wire new_AGEMA_signal_8266 ;
    wire new_AGEMA_signal_8267 ;
    wire new_AGEMA_signal_8268 ;
    wire new_AGEMA_signal_8269 ;
    wire new_AGEMA_signal_8270 ;
    wire new_AGEMA_signal_8271 ;
    wire new_AGEMA_signal_8272 ;
    wire new_AGEMA_signal_8273 ;
    wire new_AGEMA_signal_8274 ;
    wire new_AGEMA_signal_8275 ;
    wire new_AGEMA_signal_8276 ;
    wire new_AGEMA_signal_8277 ;
    wire new_AGEMA_signal_8278 ;
    wire new_AGEMA_signal_8279 ;
    wire new_AGEMA_signal_8280 ;
    wire new_AGEMA_signal_8281 ;
    wire new_AGEMA_signal_8282 ;
    wire new_AGEMA_signal_8283 ;
    wire new_AGEMA_signal_8284 ;
    wire new_AGEMA_signal_8285 ;
    wire new_AGEMA_signal_8286 ;
    wire new_AGEMA_signal_8287 ;
    wire new_AGEMA_signal_8288 ;
    wire new_AGEMA_signal_8289 ;
    wire new_AGEMA_signal_8290 ;
    wire new_AGEMA_signal_8291 ;
    wire new_AGEMA_signal_8292 ;
    wire new_AGEMA_signal_8293 ;
    wire new_AGEMA_signal_8294 ;
    wire new_AGEMA_signal_8295 ;
    wire new_AGEMA_signal_8296 ;
    wire new_AGEMA_signal_8297 ;
    wire new_AGEMA_signal_8298 ;
    wire new_AGEMA_signal_8299 ;
    wire new_AGEMA_signal_8300 ;
    wire new_AGEMA_signal_8301 ;
    wire new_AGEMA_signal_8302 ;
    wire new_AGEMA_signal_8303 ;
    wire new_AGEMA_signal_8304 ;
    wire new_AGEMA_signal_8305 ;
    wire new_AGEMA_signal_8306 ;
    wire new_AGEMA_signal_8307 ;
    wire new_AGEMA_signal_8308 ;
    wire new_AGEMA_signal_8309 ;
    wire new_AGEMA_signal_8310 ;
    wire new_AGEMA_signal_8311 ;
    wire new_AGEMA_signal_8312 ;
    wire new_AGEMA_signal_8313 ;
    wire new_AGEMA_signal_8314 ;
    wire new_AGEMA_signal_8315 ;
    wire new_AGEMA_signal_8316 ;
    wire new_AGEMA_signal_8317 ;
    wire new_AGEMA_signal_8318 ;
    wire new_AGEMA_signal_8319 ;
    wire new_AGEMA_signal_8320 ;
    wire new_AGEMA_signal_8321 ;
    wire new_AGEMA_signal_8322 ;
    wire new_AGEMA_signal_8323 ;
    wire new_AGEMA_signal_8324 ;
    wire new_AGEMA_signal_8325 ;
    wire new_AGEMA_signal_8326 ;
    wire new_AGEMA_signal_8327 ;
    wire new_AGEMA_signal_8328 ;
    wire new_AGEMA_signal_8329 ;
    wire new_AGEMA_signal_8330 ;
    wire new_AGEMA_signal_8331 ;
    wire new_AGEMA_signal_8332 ;
    wire new_AGEMA_signal_8333 ;
    wire new_AGEMA_signal_8334 ;
    wire new_AGEMA_signal_8335 ;
    wire new_AGEMA_signal_8336 ;
    wire new_AGEMA_signal_8337 ;
    wire new_AGEMA_signal_8338 ;
    wire new_AGEMA_signal_8339 ;
    wire new_AGEMA_signal_8340 ;
    wire new_AGEMA_signal_8341 ;
    wire new_AGEMA_signal_8342 ;
    wire new_AGEMA_signal_8343 ;
    wire new_AGEMA_signal_8344 ;
    wire new_AGEMA_signal_8345 ;
    wire new_AGEMA_signal_8346 ;
    wire new_AGEMA_signal_8347 ;
    wire new_AGEMA_signal_8348 ;
    wire new_AGEMA_signal_8349 ;
    wire new_AGEMA_signal_8350 ;
    wire new_AGEMA_signal_8351 ;
    wire new_AGEMA_signal_8352 ;
    wire new_AGEMA_signal_8353 ;
    wire new_AGEMA_signal_8354 ;
    wire new_AGEMA_signal_8355 ;
    wire new_AGEMA_signal_8356 ;
    wire new_AGEMA_signal_8357 ;
    wire new_AGEMA_signal_8358 ;
    wire new_AGEMA_signal_8359 ;
    wire new_AGEMA_signal_8360 ;
    wire new_AGEMA_signal_8361 ;
    wire new_AGEMA_signal_8362 ;
    wire new_AGEMA_signal_8363 ;
    wire new_AGEMA_signal_8364 ;
    wire new_AGEMA_signal_8365 ;
    wire new_AGEMA_signal_8366 ;
    wire new_AGEMA_signal_8367 ;
    wire new_AGEMA_signal_8368 ;
    wire new_AGEMA_signal_8369 ;
    wire new_AGEMA_signal_8370 ;
    wire new_AGEMA_signal_8371 ;
    wire new_AGEMA_signal_8372 ;
    wire new_AGEMA_signal_8373 ;
    wire new_AGEMA_signal_8374 ;
    wire new_AGEMA_signal_8375 ;
    wire new_AGEMA_signal_8376 ;
    wire new_AGEMA_signal_8377 ;
    wire new_AGEMA_signal_8378 ;
    wire new_AGEMA_signal_8379 ;
    wire new_AGEMA_signal_8380 ;
    wire new_AGEMA_signal_8381 ;
    wire new_AGEMA_signal_8382 ;
    wire new_AGEMA_signal_8383 ;
    wire new_AGEMA_signal_8384 ;
    wire new_AGEMA_signal_8385 ;
    wire new_AGEMA_signal_8386 ;
    wire new_AGEMA_signal_8387 ;
    wire new_AGEMA_signal_8388 ;
    wire new_AGEMA_signal_8389 ;
    wire new_AGEMA_signal_8390 ;
    wire new_AGEMA_signal_8391 ;
    wire new_AGEMA_signal_8392 ;
    wire new_AGEMA_signal_8393 ;
    wire new_AGEMA_signal_8394 ;
    wire new_AGEMA_signal_8395 ;
    wire new_AGEMA_signal_8396 ;
    wire new_AGEMA_signal_8397 ;
    wire new_AGEMA_signal_8398 ;
    wire new_AGEMA_signal_8399 ;
    wire new_AGEMA_signal_8400 ;
    wire new_AGEMA_signal_8401 ;
    wire new_AGEMA_signal_8402 ;
    wire new_AGEMA_signal_8403 ;
    wire new_AGEMA_signal_8404 ;
    wire new_AGEMA_signal_8405 ;
    wire new_AGEMA_signal_8406 ;
    wire new_AGEMA_signal_8407 ;
    wire new_AGEMA_signal_8408 ;
    wire new_AGEMA_signal_8409 ;
    wire new_AGEMA_signal_8410 ;
    wire new_AGEMA_signal_8411 ;
    wire new_AGEMA_signal_8412 ;
    wire new_AGEMA_signal_8413 ;
    wire new_AGEMA_signal_8414 ;
    wire new_AGEMA_signal_8415 ;
    wire new_AGEMA_signal_8416 ;
    wire new_AGEMA_signal_8417 ;
    wire new_AGEMA_signal_8418 ;
    wire new_AGEMA_signal_8419 ;
    wire new_AGEMA_signal_8420 ;
    wire new_AGEMA_signal_8421 ;
    wire new_AGEMA_signal_8422 ;
    wire new_AGEMA_signal_8423 ;
    wire new_AGEMA_signal_8424 ;
    wire new_AGEMA_signal_8425 ;
    wire new_AGEMA_signal_8426 ;
    wire new_AGEMA_signal_8427 ;
    wire new_AGEMA_signal_8428 ;
    wire new_AGEMA_signal_8429 ;
    wire new_AGEMA_signal_8430 ;
    wire new_AGEMA_signal_8431 ;
    wire new_AGEMA_signal_8432 ;
    wire new_AGEMA_signal_8433 ;
    wire new_AGEMA_signal_8434 ;
    wire new_AGEMA_signal_8435 ;
    wire new_AGEMA_signal_8436 ;
    wire new_AGEMA_signal_8437 ;
    wire new_AGEMA_signal_8438 ;
    wire new_AGEMA_signal_8439 ;
    wire new_AGEMA_signal_8440 ;
    wire new_AGEMA_signal_8441 ;
    wire new_AGEMA_signal_8442 ;
    wire new_AGEMA_signal_8443 ;
    wire new_AGEMA_signal_8444 ;
    wire new_AGEMA_signal_8445 ;
    wire new_AGEMA_signal_8446 ;
    wire new_AGEMA_signal_8447 ;
    wire new_AGEMA_signal_8448 ;
    wire new_AGEMA_signal_8449 ;
    wire new_AGEMA_signal_8450 ;
    wire new_AGEMA_signal_8451 ;
    wire new_AGEMA_signal_8452 ;
    wire new_AGEMA_signal_8453 ;
    wire new_AGEMA_signal_8454 ;
    wire new_AGEMA_signal_8455 ;
    wire new_AGEMA_signal_8456 ;
    wire new_AGEMA_signal_8457 ;
    wire new_AGEMA_signal_8458 ;
    wire new_AGEMA_signal_8459 ;
    wire new_AGEMA_signal_8460 ;
    wire new_AGEMA_signal_8461 ;
    wire new_AGEMA_signal_8462 ;
    wire new_AGEMA_signal_8463 ;
    wire new_AGEMA_signal_8464 ;
    wire new_AGEMA_signal_8465 ;
    wire new_AGEMA_signal_8466 ;
    wire new_AGEMA_signal_8467 ;
    wire new_AGEMA_signal_8468 ;
    wire new_AGEMA_signal_8469 ;
    wire new_AGEMA_signal_8470 ;
    wire new_AGEMA_signal_8471 ;
    wire new_AGEMA_signal_8472 ;
    wire new_AGEMA_signal_8473 ;
    wire new_AGEMA_signal_8474 ;
    wire new_AGEMA_signal_8475 ;
    wire new_AGEMA_signal_8476 ;
    wire new_AGEMA_signal_8477 ;
    wire new_AGEMA_signal_8478 ;
    wire new_AGEMA_signal_8479 ;
    wire new_AGEMA_signal_8480 ;
    wire new_AGEMA_signal_8481 ;
    wire new_AGEMA_signal_8482 ;
    wire new_AGEMA_signal_8483 ;
    wire new_AGEMA_signal_8484 ;
    wire new_AGEMA_signal_8485 ;
    wire new_AGEMA_signal_8486 ;
    wire new_AGEMA_signal_8487 ;
    wire new_AGEMA_signal_8488 ;
    wire new_AGEMA_signal_8489 ;
    wire new_AGEMA_signal_8490 ;
    wire new_AGEMA_signal_8491 ;
    wire new_AGEMA_signal_8492 ;
    wire new_AGEMA_signal_8493 ;
    wire new_AGEMA_signal_8494 ;
    wire new_AGEMA_signal_8495 ;
    wire new_AGEMA_signal_8496 ;
    wire new_AGEMA_signal_8497 ;
    wire new_AGEMA_signal_8498 ;
    wire new_AGEMA_signal_8499 ;
    wire new_AGEMA_signal_8500 ;
    wire new_AGEMA_signal_8501 ;
    wire new_AGEMA_signal_8502 ;
    wire new_AGEMA_signal_8503 ;
    wire new_AGEMA_signal_8504 ;
    wire new_AGEMA_signal_8505 ;
    wire new_AGEMA_signal_8506 ;
    wire new_AGEMA_signal_8507 ;
    wire new_AGEMA_signal_8508 ;
    wire new_AGEMA_signal_8509 ;
    wire new_AGEMA_signal_8510 ;
    wire new_AGEMA_signal_8511 ;
    wire new_AGEMA_signal_8512 ;
    wire new_AGEMA_signal_8513 ;
    wire new_AGEMA_signal_8514 ;
    wire new_AGEMA_signal_8515 ;
    wire new_AGEMA_signal_8516 ;
    wire new_AGEMA_signal_8517 ;
    wire new_AGEMA_signal_8518 ;
    wire new_AGEMA_signal_8519 ;
    wire new_AGEMA_signal_8520 ;
    wire new_AGEMA_signal_8521 ;
    wire new_AGEMA_signal_8522 ;
    wire new_AGEMA_signal_8523 ;
    wire new_AGEMA_signal_8524 ;
    wire new_AGEMA_signal_8525 ;
    wire new_AGEMA_signal_8526 ;
    wire new_AGEMA_signal_8527 ;
    wire new_AGEMA_signal_8528 ;
    wire new_AGEMA_signal_8529 ;
    wire new_AGEMA_signal_8530 ;
    wire new_AGEMA_signal_8531 ;
    wire new_AGEMA_signal_8532 ;
    wire new_AGEMA_signal_8533 ;
    wire new_AGEMA_signal_8534 ;
    wire new_AGEMA_signal_8535 ;
    wire new_AGEMA_signal_8536 ;
    wire new_AGEMA_signal_8537 ;
    wire new_AGEMA_signal_8538 ;
    wire new_AGEMA_signal_8539 ;
    wire new_AGEMA_signal_8540 ;
    wire new_AGEMA_signal_8541 ;
    wire new_AGEMA_signal_8542 ;
    wire new_AGEMA_signal_8543 ;
    wire new_AGEMA_signal_8544 ;
    wire new_AGEMA_signal_8545 ;
    wire new_AGEMA_signal_8546 ;
    wire new_AGEMA_signal_8547 ;
    wire new_AGEMA_signal_8548 ;
    wire new_AGEMA_signal_8549 ;
    wire new_AGEMA_signal_8550 ;
    wire new_AGEMA_signal_8551 ;
    wire new_AGEMA_signal_8552 ;
    wire new_AGEMA_signal_8553 ;
    wire new_AGEMA_signal_8554 ;
    wire new_AGEMA_signal_8555 ;
    wire new_AGEMA_signal_8556 ;
    wire new_AGEMA_signal_8557 ;
    wire new_AGEMA_signal_8558 ;
    wire new_AGEMA_signal_8559 ;
    wire new_AGEMA_signal_8560 ;
    wire new_AGEMA_signal_8561 ;
    wire new_AGEMA_signal_8562 ;
    wire new_AGEMA_signal_8563 ;
    wire new_AGEMA_signal_8564 ;
    wire new_AGEMA_signal_8565 ;
    wire new_AGEMA_signal_8566 ;
    wire new_AGEMA_signal_8567 ;
    wire new_AGEMA_signal_8568 ;
    wire new_AGEMA_signal_8569 ;
    wire new_AGEMA_signal_8570 ;
    wire new_AGEMA_signal_8571 ;
    wire new_AGEMA_signal_8572 ;
    wire new_AGEMA_signal_8573 ;
    wire new_AGEMA_signal_8574 ;
    wire new_AGEMA_signal_8575 ;
    wire new_AGEMA_signal_8576 ;
    wire new_AGEMA_signal_8577 ;
    wire new_AGEMA_signal_8578 ;
    wire new_AGEMA_signal_8579 ;
    wire new_AGEMA_signal_8580 ;
    wire new_AGEMA_signal_8581 ;
    wire new_AGEMA_signal_8582 ;
    wire new_AGEMA_signal_8583 ;
    wire new_AGEMA_signal_8584 ;
    wire new_AGEMA_signal_8585 ;
    wire new_AGEMA_signal_8586 ;
    wire new_AGEMA_signal_8587 ;
    wire new_AGEMA_signal_8588 ;
    wire new_AGEMA_signal_8589 ;
    wire new_AGEMA_signal_8590 ;
    wire new_AGEMA_signal_8591 ;
    wire new_AGEMA_signal_8592 ;
    wire new_AGEMA_signal_8593 ;
    wire new_AGEMA_signal_8594 ;
    wire new_AGEMA_signal_8595 ;
    wire new_AGEMA_signal_8596 ;
    wire new_AGEMA_signal_8597 ;
    wire new_AGEMA_signal_8598 ;
    wire new_AGEMA_signal_8599 ;
    wire new_AGEMA_signal_8600 ;
    wire new_AGEMA_signal_8601 ;
    wire new_AGEMA_signal_8602 ;
    wire new_AGEMA_signal_8603 ;
    wire new_AGEMA_signal_8604 ;
    wire new_AGEMA_signal_8605 ;
    wire new_AGEMA_signal_8606 ;
    wire new_AGEMA_signal_8607 ;
    wire new_AGEMA_signal_8608 ;
    wire new_AGEMA_signal_8609 ;
    wire new_AGEMA_signal_8610 ;
    wire new_AGEMA_signal_8611 ;
    wire new_AGEMA_signal_8612 ;
    wire new_AGEMA_signal_8613 ;
    wire new_AGEMA_signal_8614 ;
    wire new_AGEMA_signal_8615 ;
    wire new_AGEMA_signal_8616 ;
    wire new_AGEMA_signal_8617 ;
    wire new_AGEMA_signal_8618 ;
    wire new_AGEMA_signal_8619 ;
    wire new_AGEMA_signal_8620 ;
    wire new_AGEMA_signal_8621 ;
    wire new_AGEMA_signal_8622 ;
    wire new_AGEMA_signal_8623 ;
    wire new_AGEMA_signal_8624 ;
    wire new_AGEMA_signal_8625 ;
    wire new_AGEMA_signal_8626 ;
    wire new_AGEMA_signal_8627 ;
    wire new_AGEMA_signal_8628 ;
    wire new_AGEMA_signal_8629 ;
    wire new_AGEMA_signal_8630 ;
    wire new_AGEMA_signal_8631 ;
    wire new_AGEMA_signal_8632 ;
    wire new_AGEMA_signal_8633 ;
    wire new_AGEMA_signal_8634 ;
    wire new_AGEMA_signal_8635 ;
    wire new_AGEMA_signal_8636 ;
    wire new_AGEMA_signal_8637 ;
    wire new_AGEMA_signal_8638 ;
    wire new_AGEMA_signal_8639 ;
    wire new_AGEMA_signal_8640 ;
    wire new_AGEMA_signal_8641 ;
    wire new_AGEMA_signal_8642 ;
    wire new_AGEMA_signal_8643 ;
    wire new_AGEMA_signal_8644 ;
    wire new_AGEMA_signal_8645 ;
    wire new_AGEMA_signal_8646 ;
    wire new_AGEMA_signal_8647 ;
    wire new_AGEMA_signal_8648 ;
    wire new_AGEMA_signal_8649 ;
    wire new_AGEMA_signal_8650 ;
    wire new_AGEMA_signal_8651 ;
    wire new_AGEMA_signal_8652 ;
    wire new_AGEMA_signal_8653 ;
    wire new_AGEMA_signal_8654 ;
    wire new_AGEMA_signal_8655 ;
    wire new_AGEMA_signal_8656 ;
    wire new_AGEMA_signal_8657 ;
    wire new_AGEMA_signal_8658 ;
    wire new_AGEMA_signal_8659 ;
    wire new_AGEMA_signal_8660 ;
    wire new_AGEMA_signal_8661 ;
    wire new_AGEMA_signal_8662 ;
    wire new_AGEMA_signal_8663 ;
    wire new_AGEMA_signal_8664 ;
    wire new_AGEMA_signal_8665 ;
    wire new_AGEMA_signal_8666 ;
    wire new_AGEMA_signal_8667 ;
    wire new_AGEMA_signal_8668 ;
    wire new_AGEMA_signal_8669 ;
    wire new_AGEMA_signal_8670 ;
    wire new_AGEMA_signal_8671 ;
    wire new_AGEMA_signal_8672 ;
    wire new_AGEMA_signal_8673 ;
    wire new_AGEMA_signal_8674 ;
    wire new_AGEMA_signal_8675 ;
    wire new_AGEMA_signal_8676 ;
    wire new_AGEMA_signal_8677 ;
    wire new_AGEMA_signal_8678 ;
    wire new_AGEMA_signal_8679 ;
    wire new_AGEMA_signal_8680 ;
    wire new_AGEMA_signal_8681 ;
    wire new_AGEMA_signal_8682 ;
    wire new_AGEMA_signal_8683 ;
    wire new_AGEMA_signal_8684 ;
    wire new_AGEMA_signal_8685 ;
    wire new_AGEMA_signal_8686 ;
    wire new_AGEMA_signal_8687 ;
    wire new_AGEMA_signal_8688 ;
    wire new_AGEMA_signal_8689 ;
    wire new_AGEMA_signal_8690 ;
    wire new_AGEMA_signal_8691 ;
    wire new_AGEMA_signal_8692 ;
    wire new_AGEMA_signal_8693 ;
    wire new_AGEMA_signal_8694 ;
    wire new_AGEMA_signal_8695 ;
    wire new_AGEMA_signal_8696 ;
    wire new_AGEMA_signal_8697 ;
    wire new_AGEMA_signal_8698 ;
    wire new_AGEMA_signal_8699 ;
    wire new_AGEMA_signal_8700 ;
    wire new_AGEMA_signal_8701 ;
    wire new_AGEMA_signal_8702 ;
    wire new_AGEMA_signal_8703 ;
    wire new_AGEMA_signal_8704 ;
    wire new_AGEMA_signal_8705 ;
    wire new_AGEMA_signal_8706 ;
    wire new_AGEMA_signal_8707 ;
    wire new_AGEMA_signal_8708 ;
    wire new_AGEMA_signal_8709 ;
    wire new_AGEMA_signal_8710 ;
    wire new_AGEMA_signal_8711 ;
    wire new_AGEMA_signal_8712 ;
    wire new_AGEMA_signal_8713 ;
    wire new_AGEMA_signal_8714 ;
    wire new_AGEMA_signal_8715 ;
    wire new_AGEMA_signal_8716 ;
    wire new_AGEMA_signal_8717 ;
    wire new_AGEMA_signal_8718 ;
    wire new_AGEMA_signal_8719 ;
    wire new_AGEMA_signal_8720 ;
    wire new_AGEMA_signal_8721 ;
    wire new_AGEMA_signal_8722 ;
    wire new_AGEMA_signal_8723 ;
    wire new_AGEMA_signal_8724 ;
    wire new_AGEMA_signal_8725 ;
    wire new_AGEMA_signal_8726 ;
    wire new_AGEMA_signal_8727 ;
    wire new_AGEMA_signal_8728 ;
    wire new_AGEMA_signal_8729 ;
    wire new_AGEMA_signal_8730 ;
    wire new_AGEMA_signal_8731 ;
    wire new_AGEMA_signal_8732 ;
    wire new_AGEMA_signal_8733 ;
    wire new_AGEMA_signal_8734 ;
    wire new_AGEMA_signal_8735 ;
    wire new_AGEMA_signal_8736 ;
    wire new_AGEMA_signal_8737 ;
    wire new_AGEMA_signal_8738 ;
    wire new_AGEMA_signal_8739 ;
    wire new_AGEMA_signal_8740 ;
    wire new_AGEMA_signal_8741 ;
    wire new_AGEMA_signal_8742 ;
    wire new_AGEMA_signal_8743 ;
    wire new_AGEMA_signal_8744 ;
    wire new_AGEMA_signal_8745 ;
    wire new_AGEMA_signal_8746 ;
    wire new_AGEMA_signal_8747 ;
    wire new_AGEMA_signal_8748 ;
    wire new_AGEMA_signal_8749 ;
    wire new_AGEMA_signal_8750 ;
    wire new_AGEMA_signal_8751 ;
    wire new_AGEMA_signal_8752 ;
    wire new_AGEMA_signal_8753 ;
    wire new_AGEMA_signal_8754 ;
    wire new_AGEMA_signal_8755 ;
    wire new_AGEMA_signal_8756 ;
    wire new_AGEMA_signal_8757 ;
    wire new_AGEMA_signal_8758 ;
    wire new_AGEMA_signal_8759 ;
    wire new_AGEMA_signal_8760 ;
    wire new_AGEMA_signal_8761 ;
    wire new_AGEMA_signal_8762 ;
    wire new_AGEMA_signal_8763 ;
    wire new_AGEMA_signal_8764 ;
    wire new_AGEMA_signal_8765 ;
    wire new_AGEMA_signal_8766 ;
    wire new_AGEMA_signal_8767 ;
    wire new_AGEMA_signal_8768 ;
    wire new_AGEMA_signal_8769 ;
    wire new_AGEMA_signal_8770 ;
    wire new_AGEMA_signal_8771 ;
    wire new_AGEMA_signal_8772 ;
    wire new_AGEMA_signal_8773 ;
    wire new_AGEMA_signal_8774 ;
    wire new_AGEMA_signal_8775 ;
    wire new_AGEMA_signal_8776 ;
    wire new_AGEMA_signal_8777 ;
    wire new_AGEMA_signal_8778 ;
    wire new_AGEMA_signal_8779 ;
    wire new_AGEMA_signal_8780 ;
    wire new_AGEMA_signal_8781 ;
    wire new_AGEMA_signal_8782 ;
    wire new_AGEMA_signal_8783 ;
    wire new_AGEMA_signal_8784 ;
    wire new_AGEMA_signal_8785 ;
    wire new_AGEMA_signal_8786 ;
    wire new_AGEMA_signal_8787 ;
    wire new_AGEMA_signal_8788 ;
    wire new_AGEMA_signal_8789 ;
    wire new_AGEMA_signal_8790 ;
    wire new_AGEMA_signal_8791 ;
    wire new_AGEMA_signal_8792 ;
    wire new_AGEMA_signal_8793 ;
    wire new_AGEMA_signal_8794 ;
    wire new_AGEMA_signal_8795 ;
    wire new_AGEMA_signal_8796 ;
    wire new_AGEMA_signal_8797 ;
    wire new_AGEMA_signal_8798 ;
    wire new_AGEMA_signal_8799 ;
    wire new_AGEMA_signal_8800 ;
    wire new_AGEMA_signal_8801 ;
    wire new_AGEMA_signal_8802 ;
    wire new_AGEMA_signal_8803 ;
    wire new_AGEMA_signal_8804 ;
    wire new_AGEMA_signal_8805 ;
    wire new_AGEMA_signal_8806 ;
    wire new_AGEMA_signal_8807 ;
    wire new_AGEMA_signal_8808 ;
    wire new_AGEMA_signal_8809 ;
    wire new_AGEMA_signal_8810 ;
    wire new_AGEMA_signal_8811 ;
    wire new_AGEMA_signal_8812 ;
    wire new_AGEMA_signal_8813 ;
    wire new_AGEMA_signal_8814 ;
    wire new_AGEMA_signal_8815 ;
    wire new_AGEMA_signal_8816 ;
    wire new_AGEMA_signal_8817 ;
    wire new_AGEMA_signal_8818 ;
    wire new_AGEMA_signal_8819 ;
    wire new_AGEMA_signal_8820 ;
    wire new_AGEMA_signal_8821 ;
    wire new_AGEMA_signal_8822 ;
    wire new_AGEMA_signal_8823 ;
    wire new_AGEMA_signal_8824 ;
    wire new_AGEMA_signal_8825 ;
    wire new_AGEMA_signal_8826 ;
    wire new_AGEMA_signal_8827 ;
    wire new_AGEMA_signal_8828 ;
    wire new_AGEMA_signal_8829 ;
    wire new_AGEMA_signal_8830 ;
    wire new_AGEMA_signal_8831 ;
    wire new_AGEMA_signal_8832 ;
    wire new_AGEMA_signal_8833 ;
    wire new_AGEMA_signal_8834 ;
    wire new_AGEMA_signal_8835 ;
    wire new_AGEMA_signal_8836 ;
    wire new_AGEMA_signal_8837 ;
    wire new_AGEMA_signal_8838 ;
    wire new_AGEMA_signal_8839 ;
    wire new_AGEMA_signal_8840 ;
    wire new_AGEMA_signal_8841 ;
    wire new_AGEMA_signal_8842 ;
    wire new_AGEMA_signal_8843 ;
    wire new_AGEMA_signal_8844 ;
    wire new_AGEMA_signal_8845 ;
    wire new_AGEMA_signal_8846 ;
    wire new_AGEMA_signal_8847 ;
    wire new_AGEMA_signal_8848 ;
    wire new_AGEMA_signal_8849 ;
    wire new_AGEMA_signal_8850 ;
    wire new_AGEMA_signal_8851 ;
    wire new_AGEMA_signal_8852 ;
    wire new_AGEMA_signal_8853 ;
    wire new_AGEMA_signal_8854 ;
    wire new_AGEMA_signal_8855 ;
    wire new_AGEMA_signal_8856 ;
    wire new_AGEMA_signal_8857 ;
    wire new_AGEMA_signal_8858 ;
    wire new_AGEMA_signal_8859 ;
    wire new_AGEMA_signal_8860 ;
    wire new_AGEMA_signal_8861 ;
    wire new_AGEMA_signal_8862 ;
    wire new_AGEMA_signal_8863 ;
    wire new_AGEMA_signal_8864 ;
    wire new_AGEMA_signal_8865 ;
    wire new_AGEMA_signal_8866 ;
    wire new_AGEMA_signal_8867 ;
    wire new_AGEMA_signal_8868 ;
    wire new_AGEMA_signal_8869 ;
    wire new_AGEMA_signal_8870 ;
    wire new_AGEMA_signal_8871 ;
    wire new_AGEMA_signal_8872 ;
    wire new_AGEMA_signal_8873 ;
    wire new_AGEMA_signal_8874 ;
    wire new_AGEMA_signal_8875 ;
    wire new_AGEMA_signal_8876 ;
    wire new_AGEMA_signal_8877 ;
    wire new_AGEMA_signal_8878 ;
    wire new_AGEMA_signal_8879 ;
    wire new_AGEMA_signal_8880 ;
    wire new_AGEMA_signal_8881 ;
    wire new_AGEMA_signal_8882 ;
    wire new_AGEMA_signal_8883 ;
    wire new_AGEMA_signal_8884 ;
    wire new_AGEMA_signal_8885 ;
    wire new_AGEMA_signal_8886 ;
    wire new_AGEMA_signal_8887 ;
    wire new_AGEMA_signal_8888 ;
    wire new_AGEMA_signal_8889 ;
    wire new_AGEMA_signal_8890 ;
    wire new_AGEMA_signal_8891 ;
    wire new_AGEMA_signal_8892 ;
    wire new_AGEMA_signal_8893 ;
    wire new_AGEMA_signal_8894 ;
    wire new_AGEMA_signal_8895 ;
    wire new_AGEMA_signal_8896 ;
    wire new_AGEMA_signal_8897 ;
    wire new_AGEMA_signal_8898 ;
    wire new_AGEMA_signal_8899 ;
    wire new_AGEMA_signal_8900 ;
    wire new_AGEMA_signal_8901 ;
    wire new_AGEMA_signal_8902 ;
    wire new_AGEMA_signal_8903 ;
    wire new_AGEMA_signal_8904 ;
    wire new_AGEMA_signal_8905 ;
    wire new_AGEMA_signal_8906 ;
    wire new_AGEMA_signal_8907 ;
    wire new_AGEMA_signal_8908 ;
    wire new_AGEMA_signal_8909 ;
    wire new_AGEMA_signal_8910 ;
    wire new_AGEMA_signal_8911 ;
    wire new_AGEMA_signal_8912 ;
    wire new_AGEMA_signal_8913 ;
    wire new_AGEMA_signal_8914 ;
    wire new_AGEMA_signal_8915 ;
    wire new_AGEMA_signal_8916 ;
    wire new_AGEMA_signal_8917 ;
    wire new_AGEMA_signal_8918 ;
    wire new_AGEMA_signal_8919 ;
    wire new_AGEMA_signal_8920 ;
    wire new_AGEMA_signal_8921 ;
    wire new_AGEMA_signal_8922 ;
    wire new_AGEMA_signal_8923 ;
    wire new_AGEMA_signal_8924 ;
    wire new_AGEMA_signal_8925 ;
    wire new_AGEMA_signal_8926 ;
    wire new_AGEMA_signal_8927 ;
    wire new_AGEMA_signal_8928 ;
    wire new_AGEMA_signal_8929 ;
    wire new_AGEMA_signal_8930 ;
    wire new_AGEMA_signal_8931 ;
    wire new_AGEMA_signal_8932 ;
    wire new_AGEMA_signal_8933 ;
    wire new_AGEMA_signal_8934 ;
    wire new_AGEMA_signal_8935 ;
    wire new_AGEMA_signal_8936 ;
    wire new_AGEMA_signal_8937 ;
    wire new_AGEMA_signal_8938 ;
    wire new_AGEMA_signal_8939 ;
    wire new_AGEMA_signal_8940 ;
    wire new_AGEMA_signal_8941 ;
    wire new_AGEMA_signal_8942 ;
    wire new_AGEMA_signal_8943 ;
    wire new_AGEMA_signal_8944 ;
    wire new_AGEMA_signal_8945 ;
    wire new_AGEMA_signal_8946 ;
    wire new_AGEMA_signal_8947 ;
    wire new_AGEMA_signal_8948 ;
    wire new_AGEMA_signal_8949 ;
    wire new_AGEMA_signal_8950 ;
    wire new_AGEMA_signal_8951 ;
    wire new_AGEMA_signal_8952 ;
    wire new_AGEMA_signal_8953 ;
    wire new_AGEMA_signal_8954 ;
    wire new_AGEMA_signal_8955 ;
    wire new_AGEMA_signal_8956 ;
    wire new_AGEMA_signal_8957 ;
    wire new_AGEMA_signal_8958 ;
    wire new_AGEMA_signal_8959 ;
    wire new_AGEMA_signal_8960 ;
    wire new_AGEMA_signal_8961 ;
    wire new_AGEMA_signal_8962 ;
    wire new_AGEMA_signal_8963 ;
    wire new_AGEMA_signal_8964 ;
    wire new_AGEMA_signal_8965 ;
    wire new_AGEMA_signal_8966 ;
    wire new_AGEMA_signal_8967 ;
    wire new_AGEMA_signal_8968 ;
    wire new_AGEMA_signal_8969 ;
    wire new_AGEMA_signal_8970 ;
    wire new_AGEMA_signal_8971 ;
    wire new_AGEMA_signal_8972 ;
    wire new_AGEMA_signal_8973 ;
    wire new_AGEMA_signal_8974 ;
    wire new_AGEMA_signal_8975 ;
    wire new_AGEMA_signal_8976 ;
    wire new_AGEMA_signal_8977 ;
    wire new_AGEMA_signal_8978 ;
    wire new_AGEMA_signal_8979 ;
    wire new_AGEMA_signal_8980 ;
    wire new_AGEMA_signal_8981 ;
    wire new_AGEMA_signal_8982 ;
    wire new_AGEMA_signal_8983 ;
    wire new_AGEMA_signal_8984 ;
    wire new_AGEMA_signal_8985 ;
    wire new_AGEMA_signal_8986 ;
    wire new_AGEMA_signal_8987 ;
    wire new_AGEMA_signal_8988 ;
    wire new_AGEMA_signal_8989 ;
    wire new_AGEMA_signal_8990 ;
    wire new_AGEMA_signal_8991 ;
    wire new_AGEMA_signal_8992 ;
    wire new_AGEMA_signal_8993 ;
    wire new_AGEMA_signal_8994 ;
    wire new_AGEMA_signal_8995 ;
    wire new_AGEMA_signal_8996 ;
    wire new_AGEMA_signal_8997 ;
    wire new_AGEMA_signal_8998 ;
    wire new_AGEMA_signal_8999 ;
    wire new_AGEMA_signal_9000 ;
    wire new_AGEMA_signal_9001 ;
    wire new_AGEMA_signal_9002 ;
    wire new_AGEMA_signal_9003 ;
    wire new_AGEMA_signal_9004 ;
    wire new_AGEMA_signal_9005 ;
    wire new_AGEMA_signal_9006 ;
    wire new_AGEMA_signal_9007 ;
    wire new_AGEMA_signal_9008 ;
    wire new_AGEMA_signal_9009 ;
    wire new_AGEMA_signal_9010 ;
    wire new_AGEMA_signal_9011 ;
    wire new_AGEMA_signal_9012 ;
    wire new_AGEMA_signal_9013 ;
    wire new_AGEMA_signal_9014 ;
    wire new_AGEMA_signal_9015 ;
    wire new_AGEMA_signal_9016 ;
    wire new_AGEMA_signal_9017 ;
    wire new_AGEMA_signal_9018 ;
    wire new_AGEMA_signal_9019 ;
    wire new_AGEMA_signal_9020 ;
    wire new_AGEMA_signal_9021 ;
    wire new_AGEMA_signal_9022 ;
    wire new_AGEMA_signal_9023 ;
    wire new_AGEMA_signal_9024 ;
    wire new_AGEMA_signal_9025 ;
    wire new_AGEMA_signal_9026 ;
    wire new_AGEMA_signal_9027 ;
    wire new_AGEMA_signal_9028 ;
    wire new_AGEMA_signal_9029 ;
    wire new_AGEMA_signal_9030 ;
    wire new_AGEMA_signal_9031 ;
    wire new_AGEMA_signal_9032 ;
    wire new_AGEMA_signal_9033 ;
    wire new_AGEMA_signal_9034 ;
    wire new_AGEMA_signal_9035 ;
    wire new_AGEMA_signal_9036 ;
    wire new_AGEMA_signal_9037 ;
    wire new_AGEMA_signal_9038 ;
    wire new_AGEMA_signal_9039 ;
    wire new_AGEMA_signal_9040 ;
    wire new_AGEMA_signal_9041 ;
    wire new_AGEMA_signal_9042 ;
    wire new_AGEMA_signal_9043 ;
    wire new_AGEMA_signal_9044 ;
    wire new_AGEMA_signal_9045 ;
    wire new_AGEMA_signal_9046 ;
    wire new_AGEMA_signal_9047 ;
    wire new_AGEMA_signal_9048 ;
    wire new_AGEMA_signal_9049 ;
    wire new_AGEMA_signal_9050 ;
    wire new_AGEMA_signal_9051 ;
    wire new_AGEMA_signal_9052 ;
    wire new_AGEMA_signal_9053 ;
    wire new_AGEMA_signal_9054 ;
    wire new_AGEMA_signal_9055 ;
    wire new_AGEMA_signal_9056 ;
    wire new_AGEMA_signal_9057 ;
    wire new_AGEMA_signal_9058 ;
    wire new_AGEMA_signal_9059 ;
    wire new_AGEMA_signal_9060 ;
    wire new_AGEMA_signal_9061 ;
    wire new_AGEMA_signal_9062 ;
    wire new_AGEMA_signal_9063 ;
    wire new_AGEMA_signal_9064 ;
    wire new_AGEMA_signal_9065 ;
    wire new_AGEMA_signal_9066 ;
    wire new_AGEMA_signal_9067 ;
    wire new_AGEMA_signal_9068 ;
    wire new_AGEMA_signal_9069 ;
    wire new_AGEMA_signal_9070 ;
    wire new_AGEMA_signal_9071 ;
    wire new_AGEMA_signal_9072 ;
    wire new_AGEMA_signal_9073 ;
    wire new_AGEMA_signal_9074 ;
    wire new_AGEMA_signal_9075 ;
    wire new_AGEMA_signal_9076 ;
    wire new_AGEMA_signal_9077 ;
    wire new_AGEMA_signal_9078 ;
    wire new_AGEMA_signal_9079 ;
    wire new_AGEMA_signal_9080 ;
    wire new_AGEMA_signal_9081 ;
    wire new_AGEMA_signal_9082 ;
    wire new_AGEMA_signal_9083 ;
    wire new_AGEMA_signal_9084 ;
    wire new_AGEMA_signal_9085 ;
    wire new_AGEMA_signal_9086 ;
    wire new_AGEMA_signal_9087 ;
    wire new_AGEMA_signal_9088 ;
    wire new_AGEMA_signal_9089 ;
    wire new_AGEMA_signal_9090 ;
    wire new_AGEMA_signal_9091 ;
    wire new_AGEMA_signal_9092 ;
    wire new_AGEMA_signal_9093 ;
    wire new_AGEMA_signal_9094 ;
    wire new_AGEMA_signal_9095 ;
    wire new_AGEMA_signal_9096 ;
    wire new_AGEMA_signal_9097 ;
    wire new_AGEMA_signal_9098 ;
    wire new_AGEMA_signal_9099 ;
    wire new_AGEMA_signal_9100 ;
    wire new_AGEMA_signal_9101 ;
    wire new_AGEMA_signal_9102 ;
    wire new_AGEMA_signal_9103 ;
    wire new_AGEMA_signal_9104 ;
    wire new_AGEMA_signal_9105 ;
    wire new_AGEMA_signal_9106 ;
    wire new_AGEMA_signal_9107 ;
    wire new_AGEMA_signal_9108 ;
    wire new_AGEMA_signal_9109 ;
    wire new_AGEMA_signal_9110 ;
    wire new_AGEMA_signal_9111 ;
    wire new_AGEMA_signal_9112 ;
    wire new_AGEMA_signal_9113 ;
    wire new_AGEMA_signal_9114 ;
    wire new_AGEMA_signal_9115 ;
    wire new_AGEMA_signal_9116 ;
    wire new_AGEMA_signal_9117 ;
    wire new_AGEMA_signal_9118 ;
    wire new_AGEMA_signal_9119 ;
    wire new_AGEMA_signal_9120 ;
    wire new_AGEMA_signal_9121 ;
    wire new_AGEMA_signal_9122 ;
    wire new_AGEMA_signal_9123 ;
    wire new_AGEMA_signal_9124 ;
    wire new_AGEMA_signal_9125 ;
    wire new_AGEMA_signal_9126 ;
    wire new_AGEMA_signal_9127 ;
    wire new_AGEMA_signal_9128 ;
    wire new_AGEMA_signal_9129 ;
    wire new_AGEMA_signal_9130 ;
    wire new_AGEMA_signal_9131 ;
    wire new_AGEMA_signal_9132 ;
    wire new_AGEMA_signal_9133 ;
    wire new_AGEMA_signal_9134 ;
    wire new_AGEMA_signal_9135 ;
    wire new_AGEMA_signal_9136 ;
    wire new_AGEMA_signal_9137 ;
    wire new_AGEMA_signal_9138 ;
    wire new_AGEMA_signal_9139 ;
    wire new_AGEMA_signal_9140 ;
    wire new_AGEMA_signal_9141 ;
    wire new_AGEMA_signal_9142 ;
    wire new_AGEMA_signal_9143 ;
    wire new_AGEMA_signal_9144 ;
    wire new_AGEMA_signal_9145 ;
    wire new_AGEMA_signal_9146 ;
    wire new_AGEMA_signal_9147 ;
    wire new_AGEMA_signal_9148 ;
    wire new_AGEMA_signal_9149 ;
    wire new_AGEMA_signal_9150 ;
    wire new_AGEMA_signal_9151 ;
    wire new_AGEMA_signal_9152 ;
    wire new_AGEMA_signal_9153 ;
    wire new_AGEMA_signal_9154 ;
    wire new_AGEMA_signal_9155 ;
    wire new_AGEMA_signal_9156 ;
    wire new_AGEMA_signal_9157 ;
    wire new_AGEMA_signal_9158 ;
    wire new_AGEMA_signal_9159 ;
    wire new_AGEMA_signal_9160 ;
    wire new_AGEMA_signal_9161 ;
    wire new_AGEMA_signal_9162 ;
    wire new_AGEMA_signal_9163 ;
    wire new_AGEMA_signal_9164 ;
    wire new_AGEMA_signal_9165 ;
    wire new_AGEMA_signal_9166 ;
    wire new_AGEMA_signal_9167 ;
    wire new_AGEMA_signal_9168 ;
    wire new_AGEMA_signal_9169 ;
    wire new_AGEMA_signal_9170 ;
    wire new_AGEMA_signal_9171 ;
    wire new_AGEMA_signal_9172 ;
    wire new_AGEMA_signal_9173 ;
    wire new_AGEMA_signal_9174 ;
    wire new_AGEMA_signal_9175 ;
    wire new_AGEMA_signal_9176 ;
    wire new_AGEMA_signal_9177 ;
    wire new_AGEMA_signal_9178 ;
    wire new_AGEMA_signal_9179 ;
    wire new_AGEMA_signal_9180 ;
    wire new_AGEMA_signal_9181 ;
    wire new_AGEMA_signal_9182 ;
    wire new_AGEMA_signal_9183 ;
    wire new_AGEMA_signal_9184 ;
    wire new_AGEMA_signal_9185 ;
    wire new_AGEMA_signal_9186 ;
    wire new_AGEMA_signal_9187 ;
    wire new_AGEMA_signal_9188 ;
    wire new_AGEMA_signal_9189 ;
    wire new_AGEMA_signal_9190 ;
    wire new_AGEMA_signal_9191 ;
    wire new_AGEMA_signal_9192 ;
    wire new_AGEMA_signal_9193 ;
    wire new_AGEMA_signal_9194 ;
    wire new_AGEMA_signal_9195 ;
    wire new_AGEMA_signal_9196 ;
    wire new_AGEMA_signal_9197 ;
    wire new_AGEMA_signal_9198 ;
    wire new_AGEMA_signal_9199 ;
    wire new_AGEMA_signal_9200 ;
    wire new_AGEMA_signal_9201 ;
    wire new_AGEMA_signal_9202 ;
    wire new_AGEMA_signal_9203 ;
    wire new_AGEMA_signal_9204 ;
    wire new_AGEMA_signal_9205 ;
    wire new_AGEMA_signal_9206 ;
    wire new_AGEMA_signal_9207 ;
    wire new_AGEMA_signal_9208 ;
    wire new_AGEMA_signal_9209 ;
    wire new_AGEMA_signal_9210 ;
    wire new_AGEMA_signal_9211 ;
    wire new_AGEMA_signal_9212 ;
    wire new_AGEMA_signal_9213 ;
    wire new_AGEMA_signal_9214 ;
    wire new_AGEMA_signal_9215 ;
    wire new_AGEMA_signal_9216 ;
    wire new_AGEMA_signal_9217 ;
    wire new_AGEMA_signal_9218 ;
    wire new_AGEMA_signal_9219 ;
    wire new_AGEMA_signal_9220 ;
    wire new_AGEMA_signal_9221 ;
    wire new_AGEMA_signal_9222 ;
    wire new_AGEMA_signal_9223 ;
    wire new_AGEMA_signal_9224 ;
    wire new_AGEMA_signal_9225 ;
    wire new_AGEMA_signal_9226 ;
    wire new_AGEMA_signal_9227 ;
    wire new_AGEMA_signal_9228 ;
    wire new_AGEMA_signal_9229 ;
    wire new_AGEMA_signal_9230 ;
    wire new_AGEMA_signal_9231 ;
    wire new_AGEMA_signal_9232 ;
    wire new_AGEMA_signal_9233 ;
    wire new_AGEMA_signal_9234 ;
    wire new_AGEMA_signal_9235 ;
    wire new_AGEMA_signal_9236 ;
    wire new_AGEMA_signal_9237 ;
    wire new_AGEMA_signal_9238 ;
    wire new_AGEMA_signal_9239 ;
    wire new_AGEMA_signal_9240 ;
    wire new_AGEMA_signal_9241 ;
    wire new_AGEMA_signal_9242 ;
    wire new_AGEMA_signal_9243 ;
    wire new_AGEMA_signal_9244 ;
    wire new_AGEMA_signal_9245 ;
    wire new_AGEMA_signal_9246 ;
    wire new_AGEMA_signal_9247 ;
    wire new_AGEMA_signal_9248 ;
    wire new_AGEMA_signal_9249 ;
    wire new_AGEMA_signal_9250 ;
    wire new_AGEMA_signal_9251 ;
    wire new_AGEMA_signal_9252 ;
    wire new_AGEMA_signal_9253 ;
    wire new_AGEMA_signal_9254 ;
    wire new_AGEMA_signal_9255 ;
    wire new_AGEMA_signal_9256 ;
    wire new_AGEMA_signal_9257 ;
    wire new_AGEMA_signal_9258 ;
    wire new_AGEMA_signal_9259 ;
    wire new_AGEMA_signal_9260 ;
    wire new_AGEMA_signal_9261 ;
    wire new_AGEMA_signal_9262 ;
    wire new_AGEMA_signal_9263 ;
    wire new_AGEMA_signal_9264 ;
    wire new_AGEMA_signal_9265 ;
    wire new_AGEMA_signal_9266 ;
    wire new_AGEMA_signal_9267 ;
    wire new_AGEMA_signal_9268 ;
    wire new_AGEMA_signal_9269 ;
    wire new_AGEMA_signal_9270 ;
    wire new_AGEMA_signal_9271 ;
    wire new_AGEMA_signal_9272 ;
    wire new_AGEMA_signal_9273 ;
    wire new_AGEMA_signal_9274 ;
    wire new_AGEMA_signal_9275 ;
    wire new_AGEMA_signal_9276 ;
    wire new_AGEMA_signal_9277 ;
    wire new_AGEMA_signal_9278 ;
    wire new_AGEMA_signal_9279 ;
    wire new_AGEMA_signal_9280 ;
    wire new_AGEMA_signal_9281 ;
    wire new_AGEMA_signal_9282 ;
    wire new_AGEMA_signal_9283 ;
    wire new_AGEMA_signal_9284 ;
    wire new_AGEMA_signal_9285 ;
    wire new_AGEMA_signal_9286 ;
    wire new_AGEMA_signal_9287 ;
    wire new_AGEMA_signal_9288 ;
    wire new_AGEMA_signal_9289 ;
    wire new_AGEMA_signal_9290 ;
    wire new_AGEMA_signal_9291 ;
    wire new_AGEMA_signal_9292 ;
    wire new_AGEMA_signal_9293 ;
    wire new_AGEMA_signal_9294 ;
    wire new_AGEMA_signal_9295 ;
    wire new_AGEMA_signal_9296 ;
    wire new_AGEMA_signal_9297 ;
    wire new_AGEMA_signal_9298 ;
    wire new_AGEMA_signal_9299 ;
    wire new_AGEMA_signal_9300 ;
    wire new_AGEMA_signal_9301 ;
    wire new_AGEMA_signal_9302 ;
    wire new_AGEMA_signal_9303 ;
    wire new_AGEMA_signal_9304 ;
    wire new_AGEMA_signal_9305 ;
    wire new_AGEMA_signal_9306 ;
    wire new_AGEMA_signal_9307 ;
    wire new_AGEMA_signal_9308 ;
    wire new_AGEMA_signal_9309 ;
    wire new_AGEMA_signal_9310 ;
    wire new_AGEMA_signal_9311 ;
    wire new_AGEMA_signal_9312 ;
    wire new_AGEMA_signal_9313 ;
    wire new_AGEMA_signal_9314 ;
    wire new_AGEMA_signal_9315 ;
    wire new_AGEMA_signal_9316 ;
    wire new_AGEMA_signal_9317 ;
    wire new_AGEMA_signal_9318 ;
    wire new_AGEMA_signal_9319 ;
    wire new_AGEMA_signal_9320 ;
    wire new_AGEMA_signal_9321 ;
    wire new_AGEMA_signal_9322 ;
    wire new_AGEMA_signal_9323 ;
    wire new_AGEMA_signal_9324 ;
    wire new_AGEMA_signal_9325 ;
    wire new_AGEMA_signal_9326 ;
    wire new_AGEMA_signal_9327 ;
    wire new_AGEMA_signal_9328 ;
    wire new_AGEMA_signal_9329 ;
    wire new_AGEMA_signal_9330 ;
    wire new_AGEMA_signal_9331 ;
    wire new_AGEMA_signal_9332 ;
    wire new_AGEMA_signal_9333 ;
    wire new_AGEMA_signal_9334 ;
    wire new_AGEMA_signal_9335 ;
    wire new_AGEMA_signal_9336 ;
    wire new_AGEMA_signal_9337 ;
    wire new_AGEMA_signal_9338 ;
    wire new_AGEMA_signal_9339 ;
    wire new_AGEMA_signal_9340 ;
    wire new_AGEMA_signal_9341 ;
    wire new_AGEMA_signal_9342 ;
    wire new_AGEMA_signal_9343 ;
    wire new_AGEMA_signal_9344 ;
    wire new_AGEMA_signal_9345 ;
    wire new_AGEMA_signal_9346 ;
    wire new_AGEMA_signal_9347 ;
    wire new_AGEMA_signal_9348 ;
    wire new_AGEMA_signal_9349 ;
    wire new_AGEMA_signal_9350 ;
    wire new_AGEMA_signal_9351 ;
    wire new_AGEMA_signal_9352 ;
    wire new_AGEMA_signal_9353 ;
    wire new_AGEMA_signal_9354 ;
    wire new_AGEMA_signal_9355 ;
    wire new_AGEMA_signal_9356 ;
    wire new_AGEMA_signal_9357 ;
    wire new_AGEMA_signal_9358 ;
    wire new_AGEMA_signal_9359 ;
    wire new_AGEMA_signal_9360 ;
    wire new_AGEMA_signal_9361 ;
    wire new_AGEMA_signal_9362 ;
    wire new_AGEMA_signal_9363 ;
    wire new_AGEMA_signal_9364 ;
    wire new_AGEMA_signal_9365 ;
    wire new_AGEMA_signal_9366 ;
    wire new_AGEMA_signal_9367 ;
    wire new_AGEMA_signal_9368 ;
    wire new_AGEMA_signal_9369 ;
    wire new_AGEMA_signal_9370 ;
    wire new_AGEMA_signal_9371 ;
    wire new_AGEMA_signal_9372 ;
    wire new_AGEMA_signal_9373 ;
    wire new_AGEMA_signal_9374 ;
    wire new_AGEMA_signal_9375 ;
    wire new_AGEMA_signal_9376 ;
    wire new_AGEMA_signal_9377 ;
    wire new_AGEMA_signal_9378 ;
    wire new_AGEMA_signal_9379 ;
    wire new_AGEMA_signal_9380 ;
    wire new_AGEMA_signal_9381 ;
    wire new_AGEMA_signal_9382 ;
    wire new_AGEMA_signal_9383 ;
    wire new_AGEMA_signal_9384 ;
    wire new_AGEMA_signal_9385 ;
    wire new_AGEMA_signal_9386 ;
    wire new_AGEMA_signal_9387 ;
    wire new_AGEMA_signal_9388 ;
    wire new_AGEMA_signal_9389 ;
    wire new_AGEMA_signal_9390 ;
    wire new_AGEMA_signal_9391 ;
    wire new_AGEMA_signal_9392 ;
    wire new_AGEMA_signal_9393 ;
    wire new_AGEMA_signal_9394 ;
    wire new_AGEMA_signal_9395 ;
    wire new_AGEMA_signal_9396 ;
    wire new_AGEMA_signal_9397 ;
    wire new_AGEMA_signal_9398 ;
    wire new_AGEMA_signal_9399 ;
    wire new_AGEMA_signal_9400 ;
    wire new_AGEMA_signal_9401 ;
    wire new_AGEMA_signal_9402 ;
    wire new_AGEMA_signal_9403 ;
    wire new_AGEMA_signal_9404 ;
    wire new_AGEMA_signal_9405 ;
    wire new_AGEMA_signal_9406 ;
    wire new_AGEMA_signal_9407 ;
    wire new_AGEMA_signal_9408 ;
    wire new_AGEMA_signal_9409 ;
    wire new_AGEMA_signal_9410 ;
    wire new_AGEMA_signal_9411 ;
    wire new_AGEMA_signal_9412 ;
    wire new_AGEMA_signal_9413 ;
    wire new_AGEMA_signal_9414 ;
    wire new_AGEMA_signal_9415 ;
    wire new_AGEMA_signal_9416 ;
    wire new_AGEMA_signal_9417 ;
    wire new_AGEMA_signal_9418 ;
    wire new_AGEMA_signal_9419 ;
    wire new_AGEMA_signal_9420 ;
    wire new_AGEMA_signal_9421 ;
    wire new_AGEMA_signal_9422 ;
    wire new_AGEMA_signal_9423 ;
    wire new_AGEMA_signal_9424 ;
    wire new_AGEMA_signal_9425 ;
    wire new_AGEMA_signal_9426 ;
    wire new_AGEMA_signal_9427 ;
    wire new_AGEMA_signal_9428 ;
    wire new_AGEMA_signal_9429 ;
    wire new_AGEMA_signal_9430 ;
    wire new_AGEMA_signal_9431 ;
    wire new_AGEMA_signal_9432 ;
    wire new_AGEMA_signal_9433 ;
    wire new_AGEMA_signal_9434 ;
    wire new_AGEMA_signal_9435 ;
    wire new_AGEMA_signal_9436 ;
    wire new_AGEMA_signal_9437 ;
    wire new_AGEMA_signal_9438 ;
    wire new_AGEMA_signal_9439 ;
    wire new_AGEMA_signal_9440 ;
    wire new_AGEMA_signal_9441 ;
    wire new_AGEMA_signal_9442 ;
    wire new_AGEMA_signal_9443 ;
    wire new_AGEMA_signal_9444 ;
    wire new_AGEMA_signal_9445 ;
    wire new_AGEMA_signal_9446 ;
    wire new_AGEMA_signal_9447 ;
    wire new_AGEMA_signal_9448 ;
    wire new_AGEMA_signal_9449 ;
    wire new_AGEMA_signal_9450 ;
    wire new_AGEMA_signal_9451 ;
    wire new_AGEMA_signal_9452 ;
    wire new_AGEMA_signal_9453 ;
    wire new_AGEMA_signal_9454 ;
    wire new_AGEMA_signal_9455 ;
    wire new_AGEMA_signal_9456 ;
    wire new_AGEMA_signal_9457 ;
    wire new_AGEMA_signal_9458 ;
    wire new_AGEMA_signal_9459 ;
    wire new_AGEMA_signal_9460 ;
    wire new_AGEMA_signal_9461 ;
    wire new_AGEMA_signal_9462 ;
    wire new_AGEMA_signal_9463 ;
    wire new_AGEMA_signal_9464 ;
    wire new_AGEMA_signal_9465 ;
    wire new_AGEMA_signal_9466 ;
    wire new_AGEMA_signal_9467 ;
    wire new_AGEMA_signal_9468 ;
    wire new_AGEMA_signal_9469 ;
    wire new_AGEMA_signal_9470 ;
    wire new_AGEMA_signal_9471 ;
    wire new_AGEMA_signal_9472 ;
    wire new_AGEMA_signal_9473 ;
    wire new_AGEMA_signal_9474 ;
    wire new_AGEMA_signal_9475 ;
    wire new_AGEMA_signal_9476 ;
    wire new_AGEMA_signal_9477 ;
    wire new_AGEMA_signal_9478 ;
    wire new_AGEMA_signal_9479 ;
    wire new_AGEMA_signal_9480 ;
    wire new_AGEMA_signal_9481 ;
    wire new_AGEMA_signal_9482 ;
    wire new_AGEMA_signal_9483 ;
    wire new_AGEMA_signal_9484 ;
    wire new_AGEMA_signal_9485 ;
    wire new_AGEMA_signal_9486 ;
    wire new_AGEMA_signal_9487 ;
    wire new_AGEMA_signal_9488 ;
    wire new_AGEMA_signal_9489 ;
    wire new_AGEMA_signal_9490 ;
    wire new_AGEMA_signal_9491 ;
    wire new_AGEMA_signal_9492 ;
    wire new_AGEMA_signal_9493 ;
    wire new_AGEMA_signal_9494 ;
    wire new_AGEMA_signal_9495 ;
    wire new_AGEMA_signal_9496 ;
    wire new_AGEMA_signal_9497 ;
    wire new_AGEMA_signal_9498 ;
    wire new_AGEMA_signal_9499 ;
    wire new_AGEMA_signal_9500 ;
    wire new_AGEMA_signal_9501 ;
    wire new_AGEMA_signal_9502 ;
    wire new_AGEMA_signal_9503 ;
    wire new_AGEMA_signal_9504 ;
    wire new_AGEMA_signal_9505 ;
    wire new_AGEMA_signal_9506 ;
    wire new_AGEMA_signal_9507 ;
    wire new_AGEMA_signal_9508 ;
    wire new_AGEMA_signal_9509 ;
    wire new_AGEMA_signal_9510 ;
    wire new_AGEMA_signal_9511 ;
    wire new_AGEMA_signal_9512 ;
    wire new_AGEMA_signal_9513 ;
    wire new_AGEMA_signal_9514 ;
    wire new_AGEMA_signal_9515 ;
    wire new_AGEMA_signal_9516 ;
    wire new_AGEMA_signal_9517 ;
    wire new_AGEMA_signal_9518 ;
    wire new_AGEMA_signal_9519 ;
    wire new_AGEMA_signal_9520 ;
    wire new_AGEMA_signal_9521 ;
    wire new_AGEMA_signal_9522 ;
    wire new_AGEMA_signal_9523 ;
    wire new_AGEMA_signal_9524 ;
    wire new_AGEMA_signal_9525 ;
    wire new_AGEMA_signal_9526 ;
    wire new_AGEMA_signal_9527 ;
    wire new_AGEMA_signal_9528 ;
    wire new_AGEMA_signal_9529 ;
    wire new_AGEMA_signal_9530 ;
    wire new_AGEMA_signal_9531 ;
    wire new_AGEMA_signal_9532 ;
    wire new_AGEMA_signal_9533 ;
    wire new_AGEMA_signal_9534 ;
    wire new_AGEMA_signal_9535 ;
    wire new_AGEMA_signal_9536 ;
    wire new_AGEMA_signal_9537 ;
    wire new_AGEMA_signal_9538 ;
    wire new_AGEMA_signal_9539 ;
    wire new_AGEMA_signal_9540 ;
    wire new_AGEMA_signal_9541 ;
    wire new_AGEMA_signal_9542 ;
    wire new_AGEMA_signal_9543 ;
    wire new_AGEMA_signal_9544 ;
    wire new_AGEMA_signal_9545 ;
    wire new_AGEMA_signal_9546 ;
    wire new_AGEMA_signal_9547 ;
    wire new_AGEMA_signal_9548 ;
    wire new_AGEMA_signal_9549 ;
    wire new_AGEMA_signal_9550 ;
    wire new_AGEMA_signal_9551 ;
    wire new_AGEMA_signal_9552 ;
    wire new_AGEMA_signal_9553 ;
    wire new_AGEMA_signal_9554 ;
    wire new_AGEMA_signal_9555 ;
    wire new_AGEMA_signal_9556 ;
    wire new_AGEMA_signal_9557 ;
    wire new_AGEMA_signal_9558 ;
    wire new_AGEMA_signal_9559 ;
    wire new_AGEMA_signal_9560 ;
    wire new_AGEMA_signal_9561 ;
    wire new_AGEMA_signal_9562 ;
    wire new_AGEMA_signal_9563 ;
    wire new_AGEMA_signal_9564 ;
    wire new_AGEMA_signal_9565 ;
    wire new_AGEMA_signal_9566 ;
    wire new_AGEMA_signal_9567 ;
    wire new_AGEMA_signal_9568 ;
    wire new_AGEMA_signal_9569 ;
    wire new_AGEMA_signal_9570 ;
    wire new_AGEMA_signal_9571 ;
    wire new_AGEMA_signal_9572 ;
    wire new_AGEMA_signal_9573 ;
    wire new_AGEMA_signal_9574 ;
    wire new_AGEMA_signal_9575 ;
    wire new_AGEMA_signal_9576 ;
    wire new_AGEMA_signal_9577 ;
    wire new_AGEMA_signal_9578 ;
    wire new_AGEMA_signal_9579 ;
    wire new_AGEMA_signal_9580 ;
    wire new_AGEMA_signal_9581 ;
    wire new_AGEMA_signal_9582 ;
    wire new_AGEMA_signal_9583 ;
    wire new_AGEMA_signal_9584 ;
    wire new_AGEMA_signal_9585 ;
    wire new_AGEMA_signal_9586 ;
    wire new_AGEMA_signal_9587 ;
    wire new_AGEMA_signal_9588 ;
    wire new_AGEMA_signal_9589 ;
    wire new_AGEMA_signal_9590 ;
    wire new_AGEMA_signal_9591 ;
    wire new_AGEMA_signal_9592 ;
    wire new_AGEMA_signal_9593 ;
    wire new_AGEMA_signal_9594 ;
    wire new_AGEMA_signal_9595 ;
    wire new_AGEMA_signal_9596 ;
    wire new_AGEMA_signal_9597 ;
    wire new_AGEMA_signal_9598 ;
    wire new_AGEMA_signal_9599 ;
    wire new_AGEMA_signal_9600 ;
    wire new_AGEMA_signal_9601 ;
    wire new_AGEMA_signal_9602 ;
    wire new_AGEMA_signal_9603 ;
    wire new_AGEMA_signal_9604 ;
    wire new_AGEMA_signal_9605 ;
    wire new_AGEMA_signal_9606 ;
    wire new_AGEMA_signal_9607 ;
    wire new_AGEMA_signal_9608 ;
    wire new_AGEMA_signal_9609 ;
    wire new_AGEMA_signal_9610 ;
    wire new_AGEMA_signal_9611 ;
    wire new_AGEMA_signal_9612 ;
    wire new_AGEMA_signal_9613 ;
    wire new_AGEMA_signal_9614 ;
    wire new_AGEMA_signal_9615 ;
    wire new_AGEMA_signal_9616 ;
    wire new_AGEMA_signal_9617 ;
    wire new_AGEMA_signal_9618 ;
    wire new_AGEMA_signal_9619 ;
    wire new_AGEMA_signal_9620 ;
    wire new_AGEMA_signal_9621 ;
    wire new_AGEMA_signal_9622 ;
    wire new_AGEMA_signal_9623 ;
    wire new_AGEMA_signal_9624 ;
    wire new_AGEMA_signal_9625 ;
    wire new_AGEMA_signal_9626 ;
    wire new_AGEMA_signal_9627 ;
    wire new_AGEMA_signal_9628 ;
    wire new_AGEMA_signal_9629 ;
    wire new_AGEMA_signal_9630 ;
    wire new_AGEMA_signal_9631 ;
    wire new_AGEMA_signal_9632 ;
    wire new_AGEMA_signal_9633 ;
    wire new_AGEMA_signal_9634 ;
    wire new_AGEMA_signal_9635 ;
    wire new_AGEMA_signal_9636 ;
    wire new_AGEMA_signal_9637 ;
    wire new_AGEMA_signal_9638 ;
    wire new_AGEMA_signal_9639 ;
    wire new_AGEMA_signal_9640 ;
    wire new_AGEMA_signal_9641 ;
    wire new_AGEMA_signal_9642 ;
    wire new_AGEMA_signal_9643 ;
    wire new_AGEMA_signal_9644 ;
    wire new_AGEMA_signal_9645 ;
    wire new_AGEMA_signal_9646 ;
    wire new_AGEMA_signal_9647 ;
    wire new_AGEMA_signal_9648 ;
    wire new_AGEMA_signal_9649 ;
    wire new_AGEMA_signal_9650 ;
    wire new_AGEMA_signal_9651 ;
    wire new_AGEMA_signal_9652 ;
    wire new_AGEMA_signal_9653 ;
    wire new_AGEMA_signal_9654 ;
    wire new_AGEMA_signal_9655 ;
    wire new_AGEMA_signal_9656 ;
    wire new_AGEMA_signal_9657 ;
    wire new_AGEMA_signal_9658 ;
    wire new_AGEMA_signal_9659 ;
    wire new_AGEMA_signal_9660 ;
    wire new_AGEMA_signal_9661 ;
    wire new_AGEMA_signal_9662 ;
    wire new_AGEMA_signal_9663 ;
    wire new_AGEMA_signal_9664 ;
    wire new_AGEMA_signal_9665 ;
    wire new_AGEMA_signal_9666 ;
    wire new_AGEMA_signal_9667 ;
    wire new_AGEMA_signal_9668 ;
    wire new_AGEMA_signal_9669 ;
    wire new_AGEMA_signal_9670 ;
    wire new_AGEMA_signal_9671 ;
    wire new_AGEMA_signal_9672 ;
    wire new_AGEMA_signal_9673 ;
    wire new_AGEMA_signal_9674 ;
    wire new_AGEMA_signal_9675 ;
    wire new_AGEMA_signal_9676 ;
    wire new_AGEMA_signal_9677 ;
    wire new_AGEMA_signal_9678 ;
    wire new_AGEMA_signal_9679 ;
    wire new_AGEMA_signal_9680 ;
    wire new_AGEMA_signal_9681 ;
    wire new_AGEMA_signal_9682 ;
    wire new_AGEMA_signal_9683 ;
    wire new_AGEMA_signal_9684 ;
    wire new_AGEMA_signal_9685 ;
    wire new_AGEMA_signal_9686 ;
    wire new_AGEMA_signal_9687 ;
    wire new_AGEMA_signal_9688 ;
    wire new_AGEMA_signal_9689 ;
    wire new_AGEMA_signal_9690 ;
    wire new_AGEMA_signal_9691 ;
    wire new_AGEMA_signal_9692 ;
    wire new_AGEMA_signal_9693 ;
    wire new_AGEMA_signal_9694 ;
    wire new_AGEMA_signal_9695 ;
    wire new_AGEMA_signal_9696 ;
    wire new_AGEMA_signal_9697 ;
    wire new_AGEMA_signal_9698 ;
    wire new_AGEMA_signal_9699 ;
    wire new_AGEMA_signal_9700 ;
    wire new_AGEMA_signal_9701 ;
    wire new_AGEMA_signal_9702 ;
    wire new_AGEMA_signal_9703 ;
    wire new_AGEMA_signal_9704 ;
    wire new_AGEMA_signal_9705 ;
    wire new_AGEMA_signal_9706 ;
    wire new_AGEMA_signal_9707 ;
    wire new_AGEMA_signal_9708 ;
    wire new_AGEMA_signal_9709 ;
    wire new_AGEMA_signal_9710 ;
    wire new_AGEMA_signal_9711 ;
    wire new_AGEMA_signal_9712 ;
    wire new_AGEMA_signal_9713 ;
    wire new_AGEMA_signal_9714 ;
    wire new_AGEMA_signal_9715 ;
    wire new_AGEMA_signal_9716 ;
    wire new_AGEMA_signal_9717 ;
    wire new_AGEMA_signal_9718 ;
    wire new_AGEMA_signal_9719 ;
    wire new_AGEMA_signal_9720 ;
    wire new_AGEMA_signal_9721 ;
    wire new_AGEMA_signal_9722 ;
    wire new_AGEMA_signal_9723 ;
    wire new_AGEMA_signal_9724 ;
    wire new_AGEMA_signal_9725 ;
    wire new_AGEMA_signal_9726 ;
    wire new_AGEMA_signal_9727 ;
    wire new_AGEMA_signal_9728 ;
    wire new_AGEMA_signal_9729 ;
    wire new_AGEMA_signal_9730 ;
    wire new_AGEMA_signal_9731 ;
    wire new_AGEMA_signal_9732 ;
    wire new_AGEMA_signal_9733 ;
    wire new_AGEMA_signal_9734 ;
    wire new_AGEMA_signal_9735 ;
    wire new_AGEMA_signal_9736 ;
    wire new_AGEMA_signal_9737 ;
    wire new_AGEMA_signal_9738 ;
    wire new_AGEMA_signal_9739 ;
    wire new_AGEMA_signal_9740 ;
    wire new_AGEMA_signal_9741 ;
    wire new_AGEMA_signal_9742 ;
    wire new_AGEMA_signal_9743 ;
    wire new_AGEMA_signal_9744 ;
    wire new_AGEMA_signal_9745 ;
    wire new_AGEMA_signal_9746 ;
    wire new_AGEMA_signal_9747 ;
    wire new_AGEMA_signal_9748 ;
    wire new_AGEMA_signal_9749 ;
    wire new_AGEMA_signal_9750 ;
    wire new_AGEMA_signal_9751 ;
    wire new_AGEMA_signal_9752 ;
    wire new_AGEMA_signal_9753 ;
    wire new_AGEMA_signal_9754 ;
    wire new_AGEMA_signal_9755 ;
    wire new_AGEMA_signal_9756 ;
    wire new_AGEMA_signal_9757 ;
    wire new_AGEMA_signal_9758 ;
    wire new_AGEMA_signal_9759 ;
    wire new_AGEMA_signal_9760 ;
    wire new_AGEMA_signal_9761 ;
    wire new_AGEMA_signal_9762 ;
    wire new_AGEMA_signal_9763 ;
    wire new_AGEMA_signal_9764 ;
    wire new_AGEMA_signal_9765 ;
    wire new_AGEMA_signal_9766 ;
    wire new_AGEMA_signal_9767 ;
    wire new_AGEMA_signal_9768 ;
    wire new_AGEMA_signal_9769 ;
    wire new_AGEMA_signal_9770 ;
    wire new_AGEMA_signal_9771 ;
    wire new_AGEMA_signal_9772 ;
    wire new_AGEMA_signal_9773 ;
    wire new_AGEMA_signal_9774 ;
    wire new_AGEMA_signal_9775 ;
    wire new_AGEMA_signal_9776 ;
    wire new_AGEMA_signal_9777 ;
    wire new_AGEMA_signal_9778 ;
    wire new_AGEMA_signal_9779 ;
    wire new_AGEMA_signal_9780 ;
    wire new_AGEMA_signal_9781 ;
    wire new_AGEMA_signal_9782 ;
    wire new_AGEMA_signal_9783 ;
    wire new_AGEMA_signal_9784 ;
    wire new_AGEMA_signal_9785 ;
    wire new_AGEMA_signal_9786 ;
    wire new_AGEMA_signal_9787 ;
    wire new_AGEMA_signal_9788 ;
    wire new_AGEMA_signal_9789 ;
    wire new_AGEMA_signal_9790 ;
    wire new_AGEMA_signal_9791 ;
    wire new_AGEMA_signal_9792 ;
    wire new_AGEMA_signal_9793 ;
    wire new_AGEMA_signal_9794 ;
    wire new_AGEMA_signal_9795 ;
    wire new_AGEMA_signal_9796 ;
    wire new_AGEMA_signal_9797 ;
    wire new_AGEMA_signal_9798 ;
    wire new_AGEMA_signal_9799 ;
    wire new_AGEMA_signal_9800 ;
    wire new_AGEMA_signal_9801 ;
    wire new_AGEMA_signal_9802 ;
    wire new_AGEMA_signal_9803 ;
    wire new_AGEMA_signal_9804 ;
    wire new_AGEMA_signal_9805 ;
    wire new_AGEMA_signal_9806 ;
    wire new_AGEMA_signal_9807 ;
    wire new_AGEMA_signal_9808 ;
    wire new_AGEMA_signal_9809 ;
    wire new_AGEMA_signal_9810 ;
    wire new_AGEMA_signal_9811 ;
    wire new_AGEMA_signal_9812 ;
    wire new_AGEMA_signal_9813 ;
    wire new_AGEMA_signal_9814 ;
    wire new_AGEMA_signal_9815 ;
    wire new_AGEMA_signal_9816 ;
    wire new_AGEMA_signal_9817 ;
    wire new_AGEMA_signal_9818 ;
    wire new_AGEMA_signal_9819 ;
    wire new_AGEMA_signal_9820 ;
    wire new_AGEMA_signal_9821 ;
    wire new_AGEMA_signal_9822 ;
    wire new_AGEMA_signal_9823 ;
    wire new_AGEMA_signal_9824 ;
    wire new_AGEMA_signal_9825 ;
    wire new_AGEMA_signal_9826 ;
    wire new_AGEMA_signal_9827 ;
    wire new_AGEMA_signal_9828 ;
    wire new_AGEMA_signal_9829 ;
    wire new_AGEMA_signal_9830 ;
    wire new_AGEMA_signal_9831 ;
    wire new_AGEMA_signal_9832 ;
    wire new_AGEMA_signal_9833 ;
    wire new_AGEMA_signal_9834 ;
    wire new_AGEMA_signal_9835 ;
    wire new_AGEMA_signal_9836 ;
    wire new_AGEMA_signal_9837 ;
    wire new_AGEMA_signal_9838 ;
    wire new_AGEMA_signal_9839 ;
    wire new_AGEMA_signal_9840 ;
    wire new_AGEMA_signal_9841 ;
    wire new_AGEMA_signal_9842 ;
    wire new_AGEMA_signal_9843 ;
    wire new_AGEMA_signal_9844 ;
    wire new_AGEMA_signal_9845 ;
    wire new_AGEMA_signal_9846 ;
    wire new_AGEMA_signal_9847 ;
    wire new_AGEMA_signal_9848 ;
    wire new_AGEMA_signal_9849 ;
    wire new_AGEMA_signal_9850 ;
    wire new_AGEMA_signal_9851 ;
    wire new_AGEMA_signal_9852 ;
    wire new_AGEMA_signal_9853 ;
    wire new_AGEMA_signal_9854 ;
    wire new_AGEMA_signal_9855 ;
    wire new_AGEMA_signal_9856 ;
    wire new_AGEMA_signal_9857 ;
    wire new_AGEMA_signal_9858 ;
    wire new_AGEMA_signal_9859 ;
    wire new_AGEMA_signal_9860 ;
    wire new_AGEMA_signal_9861 ;
    wire new_AGEMA_signal_9862 ;
    wire new_AGEMA_signal_9863 ;
    wire new_AGEMA_signal_9864 ;
    wire new_AGEMA_signal_9865 ;
    wire new_AGEMA_signal_9866 ;
    wire new_AGEMA_signal_9867 ;
    wire new_AGEMA_signal_9868 ;
    wire new_AGEMA_signal_9869 ;
    wire new_AGEMA_signal_9870 ;
    wire new_AGEMA_signal_9871 ;
    wire new_AGEMA_signal_9872 ;
    wire new_AGEMA_signal_9873 ;
    wire new_AGEMA_signal_9874 ;
    wire new_AGEMA_signal_9875 ;
    wire new_AGEMA_signal_9876 ;
    wire new_AGEMA_signal_9877 ;
    wire new_AGEMA_signal_9878 ;
    wire new_AGEMA_signal_9879 ;
    wire new_AGEMA_signal_9880 ;
    wire new_AGEMA_signal_9881 ;
    wire new_AGEMA_signal_9882 ;
    wire new_AGEMA_signal_9883 ;
    wire new_AGEMA_signal_9884 ;
    wire new_AGEMA_signal_9885 ;
    wire new_AGEMA_signal_9886 ;
    wire new_AGEMA_signal_9887 ;
    wire new_AGEMA_signal_9888 ;
    wire new_AGEMA_signal_9889 ;
    wire new_AGEMA_signal_9890 ;
    wire new_AGEMA_signal_9891 ;
    wire new_AGEMA_signal_9892 ;
    wire new_AGEMA_signal_9893 ;
    wire new_AGEMA_signal_9894 ;
    wire new_AGEMA_signal_9895 ;
    wire new_AGEMA_signal_9896 ;
    wire new_AGEMA_signal_9897 ;
    wire new_AGEMA_signal_9898 ;
    wire new_AGEMA_signal_9899 ;
    wire new_AGEMA_signal_9900 ;
    wire new_AGEMA_signal_9901 ;
    wire new_AGEMA_signal_9902 ;
    wire new_AGEMA_signal_9903 ;
    wire new_AGEMA_signal_9904 ;
    wire new_AGEMA_signal_9905 ;
    wire new_AGEMA_signal_9906 ;
    wire new_AGEMA_signal_9907 ;
    wire new_AGEMA_signal_9908 ;
    wire new_AGEMA_signal_9909 ;
    wire new_AGEMA_signal_9910 ;
    wire new_AGEMA_signal_9911 ;
    wire new_AGEMA_signal_9912 ;
    wire new_AGEMA_signal_9913 ;
    wire new_AGEMA_signal_9914 ;
    wire new_AGEMA_signal_9915 ;
    wire new_AGEMA_signal_9916 ;
    wire new_AGEMA_signal_9917 ;
    wire new_AGEMA_signal_9918 ;
    wire new_AGEMA_signal_9919 ;
    wire new_AGEMA_signal_9920 ;
    wire new_AGEMA_signal_9921 ;
    wire new_AGEMA_signal_9922 ;
    wire new_AGEMA_signal_9923 ;
    wire new_AGEMA_signal_9924 ;
    wire new_AGEMA_signal_9925 ;
    wire new_AGEMA_signal_9926 ;
    wire new_AGEMA_signal_9927 ;
    wire new_AGEMA_signal_9928 ;
    wire new_AGEMA_signal_9929 ;
    wire new_AGEMA_signal_9930 ;
    wire new_AGEMA_signal_9931 ;
    wire new_AGEMA_signal_9932 ;
    wire new_AGEMA_signal_9933 ;
    wire new_AGEMA_signal_9934 ;
    wire new_AGEMA_signal_9935 ;
    wire new_AGEMA_signal_9936 ;
    wire new_AGEMA_signal_9937 ;
    wire new_AGEMA_signal_9938 ;
    wire new_AGEMA_signal_9939 ;
    wire new_AGEMA_signal_9940 ;
    wire new_AGEMA_signal_9941 ;
    wire new_AGEMA_signal_9942 ;
    wire new_AGEMA_signal_9943 ;
    wire new_AGEMA_signal_9944 ;
    wire new_AGEMA_signal_9945 ;
    wire new_AGEMA_signal_9946 ;
    wire new_AGEMA_signal_9947 ;
    wire new_AGEMA_signal_9948 ;
    wire new_AGEMA_signal_9949 ;
    wire new_AGEMA_signal_9950 ;
    wire new_AGEMA_signal_9951 ;
    wire new_AGEMA_signal_9952 ;
    wire new_AGEMA_signal_9953 ;
    wire new_AGEMA_signal_9954 ;
    wire new_AGEMA_signal_9955 ;
    wire new_AGEMA_signal_9956 ;
    wire new_AGEMA_signal_9957 ;
    wire new_AGEMA_signal_9958 ;
    wire new_AGEMA_signal_9959 ;
    wire new_AGEMA_signal_9960 ;
    wire new_AGEMA_signal_9961 ;
    wire new_AGEMA_signal_9962 ;
    wire new_AGEMA_signal_9963 ;
    wire new_AGEMA_signal_9964 ;
    wire new_AGEMA_signal_9965 ;
    wire new_AGEMA_signal_9966 ;
    wire new_AGEMA_signal_9967 ;
    wire new_AGEMA_signal_9968 ;
    wire new_AGEMA_signal_9969 ;
    wire new_AGEMA_signal_9970 ;
    wire new_AGEMA_signal_9971 ;
    wire new_AGEMA_signal_9972 ;
    wire new_AGEMA_signal_9973 ;
    wire new_AGEMA_signal_9974 ;
    wire new_AGEMA_signal_9975 ;
    wire new_AGEMA_signal_9976 ;
    wire new_AGEMA_signal_9977 ;
    wire new_AGEMA_signal_9978 ;
    wire new_AGEMA_signal_9979 ;
    wire new_AGEMA_signal_9980 ;
    wire new_AGEMA_signal_9981 ;
    wire new_AGEMA_signal_9982 ;
    wire new_AGEMA_signal_9983 ;
    wire new_AGEMA_signal_9984 ;
    wire new_AGEMA_signal_9985 ;
    wire new_AGEMA_signal_9986 ;
    wire new_AGEMA_signal_9987 ;
    wire new_AGEMA_signal_9988 ;
    wire new_AGEMA_signal_9989 ;
    wire new_AGEMA_signal_9990 ;
    wire new_AGEMA_signal_9991 ;
    wire new_AGEMA_signal_9992 ;
    wire new_AGEMA_signal_9993 ;
    wire new_AGEMA_signal_9994 ;
    wire new_AGEMA_signal_9995 ;
    wire new_AGEMA_signal_9996 ;
    wire new_AGEMA_signal_9997 ;
    wire new_AGEMA_signal_9998 ;
    wire new_AGEMA_signal_9999 ;
    wire new_AGEMA_signal_10000 ;
    wire new_AGEMA_signal_10001 ;
    wire new_AGEMA_signal_10002 ;
    wire new_AGEMA_signal_10003 ;
    wire new_AGEMA_signal_10004 ;
    wire new_AGEMA_signal_10005 ;
    wire new_AGEMA_signal_10006 ;
    wire new_AGEMA_signal_10007 ;
    wire new_AGEMA_signal_10008 ;
    wire new_AGEMA_signal_10009 ;
    wire new_AGEMA_signal_10010 ;
    wire new_AGEMA_signal_10011 ;
    wire new_AGEMA_signal_10012 ;
    wire new_AGEMA_signal_10013 ;
    wire new_AGEMA_signal_10014 ;
    wire new_AGEMA_signal_10015 ;
    wire new_AGEMA_signal_10016 ;
    wire new_AGEMA_signal_10017 ;
    wire new_AGEMA_signal_10018 ;
    wire new_AGEMA_signal_10019 ;
    wire new_AGEMA_signal_10020 ;
    wire new_AGEMA_signal_10021 ;
    wire new_AGEMA_signal_10022 ;
    wire new_AGEMA_signal_10023 ;
    wire new_AGEMA_signal_10024 ;
    wire new_AGEMA_signal_10025 ;
    wire new_AGEMA_signal_10026 ;
    wire new_AGEMA_signal_10027 ;
    wire new_AGEMA_signal_10028 ;
    wire new_AGEMA_signal_10029 ;
    wire new_AGEMA_signal_10030 ;
    wire new_AGEMA_signal_10031 ;
    wire new_AGEMA_signal_10032 ;
    wire new_AGEMA_signal_10033 ;
    wire new_AGEMA_signal_10034 ;
    wire new_AGEMA_signal_10035 ;
    wire new_AGEMA_signal_10036 ;
    wire new_AGEMA_signal_10037 ;
    wire new_AGEMA_signal_10038 ;
    wire new_AGEMA_signal_10039 ;
    wire new_AGEMA_signal_10040 ;
    wire new_AGEMA_signal_10041 ;
    wire new_AGEMA_signal_10042 ;
    wire new_AGEMA_signal_10043 ;
    wire new_AGEMA_signal_10044 ;
    wire new_AGEMA_signal_10045 ;
    wire new_AGEMA_signal_10046 ;
    wire new_AGEMA_signal_10047 ;
    wire new_AGEMA_signal_10048 ;
    wire new_AGEMA_signal_10049 ;
    wire new_AGEMA_signal_10050 ;
    wire new_AGEMA_signal_10051 ;
    wire new_AGEMA_signal_10052 ;
    wire new_AGEMA_signal_10053 ;
    wire new_AGEMA_signal_10054 ;
    wire new_AGEMA_signal_10055 ;
    wire new_AGEMA_signal_10056 ;
    wire new_AGEMA_signal_10057 ;
    wire new_AGEMA_signal_10058 ;
    wire new_AGEMA_signal_10059 ;
    wire new_AGEMA_signal_10060 ;
    wire new_AGEMA_signal_10061 ;
    wire new_AGEMA_signal_10062 ;
    wire new_AGEMA_signal_10063 ;
    wire new_AGEMA_signal_10064 ;
    wire new_AGEMA_signal_10065 ;
    wire new_AGEMA_signal_10066 ;
    wire new_AGEMA_signal_10067 ;
    wire new_AGEMA_signal_10068 ;
    wire new_AGEMA_signal_10069 ;
    wire new_AGEMA_signal_10070 ;
    wire new_AGEMA_signal_10071 ;
    wire new_AGEMA_signal_10072 ;
    wire new_AGEMA_signal_10073 ;
    wire new_AGEMA_signal_10074 ;
    wire new_AGEMA_signal_10075 ;
    wire new_AGEMA_signal_10076 ;
    wire new_AGEMA_signal_10077 ;
    wire new_AGEMA_signal_10078 ;
    wire new_AGEMA_signal_10079 ;
    wire new_AGEMA_signal_10080 ;
    wire new_AGEMA_signal_10081 ;
    wire new_AGEMA_signal_10082 ;
    wire new_AGEMA_signal_10083 ;
    wire new_AGEMA_signal_10084 ;
    wire new_AGEMA_signal_10085 ;
    wire new_AGEMA_signal_10086 ;
    wire new_AGEMA_signal_10087 ;
    wire new_AGEMA_signal_10088 ;
    wire new_AGEMA_signal_10089 ;
    wire new_AGEMA_signal_10090 ;
    wire new_AGEMA_signal_10091 ;
    wire new_AGEMA_signal_10092 ;
    wire new_AGEMA_signal_10093 ;
    wire new_AGEMA_signal_10094 ;
    wire new_AGEMA_signal_10095 ;
    wire new_AGEMA_signal_10096 ;
    wire new_AGEMA_signal_10097 ;
    wire new_AGEMA_signal_10098 ;
    wire new_AGEMA_signal_10099 ;
    wire new_AGEMA_signal_10100 ;
    wire new_AGEMA_signal_10101 ;
    wire new_AGEMA_signal_10102 ;
    wire new_AGEMA_signal_10103 ;
    wire new_AGEMA_signal_10104 ;
    wire new_AGEMA_signal_10105 ;
    wire new_AGEMA_signal_10106 ;
    wire new_AGEMA_signal_10107 ;
    wire new_AGEMA_signal_10108 ;
    wire new_AGEMA_signal_10109 ;
    wire new_AGEMA_signal_10110 ;
    wire new_AGEMA_signal_10111 ;
    wire new_AGEMA_signal_10112 ;
    wire new_AGEMA_signal_10113 ;
    wire new_AGEMA_signal_10114 ;
    wire new_AGEMA_signal_10115 ;
    wire new_AGEMA_signal_10116 ;
    wire new_AGEMA_signal_10117 ;
    wire new_AGEMA_signal_10118 ;
    wire new_AGEMA_signal_10119 ;
    wire new_AGEMA_signal_10120 ;
    wire new_AGEMA_signal_10121 ;
    wire new_AGEMA_signal_10122 ;
    wire new_AGEMA_signal_10123 ;
    wire new_AGEMA_signal_10124 ;
    wire new_AGEMA_signal_10125 ;
    wire new_AGEMA_signal_10126 ;
    wire new_AGEMA_signal_10127 ;
    wire new_AGEMA_signal_10128 ;
    wire new_AGEMA_signal_10129 ;
    wire new_AGEMA_signal_10130 ;
    wire new_AGEMA_signal_10131 ;
    wire new_AGEMA_signal_10132 ;
    wire new_AGEMA_signal_10133 ;
    wire new_AGEMA_signal_10134 ;
    wire new_AGEMA_signal_10135 ;
    wire new_AGEMA_signal_10136 ;
    wire new_AGEMA_signal_10137 ;
    wire new_AGEMA_signal_10138 ;
    wire new_AGEMA_signal_10139 ;
    wire new_AGEMA_signal_10140 ;
    wire new_AGEMA_signal_10141 ;
    wire new_AGEMA_signal_10142 ;
    wire new_AGEMA_signal_10143 ;
    wire new_AGEMA_signal_10144 ;
    wire new_AGEMA_signal_10145 ;
    wire new_AGEMA_signal_10146 ;
    wire new_AGEMA_signal_10147 ;
    wire new_AGEMA_signal_10148 ;
    wire new_AGEMA_signal_10149 ;
    wire new_AGEMA_signal_10150 ;
    wire new_AGEMA_signal_10151 ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U64 ( .a ({key_s2[73], key_s1[73], key_s0[73]}), .b ({key_s2[9], key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_1461, new_AGEMA_signal_1460, wk[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U63 ( .a ({key_s2[72], key_s1[72], key_s0[72]}), .b ({key_s2[8], key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, wk[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U62 ( .a ({key_s2[71], key_s1[71], key_s0[71]}), .b ({key_s2[7], key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, wk[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U61 ( .a ({key_s2[6], key_s1[6], key_s0[6]}), .b ({key_s2[70], key_s1[70], key_s0[70]}), .c ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, wk[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U60 ( .a ({key_s2[127], key_s1[127], key_s0[127]}), .b ({key_s2[63], key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, wk[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U59 ( .a ({key_s2[126], key_s1[126], key_s0[126]}), .b ({key_s2[62], key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, wk[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U58 ( .a ({key_s2[125], key_s1[125], key_s0[125]}), .b ({key_s2[61], key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, wk[61]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U57 ( .a ({key_s2[124], key_s1[124], key_s0[124]}), .b ({key_s2[60], key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_1503, new_AGEMA_signal_1502, wk[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U56 ( .a ({key_s2[5], key_s1[5], key_s0[5]}), .b ({key_s2[69], key_s1[69], key_s0[69]}), .c ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, wk[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U55 ( .a ({key_s2[123], key_s1[123], key_s0[123]}), .b ({key_s2[59], key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, wk[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U54 ( .a ({key_s2[122], key_s1[122], key_s0[122]}), .b ({key_s2[58], key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_1521, new_AGEMA_signal_1520, wk[58]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U53 ( .a ({key_s2[121], key_s1[121], key_s0[121]}), .b ({key_s2[57], key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, wk[57]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U52 ( .a ({key_s2[120], key_s1[120], key_s0[120]}), .b ({key_s2[56], key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_1533, new_AGEMA_signal_1532, wk[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U51 ( .a ({key_s2[119], key_s1[119], key_s0[119]}), .b ({key_s2[55], key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_1539, new_AGEMA_signal_1538, wk[55]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U50 ( .a ({key_s2[118], key_s1[118], key_s0[118]}), .b ({key_s2[54], key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, wk[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U49 ( .a ({key_s2[117], key_s1[117], key_s0[117]}), .b ({key_s2[53], key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, wk[53]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U48 ( .a ({key_s2[116], key_s1[116], key_s0[116]}), .b ({key_s2[52], key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, wk[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U47 ( .a ({key_s2[115], key_s1[115], key_s0[115]}), .b ({key_s2[51], key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_1563, new_AGEMA_signal_1562, wk[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U46 ( .a ({key_s2[114], key_s1[114], key_s0[114]}), .b ({key_s2[50], key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, wk[50]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U45 ( .a ({key_s2[4], key_s1[4], key_s0[4]}), .b ({key_s2[68], key_s1[68], key_s0[68]}), .c ({new_AGEMA_signal_1575, new_AGEMA_signal_1574, wk[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U44 ( .a ({key_s2[113], key_s1[113], key_s0[113]}), .b ({key_s2[49], key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, wk[49]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U43 ( .a ({key_s2[112], key_s1[112], key_s0[112]}), .b ({key_s2[48], key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, wk[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U42 ( .a ({key_s2[111], key_s1[111], key_s0[111]}), .b ({key_s2[47], key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_1593, new_AGEMA_signal_1592, wk[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U41 ( .a ({key_s2[110], key_s1[110], key_s0[110]}), .b ({key_s2[46], key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, wk[46]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U40 ( .a ({key_s2[109], key_s1[109], key_s0[109]}), .b ({key_s2[45], key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, wk[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U39 ( .a ({key_s2[108], key_s1[108], key_s0[108]}), .b ({key_s2[44], key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_1611, new_AGEMA_signal_1610, wk[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U38 ( .a ({key_s2[107], key_s1[107], key_s0[107]}), .b ({key_s2[43], key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, wk[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U37 ( .a ({key_s2[106], key_s1[106], key_s0[106]}), .b ({key_s2[42], key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_1623, new_AGEMA_signal_1622, wk[42]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U36 ( .a ({key_s2[105], key_s1[105], key_s0[105]}), .b ({key_s2[41], key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_1629, new_AGEMA_signal_1628, wk[41]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U35 ( .a ({key_s2[104], key_s1[104], key_s0[104]}), .b ({key_s2[40], key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, wk[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U34 ( .a ({key_s2[3], key_s1[3], key_s0[3]}), .b ({key_s2[67], key_s1[67], key_s0[67]}), .c ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, wk[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U33 ( .a ({key_s2[103], key_s1[103], key_s0[103]}), .b ({key_s2[39], key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_1647, new_AGEMA_signal_1646, wk[39]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U32 ( .a ({key_s2[102], key_s1[102], key_s0[102]}), .b ({key_s2[38], key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, wk[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U31 ( .a ({key_s2[101], key_s1[101], key_s0[101]}), .b ({key_s2[37], key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, wk[37]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U30 ( .a ({key_s2[100], key_s1[100], key_s0[100]}), .b ({key_s2[36], key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_1665, new_AGEMA_signal_1664, wk[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U29 ( .a ({key_s2[35], key_s1[35], key_s0[35]}), .b ({key_s2[99], key_s1[99], key_s0[99]}), .c ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, wk[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U28 ( .a ({key_s2[34], key_s1[34], key_s0[34]}), .b ({key_s2[98], key_s1[98], key_s0[98]}), .c ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, wk[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U27 ( .a ({key_s2[33], key_s1[33], key_s0[33]}), .b ({key_s2[97], key_s1[97], key_s0[97]}), .c ({new_AGEMA_signal_1683, new_AGEMA_signal_1682, wk[33]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U26 ( .a ({key_s2[32], key_s1[32], key_s0[32]}), .b ({key_s2[96], key_s1[96], key_s0[96]}), .c ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, wk[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U25 ( .a ({key_s2[31], key_s1[31], key_s0[31]}), .b ({key_s2[95], key_s1[95], key_s0[95]}), .c ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, wk[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U24 ( .a ({key_s2[30], key_s1[30], key_s0[30]}), .b ({key_s2[94], key_s1[94], key_s0[94]}), .c ({new_AGEMA_signal_1701, new_AGEMA_signal_1700, wk[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U23 ( .a ({key_s2[2], key_s1[2], key_s0[2]}), .b ({key_s2[66], key_s1[66], key_s0[66]}), .c ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, wk[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U22 ( .a ({key_s2[29], key_s1[29], key_s0[29]}), .b ({key_s2[93], key_s1[93], key_s0[93]}), .c ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, wk[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U21 ( .a ({key_s2[28], key_s1[28], key_s0[28]}), .b ({key_s2[92], key_s1[92], key_s0[92]}), .c ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, wk[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U20 ( .a ({key_s2[27], key_s1[27], key_s0[27]}), .b ({key_s2[91], key_s1[91], key_s0[91]}), .c ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, wk[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U19 ( .a ({key_s2[26], key_s1[26], key_s0[26]}), .b ({key_s2[90], key_s1[90], key_s0[90]}), .c ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, wk[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U18 ( .a ({key_s2[25], key_s1[25], key_s0[25]}), .b ({key_s2[89], key_s1[89], key_s0[89]}), .c ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, wk[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U17 ( .a ({key_s2[24], key_s1[24], key_s0[24]}), .b ({key_s2[88], key_s1[88], key_s0[88]}), .c ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, wk[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U16 ( .a ({key_s2[23], key_s1[23], key_s0[23]}), .b ({key_s2[87], key_s1[87], key_s0[87]}), .c ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, wk[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U15 ( .a ({key_s2[22], key_s1[22], key_s0[22]}), .b ({key_s2[86], key_s1[86], key_s0[86]}), .c ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, wk[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U14 ( .a ({key_s2[21], key_s1[21], key_s0[21]}), .b ({key_s2[85], key_s1[85], key_s0[85]}), .c ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, wk[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U13 ( .a ({key_s2[20], key_s1[20], key_s0[20]}), .b ({key_s2[84], key_s1[84], key_s0[84]}), .c ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, wk[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U12 ( .a ({key_s2[1], key_s1[1], key_s0[1]}), .b ({key_s2[65], key_s1[65], key_s0[65]}), .c ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, wk[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U11 ( .a ({key_s2[19], key_s1[19], key_s0[19]}), .b ({key_s2[83], key_s1[83], key_s0[83]}), .c ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, wk[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U10 ( .a ({key_s2[18], key_s1[18], key_s0[18]}), .b ({key_s2[82], key_s1[82], key_s0[82]}), .c ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, wk[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U9 ( .a ({key_s2[17], key_s1[17], key_s0[17]}), .b ({key_s2[81], key_s1[81], key_s0[81]}), .c ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, wk[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U8 ( .a ({key_s2[16], key_s1[16], key_s0[16]}), .b ({key_s2[80], key_s1[80], key_s0[80]}), .c ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, wk[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U7 ( .a ({key_s2[15], key_s1[15], key_s0[15]}), .b ({key_s2[79], key_s1[79], key_s0[79]}), .c ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, wk[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U6 ( .a ({key_s2[14], key_s1[14], key_s0[14]}), .b ({key_s2[78], key_s1[78], key_s0[78]}), .c ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, wk[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U5 ( .a ({key_s2[13], key_s1[13], key_s0[13]}), .b ({key_s2[77], key_s1[77], key_s0[77]}), .c ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, wk[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U4 ( .a ({key_s2[12], key_s1[12], key_s0[12]}), .b ({key_s2[76], key_s1[76], key_s0[76]}), .c ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, wk[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U3 ( .a ({key_s2[11], key_s1[11], key_s0[11]}), .b ({key_s2[75], key_s1[75], key_s0[75]}), .c ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, wk[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U2 ( .a ({key_s2[10], key_s1[10], key_s0[10]}), .b ({key_s2[74], key_s1[74], key_s0[74]}), .c ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, wk[10]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) keys_U1 ( .a ({key_s2[0], key_s1[0], key_s0[0]}), .b ({key_s2[64], key_s1[64], key_s0[64]}), .c ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, wk[0]}) ) ;
    NOR2_X1 controller_U3 ( .A1 (controller_n2), .A2 (controller_n1), .ZN (new_AGEMA_signal_4784) ) ;
    NAND2_X1 controller_U2 ( .A1 (round_Signal[0]), .A2 (round_Signal[1]), .ZN (controller_n1) ) ;
    NAND2_X1 controller_U1 ( .A1 (round_Signal[2]), .A2 (round_Signal[3]), .ZN (controller_n2) ) ;
    INV_X1 controller_roundCounter_U14 ( .A (controller_roundCounter_n13), .ZN (controller_roundCounter_n2) ) ;
    MUX2_X1 controller_roundCounter_U13 ( .S (controller_roundCounter_n6), .A (controller_roundCounter_n12), .B (controller_roundCounter_n11), .Z (controller_roundCounter_n13) ) ;
    NOR2_X1 controller_roundCounter_U12 ( .A1 (reset), .A2 (controller_roundCounter_n10), .ZN (controller_roundCounter_N8) ) ;
    XNOR2_X1 controller_roundCounter_U11 ( .A (round_Signal[0]), .B (round_Signal[1]), .ZN (controller_roundCounter_n10) ) ;
    MUX2_X1 controller_roundCounter_U10 ( .S (round_Signal[3]), .A (controller_roundCounter_n9), .B (controller_roundCounter_n8), .Z (controller_roundCounter_N10) ) ;
    NAND2_X1 controller_roundCounter_U9 ( .A1 (controller_roundCounter_n12), .A2 (controller_roundCounter_n7), .ZN (controller_roundCounter_n8) ) ;
    NAND2_X1 controller_roundCounter_U8 ( .A1 (controller_roundCounter_n6), .A2 (controller_roundCounter_n3), .ZN (controller_roundCounter_n7) ) ;
    NOR2_X1 controller_roundCounter_U7 ( .A1 (controller_roundCounter_n5), .A2 (controller_roundCounter_N7), .ZN (controller_roundCounter_n12) ) ;
    NOR2_X1 controller_roundCounter_U6 ( .A1 (round_Signal[1]), .A2 (reset), .ZN (controller_roundCounter_n5) ) ;
    NOR2_X1 controller_roundCounter_U5 ( .A1 (controller_roundCounter_n6), .A2 (controller_roundCounter_n11), .ZN (controller_roundCounter_n9) ) ;
    NAND2_X1 controller_roundCounter_U4 ( .A1 (round_Signal[1]), .A2 (controller_roundCounter_n4), .ZN (controller_roundCounter_n11) ) ;
    NOR2_X1 controller_roundCounter_U3 ( .A1 (reset), .A2 (controller_roundCounter_n1), .ZN (controller_roundCounter_n4) ) ;
    NOR2_X1 controller_roundCounter_U2 ( .A1 (reset), .A2 (round_Signal[0]), .ZN (controller_roundCounter_N7) ) ;
    INV_X1 controller_roundCounter_U1 ( .A (reset), .ZN (controller_roundCounter_n3) ) ;
    INV_X1 controller_roundCounter_count_reg_0__U1 ( .A (round_Signal[0]), .ZN (controller_roundCounter_n1) ) ;
    INV_X1 controller_roundCounter_count_reg_2__U1 ( .A (round_Signal[2]), .ZN (controller_roundCounter_n6) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U64 ( .a ({new_AGEMA_signal_1461, new_AGEMA_signal_1460, wk[9]}), .b ({DataIn_s2[9], DataIn_s1[9], DataIn_s0[9]}), .c ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, Midori_add_Result_Start[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U63 ( .a ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, wk[8]}), .b ({DataIn_s2[8], DataIn_s1[8], DataIn_s0[8]}), .c ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, Midori_add_Result_Start[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U62 ( .a ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, wk[7]}), .b ({DataIn_s2[7], DataIn_s1[7], DataIn_s0[7]}), .c ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, Midori_add_Result_Start[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U61 ( .a ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, wk[6]}), .b ({DataIn_s2[6], DataIn_s1[6], DataIn_s0[6]}), .c ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, Midori_add_Result_Start[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U60 ( .a ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, wk[63]}), .b ({DataIn_s2[63], DataIn_s1[63], DataIn_s0[63]}), .c ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, Midori_add_Result_Start[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U59 ( .a ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, wk[62]}), .b ({DataIn_s2[62], DataIn_s1[62], DataIn_s0[62]}), .c ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, Midori_add_Result_Start[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U58 ( .a ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, wk[61]}), .b ({DataIn_s2[61], DataIn_s1[61], DataIn_s0[61]}), .c ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, Midori_add_Result_Start[61]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U57 ( .a ({new_AGEMA_signal_1503, new_AGEMA_signal_1502, wk[60]}), .b ({DataIn_s2[60], DataIn_s1[60], DataIn_s0[60]}), .c ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, Midori_add_Result_Start[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U56 ( .a ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, wk[5]}), .b ({DataIn_s2[5], DataIn_s1[5], DataIn_s0[5]}), .c ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, Midori_add_Result_Start[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U55 ( .a ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, wk[59]}), .b ({DataIn_s2[59], DataIn_s1[59], DataIn_s0[59]}), .c ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, Midori_add_Result_Start[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U54 ( .a ({new_AGEMA_signal_1521, new_AGEMA_signal_1520, wk[58]}), .b ({DataIn_s2[58], DataIn_s1[58], DataIn_s0[58]}), .c ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, Midori_add_Result_Start[58]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U53 ( .a ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, wk[57]}), .b ({DataIn_s2[57], DataIn_s1[57], DataIn_s0[57]}), .c ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, Midori_add_Result_Start[57]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U52 ( .a ({new_AGEMA_signal_1533, new_AGEMA_signal_1532, wk[56]}), .b ({DataIn_s2[56], DataIn_s1[56], DataIn_s0[56]}), .c ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, Midori_add_Result_Start[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U51 ( .a ({new_AGEMA_signal_1539, new_AGEMA_signal_1538, wk[55]}), .b ({DataIn_s2[55], DataIn_s1[55], DataIn_s0[55]}), .c ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, Midori_add_Result_Start[55]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U50 ( .a ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, wk[54]}), .b ({DataIn_s2[54], DataIn_s1[54], DataIn_s0[54]}), .c ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, Midori_add_Result_Start[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U49 ( .a ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, wk[53]}), .b ({DataIn_s2[53], DataIn_s1[53], DataIn_s0[53]}), .c ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, Midori_add_Result_Start[53]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U48 ( .a ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, wk[52]}), .b ({DataIn_s2[52], DataIn_s1[52], DataIn_s0[52]}), .c ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, Midori_add_Result_Start[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U47 ( .a ({new_AGEMA_signal_1563, new_AGEMA_signal_1562, wk[51]}), .b ({DataIn_s2[51], DataIn_s1[51], DataIn_s0[51]}), .c ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, Midori_add_Result_Start[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U46 ( .a ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, wk[50]}), .b ({DataIn_s2[50], DataIn_s1[50], DataIn_s0[50]}), .c ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, Midori_add_Result_Start[50]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U45 ( .a ({new_AGEMA_signal_1575, new_AGEMA_signal_1574, wk[4]}), .b ({DataIn_s2[4], DataIn_s1[4], DataIn_s0[4]}), .c ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, Midori_add_Result_Start[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U44 ( .a ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, wk[49]}), .b ({DataIn_s2[49], DataIn_s1[49], DataIn_s0[49]}), .c ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, Midori_add_Result_Start[49]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U43 ( .a ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, wk[48]}), .b ({DataIn_s2[48], DataIn_s1[48], DataIn_s0[48]}), .c ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, Midori_add_Result_Start[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U42 ( .a ({new_AGEMA_signal_1593, new_AGEMA_signal_1592, wk[47]}), .b ({DataIn_s2[47], DataIn_s1[47], DataIn_s0[47]}), .c ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, Midori_add_Result_Start[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U41 ( .a ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, wk[46]}), .b ({DataIn_s2[46], DataIn_s1[46], DataIn_s0[46]}), .c ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, Midori_add_Result_Start[46]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U40 ( .a ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, wk[45]}), .b ({DataIn_s2[45], DataIn_s1[45], DataIn_s0[45]}), .c ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, Midori_add_Result_Start[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U39 ( .a ({new_AGEMA_signal_1611, new_AGEMA_signal_1610, wk[44]}), .b ({DataIn_s2[44], DataIn_s1[44], DataIn_s0[44]}), .c ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, Midori_add_Result_Start[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U38 ( .a ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, wk[43]}), .b ({DataIn_s2[43], DataIn_s1[43], DataIn_s0[43]}), .c ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, Midori_add_Result_Start[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U37 ( .a ({new_AGEMA_signal_1623, new_AGEMA_signal_1622, wk[42]}), .b ({DataIn_s2[42], DataIn_s1[42], DataIn_s0[42]}), .c ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, Midori_add_Result_Start[42]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U36 ( .a ({new_AGEMA_signal_1629, new_AGEMA_signal_1628, wk[41]}), .b ({DataIn_s2[41], DataIn_s1[41], DataIn_s0[41]}), .c ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, Midori_add_Result_Start[41]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U35 ( .a ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, wk[40]}), .b ({DataIn_s2[40], DataIn_s1[40], DataIn_s0[40]}), .c ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, Midori_add_Result_Start[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U34 ( .a ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, wk[3]}), .b ({DataIn_s2[3], DataIn_s1[3], DataIn_s0[3]}), .c ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, Midori_add_Result_Start[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U33 ( .a ({new_AGEMA_signal_1647, new_AGEMA_signal_1646, wk[39]}), .b ({DataIn_s2[39], DataIn_s1[39], DataIn_s0[39]}), .c ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, Midori_add_Result_Start[39]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U32 ( .a ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, wk[38]}), .b ({DataIn_s2[38], DataIn_s1[38], DataIn_s0[38]}), .c ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, Midori_add_Result_Start[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U31 ( .a ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, wk[37]}), .b ({DataIn_s2[37], DataIn_s1[37], DataIn_s0[37]}), .c ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, Midori_add_Result_Start[37]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U30 ( .a ({new_AGEMA_signal_1665, new_AGEMA_signal_1664, wk[36]}), .b ({DataIn_s2[36], DataIn_s1[36], DataIn_s0[36]}), .c ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, Midori_add_Result_Start[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U29 ( .a ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, wk[35]}), .b ({DataIn_s2[35], DataIn_s1[35], DataIn_s0[35]}), .c ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, Midori_add_Result_Start[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U28 ( .a ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, wk[34]}), .b ({DataIn_s2[34], DataIn_s1[34], DataIn_s0[34]}), .c ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, Midori_add_Result_Start[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U27 ( .a ({new_AGEMA_signal_1683, new_AGEMA_signal_1682, wk[33]}), .b ({DataIn_s2[33], DataIn_s1[33], DataIn_s0[33]}), .c ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, Midori_add_Result_Start[33]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U26 ( .a ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, wk[32]}), .b ({DataIn_s2[32], DataIn_s1[32], DataIn_s0[32]}), .c ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, Midori_add_Result_Start[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U25 ( .a ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, wk[31]}), .b ({DataIn_s2[31], DataIn_s1[31], DataIn_s0[31]}), .c ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, Midori_add_Result_Start[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U24 ( .a ({new_AGEMA_signal_1701, new_AGEMA_signal_1700, wk[30]}), .b ({DataIn_s2[30], DataIn_s1[30], DataIn_s0[30]}), .c ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, Midori_add_Result_Start[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U23 ( .a ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, wk[2]}), .b ({DataIn_s2[2], DataIn_s1[2], DataIn_s0[2]}), .c ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, Midori_add_Result_Start[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U22 ( .a ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, wk[29]}), .b ({DataIn_s2[29], DataIn_s1[29], DataIn_s0[29]}), .c ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, Midori_add_Result_Start[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U21 ( .a ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, wk[28]}), .b ({DataIn_s2[28], DataIn_s1[28], DataIn_s0[28]}), .c ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, Midori_add_Result_Start[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U20 ( .a ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, wk[27]}), .b ({DataIn_s2[27], DataIn_s1[27], DataIn_s0[27]}), .c ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, Midori_add_Result_Start[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U19 ( .a ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, wk[26]}), .b ({DataIn_s2[26], DataIn_s1[26], DataIn_s0[26]}), .c ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, Midori_add_Result_Start[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U18 ( .a ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, wk[25]}), .b ({DataIn_s2[25], DataIn_s1[25], DataIn_s0[25]}), .c ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, Midori_add_Result_Start[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U17 ( .a ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, wk[24]}), .b ({DataIn_s2[24], DataIn_s1[24], DataIn_s0[24]}), .c ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, Midori_add_Result_Start[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U16 ( .a ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, wk[23]}), .b ({DataIn_s2[23], DataIn_s1[23], DataIn_s0[23]}), .c ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, Midori_add_Result_Start[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U15 ( .a ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, wk[22]}), .b ({DataIn_s2[22], DataIn_s1[22], DataIn_s0[22]}), .c ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, Midori_add_Result_Start[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U14 ( .a ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, wk[21]}), .b ({DataIn_s2[21], DataIn_s1[21], DataIn_s0[21]}), .c ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, Midori_add_Result_Start[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U13 ( .a ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, wk[20]}), .b ({DataIn_s2[20], DataIn_s1[20], DataIn_s0[20]}), .c ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, Midori_add_Result_Start[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U12 ( .a ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, wk[1]}), .b ({DataIn_s2[1], DataIn_s1[1], DataIn_s0[1]}), .c ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, Midori_add_Result_Start[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U11 ( .a ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, wk[19]}), .b ({DataIn_s2[19], DataIn_s1[19], DataIn_s0[19]}), .c ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, Midori_add_Result_Start[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U10 ( .a ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, wk[18]}), .b ({DataIn_s2[18], DataIn_s1[18], DataIn_s0[18]}), .c ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, Midori_add_Result_Start[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U9 ( .a ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, wk[17]}), .b ({DataIn_s2[17], DataIn_s1[17], DataIn_s0[17]}), .c ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, Midori_add_Result_Start[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U8 ( .a ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, wk[16]}), .b ({DataIn_s2[16], DataIn_s1[16], DataIn_s0[16]}), .c ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, Midori_add_Result_Start[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U7 ( .a ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, wk[15]}), .b ({DataIn_s2[15], DataIn_s1[15], DataIn_s0[15]}), .c ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, Midori_add_Result_Start[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U6 ( .a ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, wk[14]}), .b ({DataIn_s2[14], DataIn_s1[14], DataIn_s0[14]}), .c ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, Midori_add_Result_Start[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U5 ( .a ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, wk[13]}), .b ({DataIn_s2[13], DataIn_s1[13], DataIn_s0[13]}), .c ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, Midori_add_Result_Start[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U4 ( .a ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, wk[12]}), .b ({DataIn_s2[12], DataIn_s1[12], DataIn_s0[12]}), .c ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, Midori_add_Result_Start[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U3 ( .a ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, wk[11]}), .b ({DataIn_s2[11], DataIn_s1[11], DataIn_s0[11]}), .c ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, Midori_add_Result_Start[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U2 ( .a ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, wk[10]}), .b ({DataIn_s2[10], DataIn_s1[10], DataIn_s0[10]}), .c ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, Midori_add_Result_Start[10]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U1 ( .a ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, wk[0]}), .b ({DataIn_s2[0], DataIn_s1[0], DataIn_s0[0]}), .c ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, Midori_add_Result_Start[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U78 ( .a ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, Midori_rounds_SelectedKey_8_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[2]}), .c ({new_AGEMA_signal_3427, new_AGEMA_signal_3426, Midori_rounds_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U71 ( .a ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, Midori_rounds_SelectedKey_60_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[15]}), .c ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, Midori_rounds_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U65 ( .a ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, Midori_rounds_SelectedKey_56_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[14]}), .c ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, Midori_rounds_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U60 ( .a ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, Midori_rounds_SelectedKey_52_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[13]}), .c ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, Midori_rounds_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U56 ( .a ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, Midori_rounds_SelectedKey_4_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[1]}), .c ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, Midori_rounds_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U53 ( .a ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, Midori_rounds_SelectedKey_48_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[12]}), .c ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, Midori_rounds_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U48 ( .a ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, Midori_rounds_SelectedKey_44_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[11]}), .c ({new_AGEMA_signal_3465, new_AGEMA_signal_3464, Midori_rounds_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U43 ( .a ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, Midori_rounds_SelectedKey_40_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[10]}), .c ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, Midori_rounds_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U37 ( .a ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, Midori_rounds_SelectedKey_36_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[9]}), .c ({new_AGEMA_signal_3481, new_AGEMA_signal_3480, Midori_rounds_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U32 ( .a ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, Midori_rounds_SelectedKey_32_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[8]}), .c ({new_AGEMA_signal_3547, new_AGEMA_signal_3546, Midori_rounds_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U26 ( .a ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, Midori_rounds_SelectedKey_28_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[7]}), .c ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, Midori_rounds_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U21 ( .a ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, Midori_rounds_SelectedKey_24_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[6]}), .c ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, Midori_rounds_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U16 ( .a ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, Midori_rounds_SelectedKey_20_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[5]}), .c ({new_AGEMA_signal_3509, new_AGEMA_signal_3508, Midori_rounds_n4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U10 ( .a ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, Midori_rounds_SelectedKey_16_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[4]}), .c ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, Midori_rounds_n3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U5 ( .a ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, Midori_rounds_SelectedKey_12_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[3]}), .c ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, Midori_rounds_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U1 ( .a ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, Midori_rounds_SelectedKey_0_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[0]}), .c ({new_AGEMA_signal_3555, new_AGEMA_signal_3554, Midori_rounds_n1}) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U106 ( .A1 (Midori_rounds_constant_MUX_n217), .A2 (Midori_rounds_constant_MUX_n216), .ZN (Midori_rounds_round_Constant[9]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U105 ( .A1 (Midori_rounds_constant_MUX_n215), .A2 (Midori_rounds_constant_MUX_n214), .ZN (Midori_rounds_constant_MUX_n217) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U104 ( .A1 (Midori_rounds_constant_MUX_n213), .A2 (Midori_rounds_constant_MUX_n212), .ZN (Midori_rounds_constant_MUX_n214) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U103 ( .A1 (Midori_rounds_constant_MUX_n211), .A2 (Midori_rounds_constant_MUX_n210), .ZN (Midori_rounds_round_Constant[8]) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U102 ( .A1 (Midori_rounds_constant_MUX_n209), .A2 (Midori_rounds_constant_MUX_n208), .ZN (Midori_rounds_round_Constant[7]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U101 ( .A1 (Midori_rounds_round_Constant[11]), .A2 (Midori_rounds_constant_MUX_n207), .ZN (Midori_rounds_constant_MUX_n208) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U100 ( .A1 (Midori_rounds_constant_MUX_n206), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n207) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U99 ( .A1 (Midori_rounds_constant_MUX_n204), .A2 (Midori_rounds_constant_MUX_n203), .ZN (Midori_rounds_constant_MUX_n206) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U98 ( .A1 (Midori_rounds_constant_MUX_n202), .A2 (Midori_rounds_constant_MUX_n201), .ZN (Midori_rounds_round_Constant[6]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U97 ( .A1 (Midori_rounds_constant_MUX_n200), .A2 (Midori_rounds_constant_MUX_n199), .ZN (Midori_rounds_constant_MUX_n201) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U96 ( .A1 (Midori_rounds_constant_MUX_n198), .A2 (Midori_rounds_constant_MUX_n197), .ZN (Midori_rounds_round_Constant[5]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U95 ( .A1 (Midori_rounds_constant_MUX_n212), .A2 (Midori_rounds_constant_MUX_n196), .ZN (Midori_rounds_constant_MUX_n197) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U94 ( .A1 (Midori_rounds_constant_MUX_n195), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n196) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U93 ( .A1 (Midori_rounds_constant_MUX_n194), .A2 (Midori_rounds_constant_MUX_n195), .ZN (Midori_rounds_round_Constant[4]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U92 ( .A1 (Midori_rounds_constant_MUX_n193), .A2 (Midori_rounds_constant_MUX_n192), .ZN (Midori_rounds_constant_MUX_n195) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U91 ( .A1 (Midori_rounds_constant_MUX_n191), .A2 (Midori_rounds_constant_MUX_n190), .ZN (Midori_rounds_round_Constant[3]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U90 ( .A1 (Midori_rounds_constant_MUX_n215), .A2 (Midori_rounds_constant_MUX_n189), .ZN (Midori_rounds_constant_MUX_n191) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U89 ( .A1 (Midori_rounds_constant_MUX_n188), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n189) ) ;
    INV_X1 Midori_rounds_constant_MUX_U88 ( .A (Midori_rounds_constant_MUX_n187), .ZN (Midori_rounds_constant_MUX_n188) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U87 ( .A1 (Midori_rounds_constant_MUX_n215), .A2 (Midori_rounds_constant_MUX_n186), .ZN (Midori_rounds_round_Constant[2]) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U86 ( .A1 (Midori_rounds_constant_MUX_n202), .A2 (Midori_rounds_constant_MUX_n185), .ZN (Midori_rounds_constant_MUX_n186) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U85 ( .A1 (Midori_rounds_constant_MUX_n184), .A2 (Midori_rounds_constant_MUX_n212), .ZN (Midori_rounds_constant_MUX_n202) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U84 ( .A1 (Midori_rounds_constant_MUX_n183), .A2 (Midori_rounds_constant_MUX_n210), .ZN (Midori_rounds_constant_MUX_n215) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U83 ( .A1 (Midori_rounds_constant_MUX_n182), .A2 (Midori_rounds_constant_MUX_n181), .ZN (Midori_rounds_round_Constant[1]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U82 ( .A1 (Midori_rounds_constant_MUX_n187), .A2 (Midori_rounds_constant_MUX_n180), .ZN (Midori_rounds_constant_MUX_n181) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U81 ( .A1 (Midori_rounds_constant_MUX_n212), .A2 (Midori_rounds_constant_MUX_n204), .ZN (Midori_rounds_constant_MUX_n180) ) ;
    INV_X1 Midori_rounds_constant_MUX_U80 ( .A (Midori_rounds_constant_MUX_n183), .ZN (Midori_rounds_constant_MUX_n204) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U79 ( .A1 (Midori_rounds_constant_MUX_n179), .A2 (Midori_rounds_constant_MUX_n178), .ZN (Midori_rounds_constant_MUX_n183) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U78 ( .A1 (Midori_rounds_constant_MUX_n177), .A2 (Midori_rounds_constant_MUX_n176), .ZN (Midori_rounds_constant_MUX_n178) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U77 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n175), .ZN (Midori_rounds_constant_MUX_n212) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U76 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n174), .B (Midori_rounds_constant_MUX_n173), .Z (Midori_rounds_constant_MUX_n175) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U75 ( .A1 (Midori_rounds_constant_MUX_n172), .A2 (Midori_rounds_constant_MUX_n171), .ZN (Midori_rounds_round_Constant[15]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U74 ( .A1 (Midori_rounds_constant_MUX_n200), .A2 (Midori_rounds_constant_MUX_n187), .ZN (Midori_rounds_constant_MUX_n172) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U73 ( .A1 (Midori_rounds_constant_MUX_n170), .A2 (Midori_rounds_constant_MUX_n194), .ZN (Midori_rounds_round_Constant[14]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U72 ( .A1 (Midori_rounds_constant_MUX_n169), .A2 (Midori_rounds_constant_MUX_n168), .ZN (Midori_rounds_constant_MUX_n194) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U71 ( .A1 (Midori_rounds_constant_MUX_n216), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n168) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U70 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n167), .ZN (Midori_rounds_constant_MUX_n205) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U69 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n166), .B (Midori_rounds_constant_MUX_n165), .Z (Midori_rounds_constant_MUX_n167) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U68 ( .A1 (Midori_rounds_constant_MUX_n185), .A2 (Midori_rounds_constant_MUX_n164), .ZN (Midori_rounds_round_Constant[13]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U67 ( .A1 (Midori_rounds_constant_MUX_n163), .A2 (Midori_rounds_constant_MUX_n162), .ZN (Midori_rounds_constant_MUX_n164) ) ;
    INV_X1 Midori_rounds_constant_MUX_U66 ( .A (Midori_rounds_constant_MUX_n170), .ZN (Midori_rounds_constant_MUX_n162) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U65 ( .A1 (Midori_rounds_constant_MUX_n161), .A2 (Midori_rounds_constant_MUX_n192), .ZN (Midori_rounds_constant_MUX_n185) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U64 ( .A1 (Midori_rounds_constant_MUX_n160), .A2 (Midori_rounds_constant_MUX_n190), .ZN (Midori_rounds_round_Constant[12]) ) ;
    INV_X1 Midori_rounds_constant_MUX_U63 ( .A (Midori_rounds_constant_MUX_n184), .ZN (Midori_rounds_constant_MUX_n190) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U62 ( .A1 (Midori_rounds_constant_MUX_n203), .A2 (Midori_rounds_constant_MUX_n159), .ZN (Midori_rounds_constant_MUX_n160) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U61 ( .A1 (Midori_rounds_constant_MUX_n211), .A2 (Midori_rounds_constant_MUX_n170), .ZN (Midori_rounds_constant_MUX_n159) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U60 ( .A1 (Midori_rounds_constant_MUX_n193), .A2 (Midori_rounds_constant_MUX_n169), .ZN (Midori_rounds_constant_MUX_n211) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U59 ( .A1 (Midori_rounds_constant_MUX_n198), .A2 (Midori_rounds_constant_MUX_n158), .ZN (Midori_rounds_constant_MUX_n169) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U58 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n157), .ZN (Midori_rounds_constant_MUX_n158) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U57 ( .A1 (Midori_rounds_constant_MUX_n165), .A2 (Midori_rounds_constant_MUX_n177), .ZN (Midori_rounds_constant_MUX_n157) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U56 ( .A1 (Midori_rounds_constant_MUX_n200), .A2 (Midori_rounds_constant_MUX_n156), .ZN (Midori_rounds_constant_MUX_n198) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U55 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n155), .ZN (Midori_rounds_constant_MUX_n156) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U54 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n176), .B (Midori_rounds_constant_MUX_n166), .Z (Midori_rounds_constant_MUX_n155) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U53 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n154), .ZN (Midori_rounds_constant_MUX_n200) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U52 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n174), .B (Midori_rounds_constant_MUX_n153), .Z (Midori_rounds_constant_MUX_n154) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U51 ( .A1 (Midori_rounds_constant_MUX_n199), .A2 (Midori_rounds_constant_MUX_n213), .ZN (Midori_rounds_round_Constant[11]) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U50 ( .A1 (Midori_rounds_constant_MUX_n170), .A2 (Midori_rounds_constant_MUX_n210), .ZN (Midori_rounds_constant_MUX_n199) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U49 ( .A1 (Midori_rounds_constant_MUX_n152), .A2 (Midori_rounds_constant_MUX_n151), .ZN (Midori_rounds_constant_MUX_n210) ) ;
    AND2_X1 Midori_rounds_constant_MUX_U48 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (round_Signal[2]), .ZN (Midori_rounds_constant_MUX_n151) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U47 ( .A1 (Midori_rounds_constant_MUX_n150), .A2 (Midori_rounds_constant_MUX_n187), .ZN (Midori_rounds_constant_MUX_n170) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U46 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n149), .ZN (Midori_rounds_constant_MUX_n187) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U45 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n165), .B (Midori_rounds_constant_MUX_n166), .Z (Midori_rounds_constant_MUX_n149) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U44 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n148), .ZN (Midori_rounds_constant_MUX_n150) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U43 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n153), .B (Midori_rounds_constant_MUX_n174), .Z (Midori_rounds_constant_MUX_n148) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U42 ( .A1 (Midori_rounds_constant_MUX_n147), .A2 (Midori_rounds_constant_MUX_n171), .ZN (Midori_rounds_round_Constant[10]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U41 ( .A1 (Midori_rounds_constant_MUX_n146), .A2 (Midori_rounds_constant_MUX_n213), .ZN (Midori_rounds_constant_MUX_n171) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U40 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n145), .ZN (Midori_rounds_constant_MUX_n213) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U39 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n165), .B (Midori_rounds_constant_MUX_n177), .Z (Midori_rounds_constant_MUX_n145) ) ;
    INV_X1 Midori_rounds_constant_MUX_U38 ( .A (Midori_rounds_constant_MUX_n144), .ZN (Midori_rounds_constant_MUX_n146) ) ;
    INV_X1 Midori_rounds_constant_MUX_U37 ( .A (Midori_rounds_constant_MUX_n193), .ZN (Midori_rounds_constant_MUX_n147) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U36 ( .A1 (Midori_rounds_constant_MUX_n182), .A2 (Midori_rounds_constant_MUX_n144), .ZN (Midori_rounds_round_Constant[0]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U35 ( .A1 (Midori_rounds_constant_MUX_n203), .A2 (Midori_rounds_constant_MUX_n192), .ZN (Midori_rounds_constant_MUX_n144) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U34 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n143), .ZN (Midori_rounds_constant_MUX_n192) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U33 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n173), .B (Midori_rounds_constant_MUX_n174), .Z (Midori_rounds_constant_MUX_n143) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U32 ( .A1 (Midori_rounds_constant_MUX_n142), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n174) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U31 ( .A1 (Midori_rounds_constant_MUX_n140), .A2 (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n173) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U30 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n139), .ZN (Midori_rounds_constant_MUX_n203) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U29 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n166), .B (Midori_rounds_constant_MUX_n176), .Z (Midori_rounds_constant_MUX_n139) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U28 ( .A1 (enc_dec), .A2 (Midori_rounds_constant_MUX_n152), .ZN (Midori_rounds_constant_MUX_n176) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U27 ( .A1 (round_Signal[3]), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n152) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U26 ( .A1 (Midori_rounds_constant_MUX_n138), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n166) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U25 ( .A1 (Midori_rounds_constant_MUX_n184), .A2 (Midori_rounds_constant_MUX_n137), .ZN (Midori_rounds_constant_MUX_n182) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U24 ( .A1 (Midori_rounds_constant_MUX_n209), .A2 (Midori_rounds_constant_MUX_n216), .ZN (Midori_rounds_constant_MUX_n137) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U23 ( .A1 (Midori_rounds_constant_MUX_n163), .A2 (Midori_rounds_constant_MUX_n136), .ZN (Midori_rounds_constant_MUX_n216) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U22 ( .A1 (Midori_rounds_constant_MUX_n140), .A2 (Midori_rounds_constant_MUX_n142), .ZN (Midori_rounds_constant_MUX_n136) ) ;
    AND2_X1 Midori_rounds_constant_MUX_U21 ( .A1 (round_Signal[1]), .A2 (Midori_rounds_constant_MUX_n179), .ZN (Midori_rounds_constant_MUX_n163) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U20 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (round_Signal[2]), .ZN (Midori_rounds_constant_MUX_n179) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U19 ( .A1 (Midori_rounds_constant_MUX_n193), .A2 (Midori_rounds_constant_MUX_n161), .ZN (Midori_rounds_constant_MUX_n209) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U18 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n135), .ZN (Midori_rounds_constant_MUX_n161) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U17 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n177), .B (Midori_rounds_constant_MUX_n165), .Z (Midori_rounds_constant_MUX_n135) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U16 ( .A1 (enc_dec), .A2 (Midori_rounds_constant_MUX_n134), .ZN (Midori_rounds_constant_MUX_n165) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U15 ( .A1 (round_Signal[3]), .A2 (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n134) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U14 ( .A1 (round_Signal[1]), .A2 (Midori_rounds_constant_MUX_n138), .ZN (Midori_rounds_constant_MUX_n177) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U13 ( .A1 (enc_dec), .A2 (Midori_rounds_constant_MUX_n133), .ZN (Midori_rounds_constant_MUX_n138) ) ;
    INV_X1 Midori_rounds_constant_MUX_U12 ( .A (round_Signal[3]), .ZN (Midori_rounds_constant_MUX_n133) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U11 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n132), .ZN (Midori_rounds_constant_MUX_n193) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U10 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n153), .B (Midori_rounds_constant_MUX_n131), .Z (Midori_rounds_constant_MUX_n132) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U9 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n130), .ZN (Midori_rounds_constant_MUX_n184) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U8 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n131), .B (Midori_rounds_constant_MUX_n153), .Z (Midori_rounds_constant_MUX_n130) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U7 ( .A1 (Midori_rounds_constant_MUX_n140), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n153) ) ;
    INV_X1 Midori_rounds_constant_MUX_U6 ( .A (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n141) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U5 ( .A1 (enc_dec), .A2 (round_Signal[3]), .ZN (Midori_rounds_constant_MUX_n140) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U4 ( .A1 (Midori_rounds_constant_MUX_n142), .A2 (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n131) ) ;
    AND2_X1 Midori_rounds_constant_MUX_U3 ( .A1 (enc_dec), .A2 (round_Signal[3]), .ZN (Midori_rounds_constant_MUX_n142) ) ;
    INV_X1 Midori_rounds_constant_MUX_U2 ( .A (Midori_rounds_constant_MUX_n129), .ZN (Midori_rounds_constant_MUX_n128) ) ;
    INV_X1 Midori_rounds_constant_MUX_U1 ( .A (round_Signal[0]), .ZN (Midori_rounds_constant_MUX_n129) ) ;
    INV_X1 Midori_rounds_MUXInst_U4 ( .A (round_Signal[0]), .ZN (Midori_rounds_MUXInst_n11) ) ;
    INV_X1 Midori_rounds_MUXInst_U3 ( .A (Midori_rounds_MUXInst_n11), .ZN (Midori_rounds_MUXInst_n8) ) ;
    INV_X1 Midori_rounds_MUXInst_U2 ( .A (Midori_rounds_MUXInst_n11), .ZN (Midori_rounds_MUXInst_n9) ) ;
    INV_X1 Midori_rounds_MUXInst_U1 ( .A (Midori_rounds_MUXInst_n11), .ZN (Midori_rounds_MUXInst_n10) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_0_U1 ( .s (round_Signal[0]), .b ({key_s2[64], key_s1[64], key_s0[64]}), .a ({key_s2[0], key_s1[0], key_s0[0]}), .c ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, Midori_rounds_SelectedKey_0_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_1_U1 ( .s (round_Signal[0]), .b ({key_s2[65], key_s1[65], key_s0[65]}), .a ({key_s2[1], key_s1[1], key_s0[1]}), .c ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, Midori_rounds_SelectedKey_1_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_2_U1 ( .s (round_Signal[0]), .b ({key_s2[66], key_s1[66], key_s0[66]}), .a ({key_s2[2], key_s1[2], key_s0[2]}), .c ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, Midori_rounds_SelectedKey_2_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_3_U1 ( .s (round_Signal[0]), .b ({key_s2[67], key_s1[67], key_s0[67]}), .a ({key_s2[3], key_s1[3], key_s0[3]}), .c ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, Midori_rounds_SelectedKey_3_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_4_U1 ( .s (round_Signal[0]), .b ({key_s2[68], key_s1[68], key_s0[68]}), .a ({key_s2[4], key_s1[4], key_s0[4]}), .c ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, Midori_rounds_SelectedKey_4_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_5_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[69], key_s1[69], key_s0[69]}), .a ({key_s2[5], key_s1[5], key_s0[5]}), .c ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, Midori_rounds_SelectedKey_5_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_6_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[70], key_s1[70], key_s0[70]}), .a ({key_s2[6], key_s1[6], key_s0[6]}), .c ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, Midori_rounds_SelectedKey_6_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_7_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[71], key_s1[71], key_s0[71]}), .a ({key_s2[7], key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, Midori_rounds_SelectedKey_7_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_8_U1 ( .s (round_Signal[0]), .b ({key_s2[72], key_s1[72], key_s0[72]}), .a ({key_s2[8], key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, Midori_rounds_SelectedKey_8_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_9_U1 ( .s (round_Signal[0]), .b ({key_s2[73], key_s1[73], key_s0[73]}), .a ({key_s2[9], key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, Midori_rounds_SelectedKey_9_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_10_U1 ( .s (round_Signal[0]), .b ({key_s2[74], key_s1[74], key_s0[74]}), .a ({key_s2[10], key_s1[10], key_s0[10]}), .c ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, Midori_rounds_SelectedKey_10_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_11_U1 ( .s (round_Signal[0]), .b ({key_s2[75], key_s1[75], key_s0[75]}), .a ({key_s2[11], key_s1[11], key_s0[11]}), .c ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, Midori_rounds_SelectedKey_11_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_12_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[76], key_s1[76], key_s0[76]}), .a ({key_s2[12], key_s1[12], key_s0[12]}), .c ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, Midori_rounds_SelectedKey_12_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_13_U1 ( .s (round_Signal[0]), .b ({key_s2[77], key_s1[77], key_s0[77]}), .a ({key_s2[13], key_s1[13], key_s0[13]}), .c ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, Midori_rounds_SelectedKey_13_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_14_U1 ( .s (round_Signal[0]), .b ({key_s2[78], key_s1[78], key_s0[78]}), .a ({key_s2[14], key_s1[14], key_s0[14]}), .c ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, Midori_rounds_SelectedKey_14_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_15_U1 ( .s (round_Signal[0]), .b ({key_s2[79], key_s1[79], key_s0[79]}), .a ({key_s2[15], key_s1[15], key_s0[15]}), .c ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, Midori_rounds_SelectedKey_15_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_16_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[80], key_s1[80], key_s0[80]}), .a ({key_s2[16], key_s1[16], key_s0[16]}), .c ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, Midori_rounds_SelectedKey_16_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_17_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[81], key_s1[81], key_s0[81]}), .a ({key_s2[17], key_s1[17], key_s0[17]}), .c ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, Midori_rounds_SelectedKey_17_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_18_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[82], key_s1[82], key_s0[82]}), .a ({key_s2[18], key_s1[18], key_s0[18]}), .c ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, Midori_rounds_SelectedKey_18_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_19_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[83], key_s1[83], key_s0[83]}), .a ({key_s2[19], key_s1[19], key_s0[19]}), .c ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, Midori_rounds_SelectedKey_19_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_20_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[84], key_s1[84], key_s0[84]}), .a ({key_s2[20], key_s1[20], key_s0[20]}), .c ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, Midori_rounds_SelectedKey_20_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_21_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[85], key_s1[85], key_s0[85]}), .a ({key_s2[21], key_s1[21], key_s0[21]}), .c ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, Midori_rounds_SelectedKey_21_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_22_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[86], key_s1[86], key_s0[86]}), .a ({key_s2[22], key_s1[22], key_s0[22]}), .c ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, Midori_rounds_SelectedKey_22_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_23_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[87], key_s1[87], key_s0[87]}), .a ({key_s2[23], key_s1[23], key_s0[23]}), .c ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, Midori_rounds_SelectedKey_23_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_24_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[88], key_s1[88], key_s0[88]}), .a ({key_s2[24], key_s1[24], key_s0[24]}), .c ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, Midori_rounds_SelectedKey_24_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_25_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[89], key_s1[89], key_s0[89]}), .a ({key_s2[25], key_s1[25], key_s0[25]}), .c ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, Midori_rounds_SelectedKey_25_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_26_U1 ( .s (round_Signal[0]), .b ({key_s2[90], key_s1[90], key_s0[90]}), .a ({key_s2[26], key_s1[26], key_s0[26]}), .c ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, Midori_rounds_SelectedKey_26_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_27_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[91], key_s1[91], key_s0[91]}), .a ({key_s2[27], key_s1[27], key_s0[27]}), .c ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, Midori_rounds_SelectedKey_27_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_28_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[92], key_s1[92], key_s0[92]}), .a ({key_s2[28], key_s1[28], key_s0[28]}), .c ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, Midori_rounds_SelectedKey_28_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_29_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[93], key_s1[93], key_s0[93]}), .a ({key_s2[29], key_s1[29], key_s0[29]}), .c ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, Midori_rounds_SelectedKey_29_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_30_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[94], key_s1[94], key_s0[94]}), .a ({key_s2[30], key_s1[30], key_s0[30]}), .c ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, Midori_rounds_SelectedKey_30_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_31_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[95], key_s1[95], key_s0[95]}), .a ({key_s2[31], key_s1[31], key_s0[31]}), .c ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, Midori_rounds_SelectedKey_31_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_32_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[96], key_s1[96], key_s0[96]}), .a ({key_s2[32], key_s1[32], key_s0[32]}), .c ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, Midori_rounds_SelectedKey_32_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_33_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[97], key_s1[97], key_s0[97]}), .a ({key_s2[33], key_s1[33], key_s0[33]}), .c ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, Midori_rounds_SelectedKey_33_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_34_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[98], key_s1[98], key_s0[98]}), .a ({key_s2[34], key_s1[34], key_s0[34]}), .c ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, Midori_rounds_SelectedKey_34_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_35_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[99], key_s1[99], key_s0[99]}), .a ({key_s2[35], key_s1[35], key_s0[35]}), .c ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, Midori_rounds_SelectedKey_35_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_36_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[100], key_s1[100], key_s0[100]}), .a ({key_s2[36], key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, Midori_rounds_SelectedKey_36_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_37_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[101], key_s1[101], key_s0[101]}), .a ({key_s2[37], key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, Midori_rounds_SelectedKey_37_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_38_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[102], key_s1[102], key_s0[102]}), .a ({key_s2[38], key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, Midori_rounds_SelectedKey_38_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_39_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[103], key_s1[103], key_s0[103]}), .a ({key_s2[39], key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, Midori_rounds_SelectedKey_39_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_40_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[104], key_s1[104], key_s0[104]}), .a ({key_s2[40], key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, Midori_rounds_SelectedKey_40_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_41_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[105], key_s1[105], key_s0[105]}), .a ({key_s2[41], key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, Midori_rounds_SelectedKey_41_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_42_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[106], key_s1[106], key_s0[106]}), .a ({key_s2[42], key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, Midori_rounds_SelectedKey_42_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_43_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[107], key_s1[107], key_s0[107]}), .a ({key_s2[43], key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, Midori_rounds_SelectedKey_43_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_44_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[108], key_s1[108], key_s0[108]}), .a ({key_s2[44], key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, Midori_rounds_SelectedKey_44_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_45_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[109], key_s1[109], key_s0[109]}), .a ({key_s2[45], key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, Midori_rounds_SelectedKey_45_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_46_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[110], key_s1[110], key_s0[110]}), .a ({key_s2[46], key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, Midori_rounds_SelectedKey_46_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_47_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[111], key_s1[111], key_s0[111]}), .a ({key_s2[47], key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, Midori_rounds_SelectedKey_47_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_48_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[112], key_s1[112], key_s0[112]}), .a ({key_s2[48], key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, Midori_rounds_SelectedKey_48_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_49_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[113], key_s1[113], key_s0[113]}), .a ({key_s2[49], key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, Midori_rounds_SelectedKey_49_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_50_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[114], key_s1[114], key_s0[114]}), .a ({key_s2[50], key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, Midori_rounds_SelectedKey_50_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_51_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[115], key_s1[115], key_s0[115]}), .a ({key_s2[51], key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, Midori_rounds_SelectedKey_51_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_52_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[116], key_s1[116], key_s0[116]}), .a ({key_s2[52], key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, Midori_rounds_SelectedKey_52_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_53_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[117], key_s1[117], key_s0[117]}), .a ({key_s2[53], key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, Midori_rounds_SelectedKey_53_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_54_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[118], key_s1[118], key_s0[118]}), .a ({key_s2[54], key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, Midori_rounds_SelectedKey_54_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_55_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[119], key_s1[119], key_s0[119]}), .a ({key_s2[55], key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, Midori_rounds_SelectedKey_55_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_56_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[120], key_s1[120], key_s0[120]}), .a ({key_s2[56], key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, Midori_rounds_SelectedKey_56_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_57_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[121], key_s1[121], key_s0[121]}), .a ({key_s2[57], key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, Midori_rounds_SelectedKey_57_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_58_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[122], key_s1[122], key_s0[122]}), .a ({key_s2[58], key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, Midori_rounds_SelectedKey_58_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_59_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[123], key_s1[123], key_s0[123]}), .a ({key_s2[59], key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, Midori_rounds_SelectedKey_59_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_60_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[124], key_s1[124], key_s0[124]}), .a ({key_s2[60], key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, Midori_rounds_SelectedKey_60_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_61_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[125], key_s1[125], key_s0[125]}), .a ({key_s2[61], key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, Midori_rounds_SelectedKey_61_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_62_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[126], key_s1[126], key_s0[126]}), .a ({key_s2[62], key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, Midori_rounds_SelectedKey_62_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_63_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[127], key_s1[127], key_s0[127]}), .a ({key_s2[63], key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, Midori_rounds_SelectedKey_63_}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U4 ( .a ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, Midori_rounds_roundReg_out[0]}), .b ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, Midori_rounds_sub_sBox_PRINCE_0_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U2 ( .a ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, Midori_rounds_roundReg_out[3]}), .b ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, Midori_rounds_sub_sBox_PRINCE_0_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U1 ( .a ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, Midori_rounds_roundReg_out[2]}), .b ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, Midori_rounds_sub_sBox_PRINCE_0_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U4 ( .a ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, Midori_rounds_roundReg_out[4]}), .b ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, Midori_rounds_sub_sBox_PRINCE_1_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U2 ( .a ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, Midori_rounds_roundReg_out[7]}), .b ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, Midori_rounds_sub_sBox_PRINCE_1_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U1 ( .a ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, Midori_rounds_roundReg_out[6]}), .b ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, Midori_rounds_sub_sBox_PRINCE_1_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U4 ( .a ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, Midori_rounds_roundReg_out[8]}), .b ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, Midori_rounds_sub_sBox_PRINCE_2_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U2 ( .a ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, Midori_rounds_roundReg_out[11]}), .b ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, Midori_rounds_sub_sBox_PRINCE_2_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U1 ( .a ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, Midori_rounds_roundReg_out[10]}), .b ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, Midori_rounds_sub_sBox_PRINCE_2_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U4 ( .a ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, Midori_rounds_roundReg_out[12]}), .b ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, Midori_rounds_sub_sBox_PRINCE_3_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U2 ( .a ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, Midori_rounds_roundReg_out[15]}), .b ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, Midori_rounds_sub_sBox_PRINCE_3_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U1 ( .a ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, Midori_rounds_roundReg_out[14]}), .b ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, Midori_rounds_sub_sBox_PRINCE_3_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U4 ( .a ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, Midori_rounds_roundReg_out[16]}), .b ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, Midori_rounds_sub_sBox_PRINCE_4_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U2 ( .a ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, Midori_rounds_roundReg_out[19]}), .b ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, Midori_rounds_sub_sBox_PRINCE_4_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U1 ( .a ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, Midori_rounds_roundReg_out[18]}), .b ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, Midori_rounds_sub_sBox_PRINCE_4_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U4 ( .a ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, Midori_rounds_roundReg_out[20]}), .b ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, Midori_rounds_sub_sBox_PRINCE_5_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U2 ( .a ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, Midori_rounds_roundReg_out[23]}), .b ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, Midori_rounds_sub_sBox_PRINCE_5_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U1 ( .a ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, Midori_rounds_roundReg_out[22]}), .b ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, Midori_rounds_sub_sBox_PRINCE_5_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U4 ( .a ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, Midori_rounds_roundReg_out[24]}), .b ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, Midori_rounds_sub_sBox_PRINCE_6_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U2 ( .a ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, Midori_rounds_roundReg_out[27]}), .b ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, Midori_rounds_sub_sBox_PRINCE_6_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U1 ( .a ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, Midori_rounds_roundReg_out[26]}), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, Midori_rounds_sub_sBox_PRINCE_6_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U4 ( .a ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, Midori_rounds_roundReg_out[28]}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, Midori_rounds_sub_sBox_PRINCE_7_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U2 ( .a ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, Midori_rounds_roundReg_out[31]}), .b ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, Midori_rounds_sub_sBox_PRINCE_7_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U1 ( .a ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, Midori_rounds_roundReg_out[30]}), .b ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, Midori_rounds_sub_sBox_PRINCE_7_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U4 ( .a ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, Midori_rounds_roundReg_out[32]}), .b ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, Midori_rounds_sub_sBox_PRINCE_8_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U2 ( .a ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, Midori_rounds_roundReg_out[35]}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, Midori_rounds_sub_sBox_PRINCE_8_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U1 ( .a ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, Midori_rounds_roundReg_out[34]}), .b ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, Midori_rounds_sub_sBox_PRINCE_8_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U4 ( .a ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, Midori_rounds_roundReg_out[36]}), .b ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, Midori_rounds_sub_sBox_PRINCE_9_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U2 ( .a ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, Midori_rounds_roundReg_out[39]}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, Midori_rounds_sub_sBox_PRINCE_9_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U1 ( .a ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, Midori_rounds_roundReg_out[38]}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, Midori_rounds_sub_sBox_PRINCE_9_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U4 ( .a ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, Midori_rounds_roundReg_out[40]}), .b ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, Midori_rounds_sub_sBox_PRINCE_10_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U2 ( .a ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, Midori_rounds_roundReg_out[43]}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, Midori_rounds_sub_sBox_PRINCE_10_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U1 ( .a ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, Midori_rounds_roundReg_out[42]}), .b ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, Midori_rounds_sub_sBox_PRINCE_10_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U4 ( .a ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, Midori_rounds_roundReg_out[44]}), .b ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, Midori_rounds_sub_sBox_PRINCE_11_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U2 ( .a ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, Midori_rounds_roundReg_out[47]}), .b ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, Midori_rounds_sub_sBox_PRINCE_11_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U1 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, Midori_rounds_roundReg_out[46]}), .b ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, Midori_rounds_sub_sBox_PRINCE_11_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U4 ( .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, Midori_rounds_roundReg_out[48]}), .b ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, Midori_rounds_sub_sBox_PRINCE_12_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U2 ( .a ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, Midori_rounds_roundReg_out[51]}), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, Midori_rounds_sub_sBox_PRINCE_12_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U1 ( .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, Midori_rounds_roundReg_out[50]}), .b ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, Midori_rounds_sub_sBox_PRINCE_12_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U4 ( .a ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, Midori_rounds_roundReg_out[52]}), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, Midori_rounds_sub_sBox_PRINCE_13_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U2 ( .a ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, Midori_rounds_roundReg_out[55]}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, Midori_rounds_sub_sBox_PRINCE_13_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U1 ( .a ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, Midori_rounds_roundReg_out[54]}), .b ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, Midori_rounds_sub_sBox_PRINCE_13_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U4 ( .a ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, Midori_rounds_roundReg_out[56]}), .b ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, Midori_rounds_sub_sBox_PRINCE_14_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U2 ( .a ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, Midori_rounds_roundReg_out[59]}), .b ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, Midori_rounds_sub_sBox_PRINCE_14_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U1 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, Midori_rounds_roundReg_out[58]}), .b ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, Midori_rounds_sub_sBox_PRINCE_14_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U4 ( .a ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, Midori_rounds_roundReg_out[60]}), .b ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, Midori_rounds_sub_sBox_PRINCE_15_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U2 ( .a ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, Midori_rounds_roundReg_out[63]}), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, Midori_rounds_sub_sBox_PRINCE_15_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U1 ( .a ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, Midori_rounds_roundReg_out[62]}), .b ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, Midori_rounds_sub_sBox_PRINCE_15_n9}) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_1319 ( .C (clk), .D (new_AGEMA_signal_4784), .Q (new_AGEMA_signal_4785) ) ;
    buf_clk new_AGEMA_reg_buffer_1455 ( .C (clk), .D (Midori_rounds_roundReg_out[1]), .Q (new_AGEMA_signal_4920) ) ;
    buf_clk new_AGEMA_reg_buffer_1457 ( .C (clk), .D (new_AGEMA_signal_2672), .Q (new_AGEMA_signal_4922) ) ;
    buf_clk new_AGEMA_reg_buffer_1459 ( .C (clk), .D (new_AGEMA_signal_2673), .Q (new_AGEMA_signal_4924) ) ;
    buf_clk new_AGEMA_reg_buffer_1461 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_0_n9), .Q (new_AGEMA_signal_4926) ) ;
    buf_clk new_AGEMA_reg_buffer_1463 ( .C (clk), .D (new_AGEMA_signal_1880), .Q (new_AGEMA_signal_4928) ) ;
    buf_clk new_AGEMA_reg_buffer_1465 ( .C (clk), .D (new_AGEMA_signal_1881), .Q (new_AGEMA_signal_4930) ) ;
    buf_clk new_AGEMA_reg_buffer_1467 ( .C (clk), .D (Midori_rounds_roundReg_out[0]), .Q (new_AGEMA_signal_4932) ) ;
    buf_clk new_AGEMA_reg_buffer_1469 ( .C (clk), .D (new_AGEMA_signal_1866), .Q (new_AGEMA_signal_4934) ) ;
    buf_clk new_AGEMA_reg_buffer_1471 ( .C (clk), .D (new_AGEMA_signal_1867), .Q (new_AGEMA_signal_4936) ) ;
    buf_clk new_AGEMA_reg_buffer_1473 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_0_n7), .Q (new_AGEMA_signal_4938) ) ;
    buf_clk new_AGEMA_reg_buffer_1475 ( .C (clk), .D (new_AGEMA_signal_1876), .Q (new_AGEMA_signal_4940) ) ;
    buf_clk new_AGEMA_reg_buffer_1477 ( .C (clk), .D (new_AGEMA_signal_1877), .Q (new_AGEMA_signal_4942) ) ;
    buf_clk new_AGEMA_reg_buffer_1479 ( .C (clk), .D (Midori_rounds_roundReg_out[5]), .Q (new_AGEMA_signal_4944) ) ;
    buf_clk new_AGEMA_reg_buffer_1481 ( .C (clk), .D (new_AGEMA_signal_2682), .Q (new_AGEMA_signal_4946) ) ;
    buf_clk new_AGEMA_reg_buffer_1483 ( .C (clk), .D (new_AGEMA_signal_2683), .Q (new_AGEMA_signal_4948) ) ;
    buf_clk new_AGEMA_reg_buffer_1485 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_1_n9), .Q (new_AGEMA_signal_4950) ) ;
    buf_clk new_AGEMA_reg_buffer_1487 ( .C (clk), .D (new_AGEMA_signal_1896), .Q (new_AGEMA_signal_4952) ) ;
    buf_clk new_AGEMA_reg_buffer_1489 ( .C (clk), .D (new_AGEMA_signal_1897), .Q (new_AGEMA_signal_4954) ) ;
    buf_clk new_AGEMA_reg_buffer_1491 ( .C (clk), .D (Midori_rounds_roundReg_out[4]), .Q (new_AGEMA_signal_4956) ) ;
    buf_clk new_AGEMA_reg_buffer_1493 ( .C (clk), .D (new_AGEMA_signal_1882), .Q (new_AGEMA_signal_4958) ) ;
    buf_clk new_AGEMA_reg_buffer_1495 ( .C (clk), .D (new_AGEMA_signal_1883), .Q (new_AGEMA_signal_4960) ) ;
    buf_clk new_AGEMA_reg_buffer_1497 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_1_n7), .Q (new_AGEMA_signal_4962) ) ;
    buf_clk new_AGEMA_reg_buffer_1499 ( .C (clk), .D (new_AGEMA_signal_1892), .Q (new_AGEMA_signal_4964) ) ;
    buf_clk new_AGEMA_reg_buffer_1501 ( .C (clk), .D (new_AGEMA_signal_1893), .Q (new_AGEMA_signal_4966) ) ;
    buf_clk new_AGEMA_reg_buffer_1503 ( .C (clk), .D (Midori_rounds_roundReg_out[9]), .Q (new_AGEMA_signal_4968) ) ;
    buf_clk new_AGEMA_reg_buffer_1505 ( .C (clk), .D (new_AGEMA_signal_2692), .Q (new_AGEMA_signal_4970) ) ;
    buf_clk new_AGEMA_reg_buffer_1507 ( .C (clk), .D (new_AGEMA_signal_2693), .Q (new_AGEMA_signal_4972) ) ;
    buf_clk new_AGEMA_reg_buffer_1509 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_2_n9), .Q (new_AGEMA_signal_4974) ) ;
    buf_clk new_AGEMA_reg_buffer_1511 ( .C (clk), .D (new_AGEMA_signal_1912), .Q (new_AGEMA_signal_4976) ) ;
    buf_clk new_AGEMA_reg_buffer_1513 ( .C (clk), .D (new_AGEMA_signal_1913), .Q (new_AGEMA_signal_4978) ) ;
    buf_clk new_AGEMA_reg_buffer_1515 ( .C (clk), .D (Midori_rounds_roundReg_out[8]), .Q (new_AGEMA_signal_4980) ) ;
    buf_clk new_AGEMA_reg_buffer_1517 ( .C (clk), .D (new_AGEMA_signal_1898), .Q (new_AGEMA_signal_4982) ) ;
    buf_clk new_AGEMA_reg_buffer_1519 ( .C (clk), .D (new_AGEMA_signal_1899), .Q (new_AGEMA_signal_4984) ) ;
    buf_clk new_AGEMA_reg_buffer_1521 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_2_n7), .Q (new_AGEMA_signal_4986) ) ;
    buf_clk new_AGEMA_reg_buffer_1523 ( .C (clk), .D (new_AGEMA_signal_1908), .Q (new_AGEMA_signal_4988) ) ;
    buf_clk new_AGEMA_reg_buffer_1525 ( .C (clk), .D (new_AGEMA_signal_1909), .Q (new_AGEMA_signal_4990) ) ;
    buf_clk new_AGEMA_reg_buffer_1527 ( .C (clk), .D (Midori_rounds_roundReg_out[13]), .Q (new_AGEMA_signal_4992) ) ;
    buf_clk new_AGEMA_reg_buffer_1529 ( .C (clk), .D (new_AGEMA_signal_2702), .Q (new_AGEMA_signal_4994) ) ;
    buf_clk new_AGEMA_reg_buffer_1531 ( .C (clk), .D (new_AGEMA_signal_2703), .Q (new_AGEMA_signal_4996) ) ;
    buf_clk new_AGEMA_reg_buffer_1533 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_3_n9), .Q (new_AGEMA_signal_4998) ) ;
    buf_clk new_AGEMA_reg_buffer_1535 ( .C (clk), .D (new_AGEMA_signal_1928), .Q (new_AGEMA_signal_5000) ) ;
    buf_clk new_AGEMA_reg_buffer_1537 ( .C (clk), .D (new_AGEMA_signal_1929), .Q (new_AGEMA_signal_5002) ) ;
    buf_clk new_AGEMA_reg_buffer_1539 ( .C (clk), .D (Midori_rounds_roundReg_out[12]), .Q (new_AGEMA_signal_5004) ) ;
    buf_clk new_AGEMA_reg_buffer_1541 ( .C (clk), .D (new_AGEMA_signal_1914), .Q (new_AGEMA_signal_5006) ) ;
    buf_clk new_AGEMA_reg_buffer_1543 ( .C (clk), .D (new_AGEMA_signal_1915), .Q (new_AGEMA_signal_5008) ) ;
    buf_clk new_AGEMA_reg_buffer_1545 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_3_n7), .Q (new_AGEMA_signal_5010) ) ;
    buf_clk new_AGEMA_reg_buffer_1547 ( .C (clk), .D (new_AGEMA_signal_1924), .Q (new_AGEMA_signal_5012) ) ;
    buf_clk new_AGEMA_reg_buffer_1549 ( .C (clk), .D (new_AGEMA_signal_1925), .Q (new_AGEMA_signal_5014) ) ;
    buf_clk new_AGEMA_reg_buffer_1551 ( .C (clk), .D (Midori_rounds_roundReg_out[17]), .Q (new_AGEMA_signal_5016) ) ;
    buf_clk new_AGEMA_reg_buffer_1553 ( .C (clk), .D (new_AGEMA_signal_2712), .Q (new_AGEMA_signal_5018) ) ;
    buf_clk new_AGEMA_reg_buffer_1555 ( .C (clk), .D (new_AGEMA_signal_2713), .Q (new_AGEMA_signal_5020) ) ;
    buf_clk new_AGEMA_reg_buffer_1557 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_4_n9), .Q (new_AGEMA_signal_5022) ) ;
    buf_clk new_AGEMA_reg_buffer_1559 ( .C (clk), .D (new_AGEMA_signal_1944), .Q (new_AGEMA_signal_5024) ) ;
    buf_clk new_AGEMA_reg_buffer_1561 ( .C (clk), .D (new_AGEMA_signal_1945), .Q (new_AGEMA_signal_5026) ) ;
    buf_clk new_AGEMA_reg_buffer_1563 ( .C (clk), .D (Midori_rounds_roundReg_out[16]), .Q (new_AGEMA_signal_5028) ) ;
    buf_clk new_AGEMA_reg_buffer_1565 ( .C (clk), .D (new_AGEMA_signal_1930), .Q (new_AGEMA_signal_5030) ) ;
    buf_clk new_AGEMA_reg_buffer_1567 ( .C (clk), .D (new_AGEMA_signal_1931), .Q (new_AGEMA_signal_5032) ) ;
    buf_clk new_AGEMA_reg_buffer_1569 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_4_n7), .Q (new_AGEMA_signal_5034) ) ;
    buf_clk new_AGEMA_reg_buffer_1571 ( .C (clk), .D (new_AGEMA_signal_1940), .Q (new_AGEMA_signal_5036) ) ;
    buf_clk new_AGEMA_reg_buffer_1573 ( .C (clk), .D (new_AGEMA_signal_1941), .Q (new_AGEMA_signal_5038) ) ;
    buf_clk new_AGEMA_reg_buffer_1575 ( .C (clk), .D (Midori_rounds_roundReg_out[21]), .Q (new_AGEMA_signal_5040) ) ;
    buf_clk new_AGEMA_reg_buffer_1577 ( .C (clk), .D (new_AGEMA_signal_2722), .Q (new_AGEMA_signal_5042) ) ;
    buf_clk new_AGEMA_reg_buffer_1579 ( .C (clk), .D (new_AGEMA_signal_2723), .Q (new_AGEMA_signal_5044) ) ;
    buf_clk new_AGEMA_reg_buffer_1581 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_5_n9), .Q (new_AGEMA_signal_5046) ) ;
    buf_clk new_AGEMA_reg_buffer_1583 ( .C (clk), .D (new_AGEMA_signal_1960), .Q (new_AGEMA_signal_5048) ) ;
    buf_clk new_AGEMA_reg_buffer_1585 ( .C (clk), .D (new_AGEMA_signal_1961), .Q (new_AGEMA_signal_5050) ) ;
    buf_clk new_AGEMA_reg_buffer_1587 ( .C (clk), .D (Midori_rounds_roundReg_out[20]), .Q (new_AGEMA_signal_5052) ) ;
    buf_clk new_AGEMA_reg_buffer_1589 ( .C (clk), .D (new_AGEMA_signal_1946), .Q (new_AGEMA_signal_5054) ) ;
    buf_clk new_AGEMA_reg_buffer_1591 ( .C (clk), .D (new_AGEMA_signal_1947), .Q (new_AGEMA_signal_5056) ) ;
    buf_clk new_AGEMA_reg_buffer_1593 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_5_n7), .Q (new_AGEMA_signal_5058) ) ;
    buf_clk new_AGEMA_reg_buffer_1595 ( .C (clk), .D (new_AGEMA_signal_1956), .Q (new_AGEMA_signal_5060) ) ;
    buf_clk new_AGEMA_reg_buffer_1597 ( .C (clk), .D (new_AGEMA_signal_1957), .Q (new_AGEMA_signal_5062) ) ;
    buf_clk new_AGEMA_reg_buffer_1599 ( .C (clk), .D (Midori_rounds_roundReg_out[25]), .Q (new_AGEMA_signal_5064) ) ;
    buf_clk new_AGEMA_reg_buffer_1601 ( .C (clk), .D (new_AGEMA_signal_2732), .Q (new_AGEMA_signal_5066) ) ;
    buf_clk new_AGEMA_reg_buffer_1603 ( .C (clk), .D (new_AGEMA_signal_2733), .Q (new_AGEMA_signal_5068) ) ;
    buf_clk new_AGEMA_reg_buffer_1605 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_6_n9), .Q (new_AGEMA_signal_5070) ) ;
    buf_clk new_AGEMA_reg_buffer_1607 ( .C (clk), .D (new_AGEMA_signal_1976), .Q (new_AGEMA_signal_5072) ) ;
    buf_clk new_AGEMA_reg_buffer_1609 ( .C (clk), .D (new_AGEMA_signal_1977), .Q (new_AGEMA_signal_5074) ) ;
    buf_clk new_AGEMA_reg_buffer_1611 ( .C (clk), .D (Midori_rounds_roundReg_out[24]), .Q (new_AGEMA_signal_5076) ) ;
    buf_clk new_AGEMA_reg_buffer_1613 ( .C (clk), .D (new_AGEMA_signal_1962), .Q (new_AGEMA_signal_5078) ) ;
    buf_clk new_AGEMA_reg_buffer_1615 ( .C (clk), .D (new_AGEMA_signal_1963), .Q (new_AGEMA_signal_5080) ) ;
    buf_clk new_AGEMA_reg_buffer_1617 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_6_n7), .Q (new_AGEMA_signal_5082) ) ;
    buf_clk new_AGEMA_reg_buffer_1619 ( .C (clk), .D (new_AGEMA_signal_1972), .Q (new_AGEMA_signal_5084) ) ;
    buf_clk new_AGEMA_reg_buffer_1621 ( .C (clk), .D (new_AGEMA_signal_1973), .Q (new_AGEMA_signal_5086) ) ;
    buf_clk new_AGEMA_reg_buffer_1623 ( .C (clk), .D (Midori_rounds_roundReg_out[29]), .Q (new_AGEMA_signal_5088) ) ;
    buf_clk new_AGEMA_reg_buffer_1625 ( .C (clk), .D (new_AGEMA_signal_2742), .Q (new_AGEMA_signal_5090) ) ;
    buf_clk new_AGEMA_reg_buffer_1627 ( .C (clk), .D (new_AGEMA_signal_2743), .Q (new_AGEMA_signal_5092) ) ;
    buf_clk new_AGEMA_reg_buffer_1629 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_7_n9), .Q (new_AGEMA_signal_5094) ) ;
    buf_clk new_AGEMA_reg_buffer_1631 ( .C (clk), .D (new_AGEMA_signal_1992), .Q (new_AGEMA_signal_5096) ) ;
    buf_clk new_AGEMA_reg_buffer_1633 ( .C (clk), .D (new_AGEMA_signal_1993), .Q (new_AGEMA_signal_5098) ) ;
    buf_clk new_AGEMA_reg_buffer_1635 ( .C (clk), .D (Midori_rounds_roundReg_out[28]), .Q (new_AGEMA_signal_5100) ) ;
    buf_clk new_AGEMA_reg_buffer_1637 ( .C (clk), .D (new_AGEMA_signal_1978), .Q (new_AGEMA_signal_5102) ) ;
    buf_clk new_AGEMA_reg_buffer_1639 ( .C (clk), .D (new_AGEMA_signal_1979), .Q (new_AGEMA_signal_5104) ) ;
    buf_clk new_AGEMA_reg_buffer_1641 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_7_n7), .Q (new_AGEMA_signal_5106) ) ;
    buf_clk new_AGEMA_reg_buffer_1643 ( .C (clk), .D (new_AGEMA_signal_1988), .Q (new_AGEMA_signal_5108) ) ;
    buf_clk new_AGEMA_reg_buffer_1645 ( .C (clk), .D (new_AGEMA_signal_1989), .Q (new_AGEMA_signal_5110) ) ;
    buf_clk new_AGEMA_reg_buffer_1647 ( .C (clk), .D (Midori_rounds_roundReg_out[33]), .Q (new_AGEMA_signal_5112) ) ;
    buf_clk new_AGEMA_reg_buffer_1649 ( .C (clk), .D (new_AGEMA_signal_2752), .Q (new_AGEMA_signal_5114) ) ;
    buf_clk new_AGEMA_reg_buffer_1651 ( .C (clk), .D (new_AGEMA_signal_2753), .Q (new_AGEMA_signal_5116) ) ;
    buf_clk new_AGEMA_reg_buffer_1653 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_8_n9), .Q (new_AGEMA_signal_5118) ) ;
    buf_clk new_AGEMA_reg_buffer_1655 ( .C (clk), .D (new_AGEMA_signal_2008), .Q (new_AGEMA_signal_5120) ) ;
    buf_clk new_AGEMA_reg_buffer_1657 ( .C (clk), .D (new_AGEMA_signal_2009), .Q (new_AGEMA_signal_5122) ) ;
    buf_clk new_AGEMA_reg_buffer_1659 ( .C (clk), .D (Midori_rounds_roundReg_out[32]), .Q (new_AGEMA_signal_5124) ) ;
    buf_clk new_AGEMA_reg_buffer_1661 ( .C (clk), .D (new_AGEMA_signal_1994), .Q (new_AGEMA_signal_5126) ) ;
    buf_clk new_AGEMA_reg_buffer_1663 ( .C (clk), .D (new_AGEMA_signal_1995), .Q (new_AGEMA_signal_5128) ) ;
    buf_clk new_AGEMA_reg_buffer_1665 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_8_n7), .Q (new_AGEMA_signal_5130) ) ;
    buf_clk new_AGEMA_reg_buffer_1667 ( .C (clk), .D (new_AGEMA_signal_2004), .Q (new_AGEMA_signal_5132) ) ;
    buf_clk new_AGEMA_reg_buffer_1669 ( .C (clk), .D (new_AGEMA_signal_2005), .Q (new_AGEMA_signal_5134) ) ;
    buf_clk new_AGEMA_reg_buffer_1671 ( .C (clk), .D (Midori_rounds_roundReg_out[37]), .Q (new_AGEMA_signal_5136) ) ;
    buf_clk new_AGEMA_reg_buffer_1673 ( .C (clk), .D (new_AGEMA_signal_2762), .Q (new_AGEMA_signal_5138) ) ;
    buf_clk new_AGEMA_reg_buffer_1675 ( .C (clk), .D (new_AGEMA_signal_2763), .Q (new_AGEMA_signal_5140) ) ;
    buf_clk new_AGEMA_reg_buffer_1677 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_9_n9), .Q (new_AGEMA_signal_5142) ) ;
    buf_clk new_AGEMA_reg_buffer_1679 ( .C (clk), .D (new_AGEMA_signal_2024), .Q (new_AGEMA_signal_5144) ) ;
    buf_clk new_AGEMA_reg_buffer_1681 ( .C (clk), .D (new_AGEMA_signal_2025), .Q (new_AGEMA_signal_5146) ) ;
    buf_clk new_AGEMA_reg_buffer_1683 ( .C (clk), .D (Midori_rounds_roundReg_out[36]), .Q (new_AGEMA_signal_5148) ) ;
    buf_clk new_AGEMA_reg_buffer_1685 ( .C (clk), .D (new_AGEMA_signal_2010), .Q (new_AGEMA_signal_5150) ) ;
    buf_clk new_AGEMA_reg_buffer_1687 ( .C (clk), .D (new_AGEMA_signal_2011), .Q (new_AGEMA_signal_5152) ) ;
    buf_clk new_AGEMA_reg_buffer_1689 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_9_n7), .Q (new_AGEMA_signal_5154) ) ;
    buf_clk new_AGEMA_reg_buffer_1691 ( .C (clk), .D (new_AGEMA_signal_2020), .Q (new_AGEMA_signal_5156) ) ;
    buf_clk new_AGEMA_reg_buffer_1693 ( .C (clk), .D (new_AGEMA_signal_2021), .Q (new_AGEMA_signal_5158) ) ;
    buf_clk new_AGEMA_reg_buffer_1695 ( .C (clk), .D (Midori_rounds_roundReg_out[41]), .Q (new_AGEMA_signal_5160) ) ;
    buf_clk new_AGEMA_reg_buffer_1697 ( .C (clk), .D (new_AGEMA_signal_2772), .Q (new_AGEMA_signal_5162) ) ;
    buf_clk new_AGEMA_reg_buffer_1699 ( .C (clk), .D (new_AGEMA_signal_2773), .Q (new_AGEMA_signal_5164) ) ;
    buf_clk new_AGEMA_reg_buffer_1701 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_10_n9), .Q (new_AGEMA_signal_5166) ) ;
    buf_clk new_AGEMA_reg_buffer_1703 ( .C (clk), .D (new_AGEMA_signal_2040), .Q (new_AGEMA_signal_5168) ) ;
    buf_clk new_AGEMA_reg_buffer_1705 ( .C (clk), .D (new_AGEMA_signal_2041), .Q (new_AGEMA_signal_5170) ) ;
    buf_clk new_AGEMA_reg_buffer_1707 ( .C (clk), .D (Midori_rounds_roundReg_out[40]), .Q (new_AGEMA_signal_5172) ) ;
    buf_clk new_AGEMA_reg_buffer_1709 ( .C (clk), .D (new_AGEMA_signal_2026), .Q (new_AGEMA_signal_5174) ) ;
    buf_clk new_AGEMA_reg_buffer_1711 ( .C (clk), .D (new_AGEMA_signal_2027), .Q (new_AGEMA_signal_5176) ) ;
    buf_clk new_AGEMA_reg_buffer_1713 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_10_n7), .Q (new_AGEMA_signal_5178) ) ;
    buf_clk new_AGEMA_reg_buffer_1715 ( .C (clk), .D (new_AGEMA_signal_2036), .Q (new_AGEMA_signal_5180) ) ;
    buf_clk new_AGEMA_reg_buffer_1717 ( .C (clk), .D (new_AGEMA_signal_2037), .Q (new_AGEMA_signal_5182) ) ;
    buf_clk new_AGEMA_reg_buffer_1719 ( .C (clk), .D (Midori_rounds_roundReg_out[45]), .Q (new_AGEMA_signal_5184) ) ;
    buf_clk new_AGEMA_reg_buffer_1721 ( .C (clk), .D (new_AGEMA_signal_2782), .Q (new_AGEMA_signal_5186) ) ;
    buf_clk new_AGEMA_reg_buffer_1723 ( .C (clk), .D (new_AGEMA_signal_2783), .Q (new_AGEMA_signal_5188) ) ;
    buf_clk new_AGEMA_reg_buffer_1725 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_11_n9), .Q (new_AGEMA_signal_5190) ) ;
    buf_clk new_AGEMA_reg_buffer_1727 ( .C (clk), .D (new_AGEMA_signal_2056), .Q (new_AGEMA_signal_5192) ) ;
    buf_clk new_AGEMA_reg_buffer_1729 ( .C (clk), .D (new_AGEMA_signal_2057), .Q (new_AGEMA_signal_5194) ) ;
    buf_clk new_AGEMA_reg_buffer_1731 ( .C (clk), .D (Midori_rounds_roundReg_out[44]), .Q (new_AGEMA_signal_5196) ) ;
    buf_clk new_AGEMA_reg_buffer_1733 ( .C (clk), .D (new_AGEMA_signal_2042), .Q (new_AGEMA_signal_5198) ) ;
    buf_clk new_AGEMA_reg_buffer_1735 ( .C (clk), .D (new_AGEMA_signal_2043), .Q (new_AGEMA_signal_5200) ) ;
    buf_clk new_AGEMA_reg_buffer_1737 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_11_n7), .Q (new_AGEMA_signal_5202) ) ;
    buf_clk new_AGEMA_reg_buffer_1739 ( .C (clk), .D (new_AGEMA_signal_2052), .Q (new_AGEMA_signal_5204) ) ;
    buf_clk new_AGEMA_reg_buffer_1741 ( .C (clk), .D (new_AGEMA_signal_2053), .Q (new_AGEMA_signal_5206) ) ;
    buf_clk new_AGEMA_reg_buffer_1743 ( .C (clk), .D (Midori_rounds_roundReg_out[49]), .Q (new_AGEMA_signal_5208) ) ;
    buf_clk new_AGEMA_reg_buffer_1745 ( .C (clk), .D (new_AGEMA_signal_2792), .Q (new_AGEMA_signal_5210) ) ;
    buf_clk new_AGEMA_reg_buffer_1747 ( .C (clk), .D (new_AGEMA_signal_2793), .Q (new_AGEMA_signal_5212) ) ;
    buf_clk new_AGEMA_reg_buffer_1749 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_12_n9), .Q (new_AGEMA_signal_5214) ) ;
    buf_clk new_AGEMA_reg_buffer_1751 ( .C (clk), .D (new_AGEMA_signal_2072), .Q (new_AGEMA_signal_5216) ) ;
    buf_clk new_AGEMA_reg_buffer_1753 ( .C (clk), .D (new_AGEMA_signal_2073), .Q (new_AGEMA_signal_5218) ) ;
    buf_clk new_AGEMA_reg_buffer_1755 ( .C (clk), .D (Midori_rounds_roundReg_out[48]), .Q (new_AGEMA_signal_5220) ) ;
    buf_clk new_AGEMA_reg_buffer_1757 ( .C (clk), .D (new_AGEMA_signal_2058), .Q (new_AGEMA_signal_5222) ) ;
    buf_clk new_AGEMA_reg_buffer_1759 ( .C (clk), .D (new_AGEMA_signal_2059), .Q (new_AGEMA_signal_5224) ) ;
    buf_clk new_AGEMA_reg_buffer_1761 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_12_n7), .Q (new_AGEMA_signal_5226) ) ;
    buf_clk new_AGEMA_reg_buffer_1763 ( .C (clk), .D (new_AGEMA_signal_2068), .Q (new_AGEMA_signal_5228) ) ;
    buf_clk new_AGEMA_reg_buffer_1765 ( .C (clk), .D (new_AGEMA_signal_2069), .Q (new_AGEMA_signal_5230) ) ;
    buf_clk new_AGEMA_reg_buffer_1767 ( .C (clk), .D (Midori_rounds_roundReg_out[53]), .Q (new_AGEMA_signal_5232) ) ;
    buf_clk new_AGEMA_reg_buffer_1769 ( .C (clk), .D (new_AGEMA_signal_2802), .Q (new_AGEMA_signal_5234) ) ;
    buf_clk new_AGEMA_reg_buffer_1771 ( .C (clk), .D (new_AGEMA_signal_2803), .Q (new_AGEMA_signal_5236) ) ;
    buf_clk new_AGEMA_reg_buffer_1773 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_13_n9), .Q (new_AGEMA_signal_5238) ) ;
    buf_clk new_AGEMA_reg_buffer_1775 ( .C (clk), .D (new_AGEMA_signal_2088), .Q (new_AGEMA_signal_5240) ) ;
    buf_clk new_AGEMA_reg_buffer_1777 ( .C (clk), .D (new_AGEMA_signal_2089), .Q (new_AGEMA_signal_5242) ) ;
    buf_clk new_AGEMA_reg_buffer_1779 ( .C (clk), .D (Midori_rounds_roundReg_out[52]), .Q (new_AGEMA_signal_5244) ) ;
    buf_clk new_AGEMA_reg_buffer_1781 ( .C (clk), .D (new_AGEMA_signal_2074), .Q (new_AGEMA_signal_5246) ) ;
    buf_clk new_AGEMA_reg_buffer_1783 ( .C (clk), .D (new_AGEMA_signal_2075), .Q (new_AGEMA_signal_5248) ) ;
    buf_clk new_AGEMA_reg_buffer_1785 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_13_n7), .Q (new_AGEMA_signal_5250) ) ;
    buf_clk new_AGEMA_reg_buffer_1787 ( .C (clk), .D (new_AGEMA_signal_2084), .Q (new_AGEMA_signal_5252) ) ;
    buf_clk new_AGEMA_reg_buffer_1789 ( .C (clk), .D (new_AGEMA_signal_2085), .Q (new_AGEMA_signal_5254) ) ;
    buf_clk new_AGEMA_reg_buffer_1791 ( .C (clk), .D (Midori_rounds_roundReg_out[57]), .Q (new_AGEMA_signal_5256) ) ;
    buf_clk new_AGEMA_reg_buffer_1793 ( .C (clk), .D (new_AGEMA_signal_2812), .Q (new_AGEMA_signal_5258) ) ;
    buf_clk new_AGEMA_reg_buffer_1795 ( .C (clk), .D (new_AGEMA_signal_2813), .Q (new_AGEMA_signal_5260) ) ;
    buf_clk new_AGEMA_reg_buffer_1797 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_14_n9), .Q (new_AGEMA_signal_5262) ) ;
    buf_clk new_AGEMA_reg_buffer_1799 ( .C (clk), .D (new_AGEMA_signal_2104), .Q (new_AGEMA_signal_5264) ) ;
    buf_clk new_AGEMA_reg_buffer_1801 ( .C (clk), .D (new_AGEMA_signal_2105), .Q (new_AGEMA_signal_5266) ) ;
    buf_clk new_AGEMA_reg_buffer_1803 ( .C (clk), .D (Midori_rounds_roundReg_out[56]), .Q (new_AGEMA_signal_5268) ) ;
    buf_clk new_AGEMA_reg_buffer_1805 ( .C (clk), .D (new_AGEMA_signal_2090), .Q (new_AGEMA_signal_5270) ) ;
    buf_clk new_AGEMA_reg_buffer_1807 ( .C (clk), .D (new_AGEMA_signal_2091), .Q (new_AGEMA_signal_5272) ) ;
    buf_clk new_AGEMA_reg_buffer_1809 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_14_n7), .Q (new_AGEMA_signal_5274) ) ;
    buf_clk new_AGEMA_reg_buffer_1811 ( .C (clk), .D (new_AGEMA_signal_2100), .Q (new_AGEMA_signal_5276) ) ;
    buf_clk new_AGEMA_reg_buffer_1813 ( .C (clk), .D (new_AGEMA_signal_2101), .Q (new_AGEMA_signal_5278) ) ;
    buf_clk new_AGEMA_reg_buffer_1815 ( .C (clk), .D (Midori_rounds_roundReg_out[61]), .Q (new_AGEMA_signal_5280) ) ;
    buf_clk new_AGEMA_reg_buffer_1817 ( .C (clk), .D (new_AGEMA_signal_2822), .Q (new_AGEMA_signal_5282) ) ;
    buf_clk new_AGEMA_reg_buffer_1819 ( .C (clk), .D (new_AGEMA_signal_2823), .Q (new_AGEMA_signal_5284) ) ;
    buf_clk new_AGEMA_reg_buffer_1821 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_15_n9), .Q (new_AGEMA_signal_5286) ) ;
    buf_clk new_AGEMA_reg_buffer_1823 ( .C (clk), .D (new_AGEMA_signal_2120), .Q (new_AGEMA_signal_5288) ) ;
    buf_clk new_AGEMA_reg_buffer_1825 ( .C (clk), .D (new_AGEMA_signal_2121), .Q (new_AGEMA_signal_5290) ) ;
    buf_clk new_AGEMA_reg_buffer_1827 ( .C (clk), .D (Midori_rounds_roundReg_out[60]), .Q (new_AGEMA_signal_5292) ) ;
    buf_clk new_AGEMA_reg_buffer_1829 ( .C (clk), .D (new_AGEMA_signal_2106), .Q (new_AGEMA_signal_5294) ) ;
    buf_clk new_AGEMA_reg_buffer_1831 ( .C (clk), .D (new_AGEMA_signal_2107), .Q (new_AGEMA_signal_5296) ) ;
    buf_clk new_AGEMA_reg_buffer_1833 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_15_n7), .Q (new_AGEMA_signal_5298) ) ;
    buf_clk new_AGEMA_reg_buffer_1835 ( .C (clk), .D (new_AGEMA_signal_2116), .Q (new_AGEMA_signal_5300) ) ;
    buf_clk new_AGEMA_reg_buffer_1837 ( .C (clk), .D (new_AGEMA_signal_2117), .Q (new_AGEMA_signal_5302) ) ;
    buf_clk new_AGEMA_reg_buffer_1839 ( .C (clk), .D (wk[9]), .Q (new_AGEMA_signal_5304) ) ;
    buf_clk new_AGEMA_reg_buffer_1845 ( .C (clk), .D (new_AGEMA_signal_1460), .Q (new_AGEMA_signal_5310) ) ;
    buf_clk new_AGEMA_reg_buffer_1851 ( .C (clk), .D (new_AGEMA_signal_1461), .Q (new_AGEMA_signal_5316) ) ;
    buf_clk new_AGEMA_reg_buffer_1857 ( .C (clk), .D (wk[7]), .Q (new_AGEMA_signal_5322) ) ;
    buf_clk new_AGEMA_reg_buffer_1863 ( .C (clk), .D (new_AGEMA_signal_1472), .Q (new_AGEMA_signal_5328) ) ;
    buf_clk new_AGEMA_reg_buffer_1869 ( .C (clk), .D (new_AGEMA_signal_1473), .Q (new_AGEMA_signal_5334) ) ;
    buf_clk new_AGEMA_reg_buffer_1875 ( .C (clk), .D (wk[63]), .Q (new_AGEMA_signal_5340) ) ;
    buf_clk new_AGEMA_reg_buffer_1881 ( .C (clk), .D (new_AGEMA_signal_1484), .Q (new_AGEMA_signal_5346) ) ;
    buf_clk new_AGEMA_reg_buffer_1887 ( .C (clk), .D (new_AGEMA_signal_1485), .Q (new_AGEMA_signal_5352) ) ;
    buf_clk new_AGEMA_reg_buffer_1893 ( .C (clk), .D (wk[61]), .Q (new_AGEMA_signal_5358) ) ;
    buf_clk new_AGEMA_reg_buffer_1899 ( .C (clk), .D (new_AGEMA_signal_1496), .Q (new_AGEMA_signal_5364) ) ;
    buf_clk new_AGEMA_reg_buffer_1905 ( .C (clk), .D (new_AGEMA_signal_1497), .Q (new_AGEMA_signal_5370) ) ;
    buf_clk new_AGEMA_reg_buffer_1911 ( .C (clk), .D (wk[5]), .Q (new_AGEMA_signal_5376) ) ;
    buf_clk new_AGEMA_reg_buffer_1917 ( .C (clk), .D (new_AGEMA_signal_1508), .Q (new_AGEMA_signal_5382) ) ;
    buf_clk new_AGEMA_reg_buffer_1923 ( .C (clk), .D (new_AGEMA_signal_1509), .Q (new_AGEMA_signal_5388) ) ;
    buf_clk new_AGEMA_reg_buffer_1929 ( .C (clk), .D (wk[59]), .Q (new_AGEMA_signal_5394) ) ;
    buf_clk new_AGEMA_reg_buffer_1935 ( .C (clk), .D (new_AGEMA_signal_1514), .Q (new_AGEMA_signal_5400) ) ;
    buf_clk new_AGEMA_reg_buffer_1941 ( .C (clk), .D (new_AGEMA_signal_1515), .Q (new_AGEMA_signal_5406) ) ;
    buf_clk new_AGEMA_reg_buffer_1947 ( .C (clk), .D (wk[57]), .Q (new_AGEMA_signal_5412) ) ;
    buf_clk new_AGEMA_reg_buffer_1953 ( .C (clk), .D (new_AGEMA_signal_1526), .Q (new_AGEMA_signal_5418) ) ;
    buf_clk new_AGEMA_reg_buffer_1959 ( .C (clk), .D (new_AGEMA_signal_1527), .Q (new_AGEMA_signal_5424) ) ;
    buf_clk new_AGEMA_reg_buffer_1965 ( .C (clk), .D (wk[55]), .Q (new_AGEMA_signal_5430) ) ;
    buf_clk new_AGEMA_reg_buffer_1971 ( .C (clk), .D (new_AGEMA_signal_1538), .Q (new_AGEMA_signal_5436) ) ;
    buf_clk new_AGEMA_reg_buffer_1977 ( .C (clk), .D (new_AGEMA_signal_1539), .Q (new_AGEMA_signal_5442) ) ;
    buf_clk new_AGEMA_reg_buffer_1983 ( .C (clk), .D (wk[53]), .Q (new_AGEMA_signal_5448) ) ;
    buf_clk new_AGEMA_reg_buffer_1989 ( .C (clk), .D (new_AGEMA_signal_1550), .Q (new_AGEMA_signal_5454) ) ;
    buf_clk new_AGEMA_reg_buffer_1995 ( .C (clk), .D (new_AGEMA_signal_1551), .Q (new_AGEMA_signal_5460) ) ;
    buf_clk new_AGEMA_reg_buffer_2001 ( .C (clk), .D (wk[51]), .Q (new_AGEMA_signal_5466) ) ;
    buf_clk new_AGEMA_reg_buffer_2007 ( .C (clk), .D (new_AGEMA_signal_1562), .Q (new_AGEMA_signal_5472) ) ;
    buf_clk new_AGEMA_reg_buffer_2013 ( .C (clk), .D (new_AGEMA_signal_1563), .Q (new_AGEMA_signal_5478) ) ;
    buf_clk new_AGEMA_reg_buffer_2019 ( .C (clk), .D (wk[49]), .Q (new_AGEMA_signal_5484) ) ;
    buf_clk new_AGEMA_reg_buffer_2025 ( .C (clk), .D (new_AGEMA_signal_1580), .Q (new_AGEMA_signal_5490) ) ;
    buf_clk new_AGEMA_reg_buffer_2031 ( .C (clk), .D (new_AGEMA_signal_1581), .Q (new_AGEMA_signal_5496) ) ;
    buf_clk new_AGEMA_reg_buffer_2037 ( .C (clk), .D (wk[47]), .Q (new_AGEMA_signal_5502) ) ;
    buf_clk new_AGEMA_reg_buffer_2043 ( .C (clk), .D (new_AGEMA_signal_1592), .Q (new_AGEMA_signal_5508) ) ;
    buf_clk new_AGEMA_reg_buffer_2049 ( .C (clk), .D (new_AGEMA_signal_1593), .Q (new_AGEMA_signal_5514) ) ;
    buf_clk new_AGEMA_reg_buffer_2055 ( .C (clk), .D (wk[45]), .Q (new_AGEMA_signal_5520) ) ;
    buf_clk new_AGEMA_reg_buffer_2061 ( .C (clk), .D (new_AGEMA_signal_1604), .Q (new_AGEMA_signal_5526) ) ;
    buf_clk new_AGEMA_reg_buffer_2067 ( .C (clk), .D (new_AGEMA_signal_1605), .Q (new_AGEMA_signal_5532) ) ;
    buf_clk new_AGEMA_reg_buffer_2073 ( .C (clk), .D (wk[43]), .Q (new_AGEMA_signal_5538) ) ;
    buf_clk new_AGEMA_reg_buffer_2079 ( .C (clk), .D (new_AGEMA_signal_1616), .Q (new_AGEMA_signal_5544) ) ;
    buf_clk new_AGEMA_reg_buffer_2085 ( .C (clk), .D (new_AGEMA_signal_1617), .Q (new_AGEMA_signal_5550) ) ;
    buf_clk new_AGEMA_reg_buffer_2091 ( .C (clk), .D (wk[41]), .Q (new_AGEMA_signal_5556) ) ;
    buf_clk new_AGEMA_reg_buffer_2097 ( .C (clk), .D (new_AGEMA_signal_1628), .Q (new_AGEMA_signal_5562) ) ;
    buf_clk new_AGEMA_reg_buffer_2103 ( .C (clk), .D (new_AGEMA_signal_1629), .Q (new_AGEMA_signal_5568) ) ;
    buf_clk new_AGEMA_reg_buffer_2109 ( .C (clk), .D (wk[3]), .Q (new_AGEMA_signal_5574) ) ;
    buf_clk new_AGEMA_reg_buffer_2115 ( .C (clk), .D (new_AGEMA_signal_1640), .Q (new_AGEMA_signal_5580) ) ;
    buf_clk new_AGEMA_reg_buffer_2121 ( .C (clk), .D (new_AGEMA_signal_1641), .Q (new_AGEMA_signal_5586) ) ;
    buf_clk new_AGEMA_reg_buffer_2127 ( .C (clk), .D (wk[39]), .Q (new_AGEMA_signal_5592) ) ;
    buf_clk new_AGEMA_reg_buffer_2133 ( .C (clk), .D (new_AGEMA_signal_1646), .Q (new_AGEMA_signal_5598) ) ;
    buf_clk new_AGEMA_reg_buffer_2139 ( .C (clk), .D (new_AGEMA_signal_1647), .Q (new_AGEMA_signal_5604) ) ;
    buf_clk new_AGEMA_reg_buffer_2145 ( .C (clk), .D (wk[37]), .Q (new_AGEMA_signal_5610) ) ;
    buf_clk new_AGEMA_reg_buffer_2151 ( .C (clk), .D (new_AGEMA_signal_1658), .Q (new_AGEMA_signal_5616) ) ;
    buf_clk new_AGEMA_reg_buffer_2157 ( .C (clk), .D (new_AGEMA_signal_1659), .Q (new_AGEMA_signal_5622) ) ;
    buf_clk new_AGEMA_reg_buffer_2163 ( .C (clk), .D (wk[35]), .Q (new_AGEMA_signal_5628) ) ;
    buf_clk new_AGEMA_reg_buffer_2169 ( .C (clk), .D (new_AGEMA_signal_1670), .Q (new_AGEMA_signal_5634) ) ;
    buf_clk new_AGEMA_reg_buffer_2175 ( .C (clk), .D (new_AGEMA_signal_1671), .Q (new_AGEMA_signal_5640) ) ;
    buf_clk new_AGEMA_reg_buffer_2181 ( .C (clk), .D (wk[33]), .Q (new_AGEMA_signal_5646) ) ;
    buf_clk new_AGEMA_reg_buffer_2187 ( .C (clk), .D (new_AGEMA_signal_1682), .Q (new_AGEMA_signal_5652) ) ;
    buf_clk new_AGEMA_reg_buffer_2193 ( .C (clk), .D (new_AGEMA_signal_1683), .Q (new_AGEMA_signal_5658) ) ;
    buf_clk new_AGEMA_reg_buffer_2199 ( .C (clk), .D (wk[31]), .Q (new_AGEMA_signal_5664) ) ;
    buf_clk new_AGEMA_reg_buffer_2205 ( .C (clk), .D (new_AGEMA_signal_1694), .Q (new_AGEMA_signal_5670) ) ;
    buf_clk new_AGEMA_reg_buffer_2211 ( .C (clk), .D (new_AGEMA_signal_1695), .Q (new_AGEMA_signal_5676) ) ;
    buf_clk new_AGEMA_reg_buffer_2217 ( .C (clk), .D (wk[29]), .Q (new_AGEMA_signal_5682) ) ;
    buf_clk new_AGEMA_reg_buffer_2223 ( .C (clk), .D (new_AGEMA_signal_1712), .Q (new_AGEMA_signal_5688) ) ;
    buf_clk new_AGEMA_reg_buffer_2229 ( .C (clk), .D (new_AGEMA_signal_1713), .Q (new_AGEMA_signal_5694) ) ;
    buf_clk new_AGEMA_reg_buffer_2235 ( .C (clk), .D (wk[27]), .Q (new_AGEMA_signal_5700) ) ;
    buf_clk new_AGEMA_reg_buffer_2241 ( .C (clk), .D (new_AGEMA_signal_1724), .Q (new_AGEMA_signal_5706) ) ;
    buf_clk new_AGEMA_reg_buffer_2247 ( .C (clk), .D (new_AGEMA_signal_1725), .Q (new_AGEMA_signal_5712) ) ;
    buf_clk new_AGEMA_reg_buffer_2253 ( .C (clk), .D (wk[25]), .Q (new_AGEMA_signal_5718) ) ;
    buf_clk new_AGEMA_reg_buffer_2259 ( .C (clk), .D (new_AGEMA_signal_1736), .Q (new_AGEMA_signal_5724) ) ;
    buf_clk new_AGEMA_reg_buffer_2265 ( .C (clk), .D (new_AGEMA_signal_1737), .Q (new_AGEMA_signal_5730) ) ;
    buf_clk new_AGEMA_reg_buffer_2271 ( .C (clk), .D (wk[23]), .Q (new_AGEMA_signal_5736) ) ;
    buf_clk new_AGEMA_reg_buffer_2277 ( .C (clk), .D (new_AGEMA_signal_1748), .Q (new_AGEMA_signal_5742) ) ;
    buf_clk new_AGEMA_reg_buffer_2283 ( .C (clk), .D (new_AGEMA_signal_1749), .Q (new_AGEMA_signal_5748) ) ;
    buf_clk new_AGEMA_reg_buffer_2289 ( .C (clk), .D (wk[21]), .Q (new_AGEMA_signal_5754) ) ;
    buf_clk new_AGEMA_reg_buffer_2295 ( .C (clk), .D (new_AGEMA_signal_1760), .Q (new_AGEMA_signal_5760) ) ;
    buf_clk new_AGEMA_reg_buffer_2301 ( .C (clk), .D (new_AGEMA_signal_1761), .Q (new_AGEMA_signal_5766) ) ;
    buf_clk new_AGEMA_reg_buffer_2307 ( .C (clk), .D (wk[1]), .Q (new_AGEMA_signal_5772) ) ;
    buf_clk new_AGEMA_reg_buffer_2313 ( .C (clk), .D (new_AGEMA_signal_1772), .Q (new_AGEMA_signal_5778) ) ;
    buf_clk new_AGEMA_reg_buffer_2319 ( .C (clk), .D (new_AGEMA_signal_1773), .Q (new_AGEMA_signal_5784) ) ;
    buf_clk new_AGEMA_reg_buffer_2325 ( .C (clk), .D (wk[19]), .Q (new_AGEMA_signal_5790) ) ;
    buf_clk new_AGEMA_reg_buffer_2331 ( .C (clk), .D (new_AGEMA_signal_1778), .Q (new_AGEMA_signal_5796) ) ;
    buf_clk new_AGEMA_reg_buffer_2337 ( .C (clk), .D (new_AGEMA_signal_1779), .Q (new_AGEMA_signal_5802) ) ;
    buf_clk new_AGEMA_reg_buffer_2343 ( .C (clk), .D (wk[17]), .Q (new_AGEMA_signal_5808) ) ;
    buf_clk new_AGEMA_reg_buffer_2349 ( .C (clk), .D (new_AGEMA_signal_1790), .Q (new_AGEMA_signal_5814) ) ;
    buf_clk new_AGEMA_reg_buffer_2355 ( .C (clk), .D (new_AGEMA_signal_1791), .Q (new_AGEMA_signal_5820) ) ;
    buf_clk new_AGEMA_reg_buffer_2361 ( .C (clk), .D (wk[15]), .Q (new_AGEMA_signal_5826) ) ;
    buf_clk new_AGEMA_reg_buffer_2367 ( .C (clk), .D (new_AGEMA_signal_1802), .Q (new_AGEMA_signal_5832) ) ;
    buf_clk new_AGEMA_reg_buffer_2373 ( .C (clk), .D (new_AGEMA_signal_1803), .Q (new_AGEMA_signal_5838) ) ;
    buf_clk new_AGEMA_reg_buffer_2379 ( .C (clk), .D (wk[13]), .Q (new_AGEMA_signal_5844) ) ;
    buf_clk new_AGEMA_reg_buffer_2385 ( .C (clk), .D (new_AGEMA_signal_1814), .Q (new_AGEMA_signal_5850) ) ;
    buf_clk new_AGEMA_reg_buffer_2391 ( .C (clk), .D (new_AGEMA_signal_1815), .Q (new_AGEMA_signal_5856) ) ;
    buf_clk new_AGEMA_reg_buffer_2397 ( .C (clk), .D (wk[11]), .Q (new_AGEMA_signal_5862) ) ;
    buf_clk new_AGEMA_reg_buffer_2403 ( .C (clk), .D (new_AGEMA_signal_1826), .Q (new_AGEMA_signal_5868) ) ;
    buf_clk new_AGEMA_reg_buffer_2409 ( .C (clk), .D (new_AGEMA_signal_1827), .Q (new_AGEMA_signal_5874) ) ;
    buf_clk new_AGEMA_reg_buffer_2415 ( .C (clk), .D (Midori_rounds_SelectedKey_9_), .Q (new_AGEMA_signal_5880) ) ;
    buf_clk new_AGEMA_reg_buffer_2421 ( .C (clk), .D (new_AGEMA_signal_1852), .Q (new_AGEMA_signal_5886) ) ;
    buf_clk new_AGEMA_reg_buffer_2427 ( .C (clk), .D (new_AGEMA_signal_1853), .Q (new_AGEMA_signal_5892) ) ;
    buf_clk new_AGEMA_reg_buffer_2433 ( .C (clk), .D (Midori_rounds_SelectedKey_7_), .Q (new_AGEMA_signal_5898) ) ;
    buf_clk new_AGEMA_reg_buffer_2439 ( .C (clk), .D (new_AGEMA_signal_2574), .Q (new_AGEMA_signal_5904) ) ;
    buf_clk new_AGEMA_reg_buffer_2445 ( .C (clk), .D (new_AGEMA_signal_2575), .Q (new_AGEMA_signal_5910) ) ;
    buf_clk new_AGEMA_reg_buffer_2451 ( .C (clk), .D (Midori_rounds_SelectedKey_63_), .Q (new_AGEMA_signal_5916) ) ;
    buf_clk new_AGEMA_reg_buffer_2457 ( .C (clk), .D (new_AGEMA_signal_2670), .Q (new_AGEMA_signal_5922) ) ;
    buf_clk new_AGEMA_reg_buffer_2463 ( .C (clk), .D (new_AGEMA_signal_2671), .Q (new_AGEMA_signal_5928) ) ;
    buf_clk new_AGEMA_reg_buffer_2469 ( .C (clk), .D (Midori_rounds_SelectedKey_61_), .Q (new_AGEMA_signal_5934) ) ;
    buf_clk new_AGEMA_reg_buffer_2475 ( .C (clk), .D (new_AGEMA_signal_2666), .Q (new_AGEMA_signal_5940) ) ;
    buf_clk new_AGEMA_reg_buffer_2481 ( .C (clk), .D (new_AGEMA_signal_2667), .Q (new_AGEMA_signal_5946) ) ;
    buf_clk new_AGEMA_reg_buffer_2487 ( .C (clk), .D (Midori_rounds_SelectedKey_5_), .Q (new_AGEMA_signal_5952) ) ;
    buf_clk new_AGEMA_reg_buffer_2493 ( .C (clk), .D (new_AGEMA_signal_2570), .Q (new_AGEMA_signal_5958) ) ;
    buf_clk new_AGEMA_reg_buffer_2499 ( .C (clk), .D (new_AGEMA_signal_2571), .Q (new_AGEMA_signal_5964) ) ;
    buf_clk new_AGEMA_reg_buffer_2505 ( .C (clk), .D (Midori_rounds_SelectedKey_59_), .Q (new_AGEMA_signal_5970) ) ;
    buf_clk new_AGEMA_reg_buffer_2511 ( .C (clk), .D (new_AGEMA_signal_2662), .Q (new_AGEMA_signal_5976) ) ;
    buf_clk new_AGEMA_reg_buffer_2517 ( .C (clk), .D (new_AGEMA_signal_2663), .Q (new_AGEMA_signal_5982) ) ;
    buf_clk new_AGEMA_reg_buffer_2523 ( .C (clk), .D (Midori_rounds_SelectedKey_57_), .Q (new_AGEMA_signal_5988) ) ;
    buf_clk new_AGEMA_reg_buffer_2529 ( .C (clk), .D (new_AGEMA_signal_2658), .Q (new_AGEMA_signal_5994) ) ;
    buf_clk new_AGEMA_reg_buffer_2535 ( .C (clk), .D (new_AGEMA_signal_2659), .Q (new_AGEMA_signal_6000) ) ;
    buf_clk new_AGEMA_reg_buffer_2541 ( .C (clk), .D (Midori_rounds_SelectedKey_55_), .Q (new_AGEMA_signal_6006) ) ;
    buf_clk new_AGEMA_reg_buffer_2547 ( .C (clk), .D (new_AGEMA_signal_2654), .Q (new_AGEMA_signal_6012) ) ;
    buf_clk new_AGEMA_reg_buffer_2553 ( .C (clk), .D (new_AGEMA_signal_2655), .Q (new_AGEMA_signal_6018) ) ;
    buf_clk new_AGEMA_reg_buffer_2559 ( .C (clk), .D (Midori_rounds_SelectedKey_53_), .Q (new_AGEMA_signal_6024) ) ;
    buf_clk new_AGEMA_reg_buffer_2565 ( .C (clk), .D (new_AGEMA_signal_2650), .Q (new_AGEMA_signal_6030) ) ;
    buf_clk new_AGEMA_reg_buffer_2571 ( .C (clk), .D (new_AGEMA_signal_2651), .Q (new_AGEMA_signal_6036) ) ;
    buf_clk new_AGEMA_reg_buffer_2577 ( .C (clk), .D (Midori_rounds_SelectedKey_51_), .Q (new_AGEMA_signal_6042) ) ;
    buf_clk new_AGEMA_reg_buffer_2583 ( .C (clk), .D (new_AGEMA_signal_2646), .Q (new_AGEMA_signal_6048) ) ;
    buf_clk new_AGEMA_reg_buffer_2589 ( .C (clk), .D (new_AGEMA_signal_2647), .Q (new_AGEMA_signal_6054) ) ;
    buf_clk new_AGEMA_reg_buffer_2595 ( .C (clk), .D (Midori_rounds_SelectedKey_49_), .Q (new_AGEMA_signal_6060) ) ;
    buf_clk new_AGEMA_reg_buffer_2601 ( .C (clk), .D (new_AGEMA_signal_2642), .Q (new_AGEMA_signal_6066) ) ;
    buf_clk new_AGEMA_reg_buffer_2607 ( .C (clk), .D (new_AGEMA_signal_2643), .Q (new_AGEMA_signal_6072) ) ;
    buf_clk new_AGEMA_reg_buffer_2613 ( .C (clk), .D (Midori_rounds_SelectedKey_47_), .Q (new_AGEMA_signal_6078) ) ;
    buf_clk new_AGEMA_reg_buffer_2619 ( .C (clk), .D (new_AGEMA_signal_2638), .Q (new_AGEMA_signal_6084) ) ;
    buf_clk new_AGEMA_reg_buffer_2625 ( .C (clk), .D (new_AGEMA_signal_2639), .Q (new_AGEMA_signal_6090) ) ;
    buf_clk new_AGEMA_reg_buffer_2631 ( .C (clk), .D (Midori_rounds_SelectedKey_45_), .Q (new_AGEMA_signal_6096) ) ;
    buf_clk new_AGEMA_reg_buffer_2637 ( .C (clk), .D (new_AGEMA_signal_2634), .Q (new_AGEMA_signal_6102) ) ;
    buf_clk new_AGEMA_reg_buffer_2643 ( .C (clk), .D (new_AGEMA_signal_2635), .Q (new_AGEMA_signal_6108) ) ;
    buf_clk new_AGEMA_reg_buffer_2649 ( .C (clk), .D (Midori_rounds_SelectedKey_43_), .Q (new_AGEMA_signal_6114) ) ;
    buf_clk new_AGEMA_reg_buffer_2655 ( .C (clk), .D (new_AGEMA_signal_2630), .Q (new_AGEMA_signal_6120) ) ;
    buf_clk new_AGEMA_reg_buffer_2661 ( .C (clk), .D (new_AGEMA_signal_2631), .Q (new_AGEMA_signal_6126) ) ;
    buf_clk new_AGEMA_reg_buffer_2667 ( .C (clk), .D (Midori_rounds_SelectedKey_41_), .Q (new_AGEMA_signal_6132) ) ;
    buf_clk new_AGEMA_reg_buffer_2673 ( .C (clk), .D (new_AGEMA_signal_2626), .Q (new_AGEMA_signal_6138) ) ;
    buf_clk new_AGEMA_reg_buffer_2679 ( .C (clk), .D (new_AGEMA_signal_2627), .Q (new_AGEMA_signal_6144) ) ;
    buf_clk new_AGEMA_reg_buffer_2685 ( .C (clk), .D (Midori_rounds_SelectedKey_3_), .Q (new_AGEMA_signal_6150) ) ;
    buf_clk new_AGEMA_reg_buffer_2691 ( .C (clk), .D (new_AGEMA_signal_1846), .Q (new_AGEMA_signal_6156) ) ;
    buf_clk new_AGEMA_reg_buffer_2697 ( .C (clk), .D (new_AGEMA_signal_1847), .Q (new_AGEMA_signal_6162) ) ;
    buf_clk new_AGEMA_reg_buffer_2703 ( .C (clk), .D (Midori_rounds_SelectedKey_39_), .Q (new_AGEMA_signal_6168) ) ;
    buf_clk new_AGEMA_reg_buffer_2709 ( .C (clk), .D (new_AGEMA_signal_2622), .Q (new_AGEMA_signal_6174) ) ;
    buf_clk new_AGEMA_reg_buffer_2715 ( .C (clk), .D (new_AGEMA_signal_2623), .Q (new_AGEMA_signal_6180) ) ;
    buf_clk new_AGEMA_reg_buffer_2721 ( .C (clk), .D (Midori_rounds_SelectedKey_37_), .Q (new_AGEMA_signal_6186) ) ;
    buf_clk new_AGEMA_reg_buffer_2727 ( .C (clk), .D (new_AGEMA_signal_2618), .Q (new_AGEMA_signal_6192) ) ;
    buf_clk new_AGEMA_reg_buffer_2733 ( .C (clk), .D (new_AGEMA_signal_2619), .Q (new_AGEMA_signal_6198) ) ;
    buf_clk new_AGEMA_reg_buffer_2739 ( .C (clk), .D (Midori_rounds_SelectedKey_35_), .Q (new_AGEMA_signal_6204) ) ;
    buf_clk new_AGEMA_reg_buffer_2745 ( .C (clk), .D (new_AGEMA_signal_2614), .Q (new_AGEMA_signal_6210) ) ;
    buf_clk new_AGEMA_reg_buffer_2751 ( .C (clk), .D (new_AGEMA_signal_2615), .Q (new_AGEMA_signal_6216) ) ;
    buf_clk new_AGEMA_reg_buffer_2757 ( .C (clk), .D (Midori_rounds_SelectedKey_33_), .Q (new_AGEMA_signal_6222) ) ;
    buf_clk new_AGEMA_reg_buffer_2763 ( .C (clk), .D (new_AGEMA_signal_2610), .Q (new_AGEMA_signal_6228) ) ;
    buf_clk new_AGEMA_reg_buffer_2769 ( .C (clk), .D (new_AGEMA_signal_2611), .Q (new_AGEMA_signal_6234) ) ;
    buf_clk new_AGEMA_reg_buffer_2775 ( .C (clk), .D (Midori_rounds_SelectedKey_31_), .Q (new_AGEMA_signal_6240) ) ;
    buf_clk new_AGEMA_reg_buffer_2781 ( .C (clk), .D (new_AGEMA_signal_2606), .Q (new_AGEMA_signal_6246) ) ;
    buf_clk new_AGEMA_reg_buffer_2787 ( .C (clk), .D (new_AGEMA_signal_2607), .Q (new_AGEMA_signal_6252) ) ;
    buf_clk new_AGEMA_reg_buffer_2793 ( .C (clk), .D (Midori_rounds_SelectedKey_29_), .Q (new_AGEMA_signal_6258) ) ;
    buf_clk new_AGEMA_reg_buffer_2799 ( .C (clk), .D (new_AGEMA_signal_2602), .Q (new_AGEMA_signal_6264) ) ;
    buf_clk new_AGEMA_reg_buffer_2805 ( .C (clk), .D (new_AGEMA_signal_2603), .Q (new_AGEMA_signal_6270) ) ;
    buf_clk new_AGEMA_reg_buffer_2811 ( .C (clk), .D (Midori_rounds_SelectedKey_27_), .Q (new_AGEMA_signal_6276) ) ;
    buf_clk new_AGEMA_reg_buffer_2817 ( .C (clk), .D (new_AGEMA_signal_2598), .Q (new_AGEMA_signal_6282) ) ;
    buf_clk new_AGEMA_reg_buffer_2823 ( .C (clk), .D (new_AGEMA_signal_2599), .Q (new_AGEMA_signal_6288) ) ;
    buf_clk new_AGEMA_reg_buffer_2829 ( .C (clk), .D (Midori_rounds_SelectedKey_25_), .Q (new_AGEMA_signal_6294) ) ;
    buf_clk new_AGEMA_reg_buffer_2835 ( .C (clk), .D (new_AGEMA_signal_2596), .Q (new_AGEMA_signal_6300) ) ;
    buf_clk new_AGEMA_reg_buffer_2841 ( .C (clk), .D (new_AGEMA_signal_2597), .Q (new_AGEMA_signal_6306) ) ;
    buf_clk new_AGEMA_reg_buffer_2847 ( .C (clk), .D (Midori_rounds_SelectedKey_23_), .Q (new_AGEMA_signal_6312) ) ;
    buf_clk new_AGEMA_reg_buffer_2853 ( .C (clk), .D (new_AGEMA_signal_2592), .Q (new_AGEMA_signal_6318) ) ;
    buf_clk new_AGEMA_reg_buffer_2859 ( .C (clk), .D (new_AGEMA_signal_2593), .Q (new_AGEMA_signal_6324) ) ;
    buf_clk new_AGEMA_reg_buffer_2865 ( .C (clk), .D (Midori_rounds_SelectedKey_21_), .Q (new_AGEMA_signal_6330) ) ;
    buf_clk new_AGEMA_reg_buffer_2871 ( .C (clk), .D (new_AGEMA_signal_2588), .Q (new_AGEMA_signal_6336) ) ;
    buf_clk new_AGEMA_reg_buffer_2877 ( .C (clk), .D (new_AGEMA_signal_2589), .Q (new_AGEMA_signal_6342) ) ;
    buf_clk new_AGEMA_reg_buffer_2883 ( .C (clk), .D (Midori_rounds_SelectedKey_1_), .Q (new_AGEMA_signal_6348) ) ;
    buf_clk new_AGEMA_reg_buffer_2889 ( .C (clk), .D (new_AGEMA_signal_1842), .Q (new_AGEMA_signal_6354) ) ;
    buf_clk new_AGEMA_reg_buffer_2895 ( .C (clk), .D (new_AGEMA_signal_1843), .Q (new_AGEMA_signal_6360) ) ;
    buf_clk new_AGEMA_reg_buffer_2901 ( .C (clk), .D (Midori_rounds_SelectedKey_19_), .Q (new_AGEMA_signal_6366) ) ;
    buf_clk new_AGEMA_reg_buffer_2907 ( .C (clk), .D (new_AGEMA_signal_2584), .Q (new_AGEMA_signal_6372) ) ;
    buf_clk new_AGEMA_reg_buffer_2913 ( .C (clk), .D (new_AGEMA_signal_2585), .Q (new_AGEMA_signal_6378) ) ;
    buf_clk new_AGEMA_reg_buffer_2919 ( .C (clk), .D (Midori_rounds_SelectedKey_17_), .Q (new_AGEMA_signal_6384) ) ;
    buf_clk new_AGEMA_reg_buffer_2925 ( .C (clk), .D (new_AGEMA_signal_2580), .Q (new_AGEMA_signal_6390) ) ;
    buf_clk new_AGEMA_reg_buffer_2931 ( .C (clk), .D (new_AGEMA_signal_2581), .Q (new_AGEMA_signal_6396) ) ;
    buf_clk new_AGEMA_reg_buffer_2937 ( .C (clk), .D (Midori_rounds_SelectedKey_15_), .Q (new_AGEMA_signal_6402) ) ;
    buf_clk new_AGEMA_reg_buffer_2943 ( .C (clk), .D (new_AGEMA_signal_1862), .Q (new_AGEMA_signal_6408) ) ;
    buf_clk new_AGEMA_reg_buffer_2949 ( .C (clk), .D (new_AGEMA_signal_1863), .Q (new_AGEMA_signal_6414) ) ;
    buf_clk new_AGEMA_reg_buffer_2955 ( .C (clk), .D (Midori_rounds_SelectedKey_13_), .Q (new_AGEMA_signal_6420) ) ;
    buf_clk new_AGEMA_reg_buffer_2961 ( .C (clk), .D (new_AGEMA_signal_1858), .Q (new_AGEMA_signal_6426) ) ;
    buf_clk new_AGEMA_reg_buffer_2967 ( .C (clk), .D (new_AGEMA_signal_1859), .Q (new_AGEMA_signal_6432) ) ;
    buf_clk new_AGEMA_reg_buffer_2973 ( .C (clk), .D (Midori_rounds_SelectedKey_11_), .Q (new_AGEMA_signal_6438) ) ;
    buf_clk new_AGEMA_reg_buffer_2979 ( .C (clk), .D (new_AGEMA_signal_1856), .Q (new_AGEMA_signal_6444) ) ;
    buf_clk new_AGEMA_reg_buffer_2985 ( .C (clk), .D (new_AGEMA_signal_1857), .Q (new_AGEMA_signal_6450) ) ;
    buf_clk new_AGEMA_reg_buffer_2991 ( .C (clk), .D (reset), .Q (new_AGEMA_signal_6456) ) ;
    buf_clk new_AGEMA_reg_buffer_2997 ( .C (clk), .D (Midori_add_Result_Start[1]), .Q (new_AGEMA_signal_6462) ) ;
    buf_clk new_AGEMA_reg_buffer_3003 ( .C (clk), .D (new_AGEMA_signal_2332), .Q (new_AGEMA_signal_6468) ) ;
    buf_clk new_AGEMA_reg_buffer_3009 ( .C (clk), .D (new_AGEMA_signal_2333), .Q (new_AGEMA_signal_6474) ) ;
    buf_clk new_AGEMA_reg_buffer_3015 ( .C (clk), .D (Midori_add_Result_Start[3]), .Q (new_AGEMA_signal_6480) ) ;
    buf_clk new_AGEMA_reg_buffer_3021 ( .C (clk), .D (new_AGEMA_signal_2244), .Q (new_AGEMA_signal_6486) ) ;
    buf_clk new_AGEMA_reg_buffer_3027 ( .C (clk), .D (new_AGEMA_signal_2245), .Q (new_AGEMA_signal_6492) ) ;
    buf_clk new_AGEMA_reg_buffer_3033 ( .C (clk), .D (Midori_add_Result_Start[5]), .Q (new_AGEMA_signal_6498) ) ;
    buf_clk new_AGEMA_reg_buffer_3039 ( .C (clk), .D (new_AGEMA_signal_2156), .Q (new_AGEMA_signal_6504) ) ;
    buf_clk new_AGEMA_reg_buffer_3045 ( .C (clk), .D (new_AGEMA_signal_2157), .Q (new_AGEMA_signal_6510) ) ;
    buf_clk new_AGEMA_reg_buffer_3051 ( .C (clk), .D (Midori_add_Result_Start[7]), .Q (new_AGEMA_signal_6516) ) ;
    buf_clk new_AGEMA_reg_buffer_3057 ( .C (clk), .D (new_AGEMA_signal_2132), .Q (new_AGEMA_signal_6522) ) ;
    buf_clk new_AGEMA_reg_buffer_3063 ( .C (clk), .D (new_AGEMA_signal_2133), .Q (new_AGEMA_signal_6528) ) ;
    buf_clk new_AGEMA_reg_buffer_3069 ( .C (clk), .D (Midori_add_Result_Start[9]), .Q (new_AGEMA_signal_6534) ) ;
    buf_clk new_AGEMA_reg_buffer_3075 ( .C (clk), .D (new_AGEMA_signal_2124), .Q (new_AGEMA_signal_6540) ) ;
    buf_clk new_AGEMA_reg_buffer_3081 ( .C (clk), .D (new_AGEMA_signal_2125), .Q (new_AGEMA_signal_6546) ) ;
    buf_clk new_AGEMA_reg_buffer_3087 ( .C (clk), .D (Midori_add_Result_Start[11]), .Q (new_AGEMA_signal_6552) ) ;
    buf_clk new_AGEMA_reg_buffer_3093 ( .C (clk), .D (new_AGEMA_signal_2368), .Q (new_AGEMA_signal_6558) ) ;
    buf_clk new_AGEMA_reg_buffer_3099 ( .C (clk), .D (new_AGEMA_signal_2369), .Q (new_AGEMA_signal_6564) ) ;
    buf_clk new_AGEMA_reg_buffer_3105 ( .C (clk), .D (Midori_add_Result_Start[13]), .Q (new_AGEMA_signal_6570) ) ;
    buf_clk new_AGEMA_reg_buffer_3111 ( .C (clk), .D (new_AGEMA_signal_2360), .Q (new_AGEMA_signal_6576) ) ;
    buf_clk new_AGEMA_reg_buffer_3117 ( .C (clk), .D (new_AGEMA_signal_2361), .Q (new_AGEMA_signal_6582) ) ;
    buf_clk new_AGEMA_reg_buffer_3123 ( .C (clk), .D (Midori_add_Result_Start[15]), .Q (new_AGEMA_signal_6588) ) ;
    buf_clk new_AGEMA_reg_buffer_3129 ( .C (clk), .D (new_AGEMA_signal_2352), .Q (new_AGEMA_signal_6594) ) ;
    buf_clk new_AGEMA_reg_buffer_3135 ( .C (clk), .D (new_AGEMA_signal_2353), .Q (new_AGEMA_signal_6600) ) ;
    buf_clk new_AGEMA_reg_buffer_3141 ( .C (clk), .D (Midori_add_Result_Start[17]), .Q (new_AGEMA_signal_6606) ) ;
    buf_clk new_AGEMA_reg_buffer_3147 ( .C (clk), .D (new_AGEMA_signal_2344), .Q (new_AGEMA_signal_6612) ) ;
    buf_clk new_AGEMA_reg_buffer_3153 ( .C (clk), .D (new_AGEMA_signal_2345), .Q (new_AGEMA_signal_6618) ) ;
    buf_clk new_AGEMA_reg_buffer_3159 ( .C (clk), .D (Midori_add_Result_Start[19]), .Q (new_AGEMA_signal_6624) ) ;
    buf_clk new_AGEMA_reg_buffer_3165 ( .C (clk), .D (new_AGEMA_signal_2336), .Q (new_AGEMA_signal_6630) ) ;
    buf_clk new_AGEMA_reg_buffer_3171 ( .C (clk), .D (new_AGEMA_signal_2337), .Q (new_AGEMA_signal_6636) ) ;
    buf_clk new_AGEMA_reg_buffer_3177 ( .C (clk), .D (Midori_add_Result_Start[21]), .Q (new_AGEMA_signal_6642) ) ;
    buf_clk new_AGEMA_reg_buffer_3183 ( .C (clk), .D (new_AGEMA_signal_2324), .Q (new_AGEMA_signal_6648) ) ;
    buf_clk new_AGEMA_reg_buffer_3189 ( .C (clk), .D (new_AGEMA_signal_2325), .Q (new_AGEMA_signal_6654) ) ;
    buf_clk new_AGEMA_reg_buffer_3195 ( .C (clk), .D (Midori_add_Result_Start[23]), .Q (new_AGEMA_signal_6660) ) ;
    buf_clk new_AGEMA_reg_buffer_3201 ( .C (clk), .D (new_AGEMA_signal_2316), .Q (new_AGEMA_signal_6666) ) ;
    buf_clk new_AGEMA_reg_buffer_3207 ( .C (clk), .D (new_AGEMA_signal_2317), .Q (new_AGEMA_signal_6672) ) ;
    buf_clk new_AGEMA_reg_buffer_3213 ( .C (clk), .D (Midori_add_Result_Start[25]), .Q (new_AGEMA_signal_6678) ) ;
    buf_clk new_AGEMA_reg_buffer_3219 ( .C (clk), .D (new_AGEMA_signal_2308), .Q (new_AGEMA_signal_6684) ) ;
    buf_clk new_AGEMA_reg_buffer_3225 ( .C (clk), .D (new_AGEMA_signal_2309), .Q (new_AGEMA_signal_6690) ) ;
    buf_clk new_AGEMA_reg_buffer_3231 ( .C (clk), .D (Midori_add_Result_Start[27]), .Q (new_AGEMA_signal_6696) ) ;
    buf_clk new_AGEMA_reg_buffer_3237 ( .C (clk), .D (new_AGEMA_signal_2300), .Q (new_AGEMA_signal_6702) ) ;
    buf_clk new_AGEMA_reg_buffer_3243 ( .C (clk), .D (new_AGEMA_signal_2301), .Q (new_AGEMA_signal_6708) ) ;
    buf_clk new_AGEMA_reg_buffer_3249 ( .C (clk), .D (Midori_add_Result_Start[29]), .Q (new_AGEMA_signal_6714) ) ;
    buf_clk new_AGEMA_reg_buffer_3255 ( .C (clk), .D (new_AGEMA_signal_2292), .Q (new_AGEMA_signal_6720) ) ;
    buf_clk new_AGEMA_reg_buffer_3261 ( .C (clk), .D (new_AGEMA_signal_2293), .Q (new_AGEMA_signal_6726) ) ;
    buf_clk new_AGEMA_reg_buffer_3267 ( .C (clk), .D (Midori_add_Result_Start[31]), .Q (new_AGEMA_signal_6732) ) ;
    buf_clk new_AGEMA_reg_buffer_3273 ( .C (clk), .D (new_AGEMA_signal_2280), .Q (new_AGEMA_signal_6738) ) ;
    buf_clk new_AGEMA_reg_buffer_3279 ( .C (clk), .D (new_AGEMA_signal_2281), .Q (new_AGEMA_signal_6744) ) ;
    buf_clk new_AGEMA_reg_buffer_3285 ( .C (clk), .D (Midori_add_Result_Start[33]), .Q (new_AGEMA_signal_6750) ) ;
    buf_clk new_AGEMA_reg_buffer_3291 ( .C (clk), .D (new_AGEMA_signal_2272), .Q (new_AGEMA_signal_6756) ) ;
    buf_clk new_AGEMA_reg_buffer_3297 ( .C (clk), .D (new_AGEMA_signal_2273), .Q (new_AGEMA_signal_6762) ) ;
    buf_clk new_AGEMA_reg_buffer_3303 ( .C (clk), .D (Midori_add_Result_Start[35]), .Q (new_AGEMA_signal_6768) ) ;
    buf_clk new_AGEMA_reg_buffer_3309 ( .C (clk), .D (new_AGEMA_signal_2264), .Q (new_AGEMA_signal_6774) ) ;
    buf_clk new_AGEMA_reg_buffer_3315 ( .C (clk), .D (new_AGEMA_signal_2265), .Q (new_AGEMA_signal_6780) ) ;
    buf_clk new_AGEMA_reg_buffer_3321 ( .C (clk), .D (Midori_add_Result_Start[37]), .Q (new_AGEMA_signal_6786) ) ;
    buf_clk new_AGEMA_reg_buffer_3327 ( .C (clk), .D (new_AGEMA_signal_2256), .Q (new_AGEMA_signal_6792) ) ;
    buf_clk new_AGEMA_reg_buffer_3333 ( .C (clk), .D (new_AGEMA_signal_2257), .Q (new_AGEMA_signal_6798) ) ;
    buf_clk new_AGEMA_reg_buffer_3339 ( .C (clk), .D (Midori_add_Result_Start[39]), .Q (new_AGEMA_signal_6804) ) ;
    buf_clk new_AGEMA_reg_buffer_3345 ( .C (clk), .D (new_AGEMA_signal_2248), .Q (new_AGEMA_signal_6810) ) ;
    buf_clk new_AGEMA_reg_buffer_3351 ( .C (clk), .D (new_AGEMA_signal_2249), .Q (new_AGEMA_signal_6816) ) ;
    buf_clk new_AGEMA_reg_buffer_3357 ( .C (clk), .D (Midori_add_Result_Start[41]), .Q (new_AGEMA_signal_6822) ) ;
    buf_clk new_AGEMA_reg_buffer_3363 ( .C (clk), .D (new_AGEMA_signal_2236), .Q (new_AGEMA_signal_6828) ) ;
    buf_clk new_AGEMA_reg_buffer_3369 ( .C (clk), .D (new_AGEMA_signal_2237), .Q (new_AGEMA_signal_6834) ) ;
    buf_clk new_AGEMA_reg_buffer_3375 ( .C (clk), .D (Midori_add_Result_Start[43]), .Q (new_AGEMA_signal_6840) ) ;
    buf_clk new_AGEMA_reg_buffer_3381 ( .C (clk), .D (new_AGEMA_signal_2228), .Q (new_AGEMA_signal_6846) ) ;
    buf_clk new_AGEMA_reg_buffer_3387 ( .C (clk), .D (new_AGEMA_signal_2229), .Q (new_AGEMA_signal_6852) ) ;
    buf_clk new_AGEMA_reg_buffer_3393 ( .C (clk), .D (Midori_add_Result_Start[45]), .Q (new_AGEMA_signal_6858) ) ;
    buf_clk new_AGEMA_reg_buffer_3399 ( .C (clk), .D (new_AGEMA_signal_2220), .Q (new_AGEMA_signal_6864) ) ;
    buf_clk new_AGEMA_reg_buffer_3405 ( .C (clk), .D (new_AGEMA_signal_2221), .Q (new_AGEMA_signal_6870) ) ;
    buf_clk new_AGEMA_reg_buffer_3411 ( .C (clk), .D (Midori_add_Result_Start[47]), .Q (new_AGEMA_signal_6876) ) ;
    buf_clk new_AGEMA_reg_buffer_3417 ( .C (clk), .D (new_AGEMA_signal_2212), .Q (new_AGEMA_signal_6882) ) ;
    buf_clk new_AGEMA_reg_buffer_3423 ( .C (clk), .D (new_AGEMA_signal_2213), .Q (new_AGEMA_signal_6888) ) ;
    buf_clk new_AGEMA_reg_buffer_3429 ( .C (clk), .D (Midori_add_Result_Start[49]), .Q (new_AGEMA_signal_6894) ) ;
    buf_clk new_AGEMA_reg_buffer_3435 ( .C (clk), .D (new_AGEMA_signal_2204), .Q (new_AGEMA_signal_6900) ) ;
    buf_clk new_AGEMA_reg_buffer_3441 ( .C (clk), .D (new_AGEMA_signal_2205), .Q (new_AGEMA_signal_6906) ) ;
    buf_clk new_AGEMA_reg_buffer_3447 ( .C (clk), .D (Midori_add_Result_Start[51]), .Q (new_AGEMA_signal_6912) ) ;
    buf_clk new_AGEMA_reg_buffer_3453 ( .C (clk), .D (new_AGEMA_signal_2192), .Q (new_AGEMA_signal_6918) ) ;
    buf_clk new_AGEMA_reg_buffer_3459 ( .C (clk), .D (new_AGEMA_signal_2193), .Q (new_AGEMA_signal_6924) ) ;
    buf_clk new_AGEMA_reg_buffer_3465 ( .C (clk), .D (Midori_add_Result_Start[53]), .Q (new_AGEMA_signal_6930) ) ;
    buf_clk new_AGEMA_reg_buffer_3471 ( .C (clk), .D (new_AGEMA_signal_2184), .Q (new_AGEMA_signal_6936) ) ;
    buf_clk new_AGEMA_reg_buffer_3477 ( .C (clk), .D (new_AGEMA_signal_2185), .Q (new_AGEMA_signal_6942) ) ;
    buf_clk new_AGEMA_reg_buffer_3483 ( .C (clk), .D (Midori_add_Result_Start[55]), .Q (new_AGEMA_signal_6948) ) ;
    buf_clk new_AGEMA_reg_buffer_3489 ( .C (clk), .D (new_AGEMA_signal_2176), .Q (new_AGEMA_signal_6954) ) ;
    buf_clk new_AGEMA_reg_buffer_3495 ( .C (clk), .D (new_AGEMA_signal_2177), .Q (new_AGEMA_signal_6960) ) ;
    buf_clk new_AGEMA_reg_buffer_3501 ( .C (clk), .D (Midori_add_Result_Start[57]), .Q (new_AGEMA_signal_6966) ) ;
    buf_clk new_AGEMA_reg_buffer_3507 ( .C (clk), .D (new_AGEMA_signal_2168), .Q (new_AGEMA_signal_6972) ) ;
    buf_clk new_AGEMA_reg_buffer_3513 ( .C (clk), .D (new_AGEMA_signal_2169), .Q (new_AGEMA_signal_6978) ) ;
    buf_clk new_AGEMA_reg_buffer_3519 ( .C (clk), .D (Midori_add_Result_Start[59]), .Q (new_AGEMA_signal_6984) ) ;
    buf_clk new_AGEMA_reg_buffer_3525 ( .C (clk), .D (new_AGEMA_signal_2160), .Q (new_AGEMA_signal_6990) ) ;
    buf_clk new_AGEMA_reg_buffer_3531 ( .C (clk), .D (new_AGEMA_signal_2161), .Q (new_AGEMA_signal_6996) ) ;
    buf_clk new_AGEMA_reg_buffer_3537 ( .C (clk), .D (Midori_add_Result_Start[61]), .Q (new_AGEMA_signal_7002) ) ;
    buf_clk new_AGEMA_reg_buffer_3543 ( .C (clk), .D (new_AGEMA_signal_2148), .Q (new_AGEMA_signal_7008) ) ;
    buf_clk new_AGEMA_reg_buffer_3549 ( .C (clk), .D (new_AGEMA_signal_2149), .Q (new_AGEMA_signal_7014) ) ;
    buf_clk new_AGEMA_reg_buffer_3555 ( .C (clk), .D (Midori_add_Result_Start[63]), .Q (new_AGEMA_signal_7020) ) ;
    buf_clk new_AGEMA_reg_buffer_3561 ( .C (clk), .D (new_AGEMA_signal_2140), .Q (new_AGEMA_signal_7026) ) ;
    buf_clk new_AGEMA_reg_buffer_3567 ( .C (clk), .D (new_AGEMA_signal_2141), .Q (new_AGEMA_signal_7032) ) ;
    buf_clk new_AGEMA_reg_buffer_3861 ( .C (clk), .D (enc_dec), .Q (new_AGEMA_signal_7326) ) ;
    buf_clk new_AGEMA_reg_buffer_3867 ( .C (clk), .D (wk[8]), .Q (new_AGEMA_signal_7332) ) ;
    buf_clk new_AGEMA_reg_buffer_3875 ( .C (clk), .D (new_AGEMA_signal_1466), .Q (new_AGEMA_signal_7340) ) ;
    buf_clk new_AGEMA_reg_buffer_3883 ( .C (clk), .D (new_AGEMA_signal_1467), .Q (new_AGEMA_signal_7348) ) ;
    buf_clk new_AGEMA_reg_buffer_3891 ( .C (clk), .D (wk[6]), .Q (new_AGEMA_signal_7356) ) ;
    buf_clk new_AGEMA_reg_buffer_3899 ( .C (clk), .D (new_AGEMA_signal_1478), .Q (new_AGEMA_signal_7364) ) ;
    buf_clk new_AGEMA_reg_buffer_3907 ( .C (clk), .D (new_AGEMA_signal_1479), .Q (new_AGEMA_signal_7372) ) ;
    buf_clk new_AGEMA_reg_buffer_3915 ( .C (clk), .D (wk[62]), .Q (new_AGEMA_signal_7380) ) ;
    buf_clk new_AGEMA_reg_buffer_3923 ( .C (clk), .D (new_AGEMA_signal_1490), .Q (new_AGEMA_signal_7388) ) ;
    buf_clk new_AGEMA_reg_buffer_3931 ( .C (clk), .D (new_AGEMA_signal_1491), .Q (new_AGEMA_signal_7396) ) ;
    buf_clk new_AGEMA_reg_buffer_3939 ( .C (clk), .D (wk[60]), .Q (new_AGEMA_signal_7404) ) ;
    buf_clk new_AGEMA_reg_buffer_3947 ( .C (clk), .D (new_AGEMA_signal_1502), .Q (new_AGEMA_signal_7412) ) ;
    buf_clk new_AGEMA_reg_buffer_3955 ( .C (clk), .D (new_AGEMA_signal_1503), .Q (new_AGEMA_signal_7420) ) ;
    buf_clk new_AGEMA_reg_buffer_3963 ( .C (clk), .D (wk[58]), .Q (new_AGEMA_signal_7428) ) ;
    buf_clk new_AGEMA_reg_buffer_3971 ( .C (clk), .D (new_AGEMA_signal_1520), .Q (new_AGEMA_signal_7436) ) ;
    buf_clk new_AGEMA_reg_buffer_3979 ( .C (clk), .D (new_AGEMA_signal_1521), .Q (new_AGEMA_signal_7444) ) ;
    buf_clk new_AGEMA_reg_buffer_3987 ( .C (clk), .D (wk[56]), .Q (new_AGEMA_signal_7452) ) ;
    buf_clk new_AGEMA_reg_buffer_3995 ( .C (clk), .D (new_AGEMA_signal_1532), .Q (new_AGEMA_signal_7460) ) ;
    buf_clk new_AGEMA_reg_buffer_4003 ( .C (clk), .D (new_AGEMA_signal_1533), .Q (new_AGEMA_signal_7468) ) ;
    buf_clk new_AGEMA_reg_buffer_4011 ( .C (clk), .D (wk[54]), .Q (new_AGEMA_signal_7476) ) ;
    buf_clk new_AGEMA_reg_buffer_4019 ( .C (clk), .D (new_AGEMA_signal_1544), .Q (new_AGEMA_signal_7484) ) ;
    buf_clk new_AGEMA_reg_buffer_4027 ( .C (clk), .D (new_AGEMA_signal_1545), .Q (new_AGEMA_signal_7492) ) ;
    buf_clk new_AGEMA_reg_buffer_4035 ( .C (clk), .D (wk[52]), .Q (new_AGEMA_signal_7500) ) ;
    buf_clk new_AGEMA_reg_buffer_4043 ( .C (clk), .D (new_AGEMA_signal_1556), .Q (new_AGEMA_signal_7508) ) ;
    buf_clk new_AGEMA_reg_buffer_4051 ( .C (clk), .D (new_AGEMA_signal_1557), .Q (new_AGEMA_signal_7516) ) ;
    buf_clk new_AGEMA_reg_buffer_4059 ( .C (clk), .D (wk[50]), .Q (new_AGEMA_signal_7524) ) ;
    buf_clk new_AGEMA_reg_buffer_4067 ( .C (clk), .D (new_AGEMA_signal_1568), .Q (new_AGEMA_signal_7532) ) ;
    buf_clk new_AGEMA_reg_buffer_4075 ( .C (clk), .D (new_AGEMA_signal_1569), .Q (new_AGEMA_signal_7540) ) ;
    buf_clk new_AGEMA_reg_buffer_4083 ( .C (clk), .D (wk[4]), .Q (new_AGEMA_signal_7548) ) ;
    buf_clk new_AGEMA_reg_buffer_4091 ( .C (clk), .D (new_AGEMA_signal_1574), .Q (new_AGEMA_signal_7556) ) ;
    buf_clk new_AGEMA_reg_buffer_4099 ( .C (clk), .D (new_AGEMA_signal_1575), .Q (new_AGEMA_signal_7564) ) ;
    buf_clk new_AGEMA_reg_buffer_4107 ( .C (clk), .D (wk[48]), .Q (new_AGEMA_signal_7572) ) ;
    buf_clk new_AGEMA_reg_buffer_4115 ( .C (clk), .D (new_AGEMA_signal_1586), .Q (new_AGEMA_signal_7580) ) ;
    buf_clk new_AGEMA_reg_buffer_4123 ( .C (clk), .D (new_AGEMA_signal_1587), .Q (new_AGEMA_signal_7588) ) ;
    buf_clk new_AGEMA_reg_buffer_4131 ( .C (clk), .D (wk[46]), .Q (new_AGEMA_signal_7596) ) ;
    buf_clk new_AGEMA_reg_buffer_4139 ( .C (clk), .D (new_AGEMA_signal_1598), .Q (new_AGEMA_signal_7604) ) ;
    buf_clk new_AGEMA_reg_buffer_4147 ( .C (clk), .D (new_AGEMA_signal_1599), .Q (new_AGEMA_signal_7612) ) ;
    buf_clk new_AGEMA_reg_buffer_4155 ( .C (clk), .D (wk[44]), .Q (new_AGEMA_signal_7620) ) ;
    buf_clk new_AGEMA_reg_buffer_4163 ( .C (clk), .D (new_AGEMA_signal_1610), .Q (new_AGEMA_signal_7628) ) ;
    buf_clk new_AGEMA_reg_buffer_4171 ( .C (clk), .D (new_AGEMA_signal_1611), .Q (new_AGEMA_signal_7636) ) ;
    buf_clk new_AGEMA_reg_buffer_4179 ( .C (clk), .D (wk[42]), .Q (new_AGEMA_signal_7644) ) ;
    buf_clk new_AGEMA_reg_buffer_4187 ( .C (clk), .D (new_AGEMA_signal_1622), .Q (new_AGEMA_signal_7652) ) ;
    buf_clk new_AGEMA_reg_buffer_4195 ( .C (clk), .D (new_AGEMA_signal_1623), .Q (new_AGEMA_signal_7660) ) ;
    buf_clk new_AGEMA_reg_buffer_4203 ( .C (clk), .D (wk[40]), .Q (new_AGEMA_signal_7668) ) ;
    buf_clk new_AGEMA_reg_buffer_4211 ( .C (clk), .D (new_AGEMA_signal_1634), .Q (new_AGEMA_signal_7676) ) ;
    buf_clk new_AGEMA_reg_buffer_4219 ( .C (clk), .D (new_AGEMA_signal_1635), .Q (new_AGEMA_signal_7684) ) ;
    buf_clk new_AGEMA_reg_buffer_4227 ( .C (clk), .D (wk[38]), .Q (new_AGEMA_signal_7692) ) ;
    buf_clk new_AGEMA_reg_buffer_4235 ( .C (clk), .D (new_AGEMA_signal_1652), .Q (new_AGEMA_signal_7700) ) ;
    buf_clk new_AGEMA_reg_buffer_4243 ( .C (clk), .D (new_AGEMA_signal_1653), .Q (new_AGEMA_signal_7708) ) ;
    buf_clk new_AGEMA_reg_buffer_4251 ( .C (clk), .D (wk[36]), .Q (new_AGEMA_signal_7716) ) ;
    buf_clk new_AGEMA_reg_buffer_4259 ( .C (clk), .D (new_AGEMA_signal_1664), .Q (new_AGEMA_signal_7724) ) ;
    buf_clk new_AGEMA_reg_buffer_4267 ( .C (clk), .D (new_AGEMA_signal_1665), .Q (new_AGEMA_signal_7732) ) ;
    buf_clk new_AGEMA_reg_buffer_4275 ( .C (clk), .D (wk[34]), .Q (new_AGEMA_signal_7740) ) ;
    buf_clk new_AGEMA_reg_buffer_4283 ( .C (clk), .D (new_AGEMA_signal_1676), .Q (new_AGEMA_signal_7748) ) ;
    buf_clk new_AGEMA_reg_buffer_4291 ( .C (clk), .D (new_AGEMA_signal_1677), .Q (new_AGEMA_signal_7756) ) ;
    buf_clk new_AGEMA_reg_buffer_4299 ( .C (clk), .D (wk[32]), .Q (new_AGEMA_signal_7764) ) ;
    buf_clk new_AGEMA_reg_buffer_4307 ( .C (clk), .D (new_AGEMA_signal_1688), .Q (new_AGEMA_signal_7772) ) ;
    buf_clk new_AGEMA_reg_buffer_4315 ( .C (clk), .D (new_AGEMA_signal_1689), .Q (new_AGEMA_signal_7780) ) ;
    buf_clk new_AGEMA_reg_buffer_4323 ( .C (clk), .D (wk[30]), .Q (new_AGEMA_signal_7788) ) ;
    buf_clk new_AGEMA_reg_buffer_4331 ( .C (clk), .D (new_AGEMA_signal_1700), .Q (new_AGEMA_signal_7796) ) ;
    buf_clk new_AGEMA_reg_buffer_4339 ( .C (clk), .D (new_AGEMA_signal_1701), .Q (new_AGEMA_signal_7804) ) ;
    buf_clk new_AGEMA_reg_buffer_4347 ( .C (clk), .D (wk[2]), .Q (new_AGEMA_signal_7812) ) ;
    buf_clk new_AGEMA_reg_buffer_4355 ( .C (clk), .D (new_AGEMA_signal_1706), .Q (new_AGEMA_signal_7820) ) ;
    buf_clk new_AGEMA_reg_buffer_4363 ( .C (clk), .D (new_AGEMA_signal_1707), .Q (new_AGEMA_signal_7828) ) ;
    buf_clk new_AGEMA_reg_buffer_4371 ( .C (clk), .D (wk[28]), .Q (new_AGEMA_signal_7836) ) ;
    buf_clk new_AGEMA_reg_buffer_4379 ( .C (clk), .D (new_AGEMA_signal_1718), .Q (new_AGEMA_signal_7844) ) ;
    buf_clk new_AGEMA_reg_buffer_4387 ( .C (clk), .D (new_AGEMA_signal_1719), .Q (new_AGEMA_signal_7852) ) ;
    buf_clk new_AGEMA_reg_buffer_4395 ( .C (clk), .D (wk[26]), .Q (new_AGEMA_signal_7860) ) ;
    buf_clk new_AGEMA_reg_buffer_4403 ( .C (clk), .D (new_AGEMA_signal_1730), .Q (new_AGEMA_signal_7868) ) ;
    buf_clk new_AGEMA_reg_buffer_4411 ( .C (clk), .D (new_AGEMA_signal_1731), .Q (new_AGEMA_signal_7876) ) ;
    buf_clk new_AGEMA_reg_buffer_4419 ( .C (clk), .D (wk[24]), .Q (new_AGEMA_signal_7884) ) ;
    buf_clk new_AGEMA_reg_buffer_4427 ( .C (clk), .D (new_AGEMA_signal_1742), .Q (new_AGEMA_signal_7892) ) ;
    buf_clk new_AGEMA_reg_buffer_4435 ( .C (clk), .D (new_AGEMA_signal_1743), .Q (new_AGEMA_signal_7900) ) ;
    buf_clk new_AGEMA_reg_buffer_4443 ( .C (clk), .D (wk[22]), .Q (new_AGEMA_signal_7908) ) ;
    buf_clk new_AGEMA_reg_buffer_4451 ( .C (clk), .D (new_AGEMA_signal_1754), .Q (new_AGEMA_signal_7916) ) ;
    buf_clk new_AGEMA_reg_buffer_4459 ( .C (clk), .D (new_AGEMA_signal_1755), .Q (new_AGEMA_signal_7924) ) ;
    buf_clk new_AGEMA_reg_buffer_4467 ( .C (clk), .D (wk[20]), .Q (new_AGEMA_signal_7932) ) ;
    buf_clk new_AGEMA_reg_buffer_4475 ( .C (clk), .D (new_AGEMA_signal_1766), .Q (new_AGEMA_signal_7940) ) ;
    buf_clk new_AGEMA_reg_buffer_4483 ( .C (clk), .D (new_AGEMA_signal_1767), .Q (new_AGEMA_signal_7948) ) ;
    buf_clk new_AGEMA_reg_buffer_4491 ( .C (clk), .D (wk[18]), .Q (new_AGEMA_signal_7956) ) ;
    buf_clk new_AGEMA_reg_buffer_4499 ( .C (clk), .D (new_AGEMA_signal_1784), .Q (new_AGEMA_signal_7964) ) ;
    buf_clk new_AGEMA_reg_buffer_4507 ( .C (clk), .D (new_AGEMA_signal_1785), .Q (new_AGEMA_signal_7972) ) ;
    buf_clk new_AGEMA_reg_buffer_4515 ( .C (clk), .D (wk[16]), .Q (new_AGEMA_signal_7980) ) ;
    buf_clk new_AGEMA_reg_buffer_4523 ( .C (clk), .D (new_AGEMA_signal_1796), .Q (new_AGEMA_signal_7988) ) ;
    buf_clk new_AGEMA_reg_buffer_4531 ( .C (clk), .D (new_AGEMA_signal_1797), .Q (new_AGEMA_signal_7996) ) ;
    buf_clk new_AGEMA_reg_buffer_4539 ( .C (clk), .D (wk[14]), .Q (new_AGEMA_signal_8004) ) ;
    buf_clk new_AGEMA_reg_buffer_4547 ( .C (clk), .D (new_AGEMA_signal_1808), .Q (new_AGEMA_signal_8012) ) ;
    buf_clk new_AGEMA_reg_buffer_4555 ( .C (clk), .D (new_AGEMA_signal_1809), .Q (new_AGEMA_signal_8020) ) ;
    buf_clk new_AGEMA_reg_buffer_4563 ( .C (clk), .D (wk[12]), .Q (new_AGEMA_signal_8028) ) ;
    buf_clk new_AGEMA_reg_buffer_4571 ( .C (clk), .D (new_AGEMA_signal_1820), .Q (new_AGEMA_signal_8036) ) ;
    buf_clk new_AGEMA_reg_buffer_4579 ( .C (clk), .D (new_AGEMA_signal_1821), .Q (new_AGEMA_signal_8044) ) ;
    buf_clk new_AGEMA_reg_buffer_4587 ( .C (clk), .D (wk[10]), .Q (new_AGEMA_signal_8052) ) ;
    buf_clk new_AGEMA_reg_buffer_4595 ( .C (clk), .D (new_AGEMA_signal_1832), .Q (new_AGEMA_signal_8060) ) ;
    buf_clk new_AGEMA_reg_buffer_4603 ( .C (clk), .D (new_AGEMA_signal_1833), .Q (new_AGEMA_signal_8068) ) ;
    buf_clk new_AGEMA_reg_buffer_4611 ( .C (clk), .D (wk[0]), .Q (new_AGEMA_signal_8076) ) ;
    buf_clk new_AGEMA_reg_buffer_4619 ( .C (clk), .D (new_AGEMA_signal_1838), .Q (new_AGEMA_signal_8084) ) ;
    buf_clk new_AGEMA_reg_buffer_4627 ( .C (clk), .D (new_AGEMA_signal_1839), .Q (new_AGEMA_signal_8092) ) ;
    buf_clk new_AGEMA_reg_buffer_4635 ( .C (clk), .D (Midori_rounds_n16), .Q (new_AGEMA_signal_8100) ) ;
    buf_clk new_AGEMA_reg_buffer_4643 ( .C (clk), .D (new_AGEMA_signal_3426), .Q (new_AGEMA_signal_8108) ) ;
    buf_clk new_AGEMA_reg_buffer_4651 ( .C (clk), .D (new_AGEMA_signal_3427), .Q (new_AGEMA_signal_8116) ) ;
    buf_clk new_AGEMA_reg_buffer_4659 ( .C (clk), .D (Midori_rounds_SelectedKey_6_), .Q (new_AGEMA_signal_8124) ) ;
    buf_clk new_AGEMA_reg_buffer_4667 ( .C (clk), .D (new_AGEMA_signal_2572), .Q (new_AGEMA_signal_8132) ) ;
    buf_clk new_AGEMA_reg_buffer_4675 ( .C (clk), .D (new_AGEMA_signal_2573), .Q (new_AGEMA_signal_8140) ) ;
    buf_clk new_AGEMA_reg_buffer_4683 ( .C (clk), .D (Midori_rounds_SelectedKey_62_), .Q (new_AGEMA_signal_8148) ) ;
    buf_clk new_AGEMA_reg_buffer_4691 ( .C (clk), .D (new_AGEMA_signal_2668), .Q (new_AGEMA_signal_8156) ) ;
    buf_clk new_AGEMA_reg_buffer_4699 ( .C (clk), .D (new_AGEMA_signal_2669), .Q (new_AGEMA_signal_8164) ) ;
    buf_clk new_AGEMA_reg_buffer_4707 ( .C (clk), .D (Midori_rounds_n15), .Q (new_AGEMA_signal_8172) ) ;
    buf_clk new_AGEMA_reg_buffer_4715 ( .C (clk), .D (new_AGEMA_signal_3536), .Q (new_AGEMA_signal_8180) ) ;
    buf_clk new_AGEMA_reg_buffer_4723 ( .C (clk), .D (new_AGEMA_signal_3537), .Q (new_AGEMA_signal_8188) ) ;
    buf_clk new_AGEMA_reg_buffer_4731 ( .C (clk), .D (Midori_rounds_SelectedKey_58_), .Q (new_AGEMA_signal_8196) ) ;
    buf_clk new_AGEMA_reg_buffer_4739 ( .C (clk), .D (new_AGEMA_signal_2660), .Q (new_AGEMA_signal_8204) ) ;
    buf_clk new_AGEMA_reg_buffer_4747 ( .C (clk), .D (new_AGEMA_signal_2661), .Q (new_AGEMA_signal_8212) ) ;
    buf_clk new_AGEMA_reg_buffer_4755 ( .C (clk), .D (Midori_rounds_n14), .Q (new_AGEMA_signal_8220) ) ;
    buf_clk new_AGEMA_reg_buffer_4763 ( .C (clk), .D (new_AGEMA_signal_3538), .Q (new_AGEMA_signal_8228) ) ;
    buf_clk new_AGEMA_reg_buffer_4771 ( .C (clk), .D (new_AGEMA_signal_3539), .Q (new_AGEMA_signal_8236) ) ;
    buf_clk new_AGEMA_reg_buffer_4779 ( .C (clk), .D (Midori_rounds_SelectedKey_54_), .Q (new_AGEMA_signal_8244) ) ;
    buf_clk new_AGEMA_reg_buffer_4787 ( .C (clk), .D (new_AGEMA_signal_2652), .Q (new_AGEMA_signal_8252) ) ;
    buf_clk new_AGEMA_reg_buffer_4795 ( .C (clk), .D (new_AGEMA_signal_2653), .Q (new_AGEMA_signal_8260) ) ;
    buf_clk new_AGEMA_reg_buffer_4803 ( .C (clk), .D (Midori_rounds_n13), .Q (new_AGEMA_signal_8268) ) ;
    buf_clk new_AGEMA_reg_buffer_4811 ( .C (clk), .D (new_AGEMA_signal_3540), .Q (new_AGEMA_signal_8276) ) ;
    buf_clk new_AGEMA_reg_buffer_4819 ( .C (clk), .D (new_AGEMA_signal_3541), .Q (new_AGEMA_signal_8284) ) ;
    buf_clk new_AGEMA_reg_buffer_4827 ( .C (clk), .D (Midori_rounds_SelectedKey_50_), .Q (new_AGEMA_signal_8292) ) ;
    buf_clk new_AGEMA_reg_buffer_4835 ( .C (clk), .D (new_AGEMA_signal_2644), .Q (new_AGEMA_signal_8300) ) ;
    buf_clk new_AGEMA_reg_buffer_4843 ( .C (clk), .D (new_AGEMA_signal_2645), .Q (new_AGEMA_signal_8308) ) ;
    buf_clk new_AGEMA_reg_buffer_4851 ( .C (clk), .D (Midori_rounds_n12), .Q (new_AGEMA_signal_8316) ) ;
    buf_clk new_AGEMA_reg_buffer_4859 ( .C (clk), .D (new_AGEMA_signal_3542), .Q (new_AGEMA_signal_8324) ) ;
    buf_clk new_AGEMA_reg_buffer_4867 ( .C (clk), .D (new_AGEMA_signal_3543), .Q (new_AGEMA_signal_8332) ) ;
    buf_clk new_AGEMA_reg_buffer_4875 ( .C (clk), .D (Midori_rounds_n11), .Q (new_AGEMA_signal_8340) ) ;
    buf_clk new_AGEMA_reg_buffer_4883 ( .C (clk), .D (new_AGEMA_signal_3780), .Q (new_AGEMA_signal_8348) ) ;
    buf_clk new_AGEMA_reg_buffer_4891 ( .C (clk), .D (new_AGEMA_signal_3781), .Q (new_AGEMA_signal_8356) ) ;
    buf_clk new_AGEMA_reg_buffer_4899 ( .C (clk), .D (Midori_rounds_SelectedKey_46_), .Q (new_AGEMA_signal_8364) ) ;
    buf_clk new_AGEMA_reg_buffer_4907 ( .C (clk), .D (new_AGEMA_signal_2636), .Q (new_AGEMA_signal_8372) ) ;
    buf_clk new_AGEMA_reg_buffer_4915 ( .C (clk), .D (new_AGEMA_signal_2637), .Q (new_AGEMA_signal_8380) ) ;
    buf_clk new_AGEMA_reg_buffer_4923 ( .C (clk), .D (Midori_rounds_n10), .Q (new_AGEMA_signal_8388) ) ;
    buf_clk new_AGEMA_reg_buffer_4931 ( .C (clk), .D (new_AGEMA_signal_3464), .Q (new_AGEMA_signal_8396) ) ;
    buf_clk new_AGEMA_reg_buffer_4939 ( .C (clk), .D (new_AGEMA_signal_3465), .Q (new_AGEMA_signal_8404) ) ;
    buf_clk new_AGEMA_reg_buffer_4947 ( .C (clk), .D (Midori_rounds_SelectedKey_42_), .Q (new_AGEMA_signal_8412) ) ;
    buf_clk new_AGEMA_reg_buffer_4955 ( .C (clk), .D (new_AGEMA_signal_2628), .Q (new_AGEMA_signal_8420) ) ;
    buf_clk new_AGEMA_reg_buffer_4963 ( .C (clk), .D (new_AGEMA_signal_2629), .Q (new_AGEMA_signal_8428) ) ;
    buf_clk new_AGEMA_reg_buffer_4971 ( .C (clk), .D (Midori_rounds_n9), .Q (new_AGEMA_signal_8436) ) ;
    buf_clk new_AGEMA_reg_buffer_4979 ( .C (clk), .D (new_AGEMA_signal_3544), .Q (new_AGEMA_signal_8444) ) ;
    buf_clk new_AGEMA_reg_buffer_4987 ( .C (clk), .D (new_AGEMA_signal_3545), .Q (new_AGEMA_signal_8452) ) ;
    buf_clk new_AGEMA_reg_buffer_4995 ( .C (clk), .D (Midori_rounds_SelectedKey_38_), .Q (new_AGEMA_signal_8460) ) ;
    buf_clk new_AGEMA_reg_buffer_5003 ( .C (clk), .D (new_AGEMA_signal_2620), .Q (new_AGEMA_signal_8468) ) ;
    buf_clk new_AGEMA_reg_buffer_5011 ( .C (clk), .D (new_AGEMA_signal_2621), .Q (new_AGEMA_signal_8476) ) ;
    buf_clk new_AGEMA_reg_buffer_5019 ( .C (clk), .D (Midori_rounds_n8), .Q (new_AGEMA_signal_8484) ) ;
    buf_clk new_AGEMA_reg_buffer_5027 ( .C (clk), .D (new_AGEMA_signal_3480), .Q (new_AGEMA_signal_8492) ) ;
    buf_clk new_AGEMA_reg_buffer_5035 ( .C (clk), .D (new_AGEMA_signal_3481), .Q (new_AGEMA_signal_8500) ) ;
    buf_clk new_AGEMA_reg_buffer_5043 ( .C (clk), .D (Midori_rounds_SelectedKey_34_), .Q (new_AGEMA_signal_8508) ) ;
    buf_clk new_AGEMA_reg_buffer_5051 ( .C (clk), .D (new_AGEMA_signal_2612), .Q (new_AGEMA_signal_8516) ) ;
    buf_clk new_AGEMA_reg_buffer_5059 ( .C (clk), .D (new_AGEMA_signal_2613), .Q (new_AGEMA_signal_8524) ) ;
    buf_clk new_AGEMA_reg_buffer_5067 ( .C (clk), .D (Midori_rounds_n7), .Q (new_AGEMA_signal_8532) ) ;
    buf_clk new_AGEMA_reg_buffer_5075 ( .C (clk), .D (new_AGEMA_signal_3546), .Q (new_AGEMA_signal_8540) ) ;
    buf_clk new_AGEMA_reg_buffer_5083 ( .C (clk), .D (new_AGEMA_signal_3547), .Q (new_AGEMA_signal_8548) ) ;
    buf_clk new_AGEMA_reg_buffer_5091 ( .C (clk), .D (Midori_rounds_SelectedKey_30_), .Q (new_AGEMA_signal_8556) ) ;
    buf_clk new_AGEMA_reg_buffer_5099 ( .C (clk), .D (new_AGEMA_signal_2604), .Q (new_AGEMA_signal_8564) ) ;
    buf_clk new_AGEMA_reg_buffer_5107 ( .C (clk), .D (new_AGEMA_signal_2605), .Q (new_AGEMA_signal_8572) ) ;
    buf_clk new_AGEMA_reg_buffer_5115 ( .C (clk), .D (Midori_rounds_SelectedKey_2_), .Q (new_AGEMA_signal_8580) ) ;
    buf_clk new_AGEMA_reg_buffer_5123 ( .C (clk), .D (new_AGEMA_signal_1844), .Q (new_AGEMA_signal_8588) ) ;
    buf_clk new_AGEMA_reg_buffer_5131 ( .C (clk), .D (new_AGEMA_signal_1845), .Q (new_AGEMA_signal_8596) ) ;
    buf_clk new_AGEMA_reg_buffer_5139 ( .C (clk), .D (Midori_rounds_n6), .Q (new_AGEMA_signal_8604) ) ;
    buf_clk new_AGEMA_reg_buffer_5147 ( .C (clk), .D (new_AGEMA_signal_3672), .Q (new_AGEMA_signal_8612) ) ;
    buf_clk new_AGEMA_reg_buffer_5155 ( .C (clk), .D (new_AGEMA_signal_3673), .Q (new_AGEMA_signal_8620) ) ;
    buf_clk new_AGEMA_reg_buffer_5163 ( .C (clk), .D (Midori_rounds_SelectedKey_26_), .Q (new_AGEMA_signal_8628) ) ;
    buf_clk new_AGEMA_reg_buffer_5171 ( .C (clk), .D (new_AGEMA_signal_1864), .Q (new_AGEMA_signal_8636) ) ;
    buf_clk new_AGEMA_reg_buffer_5179 ( .C (clk), .D (new_AGEMA_signal_1865), .Q (new_AGEMA_signal_8644) ) ;
    buf_clk new_AGEMA_reg_buffer_5187 ( .C (clk), .D (Midori_rounds_n5), .Q (new_AGEMA_signal_8652) ) ;
    buf_clk new_AGEMA_reg_buffer_5195 ( .C (clk), .D (new_AGEMA_signal_3548), .Q (new_AGEMA_signal_8660) ) ;
    buf_clk new_AGEMA_reg_buffer_5203 ( .C (clk), .D (new_AGEMA_signal_3549), .Q (new_AGEMA_signal_8668) ) ;
    buf_clk new_AGEMA_reg_buffer_5211 ( .C (clk), .D (Midori_rounds_SelectedKey_22_), .Q (new_AGEMA_signal_8676) ) ;
    buf_clk new_AGEMA_reg_buffer_5219 ( .C (clk), .D (new_AGEMA_signal_2590), .Q (new_AGEMA_signal_8684) ) ;
    buf_clk new_AGEMA_reg_buffer_5227 ( .C (clk), .D (new_AGEMA_signal_2591), .Q (new_AGEMA_signal_8692) ) ;
    buf_clk new_AGEMA_reg_buffer_5235 ( .C (clk), .D (Midori_rounds_n4), .Q (new_AGEMA_signal_8700) ) ;
    buf_clk new_AGEMA_reg_buffer_5243 ( .C (clk), .D (new_AGEMA_signal_3508), .Q (new_AGEMA_signal_8708) ) ;
    buf_clk new_AGEMA_reg_buffer_5251 ( .C (clk), .D (new_AGEMA_signal_3509), .Q (new_AGEMA_signal_8716) ) ;
    buf_clk new_AGEMA_reg_buffer_5259 ( .C (clk), .D (Midori_rounds_SelectedKey_18_), .Q (new_AGEMA_signal_8724) ) ;
    buf_clk new_AGEMA_reg_buffer_5267 ( .C (clk), .D (new_AGEMA_signal_2582), .Q (new_AGEMA_signal_8732) ) ;
    buf_clk new_AGEMA_reg_buffer_5275 ( .C (clk), .D (new_AGEMA_signal_2583), .Q (new_AGEMA_signal_8740) ) ;
    buf_clk new_AGEMA_reg_buffer_5283 ( .C (clk), .D (Midori_rounds_n3), .Q (new_AGEMA_signal_8748) ) ;
    buf_clk new_AGEMA_reg_buffer_5291 ( .C (clk), .D (new_AGEMA_signal_3550), .Q (new_AGEMA_signal_8756) ) ;
    buf_clk new_AGEMA_reg_buffer_5299 ( .C (clk), .D (new_AGEMA_signal_3551), .Q (new_AGEMA_signal_8764) ) ;
    buf_clk new_AGEMA_reg_buffer_5307 ( .C (clk), .D (Midori_rounds_SelectedKey_14_), .Q (new_AGEMA_signal_8772) ) ;
    buf_clk new_AGEMA_reg_buffer_5315 ( .C (clk), .D (new_AGEMA_signal_1860), .Q (new_AGEMA_signal_8780) ) ;
    buf_clk new_AGEMA_reg_buffer_5323 ( .C (clk), .D (new_AGEMA_signal_1861), .Q (new_AGEMA_signal_8788) ) ;
    buf_clk new_AGEMA_reg_buffer_5331 ( .C (clk), .D (Midori_rounds_n2), .Q (new_AGEMA_signal_8796) ) ;
    buf_clk new_AGEMA_reg_buffer_5339 ( .C (clk), .D (new_AGEMA_signal_3552), .Q (new_AGEMA_signal_8804) ) ;
    buf_clk new_AGEMA_reg_buffer_5347 ( .C (clk), .D (new_AGEMA_signal_3553), .Q (new_AGEMA_signal_8812) ) ;
    buf_clk new_AGEMA_reg_buffer_5355 ( .C (clk), .D (Midori_rounds_SelectedKey_10_), .Q (new_AGEMA_signal_8820) ) ;
    buf_clk new_AGEMA_reg_buffer_5363 ( .C (clk), .D (new_AGEMA_signal_1854), .Q (new_AGEMA_signal_8828) ) ;
    buf_clk new_AGEMA_reg_buffer_5371 ( .C (clk), .D (new_AGEMA_signal_1855), .Q (new_AGEMA_signal_8836) ) ;
    buf_clk new_AGEMA_reg_buffer_5379 ( .C (clk), .D (Midori_rounds_n1), .Q (new_AGEMA_signal_8844) ) ;
    buf_clk new_AGEMA_reg_buffer_5387 ( .C (clk), .D (new_AGEMA_signal_3554), .Q (new_AGEMA_signal_8852) ) ;
    buf_clk new_AGEMA_reg_buffer_5395 ( .C (clk), .D (new_AGEMA_signal_3555), .Q (new_AGEMA_signal_8860) ) ;
    buf_clk new_AGEMA_reg_buffer_5405 ( .C (clk), .D (Midori_add_Result_Start[0]), .Q (new_AGEMA_signal_8870) ) ;
    buf_clk new_AGEMA_reg_buffer_5413 ( .C (clk), .D (new_AGEMA_signal_2376), .Q (new_AGEMA_signal_8878) ) ;
    buf_clk new_AGEMA_reg_buffer_5421 ( .C (clk), .D (new_AGEMA_signal_2377), .Q (new_AGEMA_signal_8886) ) ;
    buf_clk new_AGEMA_reg_buffer_5429 ( .C (clk), .D (Midori_add_Result_Start[2]), .Q (new_AGEMA_signal_8894) ) ;
    buf_clk new_AGEMA_reg_buffer_5437 ( .C (clk), .D (new_AGEMA_signal_2288), .Q (new_AGEMA_signal_8902) ) ;
    buf_clk new_AGEMA_reg_buffer_5445 ( .C (clk), .D (new_AGEMA_signal_2289), .Q (new_AGEMA_signal_8910) ) ;
    buf_clk new_AGEMA_reg_buffer_5453 ( .C (clk), .D (Midori_add_Result_Start[4]), .Q (new_AGEMA_signal_8918) ) ;
    buf_clk new_AGEMA_reg_buffer_5461 ( .C (clk), .D (new_AGEMA_signal_2200), .Q (new_AGEMA_signal_8926) ) ;
    buf_clk new_AGEMA_reg_buffer_5469 ( .C (clk), .D (new_AGEMA_signal_2201), .Q (new_AGEMA_signal_8934) ) ;
    buf_clk new_AGEMA_reg_buffer_5477 ( .C (clk), .D (Midori_add_Result_Start[6]), .Q (new_AGEMA_signal_8942) ) ;
    buf_clk new_AGEMA_reg_buffer_5485 ( .C (clk), .D (new_AGEMA_signal_2136), .Q (new_AGEMA_signal_8950) ) ;
    buf_clk new_AGEMA_reg_buffer_5493 ( .C (clk), .D (new_AGEMA_signal_2137), .Q (new_AGEMA_signal_8958) ) ;
    buf_clk new_AGEMA_reg_buffer_5501 ( .C (clk), .D (Midori_add_Result_Start[8]), .Q (new_AGEMA_signal_8966) ) ;
    buf_clk new_AGEMA_reg_buffer_5509 ( .C (clk), .D (new_AGEMA_signal_2128), .Q (new_AGEMA_signal_8974) ) ;
    buf_clk new_AGEMA_reg_buffer_5517 ( .C (clk), .D (new_AGEMA_signal_2129), .Q (new_AGEMA_signal_8982) ) ;
    buf_clk new_AGEMA_reg_buffer_5525 ( .C (clk), .D (Midori_add_Result_Start[10]), .Q (new_AGEMA_signal_8990) ) ;
    buf_clk new_AGEMA_reg_buffer_5533 ( .C (clk), .D (new_AGEMA_signal_2372), .Q (new_AGEMA_signal_8998) ) ;
    buf_clk new_AGEMA_reg_buffer_5541 ( .C (clk), .D (new_AGEMA_signal_2373), .Q (new_AGEMA_signal_9006) ) ;
    buf_clk new_AGEMA_reg_buffer_5549 ( .C (clk), .D (Midori_add_Result_Start[12]), .Q (new_AGEMA_signal_9014) ) ;
    buf_clk new_AGEMA_reg_buffer_5557 ( .C (clk), .D (new_AGEMA_signal_2364), .Q (new_AGEMA_signal_9022) ) ;
    buf_clk new_AGEMA_reg_buffer_5565 ( .C (clk), .D (new_AGEMA_signal_2365), .Q (new_AGEMA_signal_9030) ) ;
    buf_clk new_AGEMA_reg_buffer_5573 ( .C (clk), .D (Midori_add_Result_Start[14]), .Q (new_AGEMA_signal_9038) ) ;
    buf_clk new_AGEMA_reg_buffer_5581 ( .C (clk), .D (new_AGEMA_signal_2356), .Q (new_AGEMA_signal_9046) ) ;
    buf_clk new_AGEMA_reg_buffer_5589 ( .C (clk), .D (new_AGEMA_signal_2357), .Q (new_AGEMA_signal_9054) ) ;
    buf_clk new_AGEMA_reg_buffer_5597 ( .C (clk), .D (Midori_add_Result_Start[16]), .Q (new_AGEMA_signal_9062) ) ;
    buf_clk new_AGEMA_reg_buffer_5605 ( .C (clk), .D (new_AGEMA_signal_2348), .Q (new_AGEMA_signal_9070) ) ;
    buf_clk new_AGEMA_reg_buffer_5613 ( .C (clk), .D (new_AGEMA_signal_2349), .Q (new_AGEMA_signal_9078) ) ;
    buf_clk new_AGEMA_reg_buffer_5621 ( .C (clk), .D (Midori_add_Result_Start[18]), .Q (new_AGEMA_signal_9086) ) ;
    buf_clk new_AGEMA_reg_buffer_5629 ( .C (clk), .D (new_AGEMA_signal_2340), .Q (new_AGEMA_signal_9094) ) ;
    buf_clk new_AGEMA_reg_buffer_5637 ( .C (clk), .D (new_AGEMA_signal_2341), .Q (new_AGEMA_signal_9102) ) ;
    buf_clk new_AGEMA_reg_buffer_5645 ( .C (clk), .D (Midori_add_Result_Start[20]), .Q (new_AGEMA_signal_9110) ) ;
    buf_clk new_AGEMA_reg_buffer_5653 ( .C (clk), .D (new_AGEMA_signal_2328), .Q (new_AGEMA_signal_9118) ) ;
    buf_clk new_AGEMA_reg_buffer_5661 ( .C (clk), .D (new_AGEMA_signal_2329), .Q (new_AGEMA_signal_9126) ) ;
    buf_clk new_AGEMA_reg_buffer_5669 ( .C (clk), .D (Midori_add_Result_Start[22]), .Q (new_AGEMA_signal_9134) ) ;
    buf_clk new_AGEMA_reg_buffer_5677 ( .C (clk), .D (new_AGEMA_signal_2320), .Q (new_AGEMA_signal_9142) ) ;
    buf_clk new_AGEMA_reg_buffer_5685 ( .C (clk), .D (new_AGEMA_signal_2321), .Q (new_AGEMA_signal_9150) ) ;
    buf_clk new_AGEMA_reg_buffer_5693 ( .C (clk), .D (Midori_add_Result_Start[24]), .Q (new_AGEMA_signal_9158) ) ;
    buf_clk new_AGEMA_reg_buffer_5701 ( .C (clk), .D (new_AGEMA_signal_2312), .Q (new_AGEMA_signal_9166) ) ;
    buf_clk new_AGEMA_reg_buffer_5709 ( .C (clk), .D (new_AGEMA_signal_2313), .Q (new_AGEMA_signal_9174) ) ;
    buf_clk new_AGEMA_reg_buffer_5717 ( .C (clk), .D (Midori_add_Result_Start[26]), .Q (new_AGEMA_signal_9182) ) ;
    buf_clk new_AGEMA_reg_buffer_5725 ( .C (clk), .D (new_AGEMA_signal_2304), .Q (new_AGEMA_signal_9190) ) ;
    buf_clk new_AGEMA_reg_buffer_5733 ( .C (clk), .D (new_AGEMA_signal_2305), .Q (new_AGEMA_signal_9198) ) ;
    buf_clk new_AGEMA_reg_buffer_5741 ( .C (clk), .D (Midori_add_Result_Start[28]), .Q (new_AGEMA_signal_9206) ) ;
    buf_clk new_AGEMA_reg_buffer_5749 ( .C (clk), .D (new_AGEMA_signal_2296), .Q (new_AGEMA_signal_9214) ) ;
    buf_clk new_AGEMA_reg_buffer_5757 ( .C (clk), .D (new_AGEMA_signal_2297), .Q (new_AGEMA_signal_9222) ) ;
    buf_clk new_AGEMA_reg_buffer_5765 ( .C (clk), .D (Midori_add_Result_Start[30]), .Q (new_AGEMA_signal_9230) ) ;
    buf_clk new_AGEMA_reg_buffer_5773 ( .C (clk), .D (new_AGEMA_signal_2284), .Q (new_AGEMA_signal_9238) ) ;
    buf_clk new_AGEMA_reg_buffer_5781 ( .C (clk), .D (new_AGEMA_signal_2285), .Q (new_AGEMA_signal_9246) ) ;
    buf_clk new_AGEMA_reg_buffer_5789 ( .C (clk), .D (Midori_add_Result_Start[32]), .Q (new_AGEMA_signal_9254) ) ;
    buf_clk new_AGEMA_reg_buffer_5797 ( .C (clk), .D (new_AGEMA_signal_2276), .Q (new_AGEMA_signal_9262) ) ;
    buf_clk new_AGEMA_reg_buffer_5805 ( .C (clk), .D (new_AGEMA_signal_2277), .Q (new_AGEMA_signal_9270) ) ;
    buf_clk new_AGEMA_reg_buffer_5813 ( .C (clk), .D (Midori_add_Result_Start[34]), .Q (new_AGEMA_signal_9278) ) ;
    buf_clk new_AGEMA_reg_buffer_5821 ( .C (clk), .D (new_AGEMA_signal_2268), .Q (new_AGEMA_signal_9286) ) ;
    buf_clk new_AGEMA_reg_buffer_5829 ( .C (clk), .D (new_AGEMA_signal_2269), .Q (new_AGEMA_signal_9294) ) ;
    buf_clk new_AGEMA_reg_buffer_5837 ( .C (clk), .D (Midori_add_Result_Start[36]), .Q (new_AGEMA_signal_9302) ) ;
    buf_clk new_AGEMA_reg_buffer_5845 ( .C (clk), .D (new_AGEMA_signal_2260), .Q (new_AGEMA_signal_9310) ) ;
    buf_clk new_AGEMA_reg_buffer_5853 ( .C (clk), .D (new_AGEMA_signal_2261), .Q (new_AGEMA_signal_9318) ) ;
    buf_clk new_AGEMA_reg_buffer_5861 ( .C (clk), .D (Midori_add_Result_Start[38]), .Q (new_AGEMA_signal_9326) ) ;
    buf_clk new_AGEMA_reg_buffer_5869 ( .C (clk), .D (new_AGEMA_signal_2252), .Q (new_AGEMA_signal_9334) ) ;
    buf_clk new_AGEMA_reg_buffer_5877 ( .C (clk), .D (new_AGEMA_signal_2253), .Q (new_AGEMA_signal_9342) ) ;
    buf_clk new_AGEMA_reg_buffer_5885 ( .C (clk), .D (Midori_add_Result_Start[40]), .Q (new_AGEMA_signal_9350) ) ;
    buf_clk new_AGEMA_reg_buffer_5893 ( .C (clk), .D (new_AGEMA_signal_2240), .Q (new_AGEMA_signal_9358) ) ;
    buf_clk new_AGEMA_reg_buffer_5901 ( .C (clk), .D (new_AGEMA_signal_2241), .Q (new_AGEMA_signal_9366) ) ;
    buf_clk new_AGEMA_reg_buffer_5909 ( .C (clk), .D (Midori_add_Result_Start[42]), .Q (new_AGEMA_signal_9374) ) ;
    buf_clk new_AGEMA_reg_buffer_5917 ( .C (clk), .D (new_AGEMA_signal_2232), .Q (new_AGEMA_signal_9382) ) ;
    buf_clk new_AGEMA_reg_buffer_5925 ( .C (clk), .D (new_AGEMA_signal_2233), .Q (new_AGEMA_signal_9390) ) ;
    buf_clk new_AGEMA_reg_buffer_5933 ( .C (clk), .D (Midori_add_Result_Start[44]), .Q (new_AGEMA_signal_9398) ) ;
    buf_clk new_AGEMA_reg_buffer_5941 ( .C (clk), .D (new_AGEMA_signal_2224), .Q (new_AGEMA_signal_9406) ) ;
    buf_clk new_AGEMA_reg_buffer_5949 ( .C (clk), .D (new_AGEMA_signal_2225), .Q (new_AGEMA_signal_9414) ) ;
    buf_clk new_AGEMA_reg_buffer_5957 ( .C (clk), .D (Midori_add_Result_Start[46]), .Q (new_AGEMA_signal_9422) ) ;
    buf_clk new_AGEMA_reg_buffer_5965 ( .C (clk), .D (new_AGEMA_signal_2216), .Q (new_AGEMA_signal_9430) ) ;
    buf_clk new_AGEMA_reg_buffer_5973 ( .C (clk), .D (new_AGEMA_signal_2217), .Q (new_AGEMA_signal_9438) ) ;
    buf_clk new_AGEMA_reg_buffer_5981 ( .C (clk), .D (Midori_add_Result_Start[48]), .Q (new_AGEMA_signal_9446) ) ;
    buf_clk new_AGEMA_reg_buffer_5989 ( .C (clk), .D (new_AGEMA_signal_2208), .Q (new_AGEMA_signal_9454) ) ;
    buf_clk new_AGEMA_reg_buffer_5997 ( .C (clk), .D (new_AGEMA_signal_2209), .Q (new_AGEMA_signal_9462) ) ;
    buf_clk new_AGEMA_reg_buffer_6005 ( .C (clk), .D (Midori_add_Result_Start[50]), .Q (new_AGEMA_signal_9470) ) ;
    buf_clk new_AGEMA_reg_buffer_6013 ( .C (clk), .D (new_AGEMA_signal_2196), .Q (new_AGEMA_signal_9478) ) ;
    buf_clk new_AGEMA_reg_buffer_6021 ( .C (clk), .D (new_AGEMA_signal_2197), .Q (new_AGEMA_signal_9486) ) ;
    buf_clk new_AGEMA_reg_buffer_6029 ( .C (clk), .D (Midori_add_Result_Start[52]), .Q (new_AGEMA_signal_9494) ) ;
    buf_clk new_AGEMA_reg_buffer_6037 ( .C (clk), .D (new_AGEMA_signal_2188), .Q (new_AGEMA_signal_9502) ) ;
    buf_clk new_AGEMA_reg_buffer_6045 ( .C (clk), .D (new_AGEMA_signal_2189), .Q (new_AGEMA_signal_9510) ) ;
    buf_clk new_AGEMA_reg_buffer_6053 ( .C (clk), .D (Midori_add_Result_Start[54]), .Q (new_AGEMA_signal_9518) ) ;
    buf_clk new_AGEMA_reg_buffer_6061 ( .C (clk), .D (new_AGEMA_signal_2180), .Q (new_AGEMA_signal_9526) ) ;
    buf_clk new_AGEMA_reg_buffer_6069 ( .C (clk), .D (new_AGEMA_signal_2181), .Q (new_AGEMA_signal_9534) ) ;
    buf_clk new_AGEMA_reg_buffer_6077 ( .C (clk), .D (Midori_add_Result_Start[56]), .Q (new_AGEMA_signal_9542) ) ;
    buf_clk new_AGEMA_reg_buffer_6085 ( .C (clk), .D (new_AGEMA_signal_2172), .Q (new_AGEMA_signal_9550) ) ;
    buf_clk new_AGEMA_reg_buffer_6093 ( .C (clk), .D (new_AGEMA_signal_2173), .Q (new_AGEMA_signal_9558) ) ;
    buf_clk new_AGEMA_reg_buffer_6101 ( .C (clk), .D (Midori_add_Result_Start[58]), .Q (new_AGEMA_signal_9566) ) ;
    buf_clk new_AGEMA_reg_buffer_6109 ( .C (clk), .D (new_AGEMA_signal_2164), .Q (new_AGEMA_signal_9574) ) ;
    buf_clk new_AGEMA_reg_buffer_6117 ( .C (clk), .D (new_AGEMA_signal_2165), .Q (new_AGEMA_signal_9582) ) ;
    buf_clk new_AGEMA_reg_buffer_6125 ( .C (clk), .D (Midori_add_Result_Start[60]), .Q (new_AGEMA_signal_9590) ) ;
    buf_clk new_AGEMA_reg_buffer_6133 ( .C (clk), .D (new_AGEMA_signal_2152), .Q (new_AGEMA_signal_9598) ) ;
    buf_clk new_AGEMA_reg_buffer_6141 ( .C (clk), .D (new_AGEMA_signal_2153), .Q (new_AGEMA_signal_9606) ) ;
    buf_clk new_AGEMA_reg_buffer_6149 ( .C (clk), .D (Midori_add_Result_Start[62]), .Q (new_AGEMA_signal_9614) ) ;
    buf_clk new_AGEMA_reg_buffer_6157 ( .C (clk), .D (new_AGEMA_signal_2144), .Q (new_AGEMA_signal_9622) ) ;
    buf_clk new_AGEMA_reg_buffer_6165 ( .C (clk), .D (new_AGEMA_signal_2145), .Q (new_AGEMA_signal_9630) ) ;
    buf_clk new_AGEMA_reg_buffer_6463 ( .C (clk), .D (controller_roundCounter_N7), .Q (new_AGEMA_signal_9928) ) ;
    buf_clk new_AGEMA_reg_buffer_6471 ( .C (clk), .D (controller_roundCounter_N8), .Q (new_AGEMA_signal_9936) ) ;
    buf_clk new_AGEMA_reg_buffer_6479 ( .C (clk), .D (controller_roundCounter_n2), .Q (new_AGEMA_signal_9944) ) ;
    buf_clk new_AGEMA_reg_buffer_6487 ( .C (clk), .D (controller_roundCounter_N10), .Q (new_AGEMA_signal_9952) ) ;

    /* cells in depth 2 */
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U14 ( .a ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, Midori_rounds_roundReg_out[0]}), .b ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, Midori_rounds_roundReg_out[3]}), .clk (clk), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_1871, new_AGEMA_signal_1870, Midori_rounds_sub_sBox_PRINCE_0_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U13 ( .a ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, Midori_rounds_sub_sBox_PRINCE_0_n8}), .b ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, Midori_rounds_sub_sBox_PRINCE_0_n7}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, Midori_rounds_sub_sBox_PRINCE_0_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U10 ( .a ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, Midori_rounds_roundReg_out[3]}), .b ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, Midori_rounds_sub_sBox_PRINCE_0_n9}), .clk (clk), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, Midori_rounds_sub_sBox_PRINCE_0_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U9 ( .a ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, Midori_rounds_roundReg_out[2]}), .b ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, Midori_rounds_sub_sBox_PRINCE_0_n8}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, Midori_rounds_sub_sBox_PRINCE_0_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U5 ( .a ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, Midori_rounds_roundReg_out[2]}), .b ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, Midori_rounds_roundReg_out[3]}), .clk (clk), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, Midori_rounds_sub_sBox_PRINCE_0_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U3 ( .a ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, Midori_rounds_sub_sBox_PRINCE_0_n9}), .b ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, Midori_rounds_sub_sBox_PRINCE_0_n8}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, Midori_rounds_sub_sBox_PRINCE_0_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U14 ( .a ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, Midori_rounds_roundReg_out[4]}), .b ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, Midori_rounds_roundReg_out[7]}), .clk (clk), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, Midori_rounds_sub_sBox_PRINCE_1_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U13 ( .a ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, Midori_rounds_sub_sBox_PRINCE_1_n8}), .b ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, Midori_rounds_sub_sBox_PRINCE_1_n7}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, Midori_rounds_sub_sBox_PRINCE_1_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U10 ( .a ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, Midori_rounds_roundReg_out[7]}), .b ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, Midori_rounds_sub_sBox_PRINCE_1_n9}), .clk (clk), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, Midori_rounds_sub_sBox_PRINCE_1_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U9 ( .a ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, Midori_rounds_roundReg_out[6]}), .b ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, Midori_rounds_sub_sBox_PRINCE_1_n8}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, Midori_rounds_sub_sBox_PRINCE_1_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U5 ( .a ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, Midori_rounds_roundReg_out[6]}), .b ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, Midori_rounds_roundReg_out[7]}), .clk (clk), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, Midori_rounds_sub_sBox_PRINCE_1_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U3 ( .a ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, Midori_rounds_sub_sBox_PRINCE_1_n9}), .b ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, Midori_rounds_sub_sBox_PRINCE_1_n8}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, Midori_rounds_sub_sBox_PRINCE_1_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U14 ( .a ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, Midori_rounds_roundReg_out[8]}), .b ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, Midori_rounds_roundReg_out[11]}), .clk (clk), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, Midori_rounds_sub_sBox_PRINCE_2_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U13 ( .a ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, Midori_rounds_sub_sBox_PRINCE_2_n8}), .b ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, Midori_rounds_sub_sBox_PRINCE_2_n7}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, Midori_rounds_sub_sBox_PRINCE_2_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U10 ( .a ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, Midori_rounds_roundReg_out[11]}), .b ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, Midori_rounds_sub_sBox_PRINCE_2_n9}), .clk (clk), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, Midori_rounds_sub_sBox_PRINCE_2_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U9 ( .a ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, Midori_rounds_roundReg_out[10]}), .b ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, Midori_rounds_sub_sBox_PRINCE_2_n8}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, Midori_rounds_sub_sBox_PRINCE_2_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U5 ( .a ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, Midori_rounds_roundReg_out[10]}), .b ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, Midori_rounds_roundReg_out[11]}), .clk (clk), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, Midori_rounds_sub_sBox_PRINCE_2_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U3 ( .a ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, Midori_rounds_sub_sBox_PRINCE_2_n9}), .b ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, Midori_rounds_sub_sBox_PRINCE_2_n8}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, Midori_rounds_sub_sBox_PRINCE_2_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U14 ( .a ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, Midori_rounds_roundReg_out[12]}), .b ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, Midori_rounds_roundReg_out[15]}), .clk (clk), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, Midori_rounds_sub_sBox_PRINCE_3_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U13 ( .a ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, Midori_rounds_sub_sBox_PRINCE_3_n8}), .b ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, Midori_rounds_sub_sBox_PRINCE_3_n7}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, Midori_rounds_sub_sBox_PRINCE_3_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U10 ( .a ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, Midori_rounds_roundReg_out[15]}), .b ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, Midori_rounds_sub_sBox_PRINCE_3_n9}), .clk (clk), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, Midori_rounds_sub_sBox_PRINCE_3_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U9 ( .a ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, Midori_rounds_roundReg_out[14]}), .b ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, Midori_rounds_sub_sBox_PRINCE_3_n8}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, Midori_rounds_sub_sBox_PRINCE_3_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U5 ( .a ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, Midori_rounds_roundReg_out[14]}), .b ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, Midori_rounds_roundReg_out[15]}), .clk (clk), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, Midori_rounds_sub_sBox_PRINCE_3_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U3 ( .a ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, Midori_rounds_sub_sBox_PRINCE_3_n9}), .b ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, Midori_rounds_sub_sBox_PRINCE_3_n8}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, Midori_rounds_sub_sBox_PRINCE_3_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U14 ( .a ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, Midori_rounds_roundReg_out[16]}), .b ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, Midori_rounds_roundReg_out[19]}), .clk (clk), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, Midori_rounds_sub_sBox_PRINCE_4_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U13 ( .a ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, Midori_rounds_sub_sBox_PRINCE_4_n8}), .b ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, Midori_rounds_sub_sBox_PRINCE_4_n7}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, Midori_rounds_sub_sBox_PRINCE_4_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U10 ( .a ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, Midori_rounds_roundReg_out[19]}), .b ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, Midori_rounds_sub_sBox_PRINCE_4_n9}), .clk (clk), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, Midori_rounds_sub_sBox_PRINCE_4_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U9 ( .a ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, Midori_rounds_roundReg_out[18]}), .b ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, Midori_rounds_sub_sBox_PRINCE_4_n8}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, Midori_rounds_sub_sBox_PRINCE_4_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U5 ( .a ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, Midori_rounds_roundReg_out[18]}), .b ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, Midori_rounds_roundReg_out[19]}), .clk (clk), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, Midori_rounds_sub_sBox_PRINCE_4_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U3 ( .a ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, Midori_rounds_sub_sBox_PRINCE_4_n9}), .b ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, Midori_rounds_sub_sBox_PRINCE_4_n8}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, Midori_rounds_sub_sBox_PRINCE_4_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U14 ( .a ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, Midori_rounds_roundReg_out[20]}), .b ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, Midori_rounds_roundReg_out[23]}), .clk (clk), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, Midori_rounds_sub_sBox_PRINCE_5_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U13 ( .a ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, Midori_rounds_sub_sBox_PRINCE_5_n8}), .b ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, Midori_rounds_sub_sBox_PRINCE_5_n7}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, Midori_rounds_sub_sBox_PRINCE_5_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U10 ( .a ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, Midori_rounds_roundReg_out[23]}), .b ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, Midori_rounds_sub_sBox_PRINCE_5_n9}), .clk (clk), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, Midori_rounds_sub_sBox_PRINCE_5_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U9 ( .a ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, Midori_rounds_roundReg_out[22]}), .b ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, Midori_rounds_sub_sBox_PRINCE_5_n8}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, Midori_rounds_sub_sBox_PRINCE_5_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U5 ( .a ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, Midori_rounds_roundReg_out[22]}), .b ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, Midori_rounds_roundReg_out[23]}), .clk (clk), .r ({Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, Midori_rounds_sub_sBox_PRINCE_5_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U3 ( .a ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, Midori_rounds_sub_sBox_PRINCE_5_n9}), .b ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, Midori_rounds_sub_sBox_PRINCE_5_n8}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105]}), .c ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, Midori_rounds_sub_sBox_PRINCE_5_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U14 ( .a ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, Midori_rounds_roundReg_out[24]}), .b ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, Midori_rounds_roundReg_out[27]}), .clk (clk), .r ({Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, Midori_rounds_sub_sBox_PRINCE_6_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U13 ( .a ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, Midori_rounds_sub_sBox_PRINCE_6_n8}), .b ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, Midori_rounds_sub_sBox_PRINCE_6_n7}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111]}), .c ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, Midori_rounds_sub_sBox_PRINCE_6_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U10 ( .a ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, Midori_rounds_roundReg_out[27]}), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, Midori_rounds_sub_sBox_PRINCE_6_n9}), .clk (clk), .r ({Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, Midori_rounds_sub_sBox_PRINCE_6_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U9 ( .a ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, Midori_rounds_roundReg_out[26]}), .b ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, Midori_rounds_sub_sBox_PRINCE_6_n8}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117]}), .c ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, Midori_rounds_sub_sBox_PRINCE_6_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U5 ( .a ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, Midori_rounds_roundReg_out[26]}), .b ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, Midori_rounds_roundReg_out[27]}), .clk (clk), .r ({Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, Midori_rounds_sub_sBox_PRINCE_6_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U3 ( .a ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, Midori_rounds_sub_sBox_PRINCE_6_n9}), .b ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, Midori_rounds_sub_sBox_PRINCE_6_n8}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123]}), .c ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, Midori_rounds_sub_sBox_PRINCE_6_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U14 ( .a ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, Midori_rounds_roundReg_out[28]}), .b ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, Midori_rounds_roundReg_out[31]}), .clk (clk), .r ({Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, Midori_rounds_sub_sBox_PRINCE_7_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U13 ( .a ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, Midori_rounds_sub_sBox_PRINCE_7_n8}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, Midori_rounds_sub_sBox_PRINCE_7_n7}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129]}), .c ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, Midori_rounds_sub_sBox_PRINCE_7_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U10 ( .a ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, Midori_rounds_roundReg_out[31]}), .b ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, Midori_rounds_sub_sBox_PRINCE_7_n9}), .clk (clk), .r ({Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, Midori_rounds_sub_sBox_PRINCE_7_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U9 ( .a ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, Midori_rounds_roundReg_out[30]}), .b ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, Midori_rounds_sub_sBox_PRINCE_7_n8}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135]}), .c ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, Midori_rounds_sub_sBox_PRINCE_7_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U5 ( .a ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, Midori_rounds_roundReg_out[30]}), .b ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, Midori_rounds_roundReg_out[31]}), .clk (clk), .r ({Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, Midori_rounds_sub_sBox_PRINCE_7_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U3 ( .a ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, Midori_rounds_sub_sBox_PRINCE_7_n9}), .b ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, Midori_rounds_sub_sBox_PRINCE_7_n8}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141]}), .c ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, Midori_rounds_sub_sBox_PRINCE_7_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U14 ( .a ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, Midori_rounds_roundReg_out[32]}), .b ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, Midori_rounds_roundReg_out[35]}), .clk (clk), .r ({Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, Midori_rounds_sub_sBox_PRINCE_8_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U13 ( .a ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, Midori_rounds_sub_sBox_PRINCE_8_n8}), .b ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, Midori_rounds_sub_sBox_PRINCE_8_n7}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147]}), .c ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, Midori_rounds_sub_sBox_PRINCE_8_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U10 ( .a ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, Midori_rounds_roundReg_out[35]}), .b ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, Midori_rounds_sub_sBox_PRINCE_8_n9}), .clk (clk), .r ({Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, Midori_rounds_sub_sBox_PRINCE_8_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U9 ( .a ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, Midori_rounds_roundReg_out[34]}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, Midori_rounds_sub_sBox_PRINCE_8_n8}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153]}), .c ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, Midori_rounds_sub_sBox_PRINCE_8_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U5 ( .a ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, Midori_rounds_roundReg_out[34]}), .b ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, Midori_rounds_roundReg_out[35]}), .clk (clk), .r ({Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, Midori_rounds_sub_sBox_PRINCE_8_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U3 ( .a ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, Midori_rounds_sub_sBox_PRINCE_8_n9}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, Midori_rounds_sub_sBox_PRINCE_8_n8}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159]}), .c ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, Midori_rounds_sub_sBox_PRINCE_8_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U14 ( .a ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, Midori_rounds_roundReg_out[36]}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, Midori_rounds_roundReg_out[39]}), .clk (clk), .r ({Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, Midori_rounds_sub_sBox_PRINCE_9_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U13 ( .a ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, Midori_rounds_sub_sBox_PRINCE_9_n8}), .b ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, Midori_rounds_sub_sBox_PRINCE_9_n7}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165]}), .c ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, Midori_rounds_sub_sBox_PRINCE_9_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U10 ( .a ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, Midori_rounds_roundReg_out[39]}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, Midori_rounds_sub_sBox_PRINCE_9_n9}), .clk (clk), .r ({Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, Midori_rounds_sub_sBox_PRINCE_9_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U9 ( .a ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, Midori_rounds_roundReg_out[38]}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, Midori_rounds_sub_sBox_PRINCE_9_n8}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171]}), .c ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, Midori_rounds_sub_sBox_PRINCE_9_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U5 ( .a ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, Midori_rounds_roundReg_out[38]}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, Midori_rounds_roundReg_out[39]}), .clk (clk), .r ({Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, Midori_rounds_sub_sBox_PRINCE_9_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U3 ( .a ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, Midori_rounds_sub_sBox_PRINCE_9_n9}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, Midori_rounds_sub_sBox_PRINCE_9_n8}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177]}), .c ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, Midori_rounds_sub_sBox_PRINCE_9_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U14 ( .a ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, Midori_rounds_roundReg_out[40]}), .b ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, Midori_rounds_roundReg_out[43]}), .clk (clk), .r ({Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, Midori_rounds_sub_sBox_PRINCE_10_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U13 ( .a ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, Midori_rounds_sub_sBox_PRINCE_10_n8}), .b ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, Midori_rounds_sub_sBox_PRINCE_10_n7}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183]}), .c ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, Midori_rounds_sub_sBox_PRINCE_10_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U10 ( .a ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, Midori_rounds_roundReg_out[43]}), .b ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, Midori_rounds_sub_sBox_PRINCE_10_n9}), .clk (clk), .r ({Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, Midori_rounds_sub_sBox_PRINCE_10_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U9 ( .a ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, Midori_rounds_roundReg_out[42]}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, Midori_rounds_sub_sBox_PRINCE_10_n8}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189]}), .c ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, Midori_rounds_sub_sBox_PRINCE_10_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U5 ( .a ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, Midori_rounds_roundReg_out[42]}), .b ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, Midori_rounds_roundReg_out[43]}), .clk (clk), .r ({Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, Midori_rounds_sub_sBox_PRINCE_10_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U3 ( .a ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, Midori_rounds_sub_sBox_PRINCE_10_n9}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, Midori_rounds_sub_sBox_PRINCE_10_n8}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195]}), .c ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, Midori_rounds_sub_sBox_PRINCE_10_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U14 ( .a ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, Midori_rounds_roundReg_out[44]}), .b ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, Midori_rounds_roundReg_out[47]}), .clk (clk), .r ({Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, Midori_rounds_sub_sBox_PRINCE_11_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U13 ( .a ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, Midori_rounds_sub_sBox_PRINCE_11_n8}), .b ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, Midori_rounds_sub_sBox_PRINCE_11_n7}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201]}), .c ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, Midori_rounds_sub_sBox_PRINCE_11_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U10 ( .a ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, Midori_rounds_roundReg_out[47]}), .b ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, Midori_rounds_sub_sBox_PRINCE_11_n9}), .clk (clk), .r ({Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, Midori_rounds_sub_sBox_PRINCE_11_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U9 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, Midori_rounds_roundReg_out[46]}), .b ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, Midori_rounds_sub_sBox_PRINCE_11_n8}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207]}), .c ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, Midori_rounds_sub_sBox_PRINCE_11_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U5 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, Midori_rounds_roundReg_out[46]}), .b ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, Midori_rounds_roundReg_out[47]}), .clk (clk), .r ({Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, Midori_rounds_sub_sBox_PRINCE_11_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U3 ( .a ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, Midori_rounds_sub_sBox_PRINCE_11_n9}), .b ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, Midori_rounds_sub_sBox_PRINCE_11_n8}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213]}), .c ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, Midori_rounds_sub_sBox_PRINCE_11_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U14 ( .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, Midori_rounds_roundReg_out[48]}), .b ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, Midori_rounds_roundReg_out[51]}), .clk (clk), .r ({Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, Midori_rounds_sub_sBox_PRINCE_12_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U13 ( .a ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, Midori_rounds_sub_sBox_PRINCE_12_n8}), .b ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, Midori_rounds_sub_sBox_PRINCE_12_n7}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219]}), .c ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, Midori_rounds_sub_sBox_PRINCE_12_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U10 ( .a ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, Midori_rounds_roundReg_out[51]}), .b ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, Midori_rounds_sub_sBox_PRINCE_12_n9}), .clk (clk), .r ({Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, Midori_rounds_sub_sBox_PRINCE_12_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U9 ( .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, Midori_rounds_roundReg_out[50]}), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, Midori_rounds_sub_sBox_PRINCE_12_n8}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225]}), .c ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, Midori_rounds_sub_sBox_PRINCE_12_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U5 ( .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, Midori_rounds_roundReg_out[50]}), .b ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, Midori_rounds_roundReg_out[51]}), .clk (clk), .r ({Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, Midori_rounds_sub_sBox_PRINCE_12_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U3 ( .a ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, Midori_rounds_sub_sBox_PRINCE_12_n9}), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, Midori_rounds_sub_sBox_PRINCE_12_n8}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231]}), .c ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, Midori_rounds_sub_sBox_PRINCE_12_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U14 ( .a ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, Midori_rounds_roundReg_out[52]}), .b ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, Midori_rounds_roundReg_out[55]}), .clk (clk), .r ({Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, Midori_rounds_sub_sBox_PRINCE_13_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U13 ( .a ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, Midori_rounds_sub_sBox_PRINCE_13_n8}), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, Midori_rounds_sub_sBox_PRINCE_13_n7}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237]}), .c ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, Midori_rounds_sub_sBox_PRINCE_13_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U10 ( .a ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, Midori_rounds_roundReg_out[55]}), .b ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, Midori_rounds_sub_sBox_PRINCE_13_n9}), .clk (clk), .r ({Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, Midori_rounds_sub_sBox_PRINCE_13_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U9 ( .a ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, Midori_rounds_roundReg_out[54]}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, Midori_rounds_sub_sBox_PRINCE_13_n8}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243]}), .c ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, Midori_rounds_sub_sBox_PRINCE_13_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U5 ( .a ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, Midori_rounds_roundReg_out[54]}), .b ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, Midori_rounds_roundReg_out[55]}), .clk (clk), .r ({Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, Midori_rounds_sub_sBox_PRINCE_13_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U3 ( .a ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, Midori_rounds_sub_sBox_PRINCE_13_n9}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, Midori_rounds_sub_sBox_PRINCE_13_n8}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249]}), .c ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, Midori_rounds_sub_sBox_PRINCE_13_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U14 ( .a ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, Midori_rounds_roundReg_out[56]}), .b ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, Midori_rounds_roundReg_out[59]}), .clk (clk), .r ({Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, Midori_rounds_sub_sBox_PRINCE_14_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U13 ( .a ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, Midori_rounds_sub_sBox_PRINCE_14_n8}), .b ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, Midori_rounds_sub_sBox_PRINCE_14_n7}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255]}), .c ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, Midori_rounds_sub_sBox_PRINCE_14_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U10 ( .a ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, Midori_rounds_roundReg_out[59]}), .b ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, Midori_rounds_sub_sBox_PRINCE_14_n9}), .clk (clk), .r ({Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, Midori_rounds_sub_sBox_PRINCE_14_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U9 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, Midori_rounds_roundReg_out[58]}), .b ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, Midori_rounds_sub_sBox_PRINCE_14_n8}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261]}), .c ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, Midori_rounds_sub_sBox_PRINCE_14_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U5 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, Midori_rounds_roundReg_out[58]}), .b ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, Midori_rounds_roundReg_out[59]}), .clk (clk), .r ({Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, Midori_rounds_sub_sBox_PRINCE_14_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U3 ( .a ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, Midori_rounds_sub_sBox_PRINCE_14_n9}), .b ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, Midori_rounds_sub_sBox_PRINCE_14_n8}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267]}), .c ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, Midori_rounds_sub_sBox_PRINCE_14_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U14 ( .a ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, Midori_rounds_roundReg_out[60]}), .b ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, Midori_rounds_roundReg_out[63]}), .clk (clk), .r ({Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, Midori_rounds_sub_sBox_PRINCE_15_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U13 ( .a ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, Midori_rounds_sub_sBox_PRINCE_15_n8}), .b ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, Midori_rounds_sub_sBox_PRINCE_15_n7}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273]}), .c ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, Midori_rounds_sub_sBox_PRINCE_15_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U10 ( .a ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, Midori_rounds_roundReg_out[63]}), .b ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, Midori_rounds_sub_sBox_PRINCE_15_n9}), .clk (clk), .r ({Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, Midori_rounds_sub_sBox_PRINCE_15_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U9 ( .a ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, Midori_rounds_roundReg_out[62]}), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, Midori_rounds_sub_sBox_PRINCE_15_n8}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279]}), .c ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, Midori_rounds_sub_sBox_PRINCE_15_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U5 ( .a ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, Midori_rounds_roundReg_out[62]}), .b ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, Midori_rounds_roundReg_out[63]}), .clk (clk), .r ({Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, Midori_rounds_sub_sBox_PRINCE_15_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U3 ( .a ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, Midori_rounds_sub_sBox_PRINCE_15_n9}), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, Midori_rounds_sub_sBox_PRINCE_15_n8}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285]}), .c ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, Midori_rounds_sub_sBox_PRINCE_15_n13}) ) ;
    buf_clk new_AGEMA_reg_buffer_1320 ( .C (clk), .D (new_AGEMA_signal_4785), .Q (new_AGEMA_signal_4786) ) ;
    buf_clk new_AGEMA_reg_buffer_1456 ( .C (clk), .D (new_AGEMA_signal_4920), .Q (new_AGEMA_signal_4921) ) ;
    buf_clk new_AGEMA_reg_buffer_1458 ( .C (clk), .D (new_AGEMA_signal_4922), .Q (new_AGEMA_signal_4923) ) ;
    buf_clk new_AGEMA_reg_buffer_1460 ( .C (clk), .D (new_AGEMA_signal_4924), .Q (new_AGEMA_signal_4925) ) ;
    buf_clk new_AGEMA_reg_buffer_1462 ( .C (clk), .D (new_AGEMA_signal_4926), .Q (new_AGEMA_signal_4927) ) ;
    buf_clk new_AGEMA_reg_buffer_1464 ( .C (clk), .D (new_AGEMA_signal_4928), .Q (new_AGEMA_signal_4929) ) ;
    buf_clk new_AGEMA_reg_buffer_1466 ( .C (clk), .D (new_AGEMA_signal_4930), .Q (new_AGEMA_signal_4931) ) ;
    buf_clk new_AGEMA_reg_buffer_1468 ( .C (clk), .D (new_AGEMA_signal_4932), .Q (new_AGEMA_signal_4933) ) ;
    buf_clk new_AGEMA_reg_buffer_1470 ( .C (clk), .D (new_AGEMA_signal_4934), .Q (new_AGEMA_signal_4935) ) ;
    buf_clk new_AGEMA_reg_buffer_1472 ( .C (clk), .D (new_AGEMA_signal_4936), .Q (new_AGEMA_signal_4937) ) ;
    buf_clk new_AGEMA_reg_buffer_1474 ( .C (clk), .D (new_AGEMA_signal_4938), .Q (new_AGEMA_signal_4939) ) ;
    buf_clk new_AGEMA_reg_buffer_1476 ( .C (clk), .D (new_AGEMA_signal_4940), .Q (new_AGEMA_signal_4941) ) ;
    buf_clk new_AGEMA_reg_buffer_1478 ( .C (clk), .D (new_AGEMA_signal_4942), .Q (new_AGEMA_signal_4943) ) ;
    buf_clk new_AGEMA_reg_buffer_1480 ( .C (clk), .D (new_AGEMA_signal_4944), .Q (new_AGEMA_signal_4945) ) ;
    buf_clk new_AGEMA_reg_buffer_1482 ( .C (clk), .D (new_AGEMA_signal_4946), .Q (new_AGEMA_signal_4947) ) ;
    buf_clk new_AGEMA_reg_buffer_1484 ( .C (clk), .D (new_AGEMA_signal_4948), .Q (new_AGEMA_signal_4949) ) ;
    buf_clk new_AGEMA_reg_buffer_1486 ( .C (clk), .D (new_AGEMA_signal_4950), .Q (new_AGEMA_signal_4951) ) ;
    buf_clk new_AGEMA_reg_buffer_1488 ( .C (clk), .D (new_AGEMA_signal_4952), .Q (new_AGEMA_signal_4953) ) ;
    buf_clk new_AGEMA_reg_buffer_1490 ( .C (clk), .D (new_AGEMA_signal_4954), .Q (new_AGEMA_signal_4955) ) ;
    buf_clk new_AGEMA_reg_buffer_1492 ( .C (clk), .D (new_AGEMA_signal_4956), .Q (new_AGEMA_signal_4957) ) ;
    buf_clk new_AGEMA_reg_buffer_1494 ( .C (clk), .D (new_AGEMA_signal_4958), .Q (new_AGEMA_signal_4959) ) ;
    buf_clk new_AGEMA_reg_buffer_1496 ( .C (clk), .D (new_AGEMA_signal_4960), .Q (new_AGEMA_signal_4961) ) ;
    buf_clk new_AGEMA_reg_buffer_1498 ( .C (clk), .D (new_AGEMA_signal_4962), .Q (new_AGEMA_signal_4963) ) ;
    buf_clk new_AGEMA_reg_buffer_1500 ( .C (clk), .D (new_AGEMA_signal_4964), .Q (new_AGEMA_signal_4965) ) ;
    buf_clk new_AGEMA_reg_buffer_1502 ( .C (clk), .D (new_AGEMA_signal_4966), .Q (new_AGEMA_signal_4967) ) ;
    buf_clk new_AGEMA_reg_buffer_1504 ( .C (clk), .D (new_AGEMA_signal_4968), .Q (new_AGEMA_signal_4969) ) ;
    buf_clk new_AGEMA_reg_buffer_1506 ( .C (clk), .D (new_AGEMA_signal_4970), .Q (new_AGEMA_signal_4971) ) ;
    buf_clk new_AGEMA_reg_buffer_1508 ( .C (clk), .D (new_AGEMA_signal_4972), .Q (new_AGEMA_signal_4973) ) ;
    buf_clk new_AGEMA_reg_buffer_1510 ( .C (clk), .D (new_AGEMA_signal_4974), .Q (new_AGEMA_signal_4975) ) ;
    buf_clk new_AGEMA_reg_buffer_1512 ( .C (clk), .D (new_AGEMA_signal_4976), .Q (new_AGEMA_signal_4977) ) ;
    buf_clk new_AGEMA_reg_buffer_1514 ( .C (clk), .D (new_AGEMA_signal_4978), .Q (new_AGEMA_signal_4979) ) ;
    buf_clk new_AGEMA_reg_buffer_1516 ( .C (clk), .D (new_AGEMA_signal_4980), .Q (new_AGEMA_signal_4981) ) ;
    buf_clk new_AGEMA_reg_buffer_1518 ( .C (clk), .D (new_AGEMA_signal_4982), .Q (new_AGEMA_signal_4983) ) ;
    buf_clk new_AGEMA_reg_buffer_1520 ( .C (clk), .D (new_AGEMA_signal_4984), .Q (new_AGEMA_signal_4985) ) ;
    buf_clk new_AGEMA_reg_buffer_1522 ( .C (clk), .D (new_AGEMA_signal_4986), .Q (new_AGEMA_signal_4987) ) ;
    buf_clk new_AGEMA_reg_buffer_1524 ( .C (clk), .D (new_AGEMA_signal_4988), .Q (new_AGEMA_signal_4989) ) ;
    buf_clk new_AGEMA_reg_buffer_1526 ( .C (clk), .D (new_AGEMA_signal_4990), .Q (new_AGEMA_signal_4991) ) ;
    buf_clk new_AGEMA_reg_buffer_1528 ( .C (clk), .D (new_AGEMA_signal_4992), .Q (new_AGEMA_signal_4993) ) ;
    buf_clk new_AGEMA_reg_buffer_1530 ( .C (clk), .D (new_AGEMA_signal_4994), .Q (new_AGEMA_signal_4995) ) ;
    buf_clk new_AGEMA_reg_buffer_1532 ( .C (clk), .D (new_AGEMA_signal_4996), .Q (new_AGEMA_signal_4997) ) ;
    buf_clk new_AGEMA_reg_buffer_1534 ( .C (clk), .D (new_AGEMA_signal_4998), .Q (new_AGEMA_signal_4999) ) ;
    buf_clk new_AGEMA_reg_buffer_1536 ( .C (clk), .D (new_AGEMA_signal_5000), .Q (new_AGEMA_signal_5001) ) ;
    buf_clk new_AGEMA_reg_buffer_1538 ( .C (clk), .D (new_AGEMA_signal_5002), .Q (new_AGEMA_signal_5003) ) ;
    buf_clk new_AGEMA_reg_buffer_1540 ( .C (clk), .D (new_AGEMA_signal_5004), .Q (new_AGEMA_signal_5005) ) ;
    buf_clk new_AGEMA_reg_buffer_1542 ( .C (clk), .D (new_AGEMA_signal_5006), .Q (new_AGEMA_signal_5007) ) ;
    buf_clk new_AGEMA_reg_buffer_1544 ( .C (clk), .D (new_AGEMA_signal_5008), .Q (new_AGEMA_signal_5009) ) ;
    buf_clk new_AGEMA_reg_buffer_1546 ( .C (clk), .D (new_AGEMA_signal_5010), .Q (new_AGEMA_signal_5011) ) ;
    buf_clk new_AGEMA_reg_buffer_1548 ( .C (clk), .D (new_AGEMA_signal_5012), .Q (new_AGEMA_signal_5013) ) ;
    buf_clk new_AGEMA_reg_buffer_1550 ( .C (clk), .D (new_AGEMA_signal_5014), .Q (new_AGEMA_signal_5015) ) ;
    buf_clk new_AGEMA_reg_buffer_1552 ( .C (clk), .D (new_AGEMA_signal_5016), .Q (new_AGEMA_signal_5017) ) ;
    buf_clk new_AGEMA_reg_buffer_1554 ( .C (clk), .D (new_AGEMA_signal_5018), .Q (new_AGEMA_signal_5019) ) ;
    buf_clk new_AGEMA_reg_buffer_1556 ( .C (clk), .D (new_AGEMA_signal_5020), .Q (new_AGEMA_signal_5021) ) ;
    buf_clk new_AGEMA_reg_buffer_1558 ( .C (clk), .D (new_AGEMA_signal_5022), .Q (new_AGEMA_signal_5023) ) ;
    buf_clk new_AGEMA_reg_buffer_1560 ( .C (clk), .D (new_AGEMA_signal_5024), .Q (new_AGEMA_signal_5025) ) ;
    buf_clk new_AGEMA_reg_buffer_1562 ( .C (clk), .D (new_AGEMA_signal_5026), .Q (new_AGEMA_signal_5027) ) ;
    buf_clk new_AGEMA_reg_buffer_1564 ( .C (clk), .D (new_AGEMA_signal_5028), .Q (new_AGEMA_signal_5029) ) ;
    buf_clk new_AGEMA_reg_buffer_1566 ( .C (clk), .D (new_AGEMA_signal_5030), .Q (new_AGEMA_signal_5031) ) ;
    buf_clk new_AGEMA_reg_buffer_1568 ( .C (clk), .D (new_AGEMA_signal_5032), .Q (new_AGEMA_signal_5033) ) ;
    buf_clk new_AGEMA_reg_buffer_1570 ( .C (clk), .D (new_AGEMA_signal_5034), .Q (new_AGEMA_signal_5035) ) ;
    buf_clk new_AGEMA_reg_buffer_1572 ( .C (clk), .D (new_AGEMA_signal_5036), .Q (new_AGEMA_signal_5037) ) ;
    buf_clk new_AGEMA_reg_buffer_1574 ( .C (clk), .D (new_AGEMA_signal_5038), .Q (new_AGEMA_signal_5039) ) ;
    buf_clk new_AGEMA_reg_buffer_1576 ( .C (clk), .D (new_AGEMA_signal_5040), .Q (new_AGEMA_signal_5041) ) ;
    buf_clk new_AGEMA_reg_buffer_1578 ( .C (clk), .D (new_AGEMA_signal_5042), .Q (new_AGEMA_signal_5043) ) ;
    buf_clk new_AGEMA_reg_buffer_1580 ( .C (clk), .D (new_AGEMA_signal_5044), .Q (new_AGEMA_signal_5045) ) ;
    buf_clk new_AGEMA_reg_buffer_1582 ( .C (clk), .D (new_AGEMA_signal_5046), .Q (new_AGEMA_signal_5047) ) ;
    buf_clk new_AGEMA_reg_buffer_1584 ( .C (clk), .D (new_AGEMA_signal_5048), .Q (new_AGEMA_signal_5049) ) ;
    buf_clk new_AGEMA_reg_buffer_1586 ( .C (clk), .D (new_AGEMA_signal_5050), .Q (new_AGEMA_signal_5051) ) ;
    buf_clk new_AGEMA_reg_buffer_1588 ( .C (clk), .D (new_AGEMA_signal_5052), .Q (new_AGEMA_signal_5053) ) ;
    buf_clk new_AGEMA_reg_buffer_1590 ( .C (clk), .D (new_AGEMA_signal_5054), .Q (new_AGEMA_signal_5055) ) ;
    buf_clk new_AGEMA_reg_buffer_1592 ( .C (clk), .D (new_AGEMA_signal_5056), .Q (new_AGEMA_signal_5057) ) ;
    buf_clk new_AGEMA_reg_buffer_1594 ( .C (clk), .D (new_AGEMA_signal_5058), .Q (new_AGEMA_signal_5059) ) ;
    buf_clk new_AGEMA_reg_buffer_1596 ( .C (clk), .D (new_AGEMA_signal_5060), .Q (new_AGEMA_signal_5061) ) ;
    buf_clk new_AGEMA_reg_buffer_1598 ( .C (clk), .D (new_AGEMA_signal_5062), .Q (new_AGEMA_signal_5063) ) ;
    buf_clk new_AGEMA_reg_buffer_1600 ( .C (clk), .D (new_AGEMA_signal_5064), .Q (new_AGEMA_signal_5065) ) ;
    buf_clk new_AGEMA_reg_buffer_1602 ( .C (clk), .D (new_AGEMA_signal_5066), .Q (new_AGEMA_signal_5067) ) ;
    buf_clk new_AGEMA_reg_buffer_1604 ( .C (clk), .D (new_AGEMA_signal_5068), .Q (new_AGEMA_signal_5069) ) ;
    buf_clk new_AGEMA_reg_buffer_1606 ( .C (clk), .D (new_AGEMA_signal_5070), .Q (new_AGEMA_signal_5071) ) ;
    buf_clk new_AGEMA_reg_buffer_1608 ( .C (clk), .D (new_AGEMA_signal_5072), .Q (new_AGEMA_signal_5073) ) ;
    buf_clk new_AGEMA_reg_buffer_1610 ( .C (clk), .D (new_AGEMA_signal_5074), .Q (new_AGEMA_signal_5075) ) ;
    buf_clk new_AGEMA_reg_buffer_1612 ( .C (clk), .D (new_AGEMA_signal_5076), .Q (new_AGEMA_signal_5077) ) ;
    buf_clk new_AGEMA_reg_buffer_1614 ( .C (clk), .D (new_AGEMA_signal_5078), .Q (new_AGEMA_signal_5079) ) ;
    buf_clk new_AGEMA_reg_buffer_1616 ( .C (clk), .D (new_AGEMA_signal_5080), .Q (new_AGEMA_signal_5081) ) ;
    buf_clk new_AGEMA_reg_buffer_1618 ( .C (clk), .D (new_AGEMA_signal_5082), .Q (new_AGEMA_signal_5083) ) ;
    buf_clk new_AGEMA_reg_buffer_1620 ( .C (clk), .D (new_AGEMA_signal_5084), .Q (new_AGEMA_signal_5085) ) ;
    buf_clk new_AGEMA_reg_buffer_1622 ( .C (clk), .D (new_AGEMA_signal_5086), .Q (new_AGEMA_signal_5087) ) ;
    buf_clk new_AGEMA_reg_buffer_1624 ( .C (clk), .D (new_AGEMA_signal_5088), .Q (new_AGEMA_signal_5089) ) ;
    buf_clk new_AGEMA_reg_buffer_1626 ( .C (clk), .D (new_AGEMA_signal_5090), .Q (new_AGEMA_signal_5091) ) ;
    buf_clk new_AGEMA_reg_buffer_1628 ( .C (clk), .D (new_AGEMA_signal_5092), .Q (new_AGEMA_signal_5093) ) ;
    buf_clk new_AGEMA_reg_buffer_1630 ( .C (clk), .D (new_AGEMA_signal_5094), .Q (new_AGEMA_signal_5095) ) ;
    buf_clk new_AGEMA_reg_buffer_1632 ( .C (clk), .D (new_AGEMA_signal_5096), .Q (new_AGEMA_signal_5097) ) ;
    buf_clk new_AGEMA_reg_buffer_1634 ( .C (clk), .D (new_AGEMA_signal_5098), .Q (new_AGEMA_signal_5099) ) ;
    buf_clk new_AGEMA_reg_buffer_1636 ( .C (clk), .D (new_AGEMA_signal_5100), .Q (new_AGEMA_signal_5101) ) ;
    buf_clk new_AGEMA_reg_buffer_1638 ( .C (clk), .D (new_AGEMA_signal_5102), .Q (new_AGEMA_signal_5103) ) ;
    buf_clk new_AGEMA_reg_buffer_1640 ( .C (clk), .D (new_AGEMA_signal_5104), .Q (new_AGEMA_signal_5105) ) ;
    buf_clk new_AGEMA_reg_buffer_1642 ( .C (clk), .D (new_AGEMA_signal_5106), .Q (new_AGEMA_signal_5107) ) ;
    buf_clk new_AGEMA_reg_buffer_1644 ( .C (clk), .D (new_AGEMA_signal_5108), .Q (new_AGEMA_signal_5109) ) ;
    buf_clk new_AGEMA_reg_buffer_1646 ( .C (clk), .D (new_AGEMA_signal_5110), .Q (new_AGEMA_signal_5111) ) ;
    buf_clk new_AGEMA_reg_buffer_1648 ( .C (clk), .D (new_AGEMA_signal_5112), .Q (new_AGEMA_signal_5113) ) ;
    buf_clk new_AGEMA_reg_buffer_1650 ( .C (clk), .D (new_AGEMA_signal_5114), .Q (new_AGEMA_signal_5115) ) ;
    buf_clk new_AGEMA_reg_buffer_1652 ( .C (clk), .D (new_AGEMA_signal_5116), .Q (new_AGEMA_signal_5117) ) ;
    buf_clk new_AGEMA_reg_buffer_1654 ( .C (clk), .D (new_AGEMA_signal_5118), .Q (new_AGEMA_signal_5119) ) ;
    buf_clk new_AGEMA_reg_buffer_1656 ( .C (clk), .D (new_AGEMA_signal_5120), .Q (new_AGEMA_signal_5121) ) ;
    buf_clk new_AGEMA_reg_buffer_1658 ( .C (clk), .D (new_AGEMA_signal_5122), .Q (new_AGEMA_signal_5123) ) ;
    buf_clk new_AGEMA_reg_buffer_1660 ( .C (clk), .D (new_AGEMA_signal_5124), .Q (new_AGEMA_signal_5125) ) ;
    buf_clk new_AGEMA_reg_buffer_1662 ( .C (clk), .D (new_AGEMA_signal_5126), .Q (new_AGEMA_signal_5127) ) ;
    buf_clk new_AGEMA_reg_buffer_1664 ( .C (clk), .D (new_AGEMA_signal_5128), .Q (new_AGEMA_signal_5129) ) ;
    buf_clk new_AGEMA_reg_buffer_1666 ( .C (clk), .D (new_AGEMA_signal_5130), .Q (new_AGEMA_signal_5131) ) ;
    buf_clk new_AGEMA_reg_buffer_1668 ( .C (clk), .D (new_AGEMA_signal_5132), .Q (new_AGEMA_signal_5133) ) ;
    buf_clk new_AGEMA_reg_buffer_1670 ( .C (clk), .D (new_AGEMA_signal_5134), .Q (new_AGEMA_signal_5135) ) ;
    buf_clk new_AGEMA_reg_buffer_1672 ( .C (clk), .D (new_AGEMA_signal_5136), .Q (new_AGEMA_signal_5137) ) ;
    buf_clk new_AGEMA_reg_buffer_1674 ( .C (clk), .D (new_AGEMA_signal_5138), .Q (new_AGEMA_signal_5139) ) ;
    buf_clk new_AGEMA_reg_buffer_1676 ( .C (clk), .D (new_AGEMA_signal_5140), .Q (new_AGEMA_signal_5141) ) ;
    buf_clk new_AGEMA_reg_buffer_1678 ( .C (clk), .D (new_AGEMA_signal_5142), .Q (new_AGEMA_signal_5143) ) ;
    buf_clk new_AGEMA_reg_buffer_1680 ( .C (clk), .D (new_AGEMA_signal_5144), .Q (new_AGEMA_signal_5145) ) ;
    buf_clk new_AGEMA_reg_buffer_1682 ( .C (clk), .D (new_AGEMA_signal_5146), .Q (new_AGEMA_signal_5147) ) ;
    buf_clk new_AGEMA_reg_buffer_1684 ( .C (clk), .D (new_AGEMA_signal_5148), .Q (new_AGEMA_signal_5149) ) ;
    buf_clk new_AGEMA_reg_buffer_1686 ( .C (clk), .D (new_AGEMA_signal_5150), .Q (new_AGEMA_signal_5151) ) ;
    buf_clk new_AGEMA_reg_buffer_1688 ( .C (clk), .D (new_AGEMA_signal_5152), .Q (new_AGEMA_signal_5153) ) ;
    buf_clk new_AGEMA_reg_buffer_1690 ( .C (clk), .D (new_AGEMA_signal_5154), .Q (new_AGEMA_signal_5155) ) ;
    buf_clk new_AGEMA_reg_buffer_1692 ( .C (clk), .D (new_AGEMA_signal_5156), .Q (new_AGEMA_signal_5157) ) ;
    buf_clk new_AGEMA_reg_buffer_1694 ( .C (clk), .D (new_AGEMA_signal_5158), .Q (new_AGEMA_signal_5159) ) ;
    buf_clk new_AGEMA_reg_buffer_1696 ( .C (clk), .D (new_AGEMA_signal_5160), .Q (new_AGEMA_signal_5161) ) ;
    buf_clk new_AGEMA_reg_buffer_1698 ( .C (clk), .D (new_AGEMA_signal_5162), .Q (new_AGEMA_signal_5163) ) ;
    buf_clk new_AGEMA_reg_buffer_1700 ( .C (clk), .D (new_AGEMA_signal_5164), .Q (new_AGEMA_signal_5165) ) ;
    buf_clk new_AGEMA_reg_buffer_1702 ( .C (clk), .D (new_AGEMA_signal_5166), .Q (new_AGEMA_signal_5167) ) ;
    buf_clk new_AGEMA_reg_buffer_1704 ( .C (clk), .D (new_AGEMA_signal_5168), .Q (new_AGEMA_signal_5169) ) ;
    buf_clk new_AGEMA_reg_buffer_1706 ( .C (clk), .D (new_AGEMA_signal_5170), .Q (new_AGEMA_signal_5171) ) ;
    buf_clk new_AGEMA_reg_buffer_1708 ( .C (clk), .D (new_AGEMA_signal_5172), .Q (new_AGEMA_signal_5173) ) ;
    buf_clk new_AGEMA_reg_buffer_1710 ( .C (clk), .D (new_AGEMA_signal_5174), .Q (new_AGEMA_signal_5175) ) ;
    buf_clk new_AGEMA_reg_buffer_1712 ( .C (clk), .D (new_AGEMA_signal_5176), .Q (new_AGEMA_signal_5177) ) ;
    buf_clk new_AGEMA_reg_buffer_1714 ( .C (clk), .D (new_AGEMA_signal_5178), .Q (new_AGEMA_signal_5179) ) ;
    buf_clk new_AGEMA_reg_buffer_1716 ( .C (clk), .D (new_AGEMA_signal_5180), .Q (new_AGEMA_signal_5181) ) ;
    buf_clk new_AGEMA_reg_buffer_1718 ( .C (clk), .D (new_AGEMA_signal_5182), .Q (new_AGEMA_signal_5183) ) ;
    buf_clk new_AGEMA_reg_buffer_1720 ( .C (clk), .D (new_AGEMA_signal_5184), .Q (new_AGEMA_signal_5185) ) ;
    buf_clk new_AGEMA_reg_buffer_1722 ( .C (clk), .D (new_AGEMA_signal_5186), .Q (new_AGEMA_signal_5187) ) ;
    buf_clk new_AGEMA_reg_buffer_1724 ( .C (clk), .D (new_AGEMA_signal_5188), .Q (new_AGEMA_signal_5189) ) ;
    buf_clk new_AGEMA_reg_buffer_1726 ( .C (clk), .D (new_AGEMA_signal_5190), .Q (new_AGEMA_signal_5191) ) ;
    buf_clk new_AGEMA_reg_buffer_1728 ( .C (clk), .D (new_AGEMA_signal_5192), .Q (new_AGEMA_signal_5193) ) ;
    buf_clk new_AGEMA_reg_buffer_1730 ( .C (clk), .D (new_AGEMA_signal_5194), .Q (new_AGEMA_signal_5195) ) ;
    buf_clk new_AGEMA_reg_buffer_1732 ( .C (clk), .D (new_AGEMA_signal_5196), .Q (new_AGEMA_signal_5197) ) ;
    buf_clk new_AGEMA_reg_buffer_1734 ( .C (clk), .D (new_AGEMA_signal_5198), .Q (new_AGEMA_signal_5199) ) ;
    buf_clk new_AGEMA_reg_buffer_1736 ( .C (clk), .D (new_AGEMA_signal_5200), .Q (new_AGEMA_signal_5201) ) ;
    buf_clk new_AGEMA_reg_buffer_1738 ( .C (clk), .D (new_AGEMA_signal_5202), .Q (new_AGEMA_signal_5203) ) ;
    buf_clk new_AGEMA_reg_buffer_1740 ( .C (clk), .D (new_AGEMA_signal_5204), .Q (new_AGEMA_signal_5205) ) ;
    buf_clk new_AGEMA_reg_buffer_1742 ( .C (clk), .D (new_AGEMA_signal_5206), .Q (new_AGEMA_signal_5207) ) ;
    buf_clk new_AGEMA_reg_buffer_1744 ( .C (clk), .D (new_AGEMA_signal_5208), .Q (new_AGEMA_signal_5209) ) ;
    buf_clk new_AGEMA_reg_buffer_1746 ( .C (clk), .D (new_AGEMA_signal_5210), .Q (new_AGEMA_signal_5211) ) ;
    buf_clk new_AGEMA_reg_buffer_1748 ( .C (clk), .D (new_AGEMA_signal_5212), .Q (new_AGEMA_signal_5213) ) ;
    buf_clk new_AGEMA_reg_buffer_1750 ( .C (clk), .D (new_AGEMA_signal_5214), .Q (new_AGEMA_signal_5215) ) ;
    buf_clk new_AGEMA_reg_buffer_1752 ( .C (clk), .D (new_AGEMA_signal_5216), .Q (new_AGEMA_signal_5217) ) ;
    buf_clk new_AGEMA_reg_buffer_1754 ( .C (clk), .D (new_AGEMA_signal_5218), .Q (new_AGEMA_signal_5219) ) ;
    buf_clk new_AGEMA_reg_buffer_1756 ( .C (clk), .D (new_AGEMA_signal_5220), .Q (new_AGEMA_signal_5221) ) ;
    buf_clk new_AGEMA_reg_buffer_1758 ( .C (clk), .D (new_AGEMA_signal_5222), .Q (new_AGEMA_signal_5223) ) ;
    buf_clk new_AGEMA_reg_buffer_1760 ( .C (clk), .D (new_AGEMA_signal_5224), .Q (new_AGEMA_signal_5225) ) ;
    buf_clk new_AGEMA_reg_buffer_1762 ( .C (clk), .D (new_AGEMA_signal_5226), .Q (new_AGEMA_signal_5227) ) ;
    buf_clk new_AGEMA_reg_buffer_1764 ( .C (clk), .D (new_AGEMA_signal_5228), .Q (new_AGEMA_signal_5229) ) ;
    buf_clk new_AGEMA_reg_buffer_1766 ( .C (clk), .D (new_AGEMA_signal_5230), .Q (new_AGEMA_signal_5231) ) ;
    buf_clk new_AGEMA_reg_buffer_1768 ( .C (clk), .D (new_AGEMA_signal_5232), .Q (new_AGEMA_signal_5233) ) ;
    buf_clk new_AGEMA_reg_buffer_1770 ( .C (clk), .D (new_AGEMA_signal_5234), .Q (new_AGEMA_signal_5235) ) ;
    buf_clk new_AGEMA_reg_buffer_1772 ( .C (clk), .D (new_AGEMA_signal_5236), .Q (new_AGEMA_signal_5237) ) ;
    buf_clk new_AGEMA_reg_buffer_1774 ( .C (clk), .D (new_AGEMA_signal_5238), .Q (new_AGEMA_signal_5239) ) ;
    buf_clk new_AGEMA_reg_buffer_1776 ( .C (clk), .D (new_AGEMA_signal_5240), .Q (new_AGEMA_signal_5241) ) ;
    buf_clk new_AGEMA_reg_buffer_1778 ( .C (clk), .D (new_AGEMA_signal_5242), .Q (new_AGEMA_signal_5243) ) ;
    buf_clk new_AGEMA_reg_buffer_1780 ( .C (clk), .D (new_AGEMA_signal_5244), .Q (new_AGEMA_signal_5245) ) ;
    buf_clk new_AGEMA_reg_buffer_1782 ( .C (clk), .D (new_AGEMA_signal_5246), .Q (new_AGEMA_signal_5247) ) ;
    buf_clk new_AGEMA_reg_buffer_1784 ( .C (clk), .D (new_AGEMA_signal_5248), .Q (new_AGEMA_signal_5249) ) ;
    buf_clk new_AGEMA_reg_buffer_1786 ( .C (clk), .D (new_AGEMA_signal_5250), .Q (new_AGEMA_signal_5251) ) ;
    buf_clk new_AGEMA_reg_buffer_1788 ( .C (clk), .D (new_AGEMA_signal_5252), .Q (new_AGEMA_signal_5253) ) ;
    buf_clk new_AGEMA_reg_buffer_1790 ( .C (clk), .D (new_AGEMA_signal_5254), .Q (new_AGEMA_signal_5255) ) ;
    buf_clk new_AGEMA_reg_buffer_1792 ( .C (clk), .D (new_AGEMA_signal_5256), .Q (new_AGEMA_signal_5257) ) ;
    buf_clk new_AGEMA_reg_buffer_1794 ( .C (clk), .D (new_AGEMA_signal_5258), .Q (new_AGEMA_signal_5259) ) ;
    buf_clk new_AGEMA_reg_buffer_1796 ( .C (clk), .D (new_AGEMA_signal_5260), .Q (new_AGEMA_signal_5261) ) ;
    buf_clk new_AGEMA_reg_buffer_1798 ( .C (clk), .D (new_AGEMA_signal_5262), .Q (new_AGEMA_signal_5263) ) ;
    buf_clk new_AGEMA_reg_buffer_1800 ( .C (clk), .D (new_AGEMA_signal_5264), .Q (new_AGEMA_signal_5265) ) ;
    buf_clk new_AGEMA_reg_buffer_1802 ( .C (clk), .D (new_AGEMA_signal_5266), .Q (new_AGEMA_signal_5267) ) ;
    buf_clk new_AGEMA_reg_buffer_1804 ( .C (clk), .D (new_AGEMA_signal_5268), .Q (new_AGEMA_signal_5269) ) ;
    buf_clk new_AGEMA_reg_buffer_1806 ( .C (clk), .D (new_AGEMA_signal_5270), .Q (new_AGEMA_signal_5271) ) ;
    buf_clk new_AGEMA_reg_buffer_1808 ( .C (clk), .D (new_AGEMA_signal_5272), .Q (new_AGEMA_signal_5273) ) ;
    buf_clk new_AGEMA_reg_buffer_1810 ( .C (clk), .D (new_AGEMA_signal_5274), .Q (new_AGEMA_signal_5275) ) ;
    buf_clk new_AGEMA_reg_buffer_1812 ( .C (clk), .D (new_AGEMA_signal_5276), .Q (new_AGEMA_signal_5277) ) ;
    buf_clk new_AGEMA_reg_buffer_1814 ( .C (clk), .D (new_AGEMA_signal_5278), .Q (new_AGEMA_signal_5279) ) ;
    buf_clk new_AGEMA_reg_buffer_1816 ( .C (clk), .D (new_AGEMA_signal_5280), .Q (new_AGEMA_signal_5281) ) ;
    buf_clk new_AGEMA_reg_buffer_1818 ( .C (clk), .D (new_AGEMA_signal_5282), .Q (new_AGEMA_signal_5283) ) ;
    buf_clk new_AGEMA_reg_buffer_1820 ( .C (clk), .D (new_AGEMA_signal_5284), .Q (new_AGEMA_signal_5285) ) ;
    buf_clk new_AGEMA_reg_buffer_1822 ( .C (clk), .D (new_AGEMA_signal_5286), .Q (new_AGEMA_signal_5287) ) ;
    buf_clk new_AGEMA_reg_buffer_1824 ( .C (clk), .D (new_AGEMA_signal_5288), .Q (new_AGEMA_signal_5289) ) ;
    buf_clk new_AGEMA_reg_buffer_1826 ( .C (clk), .D (new_AGEMA_signal_5290), .Q (new_AGEMA_signal_5291) ) ;
    buf_clk new_AGEMA_reg_buffer_1828 ( .C (clk), .D (new_AGEMA_signal_5292), .Q (new_AGEMA_signal_5293) ) ;
    buf_clk new_AGEMA_reg_buffer_1830 ( .C (clk), .D (new_AGEMA_signal_5294), .Q (new_AGEMA_signal_5295) ) ;
    buf_clk new_AGEMA_reg_buffer_1832 ( .C (clk), .D (new_AGEMA_signal_5296), .Q (new_AGEMA_signal_5297) ) ;
    buf_clk new_AGEMA_reg_buffer_1834 ( .C (clk), .D (new_AGEMA_signal_5298), .Q (new_AGEMA_signal_5299) ) ;
    buf_clk new_AGEMA_reg_buffer_1836 ( .C (clk), .D (new_AGEMA_signal_5300), .Q (new_AGEMA_signal_5301) ) ;
    buf_clk new_AGEMA_reg_buffer_1838 ( .C (clk), .D (new_AGEMA_signal_5302), .Q (new_AGEMA_signal_5303) ) ;
    buf_clk new_AGEMA_reg_buffer_1840 ( .C (clk), .D (new_AGEMA_signal_5304), .Q (new_AGEMA_signal_5305) ) ;
    buf_clk new_AGEMA_reg_buffer_1846 ( .C (clk), .D (new_AGEMA_signal_5310), .Q (new_AGEMA_signal_5311) ) ;
    buf_clk new_AGEMA_reg_buffer_1852 ( .C (clk), .D (new_AGEMA_signal_5316), .Q (new_AGEMA_signal_5317) ) ;
    buf_clk new_AGEMA_reg_buffer_1858 ( .C (clk), .D (new_AGEMA_signal_5322), .Q (new_AGEMA_signal_5323) ) ;
    buf_clk new_AGEMA_reg_buffer_1864 ( .C (clk), .D (new_AGEMA_signal_5328), .Q (new_AGEMA_signal_5329) ) ;
    buf_clk new_AGEMA_reg_buffer_1870 ( .C (clk), .D (new_AGEMA_signal_5334), .Q (new_AGEMA_signal_5335) ) ;
    buf_clk new_AGEMA_reg_buffer_1876 ( .C (clk), .D (new_AGEMA_signal_5340), .Q (new_AGEMA_signal_5341) ) ;
    buf_clk new_AGEMA_reg_buffer_1882 ( .C (clk), .D (new_AGEMA_signal_5346), .Q (new_AGEMA_signal_5347) ) ;
    buf_clk new_AGEMA_reg_buffer_1888 ( .C (clk), .D (new_AGEMA_signal_5352), .Q (new_AGEMA_signal_5353) ) ;
    buf_clk new_AGEMA_reg_buffer_1894 ( .C (clk), .D (new_AGEMA_signal_5358), .Q (new_AGEMA_signal_5359) ) ;
    buf_clk new_AGEMA_reg_buffer_1900 ( .C (clk), .D (new_AGEMA_signal_5364), .Q (new_AGEMA_signal_5365) ) ;
    buf_clk new_AGEMA_reg_buffer_1906 ( .C (clk), .D (new_AGEMA_signal_5370), .Q (new_AGEMA_signal_5371) ) ;
    buf_clk new_AGEMA_reg_buffer_1912 ( .C (clk), .D (new_AGEMA_signal_5376), .Q (new_AGEMA_signal_5377) ) ;
    buf_clk new_AGEMA_reg_buffer_1918 ( .C (clk), .D (new_AGEMA_signal_5382), .Q (new_AGEMA_signal_5383) ) ;
    buf_clk new_AGEMA_reg_buffer_1924 ( .C (clk), .D (new_AGEMA_signal_5388), .Q (new_AGEMA_signal_5389) ) ;
    buf_clk new_AGEMA_reg_buffer_1930 ( .C (clk), .D (new_AGEMA_signal_5394), .Q (new_AGEMA_signal_5395) ) ;
    buf_clk new_AGEMA_reg_buffer_1936 ( .C (clk), .D (new_AGEMA_signal_5400), .Q (new_AGEMA_signal_5401) ) ;
    buf_clk new_AGEMA_reg_buffer_1942 ( .C (clk), .D (new_AGEMA_signal_5406), .Q (new_AGEMA_signal_5407) ) ;
    buf_clk new_AGEMA_reg_buffer_1948 ( .C (clk), .D (new_AGEMA_signal_5412), .Q (new_AGEMA_signal_5413) ) ;
    buf_clk new_AGEMA_reg_buffer_1954 ( .C (clk), .D (new_AGEMA_signal_5418), .Q (new_AGEMA_signal_5419) ) ;
    buf_clk new_AGEMA_reg_buffer_1960 ( .C (clk), .D (new_AGEMA_signal_5424), .Q (new_AGEMA_signal_5425) ) ;
    buf_clk new_AGEMA_reg_buffer_1966 ( .C (clk), .D (new_AGEMA_signal_5430), .Q (new_AGEMA_signal_5431) ) ;
    buf_clk new_AGEMA_reg_buffer_1972 ( .C (clk), .D (new_AGEMA_signal_5436), .Q (new_AGEMA_signal_5437) ) ;
    buf_clk new_AGEMA_reg_buffer_1978 ( .C (clk), .D (new_AGEMA_signal_5442), .Q (new_AGEMA_signal_5443) ) ;
    buf_clk new_AGEMA_reg_buffer_1984 ( .C (clk), .D (new_AGEMA_signal_5448), .Q (new_AGEMA_signal_5449) ) ;
    buf_clk new_AGEMA_reg_buffer_1990 ( .C (clk), .D (new_AGEMA_signal_5454), .Q (new_AGEMA_signal_5455) ) ;
    buf_clk new_AGEMA_reg_buffer_1996 ( .C (clk), .D (new_AGEMA_signal_5460), .Q (new_AGEMA_signal_5461) ) ;
    buf_clk new_AGEMA_reg_buffer_2002 ( .C (clk), .D (new_AGEMA_signal_5466), .Q (new_AGEMA_signal_5467) ) ;
    buf_clk new_AGEMA_reg_buffer_2008 ( .C (clk), .D (new_AGEMA_signal_5472), .Q (new_AGEMA_signal_5473) ) ;
    buf_clk new_AGEMA_reg_buffer_2014 ( .C (clk), .D (new_AGEMA_signal_5478), .Q (new_AGEMA_signal_5479) ) ;
    buf_clk new_AGEMA_reg_buffer_2020 ( .C (clk), .D (new_AGEMA_signal_5484), .Q (new_AGEMA_signal_5485) ) ;
    buf_clk new_AGEMA_reg_buffer_2026 ( .C (clk), .D (new_AGEMA_signal_5490), .Q (new_AGEMA_signal_5491) ) ;
    buf_clk new_AGEMA_reg_buffer_2032 ( .C (clk), .D (new_AGEMA_signal_5496), .Q (new_AGEMA_signal_5497) ) ;
    buf_clk new_AGEMA_reg_buffer_2038 ( .C (clk), .D (new_AGEMA_signal_5502), .Q (new_AGEMA_signal_5503) ) ;
    buf_clk new_AGEMA_reg_buffer_2044 ( .C (clk), .D (new_AGEMA_signal_5508), .Q (new_AGEMA_signal_5509) ) ;
    buf_clk new_AGEMA_reg_buffer_2050 ( .C (clk), .D (new_AGEMA_signal_5514), .Q (new_AGEMA_signal_5515) ) ;
    buf_clk new_AGEMA_reg_buffer_2056 ( .C (clk), .D (new_AGEMA_signal_5520), .Q (new_AGEMA_signal_5521) ) ;
    buf_clk new_AGEMA_reg_buffer_2062 ( .C (clk), .D (new_AGEMA_signal_5526), .Q (new_AGEMA_signal_5527) ) ;
    buf_clk new_AGEMA_reg_buffer_2068 ( .C (clk), .D (new_AGEMA_signal_5532), .Q (new_AGEMA_signal_5533) ) ;
    buf_clk new_AGEMA_reg_buffer_2074 ( .C (clk), .D (new_AGEMA_signal_5538), .Q (new_AGEMA_signal_5539) ) ;
    buf_clk new_AGEMA_reg_buffer_2080 ( .C (clk), .D (new_AGEMA_signal_5544), .Q (new_AGEMA_signal_5545) ) ;
    buf_clk new_AGEMA_reg_buffer_2086 ( .C (clk), .D (new_AGEMA_signal_5550), .Q (new_AGEMA_signal_5551) ) ;
    buf_clk new_AGEMA_reg_buffer_2092 ( .C (clk), .D (new_AGEMA_signal_5556), .Q (new_AGEMA_signal_5557) ) ;
    buf_clk new_AGEMA_reg_buffer_2098 ( .C (clk), .D (new_AGEMA_signal_5562), .Q (new_AGEMA_signal_5563) ) ;
    buf_clk new_AGEMA_reg_buffer_2104 ( .C (clk), .D (new_AGEMA_signal_5568), .Q (new_AGEMA_signal_5569) ) ;
    buf_clk new_AGEMA_reg_buffer_2110 ( .C (clk), .D (new_AGEMA_signal_5574), .Q (new_AGEMA_signal_5575) ) ;
    buf_clk new_AGEMA_reg_buffer_2116 ( .C (clk), .D (new_AGEMA_signal_5580), .Q (new_AGEMA_signal_5581) ) ;
    buf_clk new_AGEMA_reg_buffer_2122 ( .C (clk), .D (new_AGEMA_signal_5586), .Q (new_AGEMA_signal_5587) ) ;
    buf_clk new_AGEMA_reg_buffer_2128 ( .C (clk), .D (new_AGEMA_signal_5592), .Q (new_AGEMA_signal_5593) ) ;
    buf_clk new_AGEMA_reg_buffer_2134 ( .C (clk), .D (new_AGEMA_signal_5598), .Q (new_AGEMA_signal_5599) ) ;
    buf_clk new_AGEMA_reg_buffer_2140 ( .C (clk), .D (new_AGEMA_signal_5604), .Q (new_AGEMA_signal_5605) ) ;
    buf_clk new_AGEMA_reg_buffer_2146 ( .C (clk), .D (new_AGEMA_signal_5610), .Q (new_AGEMA_signal_5611) ) ;
    buf_clk new_AGEMA_reg_buffer_2152 ( .C (clk), .D (new_AGEMA_signal_5616), .Q (new_AGEMA_signal_5617) ) ;
    buf_clk new_AGEMA_reg_buffer_2158 ( .C (clk), .D (new_AGEMA_signal_5622), .Q (new_AGEMA_signal_5623) ) ;
    buf_clk new_AGEMA_reg_buffer_2164 ( .C (clk), .D (new_AGEMA_signal_5628), .Q (new_AGEMA_signal_5629) ) ;
    buf_clk new_AGEMA_reg_buffer_2170 ( .C (clk), .D (new_AGEMA_signal_5634), .Q (new_AGEMA_signal_5635) ) ;
    buf_clk new_AGEMA_reg_buffer_2176 ( .C (clk), .D (new_AGEMA_signal_5640), .Q (new_AGEMA_signal_5641) ) ;
    buf_clk new_AGEMA_reg_buffer_2182 ( .C (clk), .D (new_AGEMA_signal_5646), .Q (new_AGEMA_signal_5647) ) ;
    buf_clk new_AGEMA_reg_buffer_2188 ( .C (clk), .D (new_AGEMA_signal_5652), .Q (new_AGEMA_signal_5653) ) ;
    buf_clk new_AGEMA_reg_buffer_2194 ( .C (clk), .D (new_AGEMA_signal_5658), .Q (new_AGEMA_signal_5659) ) ;
    buf_clk new_AGEMA_reg_buffer_2200 ( .C (clk), .D (new_AGEMA_signal_5664), .Q (new_AGEMA_signal_5665) ) ;
    buf_clk new_AGEMA_reg_buffer_2206 ( .C (clk), .D (new_AGEMA_signal_5670), .Q (new_AGEMA_signal_5671) ) ;
    buf_clk new_AGEMA_reg_buffer_2212 ( .C (clk), .D (new_AGEMA_signal_5676), .Q (new_AGEMA_signal_5677) ) ;
    buf_clk new_AGEMA_reg_buffer_2218 ( .C (clk), .D (new_AGEMA_signal_5682), .Q (new_AGEMA_signal_5683) ) ;
    buf_clk new_AGEMA_reg_buffer_2224 ( .C (clk), .D (new_AGEMA_signal_5688), .Q (new_AGEMA_signal_5689) ) ;
    buf_clk new_AGEMA_reg_buffer_2230 ( .C (clk), .D (new_AGEMA_signal_5694), .Q (new_AGEMA_signal_5695) ) ;
    buf_clk new_AGEMA_reg_buffer_2236 ( .C (clk), .D (new_AGEMA_signal_5700), .Q (new_AGEMA_signal_5701) ) ;
    buf_clk new_AGEMA_reg_buffer_2242 ( .C (clk), .D (new_AGEMA_signal_5706), .Q (new_AGEMA_signal_5707) ) ;
    buf_clk new_AGEMA_reg_buffer_2248 ( .C (clk), .D (new_AGEMA_signal_5712), .Q (new_AGEMA_signal_5713) ) ;
    buf_clk new_AGEMA_reg_buffer_2254 ( .C (clk), .D (new_AGEMA_signal_5718), .Q (new_AGEMA_signal_5719) ) ;
    buf_clk new_AGEMA_reg_buffer_2260 ( .C (clk), .D (new_AGEMA_signal_5724), .Q (new_AGEMA_signal_5725) ) ;
    buf_clk new_AGEMA_reg_buffer_2266 ( .C (clk), .D (new_AGEMA_signal_5730), .Q (new_AGEMA_signal_5731) ) ;
    buf_clk new_AGEMA_reg_buffer_2272 ( .C (clk), .D (new_AGEMA_signal_5736), .Q (new_AGEMA_signal_5737) ) ;
    buf_clk new_AGEMA_reg_buffer_2278 ( .C (clk), .D (new_AGEMA_signal_5742), .Q (new_AGEMA_signal_5743) ) ;
    buf_clk new_AGEMA_reg_buffer_2284 ( .C (clk), .D (new_AGEMA_signal_5748), .Q (new_AGEMA_signal_5749) ) ;
    buf_clk new_AGEMA_reg_buffer_2290 ( .C (clk), .D (new_AGEMA_signal_5754), .Q (new_AGEMA_signal_5755) ) ;
    buf_clk new_AGEMA_reg_buffer_2296 ( .C (clk), .D (new_AGEMA_signal_5760), .Q (new_AGEMA_signal_5761) ) ;
    buf_clk new_AGEMA_reg_buffer_2302 ( .C (clk), .D (new_AGEMA_signal_5766), .Q (new_AGEMA_signal_5767) ) ;
    buf_clk new_AGEMA_reg_buffer_2308 ( .C (clk), .D (new_AGEMA_signal_5772), .Q (new_AGEMA_signal_5773) ) ;
    buf_clk new_AGEMA_reg_buffer_2314 ( .C (clk), .D (new_AGEMA_signal_5778), .Q (new_AGEMA_signal_5779) ) ;
    buf_clk new_AGEMA_reg_buffer_2320 ( .C (clk), .D (new_AGEMA_signal_5784), .Q (new_AGEMA_signal_5785) ) ;
    buf_clk new_AGEMA_reg_buffer_2326 ( .C (clk), .D (new_AGEMA_signal_5790), .Q (new_AGEMA_signal_5791) ) ;
    buf_clk new_AGEMA_reg_buffer_2332 ( .C (clk), .D (new_AGEMA_signal_5796), .Q (new_AGEMA_signal_5797) ) ;
    buf_clk new_AGEMA_reg_buffer_2338 ( .C (clk), .D (new_AGEMA_signal_5802), .Q (new_AGEMA_signal_5803) ) ;
    buf_clk new_AGEMA_reg_buffer_2344 ( .C (clk), .D (new_AGEMA_signal_5808), .Q (new_AGEMA_signal_5809) ) ;
    buf_clk new_AGEMA_reg_buffer_2350 ( .C (clk), .D (new_AGEMA_signal_5814), .Q (new_AGEMA_signal_5815) ) ;
    buf_clk new_AGEMA_reg_buffer_2356 ( .C (clk), .D (new_AGEMA_signal_5820), .Q (new_AGEMA_signal_5821) ) ;
    buf_clk new_AGEMA_reg_buffer_2362 ( .C (clk), .D (new_AGEMA_signal_5826), .Q (new_AGEMA_signal_5827) ) ;
    buf_clk new_AGEMA_reg_buffer_2368 ( .C (clk), .D (new_AGEMA_signal_5832), .Q (new_AGEMA_signal_5833) ) ;
    buf_clk new_AGEMA_reg_buffer_2374 ( .C (clk), .D (new_AGEMA_signal_5838), .Q (new_AGEMA_signal_5839) ) ;
    buf_clk new_AGEMA_reg_buffer_2380 ( .C (clk), .D (new_AGEMA_signal_5844), .Q (new_AGEMA_signal_5845) ) ;
    buf_clk new_AGEMA_reg_buffer_2386 ( .C (clk), .D (new_AGEMA_signal_5850), .Q (new_AGEMA_signal_5851) ) ;
    buf_clk new_AGEMA_reg_buffer_2392 ( .C (clk), .D (new_AGEMA_signal_5856), .Q (new_AGEMA_signal_5857) ) ;
    buf_clk new_AGEMA_reg_buffer_2398 ( .C (clk), .D (new_AGEMA_signal_5862), .Q (new_AGEMA_signal_5863) ) ;
    buf_clk new_AGEMA_reg_buffer_2404 ( .C (clk), .D (new_AGEMA_signal_5868), .Q (new_AGEMA_signal_5869) ) ;
    buf_clk new_AGEMA_reg_buffer_2410 ( .C (clk), .D (new_AGEMA_signal_5874), .Q (new_AGEMA_signal_5875) ) ;
    buf_clk new_AGEMA_reg_buffer_2416 ( .C (clk), .D (new_AGEMA_signal_5880), .Q (new_AGEMA_signal_5881) ) ;
    buf_clk new_AGEMA_reg_buffer_2422 ( .C (clk), .D (new_AGEMA_signal_5886), .Q (new_AGEMA_signal_5887) ) ;
    buf_clk new_AGEMA_reg_buffer_2428 ( .C (clk), .D (new_AGEMA_signal_5892), .Q (new_AGEMA_signal_5893) ) ;
    buf_clk new_AGEMA_reg_buffer_2434 ( .C (clk), .D (new_AGEMA_signal_5898), .Q (new_AGEMA_signal_5899) ) ;
    buf_clk new_AGEMA_reg_buffer_2440 ( .C (clk), .D (new_AGEMA_signal_5904), .Q (new_AGEMA_signal_5905) ) ;
    buf_clk new_AGEMA_reg_buffer_2446 ( .C (clk), .D (new_AGEMA_signal_5910), .Q (new_AGEMA_signal_5911) ) ;
    buf_clk new_AGEMA_reg_buffer_2452 ( .C (clk), .D (new_AGEMA_signal_5916), .Q (new_AGEMA_signal_5917) ) ;
    buf_clk new_AGEMA_reg_buffer_2458 ( .C (clk), .D (new_AGEMA_signal_5922), .Q (new_AGEMA_signal_5923) ) ;
    buf_clk new_AGEMA_reg_buffer_2464 ( .C (clk), .D (new_AGEMA_signal_5928), .Q (new_AGEMA_signal_5929) ) ;
    buf_clk new_AGEMA_reg_buffer_2470 ( .C (clk), .D (new_AGEMA_signal_5934), .Q (new_AGEMA_signal_5935) ) ;
    buf_clk new_AGEMA_reg_buffer_2476 ( .C (clk), .D (new_AGEMA_signal_5940), .Q (new_AGEMA_signal_5941) ) ;
    buf_clk new_AGEMA_reg_buffer_2482 ( .C (clk), .D (new_AGEMA_signal_5946), .Q (new_AGEMA_signal_5947) ) ;
    buf_clk new_AGEMA_reg_buffer_2488 ( .C (clk), .D (new_AGEMA_signal_5952), .Q (new_AGEMA_signal_5953) ) ;
    buf_clk new_AGEMA_reg_buffer_2494 ( .C (clk), .D (new_AGEMA_signal_5958), .Q (new_AGEMA_signal_5959) ) ;
    buf_clk new_AGEMA_reg_buffer_2500 ( .C (clk), .D (new_AGEMA_signal_5964), .Q (new_AGEMA_signal_5965) ) ;
    buf_clk new_AGEMA_reg_buffer_2506 ( .C (clk), .D (new_AGEMA_signal_5970), .Q (new_AGEMA_signal_5971) ) ;
    buf_clk new_AGEMA_reg_buffer_2512 ( .C (clk), .D (new_AGEMA_signal_5976), .Q (new_AGEMA_signal_5977) ) ;
    buf_clk new_AGEMA_reg_buffer_2518 ( .C (clk), .D (new_AGEMA_signal_5982), .Q (new_AGEMA_signal_5983) ) ;
    buf_clk new_AGEMA_reg_buffer_2524 ( .C (clk), .D (new_AGEMA_signal_5988), .Q (new_AGEMA_signal_5989) ) ;
    buf_clk new_AGEMA_reg_buffer_2530 ( .C (clk), .D (new_AGEMA_signal_5994), .Q (new_AGEMA_signal_5995) ) ;
    buf_clk new_AGEMA_reg_buffer_2536 ( .C (clk), .D (new_AGEMA_signal_6000), .Q (new_AGEMA_signal_6001) ) ;
    buf_clk new_AGEMA_reg_buffer_2542 ( .C (clk), .D (new_AGEMA_signal_6006), .Q (new_AGEMA_signal_6007) ) ;
    buf_clk new_AGEMA_reg_buffer_2548 ( .C (clk), .D (new_AGEMA_signal_6012), .Q (new_AGEMA_signal_6013) ) ;
    buf_clk new_AGEMA_reg_buffer_2554 ( .C (clk), .D (new_AGEMA_signal_6018), .Q (new_AGEMA_signal_6019) ) ;
    buf_clk new_AGEMA_reg_buffer_2560 ( .C (clk), .D (new_AGEMA_signal_6024), .Q (new_AGEMA_signal_6025) ) ;
    buf_clk new_AGEMA_reg_buffer_2566 ( .C (clk), .D (new_AGEMA_signal_6030), .Q (new_AGEMA_signal_6031) ) ;
    buf_clk new_AGEMA_reg_buffer_2572 ( .C (clk), .D (new_AGEMA_signal_6036), .Q (new_AGEMA_signal_6037) ) ;
    buf_clk new_AGEMA_reg_buffer_2578 ( .C (clk), .D (new_AGEMA_signal_6042), .Q (new_AGEMA_signal_6043) ) ;
    buf_clk new_AGEMA_reg_buffer_2584 ( .C (clk), .D (new_AGEMA_signal_6048), .Q (new_AGEMA_signal_6049) ) ;
    buf_clk new_AGEMA_reg_buffer_2590 ( .C (clk), .D (new_AGEMA_signal_6054), .Q (new_AGEMA_signal_6055) ) ;
    buf_clk new_AGEMA_reg_buffer_2596 ( .C (clk), .D (new_AGEMA_signal_6060), .Q (new_AGEMA_signal_6061) ) ;
    buf_clk new_AGEMA_reg_buffer_2602 ( .C (clk), .D (new_AGEMA_signal_6066), .Q (new_AGEMA_signal_6067) ) ;
    buf_clk new_AGEMA_reg_buffer_2608 ( .C (clk), .D (new_AGEMA_signal_6072), .Q (new_AGEMA_signal_6073) ) ;
    buf_clk new_AGEMA_reg_buffer_2614 ( .C (clk), .D (new_AGEMA_signal_6078), .Q (new_AGEMA_signal_6079) ) ;
    buf_clk new_AGEMA_reg_buffer_2620 ( .C (clk), .D (new_AGEMA_signal_6084), .Q (new_AGEMA_signal_6085) ) ;
    buf_clk new_AGEMA_reg_buffer_2626 ( .C (clk), .D (new_AGEMA_signal_6090), .Q (new_AGEMA_signal_6091) ) ;
    buf_clk new_AGEMA_reg_buffer_2632 ( .C (clk), .D (new_AGEMA_signal_6096), .Q (new_AGEMA_signal_6097) ) ;
    buf_clk new_AGEMA_reg_buffer_2638 ( .C (clk), .D (new_AGEMA_signal_6102), .Q (new_AGEMA_signal_6103) ) ;
    buf_clk new_AGEMA_reg_buffer_2644 ( .C (clk), .D (new_AGEMA_signal_6108), .Q (new_AGEMA_signal_6109) ) ;
    buf_clk new_AGEMA_reg_buffer_2650 ( .C (clk), .D (new_AGEMA_signal_6114), .Q (new_AGEMA_signal_6115) ) ;
    buf_clk new_AGEMA_reg_buffer_2656 ( .C (clk), .D (new_AGEMA_signal_6120), .Q (new_AGEMA_signal_6121) ) ;
    buf_clk new_AGEMA_reg_buffer_2662 ( .C (clk), .D (new_AGEMA_signal_6126), .Q (new_AGEMA_signal_6127) ) ;
    buf_clk new_AGEMA_reg_buffer_2668 ( .C (clk), .D (new_AGEMA_signal_6132), .Q (new_AGEMA_signal_6133) ) ;
    buf_clk new_AGEMA_reg_buffer_2674 ( .C (clk), .D (new_AGEMA_signal_6138), .Q (new_AGEMA_signal_6139) ) ;
    buf_clk new_AGEMA_reg_buffer_2680 ( .C (clk), .D (new_AGEMA_signal_6144), .Q (new_AGEMA_signal_6145) ) ;
    buf_clk new_AGEMA_reg_buffer_2686 ( .C (clk), .D (new_AGEMA_signal_6150), .Q (new_AGEMA_signal_6151) ) ;
    buf_clk new_AGEMA_reg_buffer_2692 ( .C (clk), .D (new_AGEMA_signal_6156), .Q (new_AGEMA_signal_6157) ) ;
    buf_clk new_AGEMA_reg_buffer_2698 ( .C (clk), .D (new_AGEMA_signal_6162), .Q (new_AGEMA_signal_6163) ) ;
    buf_clk new_AGEMA_reg_buffer_2704 ( .C (clk), .D (new_AGEMA_signal_6168), .Q (new_AGEMA_signal_6169) ) ;
    buf_clk new_AGEMA_reg_buffer_2710 ( .C (clk), .D (new_AGEMA_signal_6174), .Q (new_AGEMA_signal_6175) ) ;
    buf_clk new_AGEMA_reg_buffer_2716 ( .C (clk), .D (new_AGEMA_signal_6180), .Q (new_AGEMA_signal_6181) ) ;
    buf_clk new_AGEMA_reg_buffer_2722 ( .C (clk), .D (new_AGEMA_signal_6186), .Q (new_AGEMA_signal_6187) ) ;
    buf_clk new_AGEMA_reg_buffer_2728 ( .C (clk), .D (new_AGEMA_signal_6192), .Q (new_AGEMA_signal_6193) ) ;
    buf_clk new_AGEMA_reg_buffer_2734 ( .C (clk), .D (new_AGEMA_signal_6198), .Q (new_AGEMA_signal_6199) ) ;
    buf_clk new_AGEMA_reg_buffer_2740 ( .C (clk), .D (new_AGEMA_signal_6204), .Q (new_AGEMA_signal_6205) ) ;
    buf_clk new_AGEMA_reg_buffer_2746 ( .C (clk), .D (new_AGEMA_signal_6210), .Q (new_AGEMA_signal_6211) ) ;
    buf_clk new_AGEMA_reg_buffer_2752 ( .C (clk), .D (new_AGEMA_signal_6216), .Q (new_AGEMA_signal_6217) ) ;
    buf_clk new_AGEMA_reg_buffer_2758 ( .C (clk), .D (new_AGEMA_signal_6222), .Q (new_AGEMA_signal_6223) ) ;
    buf_clk new_AGEMA_reg_buffer_2764 ( .C (clk), .D (new_AGEMA_signal_6228), .Q (new_AGEMA_signal_6229) ) ;
    buf_clk new_AGEMA_reg_buffer_2770 ( .C (clk), .D (new_AGEMA_signal_6234), .Q (new_AGEMA_signal_6235) ) ;
    buf_clk new_AGEMA_reg_buffer_2776 ( .C (clk), .D (new_AGEMA_signal_6240), .Q (new_AGEMA_signal_6241) ) ;
    buf_clk new_AGEMA_reg_buffer_2782 ( .C (clk), .D (new_AGEMA_signal_6246), .Q (new_AGEMA_signal_6247) ) ;
    buf_clk new_AGEMA_reg_buffer_2788 ( .C (clk), .D (new_AGEMA_signal_6252), .Q (new_AGEMA_signal_6253) ) ;
    buf_clk new_AGEMA_reg_buffer_2794 ( .C (clk), .D (new_AGEMA_signal_6258), .Q (new_AGEMA_signal_6259) ) ;
    buf_clk new_AGEMA_reg_buffer_2800 ( .C (clk), .D (new_AGEMA_signal_6264), .Q (new_AGEMA_signal_6265) ) ;
    buf_clk new_AGEMA_reg_buffer_2806 ( .C (clk), .D (new_AGEMA_signal_6270), .Q (new_AGEMA_signal_6271) ) ;
    buf_clk new_AGEMA_reg_buffer_2812 ( .C (clk), .D (new_AGEMA_signal_6276), .Q (new_AGEMA_signal_6277) ) ;
    buf_clk new_AGEMA_reg_buffer_2818 ( .C (clk), .D (new_AGEMA_signal_6282), .Q (new_AGEMA_signal_6283) ) ;
    buf_clk new_AGEMA_reg_buffer_2824 ( .C (clk), .D (new_AGEMA_signal_6288), .Q (new_AGEMA_signal_6289) ) ;
    buf_clk new_AGEMA_reg_buffer_2830 ( .C (clk), .D (new_AGEMA_signal_6294), .Q (new_AGEMA_signal_6295) ) ;
    buf_clk new_AGEMA_reg_buffer_2836 ( .C (clk), .D (new_AGEMA_signal_6300), .Q (new_AGEMA_signal_6301) ) ;
    buf_clk new_AGEMA_reg_buffer_2842 ( .C (clk), .D (new_AGEMA_signal_6306), .Q (new_AGEMA_signal_6307) ) ;
    buf_clk new_AGEMA_reg_buffer_2848 ( .C (clk), .D (new_AGEMA_signal_6312), .Q (new_AGEMA_signal_6313) ) ;
    buf_clk new_AGEMA_reg_buffer_2854 ( .C (clk), .D (new_AGEMA_signal_6318), .Q (new_AGEMA_signal_6319) ) ;
    buf_clk new_AGEMA_reg_buffer_2860 ( .C (clk), .D (new_AGEMA_signal_6324), .Q (new_AGEMA_signal_6325) ) ;
    buf_clk new_AGEMA_reg_buffer_2866 ( .C (clk), .D (new_AGEMA_signal_6330), .Q (new_AGEMA_signal_6331) ) ;
    buf_clk new_AGEMA_reg_buffer_2872 ( .C (clk), .D (new_AGEMA_signal_6336), .Q (new_AGEMA_signal_6337) ) ;
    buf_clk new_AGEMA_reg_buffer_2878 ( .C (clk), .D (new_AGEMA_signal_6342), .Q (new_AGEMA_signal_6343) ) ;
    buf_clk new_AGEMA_reg_buffer_2884 ( .C (clk), .D (new_AGEMA_signal_6348), .Q (new_AGEMA_signal_6349) ) ;
    buf_clk new_AGEMA_reg_buffer_2890 ( .C (clk), .D (new_AGEMA_signal_6354), .Q (new_AGEMA_signal_6355) ) ;
    buf_clk new_AGEMA_reg_buffer_2896 ( .C (clk), .D (new_AGEMA_signal_6360), .Q (new_AGEMA_signal_6361) ) ;
    buf_clk new_AGEMA_reg_buffer_2902 ( .C (clk), .D (new_AGEMA_signal_6366), .Q (new_AGEMA_signal_6367) ) ;
    buf_clk new_AGEMA_reg_buffer_2908 ( .C (clk), .D (new_AGEMA_signal_6372), .Q (new_AGEMA_signal_6373) ) ;
    buf_clk new_AGEMA_reg_buffer_2914 ( .C (clk), .D (new_AGEMA_signal_6378), .Q (new_AGEMA_signal_6379) ) ;
    buf_clk new_AGEMA_reg_buffer_2920 ( .C (clk), .D (new_AGEMA_signal_6384), .Q (new_AGEMA_signal_6385) ) ;
    buf_clk new_AGEMA_reg_buffer_2926 ( .C (clk), .D (new_AGEMA_signal_6390), .Q (new_AGEMA_signal_6391) ) ;
    buf_clk new_AGEMA_reg_buffer_2932 ( .C (clk), .D (new_AGEMA_signal_6396), .Q (new_AGEMA_signal_6397) ) ;
    buf_clk new_AGEMA_reg_buffer_2938 ( .C (clk), .D (new_AGEMA_signal_6402), .Q (new_AGEMA_signal_6403) ) ;
    buf_clk new_AGEMA_reg_buffer_2944 ( .C (clk), .D (new_AGEMA_signal_6408), .Q (new_AGEMA_signal_6409) ) ;
    buf_clk new_AGEMA_reg_buffer_2950 ( .C (clk), .D (new_AGEMA_signal_6414), .Q (new_AGEMA_signal_6415) ) ;
    buf_clk new_AGEMA_reg_buffer_2956 ( .C (clk), .D (new_AGEMA_signal_6420), .Q (new_AGEMA_signal_6421) ) ;
    buf_clk new_AGEMA_reg_buffer_2962 ( .C (clk), .D (new_AGEMA_signal_6426), .Q (new_AGEMA_signal_6427) ) ;
    buf_clk new_AGEMA_reg_buffer_2968 ( .C (clk), .D (new_AGEMA_signal_6432), .Q (new_AGEMA_signal_6433) ) ;
    buf_clk new_AGEMA_reg_buffer_2974 ( .C (clk), .D (new_AGEMA_signal_6438), .Q (new_AGEMA_signal_6439) ) ;
    buf_clk new_AGEMA_reg_buffer_2980 ( .C (clk), .D (new_AGEMA_signal_6444), .Q (new_AGEMA_signal_6445) ) ;
    buf_clk new_AGEMA_reg_buffer_2986 ( .C (clk), .D (new_AGEMA_signal_6450), .Q (new_AGEMA_signal_6451) ) ;
    buf_clk new_AGEMA_reg_buffer_2992 ( .C (clk), .D (new_AGEMA_signal_6456), .Q (new_AGEMA_signal_6457) ) ;
    buf_clk new_AGEMA_reg_buffer_2998 ( .C (clk), .D (new_AGEMA_signal_6462), .Q (new_AGEMA_signal_6463) ) ;
    buf_clk new_AGEMA_reg_buffer_3004 ( .C (clk), .D (new_AGEMA_signal_6468), .Q (new_AGEMA_signal_6469) ) ;
    buf_clk new_AGEMA_reg_buffer_3010 ( .C (clk), .D (new_AGEMA_signal_6474), .Q (new_AGEMA_signal_6475) ) ;
    buf_clk new_AGEMA_reg_buffer_3016 ( .C (clk), .D (new_AGEMA_signal_6480), .Q (new_AGEMA_signal_6481) ) ;
    buf_clk new_AGEMA_reg_buffer_3022 ( .C (clk), .D (new_AGEMA_signal_6486), .Q (new_AGEMA_signal_6487) ) ;
    buf_clk new_AGEMA_reg_buffer_3028 ( .C (clk), .D (new_AGEMA_signal_6492), .Q (new_AGEMA_signal_6493) ) ;
    buf_clk new_AGEMA_reg_buffer_3034 ( .C (clk), .D (new_AGEMA_signal_6498), .Q (new_AGEMA_signal_6499) ) ;
    buf_clk new_AGEMA_reg_buffer_3040 ( .C (clk), .D (new_AGEMA_signal_6504), .Q (new_AGEMA_signal_6505) ) ;
    buf_clk new_AGEMA_reg_buffer_3046 ( .C (clk), .D (new_AGEMA_signal_6510), .Q (new_AGEMA_signal_6511) ) ;
    buf_clk new_AGEMA_reg_buffer_3052 ( .C (clk), .D (new_AGEMA_signal_6516), .Q (new_AGEMA_signal_6517) ) ;
    buf_clk new_AGEMA_reg_buffer_3058 ( .C (clk), .D (new_AGEMA_signal_6522), .Q (new_AGEMA_signal_6523) ) ;
    buf_clk new_AGEMA_reg_buffer_3064 ( .C (clk), .D (new_AGEMA_signal_6528), .Q (new_AGEMA_signal_6529) ) ;
    buf_clk new_AGEMA_reg_buffer_3070 ( .C (clk), .D (new_AGEMA_signal_6534), .Q (new_AGEMA_signal_6535) ) ;
    buf_clk new_AGEMA_reg_buffer_3076 ( .C (clk), .D (new_AGEMA_signal_6540), .Q (new_AGEMA_signal_6541) ) ;
    buf_clk new_AGEMA_reg_buffer_3082 ( .C (clk), .D (new_AGEMA_signal_6546), .Q (new_AGEMA_signal_6547) ) ;
    buf_clk new_AGEMA_reg_buffer_3088 ( .C (clk), .D (new_AGEMA_signal_6552), .Q (new_AGEMA_signal_6553) ) ;
    buf_clk new_AGEMA_reg_buffer_3094 ( .C (clk), .D (new_AGEMA_signal_6558), .Q (new_AGEMA_signal_6559) ) ;
    buf_clk new_AGEMA_reg_buffer_3100 ( .C (clk), .D (new_AGEMA_signal_6564), .Q (new_AGEMA_signal_6565) ) ;
    buf_clk new_AGEMA_reg_buffer_3106 ( .C (clk), .D (new_AGEMA_signal_6570), .Q (new_AGEMA_signal_6571) ) ;
    buf_clk new_AGEMA_reg_buffer_3112 ( .C (clk), .D (new_AGEMA_signal_6576), .Q (new_AGEMA_signal_6577) ) ;
    buf_clk new_AGEMA_reg_buffer_3118 ( .C (clk), .D (new_AGEMA_signal_6582), .Q (new_AGEMA_signal_6583) ) ;
    buf_clk new_AGEMA_reg_buffer_3124 ( .C (clk), .D (new_AGEMA_signal_6588), .Q (new_AGEMA_signal_6589) ) ;
    buf_clk new_AGEMA_reg_buffer_3130 ( .C (clk), .D (new_AGEMA_signal_6594), .Q (new_AGEMA_signal_6595) ) ;
    buf_clk new_AGEMA_reg_buffer_3136 ( .C (clk), .D (new_AGEMA_signal_6600), .Q (new_AGEMA_signal_6601) ) ;
    buf_clk new_AGEMA_reg_buffer_3142 ( .C (clk), .D (new_AGEMA_signal_6606), .Q (new_AGEMA_signal_6607) ) ;
    buf_clk new_AGEMA_reg_buffer_3148 ( .C (clk), .D (new_AGEMA_signal_6612), .Q (new_AGEMA_signal_6613) ) ;
    buf_clk new_AGEMA_reg_buffer_3154 ( .C (clk), .D (new_AGEMA_signal_6618), .Q (new_AGEMA_signal_6619) ) ;
    buf_clk new_AGEMA_reg_buffer_3160 ( .C (clk), .D (new_AGEMA_signal_6624), .Q (new_AGEMA_signal_6625) ) ;
    buf_clk new_AGEMA_reg_buffer_3166 ( .C (clk), .D (new_AGEMA_signal_6630), .Q (new_AGEMA_signal_6631) ) ;
    buf_clk new_AGEMA_reg_buffer_3172 ( .C (clk), .D (new_AGEMA_signal_6636), .Q (new_AGEMA_signal_6637) ) ;
    buf_clk new_AGEMA_reg_buffer_3178 ( .C (clk), .D (new_AGEMA_signal_6642), .Q (new_AGEMA_signal_6643) ) ;
    buf_clk new_AGEMA_reg_buffer_3184 ( .C (clk), .D (new_AGEMA_signal_6648), .Q (new_AGEMA_signal_6649) ) ;
    buf_clk new_AGEMA_reg_buffer_3190 ( .C (clk), .D (new_AGEMA_signal_6654), .Q (new_AGEMA_signal_6655) ) ;
    buf_clk new_AGEMA_reg_buffer_3196 ( .C (clk), .D (new_AGEMA_signal_6660), .Q (new_AGEMA_signal_6661) ) ;
    buf_clk new_AGEMA_reg_buffer_3202 ( .C (clk), .D (new_AGEMA_signal_6666), .Q (new_AGEMA_signal_6667) ) ;
    buf_clk new_AGEMA_reg_buffer_3208 ( .C (clk), .D (new_AGEMA_signal_6672), .Q (new_AGEMA_signal_6673) ) ;
    buf_clk new_AGEMA_reg_buffer_3214 ( .C (clk), .D (new_AGEMA_signal_6678), .Q (new_AGEMA_signal_6679) ) ;
    buf_clk new_AGEMA_reg_buffer_3220 ( .C (clk), .D (new_AGEMA_signal_6684), .Q (new_AGEMA_signal_6685) ) ;
    buf_clk new_AGEMA_reg_buffer_3226 ( .C (clk), .D (new_AGEMA_signal_6690), .Q (new_AGEMA_signal_6691) ) ;
    buf_clk new_AGEMA_reg_buffer_3232 ( .C (clk), .D (new_AGEMA_signal_6696), .Q (new_AGEMA_signal_6697) ) ;
    buf_clk new_AGEMA_reg_buffer_3238 ( .C (clk), .D (new_AGEMA_signal_6702), .Q (new_AGEMA_signal_6703) ) ;
    buf_clk new_AGEMA_reg_buffer_3244 ( .C (clk), .D (new_AGEMA_signal_6708), .Q (new_AGEMA_signal_6709) ) ;
    buf_clk new_AGEMA_reg_buffer_3250 ( .C (clk), .D (new_AGEMA_signal_6714), .Q (new_AGEMA_signal_6715) ) ;
    buf_clk new_AGEMA_reg_buffer_3256 ( .C (clk), .D (new_AGEMA_signal_6720), .Q (new_AGEMA_signal_6721) ) ;
    buf_clk new_AGEMA_reg_buffer_3262 ( .C (clk), .D (new_AGEMA_signal_6726), .Q (new_AGEMA_signal_6727) ) ;
    buf_clk new_AGEMA_reg_buffer_3268 ( .C (clk), .D (new_AGEMA_signal_6732), .Q (new_AGEMA_signal_6733) ) ;
    buf_clk new_AGEMA_reg_buffer_3274 ( .C (clk), .D (new_AGEMA_signal_6738), .Q (new_AGEMA_signal_6739) ) ;
    buf_clk new_AGEMA_reg_buffer_3280 ( .C (clk), .D (new_AGEMA_signal_6744), .Q (new_AGEMA_signal_6745) ) ;
    buf_clk new_AGEMA_reg_buffer_3286 ( .C (clk), .D (new_AGEMA_signal_6750), .Q (new_AGEMA_signal_6751) ) ;
    buf_clk new_AGEMA_reg_buffer_3292 ( .C (clk), .D (new_AGEMA_signal_6756), .Q (new_AGEMA_signal_6757) ) ;
    buf_clk new_AGEMA_reg_buffer_3298 ( .C (clk), .D (new_AGEMA_signal_6762), .Q (new_AGEMA_signal_6763) ) ;
    buf_clk new_AGEMA_reg_buffer_3304 ( .C (clk), .D (new_AGEMA_signal_6768), .Q (new_AGEMA_signal_6769) ) ;
    buf_clk new_AGEMA_reg_buffer_3310 ( .C (clk), .D (new_AGEMA_signal_6774), .Q (new_AGEMA_signal_6775) ) ;
    buf_clk new_AGEMA_reg_buffer_3316 ( .C (clk), .D (new_AGEMA_signal_6780), .Q (new_AGEMA_signal_6781) ) ;
    buf_clk new_AGEMA_reg_buffer_3322 ( .C (clk), .D (new_AGEMA_signal_6786), .Q (new_AGEMA_signal_6787) ) ;
    buf_clk new_AGEMA_reg_buffer_3328 ( .C (clk), .D (new_AGEMA_signal_6792), .Q (new_AGEMA_signal_6793) ) ;
    buf_clk new_AGEMA_reg_buffer_3334 ( .C (clk), .D (new_AGEMA_signal_6798), .Q (new_AGEMA_signal_6799) ) ;
    buf_clk new_AGEMA_reg_buffer_3340 ( .C (clk), .D (new_AGEMA_signal_6804), .Q (new_AGEMA_signal_6805) ) ;
    buf_clk new_AGEMA_reg_buffer_3346 ( .C (clk), .D (new_AGEMA_signal_6810), .Q (new_AGEMA_signal_6811) ) ;
    buf_clk new_AGEMA_reg_buffer_3352 ( .C (clk), .D (new_AGEMA_signal_6816), .Q (new_AGEMA_signal_6817) ) ;
    buf_clk new_AGEMA_reg_buffer_3358 ( .C (clk), .D (new_AGEMA_signal_6822), .Q (new_AGEMA_signal_6823) ) ;
    buf_clk new_AGEMA_reg_buffer_3364 ( .C (clk), .D (new_AGEMA_signal_6828), .Q (new_AGEMA_signal_6829) ) ;
    buf_clk new_AGEMA_reg_buffer_3370 ( .C (clk), .D (new_AGEMA_signal_6834), .Q (new_AGEMA_signal_6835) ) ;
    buf_clk new_AGEMA_reg_buffer_3376 ( .C (clk), .D (new_AGEMA_signal_6840), .Q (new_AGEMA_signal_6841) ) ;
    buf_clk new_AGEMA_reg_buffer_3382 ( .C (clk), .D (new_AGEMA_signal_6846), .Q (new_AGEMA_signal_6847) ) ;
    buf_clk new_AGEMA_reg_buffer_3388 ( .C (clk), .D (new_AGEMA_signal_6852), .Q (new_AGEMA_signal_6853) ) ;
    buf_clk new_AGEMA_reg_buffer_3394 ( .C (clk), .D (new_AGEMA_signal_6858), .Q (new_AGEMA_signal_6859) ) ;
    buf_clk new_AGEMA_reg_buffer_3400 ( .C (clk), .D (new_AGEMA_signal_6864), .Q (new_AGEMA_signal_6865) ) ;
    buf_clk new_AGEMA_reg_buffer_3406 ( .C (clk), .D (new_AGEMA_signal_6870), .Q (new_AGEMA_signal_6871) ) ;
    buf_clk new_AGEMA_reg_buffer_3412 ( .C (clk), .D (new_AGEMA_signal_6876), .Q (new_AGEMA_signal_6877) ) ;
    buf_clk new_AGEMA_reg_buffer_3418 ( .C (clk), .D (new_AGEMA_signal_6882), .Q (new_AGEMA_signal_6883) ) ;
    buf_clk new_AGEMA_reg_buffer_3424 ( .C (clk), .D (new_AGEMA_signal_6888), .Q (new_AGEMA_signal_6889) ) ;
    buf_clk new_AGEMA_reg_buffer_3430 ( .C (clk), .D (new_AGEMA_signal_6894), .Q (new_AGEMA_signal_6895) ) ;
    buf_clk new_AGEMA_reg_buffer_3436 ( .C (clk), .D (new_AGEMA_signal_6900), .Q (new_AGEMA_signal_6901) ) ;
    buf_clk new_AGEMA_reg_buffer_3442 ( .C (clk), .D (new_AGEMA_signal_6906), .Q (new_AGEMA_signal_6907) ) ;
    buf_clk new_AGEMA_reg_buffer_3448 ( .C (clk), .D (new_AGEMA_signal_6912), .Q (new_AGEMA_signal_6913) ) ;
    buf_clk new_AGEMA_reg_buffer_3454 ( .C (clk), .D (new_AGEMA_signal_6918), .Q (new_AGEMA_signal_6919) ) ;
    buf_clk new_AGEMA_reg_buffer_3460 ( .C (clk), .D (new_AGEMA_signal_6924), .Q (new_AGEMA_signal_6925) ) ;
    buf_clk new_AGEMA_reg_buffer_3466 ( .C (clk), .D (new_AGEMA_signal_6930), .Q (new_AGEMA_signal_6931) ) ;
    buf_clk new_AGEMA_reg_buffer_3472 ( .C (clk), .D (new_AGEMA_signal_6936), .Q (new_AGEMA_signal_6937) ) ;
    buf_clk new_AGEMA_reg_buffer_3478 ( .C (clk), .D (new_AGEMA_signal_6942), .Q (new_AGEMA_signal_6943) ) ;
    buf_clk new_AGEMA_reg_buffer_3484 ( .C (clk), .D (new_AGEMA_signal_6948), .Q (new_AGEMA_signal_6949) ) ;
    buf_clk new_AGEMA_reg_buffer_3490 ( .C (clk), .D (new_AGEMA_signal_6954), .Q (new_AGEMA_signal_6955) ) ;
    buf_clk new_AGEMA_reg_buffer_3496 ( .C (clk), .D (new_AGEMA_signal_6960), .Q (new_AGEMA_signal_6961) ) ;
    buf_clk new_AGEMA_reg_buffer_3502 ( .C (clk), .D (new_AGEMA_signal_6966), .Q (new_AGEMA_signal_6967) ) ;
    buf_clk new_AGEMA_reg_buffer_3508 ( .C (clk), .D (new_AGEMA_signal_6972), .Q (new_AGEMA_signal_6973) ) ;
    buf_clk new_AGEMA_reg_buffer_3514 ( .C (clk), .D (new_AGEMA_signal_6978), .Q (new_AGEMA_signal_6979) ) ;
    buf_clk new_AGEMA_reg_buffer_3520 ( .C (clk), .D (new_AGEMA_signal_6984), .Q (new_AGEMA_signal_6985) ) ;
    buf_clk new_AGEMA_reg_buffer_3526 ( .C (clk), .D (new_AGEMA_signal_6990), .Q (new_AGEMA_signal_6991) ) ;
    buf_clk new_AGEMA_reg_buffer_3532 ( .C (clk), .D (new_AGEMA_signal_6996), .Q (new_AGEMA_signal_6997) ) ;
    buf_clk new_AGEMA_reg_buffer_3538 ( .C (clk), .D (new_AGEMA_signal_7002), .Q (new_AGEMA_signal_7003) ) ;
    buf_clk new_AGEMA_reg_buffer_3544 ( .C (clk), .D (new_AGEMA_signal_7008), .Q (new_AGEMA_signal_7009) ) ;
    buf_clk new_AGEMA_reg_buffer_3550 ( .C (clk), .D (new_AGEMA_signal_7014), .Q (new_AGEMA_signal_7015) ) ;
    buf_clk new_AGEMA_reg_buffer_3556 ( .C (clk), .D (new_AGEMA_signal_7020), .Q (new_AGEMA_signal_7021) ) ;
    buf_clk new_AGEMA_reg_buffer_3562 ( .C (clk), .D (new_AGEMA_signal_7026), .Q (new_AGEMA_signal_7027) ) ;
    buf_clk new_AGEMA_reg_buffer_3568 ( .C (clk), .D (new_AGEMA_signal_7032), .Q (new_AGEMA_signal_7033) ) ;
    buf_clk new_AGEMA_reg_buffer_3862 ( .C (clk), .D (new_AGEMA_signal_7326), .Q (new_AGEMA_signal_7327) ) ;
    buf_clk new_AGEMA_reg_buffer_3868 ( .C (clk), .D (new_AGEMA_signal_7332), .Q (new_AGEMA_signal_7333) ) ;
    buf_clk new_AGEMA_reg_buffer_3876 ( .C (clk), .D (new_AGEMA_signal_7340), .Q (new_AGEMA_signal_7341) ) ;
    buf_clk new_AGEMA_reg_buffer_3884 ( .C (clk), .D (new_AGEMA_signal_7348), .Q (new_AGEMA_signal_7349) ) ;
    buf_clk new_AGEMA_reg_buffer_3892 ( .C (clk), .D (new_AGEMA_signal_7356), .Q (new_AGEMA_signal_7357) ) ;
    buf_clk new_AGEMA_reg_buffer_3900 ( .C (clk), .D (new_AGEMA_signal_7364), .Q (new_AGEMA_signal_7365) ) ;
    buf_clk new_AGEMA_reg_buffer_3908 ( .C (clk), .D (new_AGEMA_signal_7372), .Q (new_AGEMA_signal_7373) ) ;
    buf_clk new_AGEMA_reg_buffer_3916 ( .C (clk), .D (new_AGEMA_signal_7380), .Q (new_AGEMA_signal_7381) ) ;
    buf_clk new_AGEMA_reg_buffer_3924 ( .C (clk), .D (new_AGEMA_signal_7388), .Q (new_AGEMA_signal_7389) ) ;
    buf_clk new_AGEMA_reg_buffer_3932 ( .C (clk), .D (new_AGEMA_signal_7396), .Q (new_AGEMA_signal_7397) ) ;
    buf_clk new_AGEMA_reg_buffer_3940 ( .C (clk), .D (new_AGEMA_signal_7404), .Q (new_AGEMA_signal_7405) ) ;
    buf_clk new_AGEMA_reg_buffer_3948 ( .C (clk), .D (new_AGEMA_signal_7412), .Q (new_AGEMA_signal_7413) ) ;
    buf_clk new_AGEMA_reg_buffer_3956 ( .C (clk), .D (new_AGEMA_signal_7420), .Q (new_AGEMA_signal_7421) ) ;
    buf_clk new_AGEMA_reg_buffer_3964 ( .C (clk), .D (new_AGEMA_signal_7428), .Q (new_AGEMA_signal_7429) ) ;
    buf_clk new_AGEMA_reg_buffer_3972 ( .C (clk), .D (new_AGEMA_signal_7436), .Q (new_AGEMA_signal_7437) ) ;
    buf_clk new_AGEMA_reg_buffer_3980 ( .C (clk), .D (new_AGEMA_signal_7444), .Q (new_AGEMA_signal_7445) ) ;
    buf_clk new_AGEMA_reg_buffer_3988 ( .C (clk), .D (new_AGEMA_signal_7452), .Q (new_AGEMA_signal_7453) ) ;
    buf_clk new_AGEMA_reg_buffer_3996 ( .C (clk), .D (new_AGEMA_signal_7460), .Q (new_AGEMA_signal_7461) ) ;
    buf_clk new_AGEMA_reg_buffer_4004 ( .C (clk), .D (new_AGEMA_signal_7468), .Q (new_AGEMA_signal_7469) ) ;
    buf_clk new_AGEMA_reg_buffer_4012 ( .C (clk), .D (new_AGEMA_signal_7476), .Q (new_AGEMA_signal_7477) ) ;
    buf_clk new_AGEMA_reg_buffer_4020 ( .C (clk), .D (new_AGEMA_signal_7484), .Q (new_AGEMA_signal_7485) ) ;
    buf_clk new_AGEMA_reg_buffer_4028 ( .C (clk), .D (new_AGEMA_signal_7492), .Q (new_AGEMA_signal_7493) ) ;
    buf_clk new_AGEMA_reg_buffer_4036 ( .C (clk), .D (new_AGEMA_signal_7500), .Q (new_AGEMA_signal_7501) ) ;
    buf_clk new_AGEMA_reg_buffer_4044 ( .C (clk), .D (new_AGEMA_signal_7508), .Q (new_AGEMA_signal_7509) ) ;
    buf_clk new_AGEMA_reg_buffer_4052 ( .C (clk), .D (new_AGEMA_signal_7516), .Q (new_AGEMA_signal_7517) ) ;
    buf_clk new_AGEMA_reg_buffer_4060 ( .C (clk), .D (new_AGEMA_signal_7524), .Q (new_AGEMA_signal_7525) ) ;
    buf_clk new_AGEMA_reg_buffer_4068 ( .C (clk), .D (new_AGEMA_signal_7532), .Q (new_AGEMA_signal_7533) ) ;
    buf_clk new_AGEMA_reg_buffer_4076 ( .C (clk), .D (new_AGEMA_signal_7540), .Q (new_AGEMA_signal_7541) ) ;
    buf_clk new_AGEMA_reg_buffer_4084 ( .C (clk), .D (new_AGEMA_signal_7548), .Q (new_AGEMA_signal_7549) ) ;
    buf_clk new_AGEMA_reg_buffer_4092 ( .C (clk), .D (new_AGEMA_signal_7556), .Q (new_AGEMA_signal_7557) ) ;
    buf_clk new_AGEMA_reg_buffer_4100 ( .C (clk), .D (new_AGEMA_signal_7564), .Q (new_AGEMA_signal_7565) ) ;
    buf_clk new_AGEMA_reg_buffer_4108 ( .C (clk), .D (new_AGEMA_signal_7572), .Q (new_AGEMA_signal_7573) ) ;
    buf_clk new_AGEMA_reg_buffer_4116 ( .C (clk), .D (new_AGEMA_signal_7580), .Q (new_AGEMA_signal_7581) ) ;
    buf_clk new_AGEMA_reg_buffer_4124 ( .C (clk), .D (new_AGEMA_signal_7588), .Q (new_AGEMA_signal_7589) ) ;
    buf_clk new_AGEMA_reg_buffer_4132 ( .C (clk), .D (new_AGEMA_signal_7596), .Q (new_AGEMA_signal_7597) ) ;
    buf_clk new_AGEMA_reg_buffer_4140 ( .C (clk), .D (new_AGEMA_signal_7604), .Q (new_AGEMA_signal_7605) ) ;
    buf_clk new_AGEMA_reg_buffer_4148 ( .C (clk), .D (new_AGEMA_signal_7612), .Q (new_AGEMA_signal_7613) ) ;
    buf_clk new_AGEMA_reg_buffer_4156 ( .C (clk), .D (new_AGEMA_signal_7620), .Q (new_AGEMA_signal_7621) ) ;
    buf_clk new_AGEMA_reg_buffer_4164 ( .C (clk), .D (new_AGEMA_signal_7628), .Q (new_AGEMA_signal_7629) ) ;
    buf_clk new_AGEMA_reg_buffer_4172 ( .C (clk), .D (new_AGEMA_signal_7636), .Q (new_AGEMA_signal_7637) ) ;
    buf_clk new_AGEMA_reg_buffer_4180 ( .C (clk), .D (new_AGEMA_signal_7644), .Q (new_AGEMA_signal_7645) ) ;
    buf_clk new_AGEMA_reg_buffer_4188 ( .C (clk), .D (new_AGEMA_signal_7652), .Q (new_AGEMA_signal_7653) ) ;
    buf_clk new_AGEMA_reg_buffer_4196 ( .C (clk), .D (new_AGEMA_signal_7660), .Q (new_AGEMA_signal_7661) ) ;
    buf_clk new_AGEMA_reg_buffer_4204 ( .C (clk), .D (new_AGEMA_signal_7668), .Q (new_AGEMA_signal_7669) ) ;
    buf_clk new_AGEMA_reg_buffer_4212 ( .C (clk), .D (new_AGEMA_signal_7676), .Q (new_AGEMA_signal_7677) ) ;
    buf_clk new_AGEMA_reg_buffer_4220 ( .C (clk), .D (new_AGEMA_signal_7684), .Q (new_AGEMA_signal_7685) ) ;
    buf_clk new_AGEMA_reg_buffer_4228 ( .C (clk), .D (new_AGEMA_signal_7692), .Q (new_AGEMA_signal_7693) ) ;
    buf_clk new_AGEMA_reg_buffer_4236 ( .C (clk), .D (new_AGEMA_signal_7700), .Q (new_AGEMA_signal_7701) ) ;
    buf_clk new_AGEMA_reg_buffer_4244 ( .C (clk), .D (new_AGEMA_signal_7708), .Q (new_AGEMA_signal_7709) ) ;
    buf_clk new_AGEMA_reg_buffer_4252 ( .C (clk), .D (new_AGEMA_signal_7716), .Q (new_AGEMA_signal_7717) ) ;
    buf_clk new_AGEMA_reg_buffer_4260 ( .C (clk), .D (new_AGEMA_signal_7724), .Q (new_AGEMA_signal_7725) ) ;
    buf_clk new_AGEMA_reg_buffer_4268 ( .C (clk), .D (new_AGEMA_signal_7732), .Q (new_AGEMA_signal_7733) ) ;
    buf_clk new_AGEMA_reg_buffer_4276 ( .C (clk), .D (new_AGEMA_signal_7740), .Q (new_AGEMA_signal_7741) ) ;
    buf_clk new_AGEMA_reg_buffer_4284 ( .C (clk), .D (new_AGEMA_signal_7748), .Q (new_AGEMA_signal_7749) ) ;
    buf_clk new_AGEMA_reg_buffer_4292 ( .C (clk), .D (new_AGEMA_signal_7756), .Q (new_AGEMA_signal_7757) ) ;
    buf_clk new_AGEMA_reg_buffer_4300 ( .C (clk), .D (new_AGEMA_signal_7764), .Q (new_AGEMA_signal_7765) ) ;
    buf_clk new_AGEMA_reg_buffer_4308 ( .C (clk), .D (new_AGEMA_signal_7772), .Q (new_AGEMA_signal_7773) ) ;
    buf_clk new_AGEMA_reg_buffer_4316 ( .C (clk), .D (new_AGEMA_signal_7780), .Q (new_AGEMA_signal_7781) ) ;
    buf_clk new_AGEMA_reg_buffer_4324 ( .C (clk), .D (new_AGEMA_signal_7788), .Q (new_AGEMA_signal_7789) ) ;
    buf_clk new_AGEMA_reg_buffer_4332 ( .C (clk), .D (new_AGEMA_signal_7796), .Q (new_AGEMA_signal_7797) ) ;
    buf_clk new_AGEMA_reg_buffer_4340 ( .C (clk), .D (new_AGEMA_signal_7804), .Q (new_AGEMA_signal_7805) ) ;
    buf_clk new_AGEMA_reg_buffer_4348 ( .C (clk), .D (new_AGEMA_signal_7812), .Q (new_AGEMA_signal_7813) ) ;
    buf_clk new_AGEMA_reg_buffer_4356 ( .C (clk), .D (new_AGEMA_signal_7820), .Q (new_AGEMA_signal_7821) ) ;
    buf_clk new_AGEMA_reg_buffer_4364 ( .C (clk), .D (new_AGEMA_signal_7828), .Q (new_AGEMA_signal_7829) ) ;
    buf_clk new_AGEMA_reg_buffer_4372 ( .C (clk), .D (new_AGEMA_signal_7836), .Q (new_AGEMA_signal_7837) ) ;
    buf_clk new_AGEMA_reg_buffer_4380 ( .C (clk), .D (new_AGEMA_signal_7844), .Q (new_AGEMA_signal_7845) ) ;
    buf_clk new_AGEMA_reg_buffer_4388 ( .C (clk), .D (new_AGEMA_signal_7852), .Q (new_AGEMA_signal_7853) ) ;
    buf_clk new_AGEMA_reg_buffer_4396 ( .C (clk), .D (new_AGEMA_signal_7860), .Q (new_AGEMA_signal_7861) ) ;
    buf_clk new_AGEMA_reg_buffer_4404 ( .C (clk), .D (new_AGEMA_signal_7868), .Q (new_AGEMA_signal_7869) ) ;
    buf_clk new_AGEMA_reg_buffer_4412 ( .C (clk), .D (new_AGEMA_signal_7876), .Q (new_AGEMA_signal_7877) ) ;
    buf_clk new_AGEMA_reg_buffer_4420 ( .C (clk), .D (new_AGEMA_signal_7884), .Q (new_AGEMA_signal_7885) ) ;
    buf_clk new_AGEMA_reg_buffer_4428 ( .C (clk), .D (new_AGEMA_signal_7892), .Q (new_AGEMA_signal_7893) ) ;
    buf_clk new_AGEMA_reg_buffer_4436 ( .C (clk), .D (new_AGEMA_signal_7900), .Q (new_AGEMA_signal_7901) ) ;
    buf_clk new_AGEMA_reg_buffer_4444 ( .C (clk), .D (new_AGEMA_signal_7908), .Q (new_AGEMA_signal_7909) ) ;
    buf_clk new_AGEMA_reg_buffer_4452 ( .C (clk), .D (new_AGEMA_signal_7916), .Q (new_AGEMA_signal_7917) ) ;
    buf_clk new_AGEMA_reg_buffer_4460 ( .C (clk), .D (new_AGEMA_signal_7924), .Q (new_AGEMA_signal_7925) ) ;
    buf_clk new_AGEMA_reg_buffer_4468 ( .C (clk), .D (new_AGEMA_signal_7932), .Q (new_AGEMA_signal_7933) ) ;
    buf_clk new_AGEMA_reg_buffer_4476 ( .C (clk), .D (new_AGEMA_signal_7940), .Q (new_AGEMA_signal_7941) ) ;
    buf_clk new_AGEMA_reg_buffer_4484 ( .C (clk), .D (new_AGEMA_signal_7948), .Q (new_AGEMA_signal_7949) ) ;
    buf_clk new_AGEMA_reg_buffer_4492 ( .C (clk), .D (new_AGEMA_signal_7956), .Q (new_AGEMA_signal_7957) ) ;
    buf_clk new_AGEMA_reg_buffer_4500 ( .C (clk), .D (new_AGEMA_signal_7964), .Q (new_AGEMA_signal_7965) ) ;
    buf_clk new_AGEMA_reg_buffer_4508 ( .C (clk), .D (new_AGEMA_signal_7972), .Q (new_AGEMA_signal_7973) ) ;
    buf_clk new_AGEMA_reg_buffer_4516 ( .C (clk), .D (new_AGEMA_signal_7980), .Q (new_AGEMA_signal_7981) ) ;
    buf_clk new_AGEMA_reg_buffer_4524 ( .C (clk), .D (new_AGEMA_signal_7988), .Q (new_AGEMA_signal_7989) ) ;
    buf_clk new_AGEMA_reg_buffer_4532 ( .C (clk), .D (new_AGEMA_signal_7996), .Q (new_AGEMA_signal_7997) ) ;
    buf_clk new_AGEMA_reg_buffer_4540 ( .C (clk), .D (new_AGEMA_signal_8004), .Q (new_AGEMA_signal_8005) ) ;
    buf_clk new_AGEMA_reg_buffer_4548 ( .C (clk), .D (new_AGEMA_signal_8012), .Q (new_AGEMA_signal_8013) ) ;
    buf_clk new_AGEMA_reg_buffer_4556 ( .C (clk), .D (new_AGEMA_signal_8020), .Q (new_AGEMA_signal_8021) ) ;
    buf_clk new_AGEMA_reg_buffer_4564 ( .C (clk), .D (new_AGEMA_signal_8028), .Q (new_AGEMA_signal_8029) ) ;
    buf_clk new_AGEMA_reg_buffer_4572 ( .C (clk), .D (new_AGEMA_signal_8036), .Q (new_AGEMA_signal_8037) ) ;
    buf_clk new_AGEMA_reg_buffer_4580 ( .C (clk), .D (new_AGEMA_signal_8044), .Q (new_AGEMA_signal_8045) ) ;
    buf_clk new_AGEMA_reg_buffer_4588 ( .C (clk), .D (new_AGEMA_signal_8052), .Q (new_AGEMA_signal_8053) ) ;
    buf_clk new_AGEMA_reg_buffer_4596 ( .C (clk), .D (new_AGEMA_signal_8060), .Q (new_AGEMA_signal_8061) ) ;
    buf_clk new_AGEMA_reg_buffer_4604 ( .C (clk), .D (new_AGEMA_signal_8068), .Q (new_AGEMA_signal_8069) ) ;
    buf_clk new_AGEMA_reg_buffer_4612 ( .C (clk), .D (new_AGEMA_signal_8076), .Q (new_AGEMA_signal_8077) ) ;
    buf_clk new_AGEMA_reg_buffer_4620 ( .C (clk), .D (new_AGEMA_signal_8084), .Q (new_AGEMA_signal_8085) ) ;
    buf_clk new_AGEMA_reg_buffer_4628 ( .C (clk), .D (new_AGEMA_signal_8092), .Q (new_AGEMA_signal_8093) ) ;
    buf_clk new_AGEMA_reg_buffer_4636 ( .C (clk), .D (new_AGEMA_signal_8100), .Q (new_AGEMA_signal_8101) ) ;
    buf_clk new_AGEMA_reg_buffer_4644 ( .C (clk), .D (new_AGEMA_signal_8108), .Q (new_AGEMA_signal_8109) ) ;
    buf_clk new_AGEMA_reg_buffer_4652 ( .C (clk), .D (new_AGEMA_signal_8116), .Q (new_AGEMA_signal_8117) ) ;
    buf_clk new_AGEMA_reg_buffer_4660 ( .C (clk), .D (new_AGEMA_signal_8124), .Q (new_AGEMA_signal_8125) ) ;
    buf_clk new_AGEMA_reg_buffer_4668 ( .C (clk), .D (new_AGEMA_signal_8132), .Q (new_AGEMA_signal_8133) ) ;
    buf_clk new_AGEMA_reg_buffer_4676 ( .C (clk), .D (new_AGEMA_signal_8140), .Q (new_AGEMA_signal_8141) ) ;
    buf_clk new_AGEMA_reg_buffer_4684 ( .C (clk), .D (new_AGEMA_signal_8148), .Q (new_AGEMA_signal_8149) ) ;
    buf_clk new_AGEMA_reg_buffer_4692 ( .C (clk), .D (new_AGEMA_signal_8156), .Q (new_AGEMA_signal_8157) ) ;
    buf_clk new_AGEMA_reg_buffer_4700 ( .C (clk), .D (new_AGEMA_signal_8164), .Q (new_AGEMA_signal_8165) ) ;
    buf_clk new_AGEMA_reg_buffer_4708 ( .C (clk), .D (new_AGEMA_signal_8172), .Q (new_AGEMA_signal_8173) ) ;
    buf_clk new_AGEMA_reg_buffer_4716 ( .C (clk), .D (new_AGEMA_signal_8180), .Q (new_AGEMA_signal_8181) ) ;
    buf_clk new_AGEMA_reg_buffer_4724 ( .C (clk), .D (new_AGEMA_signal_8188), .Q (new_AGEMA_signal_8189) ) ;
    buf_clk new_AGEMA_reg_buffer_4732 ( .C (clk), .D (new_AGEMA_signal_8196), .Q (new_AGEMA_signal_8197) ) ;
    buf_clk new_AGEMA_reg_buffer_4740 ( .C (clk), .D (new_AGEMA_signal_8204), .Q (new_AGEMA_signal_8205) ) ;
    buf_clk new_AGEMA_reg_buffer_4748 ( .C (clk), .D (new_AGEMA_signal_8212), .Q (new_AGEMA_signal_8213) ) ;
    buf_clk new_AGEMA_reg_buffer_4756 ( .C (clk), .D (new_AGEMA_signal_8220), .Q (new_AGEMA_signal_8221) ) ;
    buf_clk new_AGEMA_reg_buffer_4764 ( .C (clk), .D (new_AGEMA_signal_8228), .Q (new_AGEMA_signal_8229) ) ;
    buf_clk new_AGEMA_reg_buffer_4772 ( .C (clk), .D (new_AGEMA_signal_8236), .Q (new_AGEMA_signal_8237) ) ;
    buf_clk new_AGEMA_reg_buffer_4780 ( .C (clk), .D (new_AGEMA_signal_8244), .Q (new_AGEMA_signal_8245) ) ;
    buf_clk new_AGEMA_reg_buffer_4788 ( .C (clk), .D (new_AGEMA_signal_8252), .Q (new_AGEMA_signal_8253) ) ;
    buf_clk new_AGEMA_reg_buffer_4796 ( .C (clk), .D (new_AGEMA_signal_8260), .Q (new_AGEMA_signal_8261) ) ;
    buf_clk new_AGEMA_reg_buffer_4804 ( .C (clk), .D (new_AGEMA_signal_8268), .Q (new_AGEMA_signal_8269) ) ;
    buf_clk new_AGEMA_reg_buffer_4812 ( .C (clk), .D (new_AGEMA_signal_8276), .Q (new_AGEMA_signal_8277) ) ;
    buf_clk new_AGEMA_reg_buffer_4820 ( .C (clk), .D (new_AGEMA_signal_8284), .Q (new_AGEMA_signal_8285) ) ;
    buf_clk new_AGEMA_reg_buffer_4828 ( .C (clk), .D (new_AGEMA_signal_8292), .Q (new_AGEMA_signal_8293) ) ;
    buf_clk new_AGEMA_reg_buffer_4836 ( .C (clk), .D (new_AGEMA_signal_8300), .Q (new_AGEMA_signal_8301) ) ;
    buf_clk new_AGEMA_reg_buffer_4844 ( .C (clk), .D (new_AGEMA_signal_8308), .Q (new_AGEMA_signal_8309) ) ;
    buf_clk new_AGEMA_reg_buffer_4852 ( .C (clk), .D (new_AGEMA_signal_8316), .Q (new_AGEMA_signal_8317) ) ;
    buf_clk new_AGEMA_reg_buffer_4860 ( .C (clk), .D (new_AGEMA_signal_8324), .Q (new_AGEMA_signal_8325) ) ;
    buf_clk new_AGEMA_reg_buffer_4868 ( .C (clk), .D (new_AGEMA_signal_8332), .Q (new_AGEMA_signal_8333) ) ;
    buf_clk new_AGEMA_reg_buffer_4876 ( .C (clk), .D (new_AGEMA_signal_8340), .Q (new_AGEMA_signal_8341) ) ;
    buf_clk new_AGEMA_reg_buffer_4884 ( .C (clk), .D (new_AGEMA_signal_8348), .Q (new_AGEMA_signal_8349) ) ;
    buf_clk new_AGEMA_reg_buffer_4892 ( .C (clk), .D (new_AGEMA_signal_8356), .Q (new_AGEMA_signal_8357) ) ;
    buf_clk new_AGEMA_reg_buffer_4900 ( .C (clk), .D (new_AGEMA_signal_8364), .Q (new_AGEMA_signal_8365) ) ;
    buf_clk new_AGEMA_reg_buffer_4908 ( .C (clk), .D (new_AGEMA_signal_8372), .Q (new_AGEMA_signal_8373) ) ;
    buf_clk new_AGEMA_reg_buffer_4916 ( .C (clk), .D (new_AGEMA_signal_8380), .Q (new_AGEMA_signal_8381) ) ;
    buf_clk new_AGEMA_reg_buffer_4924 ( .C (clk), .D (new_AGEMA_signal_8388), .Q (new_AGEMA_signal_8389) ) ;
    buf_clk new_AGEMA_reg_buffer_4932 ( .C (clk), .D (new_AGEMA_signal_8396), .Q (new_AGEMA_signal_8397) ) ;
    buf_clk new_AGEMA_reg_buffer_4940 ( .C (clk), .D (new_AGEMA_signal_8404), .Q (new_AGEMA_signal_8405) ) ;
    buf_clk new_AGEMA_reg_buffer_4948 ( .C (clk), .D (new_AGEMA_signal_8412), .Q (new_AGEMA_signal_8413) ) ;
    buf_clk new_AGEMA_reg_buffer_4956 ( .C (clk), .D (new_AGEMA_signal_8420), .Q (new_AGEMA_signal_8421) ) ;
    buf_clk new_AGEMA_reg_buffer_4964 ( .C (clk), .D (new_AGEMA_signal_8428), .Q (new_AGEMA_signal_8429) ) ;
    buf_clk new_AGEMA_reg_buffer_4972 ( .C (clk), .D (new_AGEMA_signal_8436), .Q (new_AGEMA_signal_8437) ) ;
    buf_clk new_AGEMA_reg_buffer_4980 ( .C (clk), .D (new_AGEMA_signal_8444), .Q (new_AGEMA_signal_8445) ) ;
    buf_clk new_AGEMA_reg_buffer_4988 ( .C (clk), .D (new_AGEMA_signal_8452), .Q (new_AGEMA_signal_8453) ) ;
    buf_clk new_AGEMA_reg_buffer_4996 ( .C (clk), .D (new_AGEMA_signal_8460), .Q (new_AGEMA_signal_8461) ) ;
    buf_clk new_AGEMA_reg_buffer_5004 ( .C (clk), .D (new_AGEMA_signal_8468), .Q (new_AGEMA_signal_8469) ) ;
    buf_clk new_AGEMA_reg_buffer_5012 ( .C (clk), .D (new_AGEMA_signal_8476), .Q (new_AGEMA_signal_8477) ) ;
    buf_clk new_AGEMA_reg_buffer_5020 ( .C (clk), .D (new_AGEMA_signal_8484), .Q (new_AGEMA_signal_8485) ) ;
    buf_clk new_AGEMA_reg_buffer_5028 ( .C (clk), .D (new_AGEMA_signal_8492), .Q (new_AGEMA_signal_8493) ) ;
    buf_clk new_AGEMA_reg_buffer_5036 ( .C (clk), .D (new_AGEMA_signal_8500), .Q (new_AGEMA_signal_8501) ) ;
    buf_clk new_AGEMA_reg_buffer_5044 ( .C (clk), .D (new_AGEMA_signal_8508), .Q (new_AGEMA_signal_8509) ) ;
    buf_clk new_AGEMA_reg_buffer_5052 ( .C (clk), .D (new_AGEMA_signal_8516), .Q (new_AGEMA_signal_8517) ) ;
    buf_clk new_AGEMA_reg_buffer_5060 ( .C (clk), .D (new_AGEMA_signal_8524), .Q (new_AGEMA_signal_8525) ) ;
    buf_clk new_AGEMA_reg_buffer_5068 ( .C (clk), .D (new_AGEMA_signal_8532), .Q (new_AGEMA_signal_8533) ) ;
    buf_clk new_AGEMA_reg_buffer_5076 ( .C (clk), .D (new_AGEMA_signal_8540), .Q (new_AGEMA_signal_8541) ) ;
    buf_clk new_AGEMA_reg_buffer_5084 ( .C (clk), .D (new_AGEMA_signal_8548), .Q (new_AGEMA_signal_8549) ) ;
    buf_clk new_AGEMA_reg_buffer_5092 ( .C (clk), .D (new_AGEMA_signal_8556), .Q (new_AGEMA_signal_8557) ) ;
    buf_clk new_AGEMA_reg_buffer_5100 ( .C (clk), .D (new_AGEMA_signal_8564), .Q (new_AGEMA_signal_8565) ) ;
    buf_clk new_AGEMA_reg_buffer_5108 ( .C (clk), .D (new_AGEMA_signal_8572), .Q (new_AGEMA_signal_8573) ) ;
    buf_clk new_AGEMA_reg_buffer_5116 ( .C (clk), .D (new_AGEMA_signal_8580), .Q (new_AGEMA_signal_8581) ) ;
    buf_clk new_AGEMA_reg_buffer_5124 ( .C (clk), .D (new_AGEMA_signal_8588), .Q (new_AGEMA_signal_8589) ) ;
    buf_clk new_AGEMA_reg_buffer_5132 ( .C (clk), .D (new_AGEMA_signal_8596), .Q (new_AGEMA_signal_8597) ) ;
    buf_clk new_AGEMA_reg_buffer_5140 ( .C (clk), .D (new_AGEMA_signal_8604), .Q (new_AGEMA_signal_8605) ) ;
    buf_clk new_AGEMA_reg_buffer_5148 ( .C (clk), .D (new_AGEMA_signal_8612), .Q (new_AGEMA_signal_8613) ) ;
    buf_clk new_AGEMA_reg_buffer_5156 ( .C (clk), .D (new_AGEMA_signal_8620), .Q (new_AGEMA_signal_8621) ) ;
    buf_clk new_AGEMA_reg_buffer_5164 ( .C (clk), .D (new_AGEMA_signal_8628), .Q (new_AGEMA_signal_8629) ) ;
    buf_clk new_AGEMA_reg_buffer_5172 ( .C (clk), .D (new_AGEMA_signal_8636), .Q (new_AGEMA_signal_8637) ) ;
    buf_clk new_AGEMA_reg_buffer_5180 ( .C (clk), .D (new_AGEMA_signal_8644), .Q (new_AGEMA_signal_8645) ) ;
    buf_clk new_AGEMA_reg_buffer_5188 ( .C (clk), .D (new_AGEMA_signal_8652), .Q (new_AGEMA_signal_8653) ) ;
    buf_clk new_AGEMA_reg_buffer_5196 ( .C (clk), .D (new_AGEMA_signal_8660), .Q (new_AGEMA_signal_8661) ) ;
    buf_clk new_AGEMA_reg_buffer_5204 ( .C (clk), .D (new_AGEMA_signal_8668), .Q (new_AGEMA_signal_8669) ) ;
    buf_clk new_AGEMA_reg_buffer_5212 ( .C (clk), .D (new_AGEMA_signal_8676), .Q (new_AGEMA_signal_8677) ) ;
    buf_clk new_AGEMA_reg_buffer_5220 ( .C (clk), .D (new_AGEMA_signal_8684), .Q (new_AGEMA_signal_8685) ) ;
    buf_clk new_AGEMA_reg_buffer_5228 ( .C (clk), .D (new_AGEMA_signal_8692), .Q (new_AGEMA_signal_8693) ) ;
    buf_clk new_AGEMA_reg_buffer_5236 ( .C (clk), .D (new_AGEMA_signal_8700), .Q (new_AGEMA_signal_8701) ) ;
    buf_clk new_AGEMA_reg_buffer_5244 ( .C (clk), .D (new_AGEMA_signal_8708), .Q (new_AGEMA_signal_8709) ) ;
    buf_clk new_AGEMA_reg_buffer_5252 ( .C (clk), .D (new_AGEMA_signal_8716), .Q (new_AGEMA_signal_8717) ) ;
    buf_clk new_AGEMA_reg_buffer_5260 ( .C (clk), .D (new_AGEMA_signal_8724), .Q (new_AGEMA_signal_8725) ) ;
    buf_clk new_AGEMA_reg_buffer_5268 ( .C (clk), .D (new_AGEMA_signal_8732), .Q (new_AGEMA_signal_8733) ) ;
    buf_clk new_AGEMA_reg_buffer_5276 ( .C (clk), .D (new_AGEMA_signal_8740), .Q (new_AGEMA_signal_8741) ) ;
    buf_clk new_AGEMA_reg_buffer_5284 ( .C (clk), .D (new_AGEMA_signal_8748), .Q (new_AGEMA_signal_8749) ) ;
    buf_clk new_AGEMA_reg_buffer_5292 ( .C (clk), .D (new_AGEMA_signal_8756), .Q (new_AGEMA_signal_8757) ) ;
    buf_clk new_AGEMA_reg_buffer_5300 ( .C (clk), .D (new_AGEMA_signal_8764), .Q (new_AGEMA_signal_8765) ) ;
    buf_clk new_AGEMA_reg_buffer_5308 ( .C (clk), .D (new_AGEMA_signal_8772), .Q (new_AGEMA_signal_8773) ) ;
    buf_clk new_AGEMA_reg_buffer_5316 ( .C (clk), .D (new_AGEMA_signal_8780), .Q (new_AGEMA_signal_8781) ) ;
    buf_clk new_AGEMA_reg_buffer_5324 ( .C (clk), .D (new_AGEMA_signal_8788), .Q (new_AGEMA_signal_8789) ) ;
    buf_clk new_AGEMA_reg_buffer_5332 ( .C (clk), .D (new_AGEMA_signal_8796), .Q (new_AGEMA_signal_8797) ) ;
    buf_clk new_AGEMA_reg_buffer_5340 ( .C (clk), .D (new_AGEMA_signal_8804), .Q (new_AGEMA_signal_8805) ) ;
    buf_clk new_AGEMA_reg_buffer_5348 ( .C (clk), .D (new_AGEMA_signal_8812), .Q (new_AGEMA_signal_8813) ) ;
    buf_clk new_AGEMA_reg_buffer_5356 ( .C (clk), .D (new_AGEMA_signal_8820), .Q (new_AGEMA_signal_8821) ) ;
    buf_clk new_AGEMA_reg_buffer_5364 ( .C (clk), .D (new_AGEMA_signal_8828), .Q (new_AGEMA_signal_8829) ) ;
    buf_clk new_AGEMA_reg_buffer_5372 ( .C (clk), .D (new_AGEMA_signal_8836), .Q (new_AGEMA_signal_8837) ) ;
    buf_clk new_AGEMA_reg_buffer_5380 ( .C (clk), .D (new_AGEMA_signal_8844), .Q (new_AGEMA_signal_8845) ) ;
    buf_clk new_AGEMA_reg_buffer_5388 ( .C (clk), .D (new_AGEMA_signal_8852), .Q (new_AGEMA_signal_8853) ) ;
    buf_clk new_AGEMA_reg_buffer_5396 ( .C (clk), .D (new_AGEMA_signal_8860), .Q (new_AGEMA_signal_8861) ) ;
    buf_clk new_AGEMA_reg_buffer_5406 ( .C (clk), .D (new_AGEMA_signal_8870), .Q (new_AGEMA_signal_8871) ) ;
    buf_clk new_AGEMA_reg_buffer_5414 ( .C (clk), .D (new_AGEMA_signal_8878), .Q (new_AGEMA_signal_8879) ) ;
    buf_clk new_AGEMA_reg_buffer_5422 ( .C (clk), .D (new_AGEMA_signal_8886), .Q (new_AGEMA_signal_8887) ) ;
    buf_clk new_AGEMA_reg_buffer_5430 ( .C (clk), .D (new_AGEMA_signal_8894), .Q (new_AGEMA_signal_8895) ) ;
    buf_clk new_AGEMA_reg_buffer_5438 ( .C (clk), .D (new_AGEMA_signal_8902), .Q (new_AGEMA_signal_8903) ) ;
    buf_clk new_AGEMA_reg_buffer_5446 ( .C (clk), .D (new_AGEMA_signal_8910), .Q (new_AGEMA_signal_8911) ) ;
    buf_clk new_AGEMA_reg_buffer_5454 ( .C (clk), .D (new_AGEMA_signal_8918), .Q (new_AGEMA_signal_8919) ) ;
    buf_clk new_AGEMA_reg_buffer_5462 ( .C (clk), .D (new_AGEMA_signal_8926), .Q (new_AGEMA_signal_8927) ) ;
    buf_clk new_AGEMA_reg_buffer_5470 ( .C (clk), .D (new_AGEMA_signal_8934), .Q (new_AGEMA_signal_8935) ) ;
    buf_clk new_AGEMA_reg_buffer_5478 ( .C (clk), .D (new_AGEMA_signal_8942), .Q (new_AGEMA_signal_8943) ) ;
    buf_clk new_AGEMA_reg_buffer_5486 ( .C (clk), .D (new_AGEMA_signal_8950), .Q (new_AGEMA_signal_8951) ) ;
    buf_clk new_AGEMA_reg_buffer_5494 ( .C (clk), .D (new_AGEMA_signal_8958), .Q (new_AGEMA_signal_8959) ) ;
    buf_clk new_AGEMA_reg_buffer_5502 ( .C (clk), .D (new_AGEMA_signal_8966), .Q (new_AGEMA_signal_8967) ) ;
    buf_clk new_AGEMA_reg_buffer_5510 ( .C (clk), .D (new_AGEMA_signal_8974), .Q (new_AGEMA_signal_8975) ) ;
    buf_clk new_AGEMA_reg_buffer_5518 ( .C (clk), .D (new_AGEMA_signal_8982), .Q (new_AGEMA_signal_8983) ) ;
    buf_clk new_AGEMA_reg_buffer_5526 ( .C (clk), .D (new_AGEMA_signal_8990), .Q (new_AGEMA_signal_8991) ) ;
    buf_clk new_AGEMA_reg_buffer_5534 ( .C (clk), .D (new_AGEMA_signal_8998), .Q (new_AGEMA_signal_8999) ) ;
    buf_clk new_AGEMA_reg_buffer_5542 ( .C (clk), .D (new_AGEMA_signal_9006), .Q (new_AGEMA_signal_9007) ) ;
    buf_clk new_AGEMA_reg_buffer_5550 ( .C (clk), .D (new_AGEMA_signal_9014), .Q (new_AGEMA_signal_9015) ) ;
    buf_clk new_AGEMA_reg_buffer_5558 ( .C (clk), .D (new_AGEMA_signal_9022), .Q (new_AGEMA_signal_9023) ) ;
    buf_clk new_AGEMA_reg_buffer_5566 ( .C (clk), .D (new_AGEMA_signal_9030), .Q (new_AGEMA_signal_9031) ) ;
    buf_clk new_AGEMA_reg_buffer_5574 ( .C (clk), .D (new_AGEMA_signal_9038), .Q (new_AGEMA_signal_9039) ) ;
    buf_clk new_AGEMA_reg_buffer_5582 ( .C (clk), .D (new_AGEMA_signal_9046), .Q (new_AGEMA_signal_9047) ) ;
    buf_clk new_AGEMA_reg_buffer_5590 ( .C (clk), .D (new_AGEMA_signal_9054), .Q (new_AGEMA_signal_9055) ) ;
    buf_clk new_AGEMA_reg_buffer_5598 ( .C (clk), .D (new_AGEMA_signal_9062), .Q (new_AGEMA_signal_9063) ) ;
    buf_clk new_AGEMA_reg_buffer_5606 ( .C (clk), .D (new_AGEMA_signal_9070), .Q (new_AGEMA_signal_9071) ) ;
    buf_clk new_AGEMA_reg_buffer_5614 ( .C (clk), .D (new_AGEMA_signal_9078), .Q (new_AGEMA_signal_9079) ) ;
    buf_clk new_AGEMA_reg_buffer_5622 ( .C (clk), .D (new_AGEMA_signal_9086), .Q (new_AGEMA_signal_9087) ) ;
    buf_clk new_AGEMA_reg_buffer_5630 ( .C (clk), .D (new_AGEMA_signal_9094), .Q (new_AGEMA_signal_9095) ) ;
    buf_clk new_AGEMA_reg_buffer_5638 ( .C (clk), .D (new_AGEMA_signal_9102), .Q (new_AGEMA_signal_9103) ) ;
    buf_clk new_AGEMA_reg_buffer_5646 ( .C (clk), .D (new_AGEMA_signal_9110), .Q (new_AGEMA_signal_9111) ) ;
    buf_clk new_AGEMA_reg_buffer_5654 ( .C (clk), .D (new_AGEMA_signal_9118), .Q (new_AGEMA_signal_9119) ) ;
    buf_clk new_AGEMA_reg_buffer_5662 ( .C (clk), .D (new_AGEMA_signal_9126), .Q (new_AGEMA_signal_9127) ) ;
    buf_clk new_AGEMA_reg_buffer_5670 ( .C (clk), .D (new_AGEMA_signal_9134), .Q (new_AGEMA_signal_9135) ) ;
    buf_clk new_AGEMA_reg_buffer_5678 ( .C (clk), .D (new_AGEMA_signal_9142), .Q (new_AGEMA_signal_9143) ) ;
    buf_clk new_AGEMA_reg_buffer_5686 ( .C (clk), .D (new_AGEMA_signal_9150), .Q (new_AGEMA_signal_9151) ) ;
    buf_clk new_AGEMA_reg_buffer_5694 ( .C (clk), .D (new_AGEMA_signal_9158), .Q (new_AGEMA_signal_9159) ) ;
    buf_clk new_AGEMA_reg_buffer_5702 ( .C (clk), .D (new_AGEMA_signal_9166), .Q (new_AGEMA_signal_9167) ) ;
    buf_clk new_AGEMA_reg_buffer_5710 ( .C (clk), .D (new_AGEMA_signal_9174), .Q (new_AGEMA_signal_9175) ) ;
    buf_clk new_AGEMA_reg_buffer_5718 ( .C (clk), .D (new_AGEMA_signal_9182), .Q (new_AGEMA_signal_9183) ) ;
    buf_clk new_AGEMA_reg_buffer_5726 ( .C (clk), .D (new_AGEMA_signal_9190), .Q (new_AGEMA_signal_9191) ) ;
    buf_clk new_AGEMA_reg_buffer_5734 ( .C (clk), .D (new_AGEMA_signal_9198), .Q (new_AGEMA_signal_9199) ) ;
    buf_clk new_AGEMA_reg_buffer_5742 ( .C (clk), .D (new_AGEMA_signal_9206), .Q (new_AGEMA_signal_9207) ) ;
    buf_clk new_AGEMA_reg_buffer_5750 ( .C (clk), .D (new_AGEMA_signal_9214), .Q (new_AGEMA_signal_9215) ) ;
    buf_clk new_AGEMA_reg_buffer_5758 ( .C (clk), .D (new_AGEMA_signal_9222), .Q (new_AGEMA_signal_9223) ) ;
    buf_clk new_AGEMA_reg_buffer_5766 ( .C (clk), .D (new_AGEMA_signal_9230), .Q (new_AGEMA_signal_9231) ) ;
    buf_clk new_AGEMA_reg_buffer_5774 ( .C (clk), .D (new_AGEMA_signal_9238), .Q (new_AGEMA_signal_9239) ) ;
    buf_clk new_AGEMA_reg_buffer_5782 ( .C (clk), .D (new_AGEMA_signal_9246), .Q (new_AGEMA_signal_9247) ) ;
    buf_clk new_AGEMA_reg_buffer_5790 ( .C (clk), .D (new_AGEMA_signal_9254), .Q (new_AGEMA_signal_9255) ) ;
    buf_clk new_AGEMA_reg_buffer_5798 ( .C (clk), .D (new_AGEMA_signal_9262), .Q (new_AGEMA_signal_9263) ) ;
    buf_clk new_AGEMA_reg_buffer_5806 ( .C (clk), .D (new_AGEMA_signal_9270), .Q (new_AGEMA_signal_9271) ) ;
    buf_clk new_AGEMA_reg_buffer_5814 ( .C (clk), .D (new_AGEMA_signal_9278), .Q (new_AGEMA_signal_9279) ) ;
    buf_clk new_AGEMA_reg_buffer_5822 ( .C (clk), .D (new_AGEMA_signal_9286), .Q (new_AGEMA_signal_9287) ) ;
    buf_clk new_AGEMA_reg_buffer_5830 ( .C (clk), .D (new_AGEMA_signal_9294), .Q (new_AGEMA_signal_9295) ) ;
    buf_clk new_AGEMA_reg_buffer_5838 ( .C (clk), .D (new_AGEMA_signal_9302), .Q (new_AGEMA_signal_9303) ) ;
    buf_clk new_AGEMA_reg_buffer_5846 ( .C (clk), .D (new_AGEMA_signal_9310), .Q (new_AGEMA_signal_9311) ) ;
    buf_clk new_AGEMA_reg_buffer_5854 ( .C (clk), .D (new_AGEMA_signal_9318), .Q (new_AGEMA_signal_9319) ) ;
    buf_clk new_AGEMA_reg_buffer_5862 ( .C (clk), .D (new_AGEMA_signal_9326), .Q (new_AGEMA_signal_9327) ) ;
    buf_clk new_AGEMA_reg_buffer_5870 ( .C (clk), .D (new_AGEMA_signal_9334), .Q (new_AGEMA_signal_9335) ) ;
    buf_clk new_AGEMA_reg_buffer_5878 ( .C (clk), .D (new_AGEMA_signal_9342), .Q (new_AGEMA_signal_9343) ) ;
    buf_clk new_AGEMA_reg_buffer_5886 ( .C (clk), .D (new_AGEMA_signal_9350), .Q (new_AGEMA_signal_9351) ) ;
    buf_clk new_AGEMA_reg_buffer_5894 ( .C (clk), .D (new_AGEMA_signal_9358), .Q (new_AGEMA_signal_9359) ) ;
    buf_clk new_AGEMA_reg_buffer_5902 ( .C (clk), .D (new_AGEMA_signal_9366), .Q (new_AGEMA_signal_9367) ) ;
    buf_clk new_AGEMA_reg_buffer_5910 ( .C (clk), .D (new_AGEMA_signal_9374), .Q (new_AGEMA_signal_9375) ) ;
    buf_clk new_AGEMA_reg_buffer_5918 ( .C (clk), .D (new_AGEMA_signal_9382), .Q (new_AGEMA_signal_9383) ) ;
    buf_clk new_AGEMA_reg_buffer_5926 ( .C (clk), .D (new_AGEMA_signal_9390), .Q (new_AGEMA_signal_9391) ) ;
    buf_clk new_AGEMA_reg_buffer_5934 ( .C (clk), .D (new_AGEMA_signal_9398), .Q (new_AGEMA_signal_9399) ) ;
    buf_clk new_AGEMA_reg_buffer_5942 ( .C (clk), .D (new_AGEMA_signal_9406), .Q (new_AGEMA_signal_9407) ) ;
    buf_clk new_AGEMA_reg_buffer_5950 ( .C (clk), .D (new_AGEMA_signal_9414), .Q (new_AGEMA_signal_9415) ) ;
    buf_clk new_AGEMA_reg_buffer_5958 ( .C (clk), .D (new_AGEMA_signal_9422), .Q (new_AGEMA_signal_9423) ) ;
    buf_clk new_AGEMA_reg_buffer_5966 ( .C (clk), .D (new_AGEMA_signal_9430), .Q (new_AGEMA_signal_9431) ) ;
    buf_clk new_AGEMA_reg_buffer_5974 ( .C (clk), .D (new_AGEMA_signal_9438), .Q (new_AGEMA_signal_9439) ) ;
    buf_clk new_AGEMA_reg_buffer_5982 ( .C (clk), .D (new_AGEMA_signal_9446), .Q (new_AGEMA_signal_9447) ) ;
    buf_clk new_AGEMA_reg_buffer_5990 ( .C (clk), .D (new_AGEMA_signal_9454), .Q (new_AGEMA_signal_9455) ) ;
    buf_clk new_AGEMA_reg_buffer_5998 ( .C (clk), .D (new_AGEMA_signal_9462), .Q (new_AGEMA_signal_9463) ) ;
    buf_clk new_AGEMA_reg_buffer_6006 ( .C (clk), .D (new_AGEMA_signal_9470), .Q (new_AGEMA_signal_9471) ) ;
    buf_clk new_AGEMA_reg_buffer_6014 ( .C (clk), .D (new_AGEMA_signal_9478), .Q (new_AGEMA_signal_9479) ) ;
    buf_clk new_AGEMA_reg_buffer_6022 ( .C (clk), .D (new_AGEMA_signal_9486), .Q (new_AGEMA_signal_9487) ) ;
    buf_clk new_AGEMA_reg_buffer_6030 ( .C (clk), .D (new_AGEMA_signal_9494), .Q (new_AGEMA_signal_9495) ) ;
    buf_clk new_AGEMA_reg_buffer_6038 ( .C (clk), .D (new_AGEMA_signal_9502), .Q (new_AGEMA_signal_9503) ) ;
    buf_clk new_AGEMA_reg_buffer_6046 ( .C (clk), .D (new_AGEMA_signal_9510), .Q (new_AGEMA_signal_9511) ) ;
    buf_clk new_AGEMA_reg_buffer_6054 ( .C (clk), .D (new_AGEMA_signal_9518), .Q (new_AGEMA_signal_9519) ) ;
    buf_clk new_AGEMA_reg_buffer_6062 ( .C (clk), .D (new_AGEMA_signal_9526), .Q (new_AGEMA_signal_9527) ) ;
    buf_clk new_AGEMA_reg_buffer_6070 ( .C (clk), .D (new_AGEMA_signal_9534), .Q (new_AGEMA_signal_9535) ) ;
    buf_clk new_AGEMA_reg_buffer_6078 ( .C (clk), .D (new_AGEMA_signal_9542), .Q (new_AGEMA_signal_9543) ) ;
    buf_clk new_AGEMA_reg_buffer_6086 ( .C (clk), .D (new_AGEMA_signal_9550), .Q (new_AGEMA_signal_9551) ) ;
    buf_clk new_AGEMA_reg_buffer_6094 ( .C (clk), .D (new_AGEMA_signal_9558), .Q (new_AGEMA_signal_9559) ) ;
    buf_clk new_AGEMA_reg_buffer_6102 ( .C (clk), .D (new_AGEMA_signal_9566), .Q (new_AGEMA_signal_9567) ) ;
    buf_clk new_AGEMA_reg_buffer_6110 ( .C (clk), .D (new_AGEMA_signal_9574), .Q (new_AGEMA_signal_9575) ) ;
    buf_clk new_AGEMA_reg_buffer_6118 ( .C (clk), .D (new_AGEMA_signal_9582), .Q (new_AGEMA_signal_9583) ) ;
    buf_clk new_AGEMA_reg_buffer_6126 ( .C (clk), .D (new_AGEMA_signal_9590), .Q (new_AGEMA_signal_9591) ) ;
    buf_clk new_AGEMA_reg_buffer_6134 ( .C (clk), .D (new_AGEMA_signal_9598), .Q (new_AGEMA_signal_9599) ) ;
    buf_clk new_AGEMA_reg_buffer_6142 ( .C (clk), .D (new_AGEMA_signal_9606), .Q (new_AGEMA_signal_9607) ) ;
    buf_clk new_AGEMA_reg_buffer_6150 ( .C (clk), .D (new_AGEMA_signal_9614), .Q (new_AGEMA_signal_9615) ) ;
    buf_clk new_AGEMA_reg_buffer_6158 ( .C (clk), .D (new_AGEMA_signal_9622), .Q (new_AGEMA_signal_9623) ) ;
    buf_clk new_AGEMA_reg_buffer_6166 ( .C (clk), .D (new_AGEMA_signal_9630), .Q (new_AGEMA_signal_9631) ) ;
    buf_clk new_AGEMA_reg_buffer_6464 ( .C (clk), .D (new_AGEMA_signal_9928), .Q (new_AGEMA_signal_9929) ) ;
    buf_clk new_AGEMA_reg_buffer_6472 ( .C (clk), .D (new_AGEMA_signal_9936), .Q (new_AGEMA_signal_9937) ) ;
    buf_clk new_AGEMA_reg_buffer_6480 ( .C (clk), .D (new_AGEMA_signal_9944), .Q (new_AGEMA_signal_9945) ) ;
    buf_clk new_AGEMA_reg_buffer_6488 ( .C (clk), .D (new_AGEMA_signal_9952), .Q (new_AGEMA_signal_9953) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_1321 ( .C (clk), .D (new_AGEMA_signal_4786), .Q (new_AGEMA_signal_4787) ) ;
    buf_clk new_AGEMA_reg_buffer_1841 ( .C (clk), .D (new_AGEMA_signal_5305), .Q (new_AGEMA_signal_5306) ) ;
    buf_clk new_AGEMA_reg_buffer_1847 ( .C (clk), .D (new_AGEMA_signal_5311), .Q (new_AGEMA_signal_5312) ) ;
    buf_clk new_AGEMA_reg_buffer_1853 ( .C (clk), .D (new_AGEMA_signal_5317), .Q (new_AGEMA_signal_5318) ) ;
    buf_clk new_AGEMA_reg_buffer_1859 ( .C (clk), .D (new_AGEMA_signal_5323), .Q (new_AGEMA_signal_5324) ) ;
    buf_clk new_AGEMA_reg_buffer_1865 ( .C (clk), .D (new_AGEMA_signal_5329), .Q (new_AGEMA_signal_5330) ) ;
    buf_clk new_AGEMA_reg_buffer_1871 ( .C (clk), .D (new_AGEMA_signal_5335), .Q (new_AGEMA_signal_5336) ) ;
    buf_clk new_AGEMA_reg_buffer_1877 ( .C (clk), .D (new_AGEMA_signal_5341), .Q (new_AGEMA_signal_5342) ) ;
    buf_clk new_AGEMA_reg_buffer_1883 ( .C (clk), .D (new_AGEMA_signal_5347), .Q (new_AGEMA_signal_5348) ) ;
    buf_clk new_AGEMA_reg_buffer_1889 ( .C (clk), .D (new_AGEMA_signal_5353), .Q (new_AGEMA_signal_5354) ) ;
    buf_clk new_AGEMA_reg_buffer_1895 ( .C (clk), .D (new_AGEMA_signal_5359), .Q (new_AGEMA_signal_5360) ) ;
    buf_clk new_AGEMA_reg_buffer_1901 ( .C (clk), .D (new_AGEMA_signal_5365), .Q (new_AGEMA_signal_5366) ) ;
    buf_clk new_AGEMA_reg_buffer_1907 ( .C (clk), .D (new_AGEMA_signal_5371), .Q (new_AGEMA_signal_5372) ) ;
    buf_clk new_AGEMA_reg_buffer_1913 ( .C (clk), .D (new_AGEMA_signal_5377), .Q (new_AGEMA_signal_5378) ) ;
    buf_clk new_AGEMA_reg_buffer_1919 ( .C (clk), .D (new_AGEMA_signal_5383), .Q (new_AGEMA_signal_5384) ) ;
    buf_clk new_AGEMA_reg_buffer_1925 ( .C (clk), .D (new_AGEMA_signal_5389), .Q (new_AGEMA_signal_5390) ) ;
    buf_clk new_AGEMA_reg_buffer_1931 ( .C (clk), .D (new_AGEMA_signal_5395), .Q (new_AGEMA_signal_5396) ) ;
    buf_clk new_AGEMA_reg_buffer_1937 ( .C (clk), .D (new_AGEMA_signal_5401), .Q (new_AGEMA_signal_5402) ) ;
    buf_clk new_AGEMA_reg_buffer_1943 ( .C (clk), .D (new_AGEMA_signal_5407), .Q (new_AGEMA_signal_5408) ) ;
    buf_clk new_AGEMA_reg_buffer_1949 ( .C (clk), .D (new_AGEMA_signal_5413), .Q (new_AGEMA_signal_5414) ) ;
    buf_clk new_AGEMA_reg_buffer_1955 ( .C (clk), .D (new_AGEMA_signal_5419), .Q (new_AGEMA_signal_5420) ) ;
    buf_clk new_AGEMA_reg_buffer_1961 ( .C (clk), .D (new_AGEMA_signal_5425), .Q (new_AGEMA_signal_5426) ) ;
    buf_clk new_AGEMA_reg_buffer_1967 ( .C (clk), .D (new_AGEMA_signal_5431), .Q (new_AGEMA_signal_5432) ) ;
    buf_clk new_AGEMA_reg_buffer_1973 ( .C (clk), .D (new_AGEMA_signal_5437), .Q (new_AGEMA_signal_5438) ) ;
    buf_clk new_AGEMA_reg_buffer_1979 ( .C (clk), .D (new_AGEMA_signal_5443), .Q (new_AGEMA_signal_5444) ) ;
    buf_clk new_AGEMA_reg_buffer_1985 ( .C (clk), .D (new_AGEMA_signal_5449), .Q (new_AGEMA_signal_5450) ) ;
    buf_clk new_AGEMA_reg_buffer_1991 ( .C (clk), .D (new_AGEMA_signal_5455), .Q (new_AGEMA_signal_5456) ) ;
    buf_clk new_AGEMA_reg_buffer_1997 ( .C (clk), .D (new_AGEMA_signal_5461), .Q (new_AGEMA_signal_5462) ) ;
    buf_clk new_AGEMA_reg_buffer_2003 ( .C (clk), .D (new_AGEMA_signal_5467), .Q (new_AGEMA_signal_5468) ) ;
    buf_clk new_AGEMA_reg_buffer_2009 ( .C (clk), .D (new_AGEMA_signal_5473), .Q (new_AGEMA_signal_5474) ) ;
    buf_clk new_AGEMA_reg_buffer_2015 ( .C (clk), .D (new_AGEMA_signal_5479), .Q (new_AGEMA_signal_5480) ) ;
    buf_clk new_AGEMA_reg_buffer_2021 ( .C (clk), .D (new_AGEMA_signal_5485), .Q (new_AGEMA_signal_5486) ) ;
    buf_clk new_AGEMA_reg_buffer_2027 ( .C (clk), .D (new_AGEMA_signal_5491), .Q (new_AGEMA_signal_5492) ) ;
    buf_clk new_AGEMA_reg_buffer_2033 ( .C (clk), .D (new_AGEMA_signal_5497), .Q (new_AGEMA_signal_5498) ) ;
    buf_clk new_AGEMA_reg_buffer_2039 ( .C (clk), .D (new_AGEMA_signal_5503), .Q (new_AGEMA_signal_5504) ) ;
    buf_clk new_AGEMA_reg_buffer_2045 ( .C (clk), .D (new_AGEMA_signal_5509), .Q (new_AGEMA_signal_5510) ) ;
    buf_clk new_AGEMA_reg_buffer_2051 ( .C (clk), .D (new_AGEMA_signal_5515), .Q (new_AGEMA_signal_5516) ) ;
    buf_clk new_AGEMA_reg_buffer_2057 ( .C (clk), .D (new_AGEMA_signal_5521), .Q (new_AGEMA_signal_5522) ) ;
    buf_clk new_AGEMA_reg_buffer_2063 ( .C (clk), .D (new_AGEMA_signal_5527), .Q (new_AGEMA_signal_5528) ) ;
    buf_clk new_AGEMA_reg_buffer_2069 ( .C (clk), .D (new_AGEMA_signal_5533), .Q (new_AGEMA_signal_5534) ) ;
    buf_clk new_AGEMA_reg_buffer_2075 ( .C (clk), .D (new_AGEMA_signal_5539), .Q (new_AGEMA_signal_5540) ) ;
    buf_clk new_AGEMA_reg_buffer_2081 ( .C (clk), .D (new_AGEMA_signal_5545), .Q (new_AGEMA_signal_5546) ) ;
    buf_clk new_AGEMA_reg_buffer_2087 ( .C (clk), .D (new_AGEMA_signal_5551), .Q (new_AGEMA_signal_5552) ) ;
    buf_clk new_AGEMA_reg_buffer_2093 ( .C (clk), .D (new_AGEMA_signal_5557), .Q (new_AGEMA_signal_5558) ) ;
    buf_clk new_AGEMA_reg_buffer_2099 ( .C (clk), .D (new_AGEMA_signal_5563), .Q (new_AGEMA_signal_5564) ) ;
    buf_clk new_AGEMA_reg_buffer_2105 ( .C (clk), .D (new_AGEMA_signal_5569), .Q (new_AGEMA_signal_5570) ) ;
    buf_clk new_AGEMA_reg_buffer_2111 ( .C (clk), .D (new_AGEMA_signal_5575), .Q (new_AGEMA_signal_5576) ) ;
    buf_clk new_AGEMA_reg_buffer_2117 ( .C (clk), .D (new_AGEMA_signal_5581), .Q (new_AGEMA_signal_5582) ) ;
    buf_clk new_AGEMA_reg_buffer_2123 ( .C (clk), .D (new_AGEMA_signal_5587), .Q (new_AGEMA_signal_5588) ) ;
    buf_clk new_AGEMA_reg_buffer_2129 ( .C (clk), .D (new_AGEMA_signal_5593), .Q (new_AGEMA_signal_5594) ) ;
    buf_clk new_AGEMA_reg_buffer_2135 ( .C (clk), .D (new_AGEMA_signal_5599), .Q (new_AGEMA_signal_5600) ) ;
    buf_clk new_AGEMA_reg_buffer_2141 ( .C (clk), .D (new_AGEMA_signal_5605), .Q (new_AGEMA_signal_5606) ) ;
    buf_clk new_AGEMA_reg_buffer_2147 ( .C (clk), .D (new_AGEMA_signal_5611), .Q (new_AGEMA_signal_5612) ) ;
    buf_clk new_AGEMA_reg_buffer_2153 ( .C (clk), .D (new_AGEMA_signal_5617), .Q (new_AGEMA_signal_5618) ) ;
    buf_clk new_AGEMA_reg_buffer_2159 ( .C (clk), .D (new_AGEMA_signal_5623), .Q (new_AGEMA_signal_5624) ) ;
    buf_clk new_AGEMA_reg_buffer_2165 ( .C (clk), .D (new_AGEMA_signal_5629), .Q (new_AGEMA_signal_5630) ) ;
    buf_clk new_AGEMA_reg_buffer_2171 ( .C (clk), .D (new_AGEMA_signal_5635), .Q (new_AGEMA_signal_5636) ) ;
    buf_clk new_AGEMA_reg_buffer_2177 ( .C (clk), .D (new_AGEMA_signal_5641), .Q (new_AGEMA_signal_5642) ) ;
    buf_clk new_AGEMA_reg_buffer_2183 ( .C (clk), .D (new_AGEMA_signal_5647), .Q (new_AGEMA_signal_5648) ) ;
    buf_clk new_AGEMA_reg_buffer_2189 ( .C (clk), .D (new_AGEMA_signal_5653), .Q (new_AGEMA_signal_5654) ) ;
    buf_clk new_AGEMA_reg_buffer_2195 ( .C (clk), .D (new_AGEMA_signal_5659), .Q (new_AGEMA_signal_5660) ) ;
    buf_clk new_AGEMA_reg_buffer_2201 ( .C (clk), .D (new_AGEMA_signal_5665), .Q (new_AGEMA_signal_5666) ) ;
    buf_clk new_AGEMA_reg_buffer_2207 ( .C (clk), .D (new_AGEMA_signal_5671), .Q (new_AGEMA_signal_5672) ) ;
    buf_clk new_AGEMA_reg_buffer_2213 ( .C (clk), .D (new_AGEMA_signal_5677), .Q (new_AGEMA_signal_5678) ) ;
    buf_clk new_AGEMA_reg_buffer_2219 ( .C (clk), .D (new_AGEMA_signal_5683), .Q (new_AGEMA_signal_5684) ) ;
    buf_clk new_AGEMA_reg_buffer_2225 ( .C (clk), .D (new_AGEMA_signal_5689), .Q (new_AGEMA_signal_5690) ) ;
    buf_clk new_AGEMA_reg_buffer_2231 ( .C (clk), .D (new_AGEMA_signal_5695), .Q (new_AGEMA_signal_5696) ) ;
    buf_clk new_AGEMA_reg_buffer_2237 ( .C (clk), .D (new_AGEMA_signal_5701), .Q (new_AGEMA_signal_5702) ) ;
    buf_clk new_AGEMA_reg_buffer_2243 ( .C (clk), .D (new_AGEMA_signal_5707), .Q (new_AGEMA_signal_5708) ) ;
    buf_clk new_AGEMA_reg_buffer_2249 ( .C (clk), .D (new_AGEMA_signal_5713), .Q (new_AGEMA_signal_5714) ) ;
    buf_clk new_AGEMA_reg_buffer_2255 ( .C (clk), .D (new_AGEMA_signal_5719), .Q (new_AGEMA_signal_5720) ) ;
    buf_clk new_AGEMA_reg_buffer_2261 ( .C (clk), .D (new_AGEMA_signal_5725), .Q (new_AGEMA_signal_5726) ) ;
    buf_clk new_AGEMA_reg_buffer_2267 ( .C (clk), .D (new_AGEMA_signal_5731), .Q (new_AGEMA_signal_5732) ) ;
    buf_clk new_AGEMA_reg_buffer_2273 ( .C (clk), .D (new_AGEMA_signal_5737), .Q (new_AGEMA_signal_5738) ) ;
    buf_clk new_AGEMA_reg_buffer_2279 ( .C (clk), .D (new_AGEMA_signal_5743), .Q (new_AGEMA_signal_5744) ) ;
    buf_clk new_AGEMA_reg_buffer_2285 ( .C (clk), .D (new_AGEMA_signal_5749), .Q (new_AGEMA_signal_5750) ) ;
    buf_clk new_AGEMA_reg_buffer_2291 ( .C (clk), .D (new_AGEMA_signal_5755), .Q (new_AGEMA_signal_5756) ) ;
    buf_clk new_AGEMA_reg_buffer_2297 ( .C (clk), .D (new_AGEMA_signal_5761), .Q (new_AGEMA_signal_5762) ) ;
    buf_clk new_AGEMA_reg_buffer_2303 ( .C (clk), .D (new_AGEMA_signal_5767), .Q (new_AGEMA_signal_5768) ) ;
    buf_clk new_AGEMA_reg_buffer_2309 ( .C (clk), .D (new_AGEMA_signal_5773), .Q (new_AGEMA_signal_5774) ) ;
    buf_clk new_AGEMA_reg_buffer_2315 ( .C (clk), .D (new_AGEMA_signal_5779), .Q (new_AGEMA_signal_5780) ) ;
    buf_clk new_AGEMA_reg_buffer_2321 ( .C (clk), .D (new_AGEMA_signal_5785), .Q (new_AGEMA_signal_5786) ) ;
    buf_clk new_AGEMA_reg_buffer_2327 ( .C (clk), .D (new_AGEMA_signal_5791), .Q (new_AGEMA_signal_5792) ) ;
    buf_clk new_AGEMA_reg_buffer_2333 ( .C (clk), .D (new_AGEMA_signal_5797), .Q (new_AGEMA_signal_5798) ) ;
    buf_clk new_AGEMA_reg_buffer_2339 ( .C (clk), .D (new_AGEMA_signal_5803), .Q (new_AGEMA_signal_5804) ) ;
    buf_clk new_AGEMA_reg_buffer_2345 ( .C (clk), .D (new_AGEMA_signal_5809), .Q (new_AGEMA_signal_5810) ) ;
    buf_clk new_AGEMA_reg_buffer_2351 ( .C (clk), .D (new_AGEMA_signal_5815), .Q (new_AGEMA_signal_5816) ) ;
    buf_clk new_AGEMA_reg_buffer_2357 ( .C (clk), .D (new_AGEMA_signal_5821), .Q (new_AGEMA_signal_5822) ) ;
    buf_clk new_AGEMA_reg_buffer_2363 ( .C (clk), .D (new_AGEMA_signal_5827), .Q (new_AGEMA_signal_5828) ) ;
    buf_clk new_AGEMA_reg_buffer_2369 ( .C (clk), .D (new_AGEMA_signal_5833), .Q (new_AGEMA_signal_5834) ) ;
    buf_clk new_AGEMA_reg_buffer_2375 ( .C (clk), .D (new_AGEMA_signal_5839), .Q (new_AGEMA_signal_5840) ) ;
    buf_clk new_AGEMA_reg_buffer_2381 ( .C (clk), .D (new_AGEMA_signal_5845), .Q (new_AGEMA_signal_5846) ) ;
    buf_clk new_AGEMA_reg_buffer_2387 ( .C (clk), .D (new_AGEMA_signal_5851), .Q (new_AGEMA_signal_5852) ) ;
    buf_clk new_AGEMA_reg_buffer_2393 ( .C (clk), .D (new_AGEMA_signal_5857), .Q (new_AGEMA_signal_5858) ) ;
    buf_clk new_AGEMA_reg_buffer_2399 ( .C (clk), .D (new_AGEMA_signal_5863), .Q (new_AGEMA_signal_5864) ) ;
    buf_clk new_AGEMA_reg_buffer_2405 ( .C (clk), .D (new_AGEMA_signal_5869), .Q (new_AGEMA_signal_5870) ) ;
    buf_clk new_AGEMA_reg_buffer_2411 ( .C (clk), .D (new_AGEMA_signal_5875), .Q (new_AGEMA_signal_5876) ) ;
    buf_clk new_AGEMA_reg_buffer_2417 ( .C (clk), .D (new_AGEMA_signal_5881), .Q (new_AGEMA_signal_5882) ) ;
    buf_clk new_AGEMA_reg_buffer_2423 ( .C (clk), .D (new_AGEMA_signal_5887), .Q (new_AGEMA_signal_5888) ) ;
    buf_clk new_AGEMA_reg_buffer_2429 ( .C (clk), .D (new_AGEMA_signal_5893), .Q (new_AGEMA_signal_5894) ) ;
    buf_clk new_AGEMA_reg_buffer_2435 ( .C (clk), .D (new_AGEMA_signal_5899), .Q (new_AGEMA_signal_5900) ) ;
    buf_clk new_AGEMA_reg_buffer_2441 ( .C (clk), .D (new_AGEMA_signal_5905), .Q (new_AGEMA_signal_5906) ) ;
    buf_clk new_AGEMA_reg_buffer_2447 ( .C (clk), .D (new_AGEMA_signal_5911), .Q (new_AGEMA_signal_5912) ) ;
    buf_clk new_AGEMA_reg_buffer_2453 ( .C (clk), .D (new_AGEMA_signal_5917), .Q (new_AGEMA_signal_5918) ) ;
    buf_clk new_AGEMA_reg_buffer_2459 ( .C (clk), .D (new_AGEMA_signal_5923), .Q (new_AGEMA_signal_5924) ) ;
    buf_clk new_AGEMA_reg_buffer_2465 ( .C (clk), .D (new_AGEMA_signal_5929), .Q (new_AGEMA_signal_5930) ) ;
    buf_clk new_AGEMA_reg_buffer_2471 ( .C (clk), .D (new_AGEMA_signal_5935), .Q (new_AGEMA_signal_5936) ) ;
    buf_clk new_AGEMA_reg_buffer_2477 ( .C (clk), .D (new_AGEMA_signal_5941), .Q (new_AGEMA_signal_5942) ) ;
    buf_clk new_AGEMA_reg_buffer_2483 ( .C (clk), .D (new_AGEMA_signal_5947), .Q (new_AGEMA_signal_5948) ) ;
    buf_clk new_AGEMA_reg_buffer_2489 ( .C (clk), .D (new_AGEMA_signal_5953), .Q (new_AGEMA_signal_5954) ) ;
    buf_clk new_AGEMA_reg_buffer_2495 ( .C (clk), .D (new_AGEMA_signal_5959), .Q (new_AGEMA_signal_5960) ) ;
    buf_clk new_AGEMA_reg_buffer_2501 ( .C (clk), .D (new_AGEMA_signal_5965), .Q (new_AGEMA_signal_5966) ) ;
    buf_clk new_AGEMA_reg_buffer_2507 ( .C (clk), .D (new_AGEMA_signal_5971), .Q (new_AGEMA_signal_5972) ) ;
    buf_clk new_AGEMA_reg_buffer_2513 ( .C (clk), .D (new_AGEMA_signal_5977), .Q (new_AGEMA_signal_5978) ) ;
    buf_clk new_AGEMA_reg_buffer_2519 ( .C (clk), .D (new_AGEMA_signal_5983), .Q (new_AGEMA_signal_5984) ) ;
    buf_clk new_AGEMA_reg_buffer_2525 ( .C (clk), .D (new_AGEMA_signal_5989), .Q (new_AGEMA_signal_5990) ) ;
    buf_clk new_AGEMA_reg_buffer_2531 ( .C (clk), .D (new_AGEMA_signal_5995), .Q (new_AGEMA_signal_5996) ) ;
    buf_clk new_AGEMA_reg_buffer_2537 ( .C (clk), .D (new_AGEMA_signal_6001), .Q (new_AGEMA_signal_6002) ) ;
    buf_clk new_AGEMA_reg_buffer_2543 ( .C (clk), .D (new_AGEMA_signal_6007), .Q (new_AGEMA_signal_6008) ) ;
    buf_clk new_AGEMA_reg_buffer_2549 ( .C (clk), .D (new_AGEMA_signal_6013), .Q (new_AGEMA_signal_6014) ) ;
    buf_clk new_AGEMA_reg_buffer_2555 ( .C (clk), .D (new_AGEMA_signal_6019), .Q (new_AGEMA_signal_6020) ) ;
    buf_clk new_AGEMA_reg_buffer_2561 ( .C (clk), .D (new_AGEMA_signal_6025), .Q (new_AGEMA_signal_6026) ) ;
    buf_clk new_AGEMA_reg_buffer_2567 ( .C (clk), .D (new_AGEMA_signal_6031), .Q (new_AGEMA_signal_6032) ) ;
    buf_clk new_AGEMA_reg_buffer_2573 ( .C (clk), .D (new_AGEMA_signal_6037), .Q (new_AGEMA_signal_6038) ) ;
    buf_clk new_AGEMA_reg_buffer_2579 ( .C (clk), .D (new_AGEMA_signal_6043), .Q (new_AGEMA_signal_6044) ) ;
    buf_clk new_AGEMA_reg_buffer_2585 ( .C (clk), .D (new_AGEMA_signal_6049), .Q (new_AGEMA_signal_6050) ) ;
    buf_clk new_AGEMA_reg_buffer_2591 ( .C (clk), .D (new_AGEMA_signal_6055), .Q (new_AGEMA_signal_6056) ) ;
    buf_clk new_AGEMA_reg_buffer_2597 ( .C (clk), .D (new_AGEMA_signal_6061), .Q (new_AGEMA_signal_6062) ) ;
    buf_clk new_AGEMA_reg_buffer_2603 ( .C (clk), .D (new_AGEMA_signal_6067), .Q (new_AGEMA_signal_6068) ) ;
    buf_clk new_AGEMA_reg_buffer_2609 ( .C (clk), .D (new_AGEMA_signal_6073), .Q (new_AGEMA_signal_6074) ) ;
    buf_clk new_AGEMA_reg_buffer_2615 ( .C (clk), .D (new_AGEMA_signal_6079), .Q (new_AGEMA_signal_6080) ) ;
    buf_clk new_AGEMA_reg_buffer_2621 ( .C (clk), .D (new_AGEMA_signal_6085), .Q (new_AGEMA_signal_6086) ) ;
    buf_clk new_AGEMA_reg_buffer_2627 ( .C (clk), .D (new_AGEMA_signal_6091), .Q (new_AGEMA_signal_6092) ) ;
    buf_clk new_AGEMA_reg_buffer_2633 ( .C (clk), .D (new_AGEMA_signal_6097), .Q (new_AGEMA_signal_6098) ) ;
    buf_clk new_AGEMA_reg_buffer_2639 ( .C (clk), .D (new_AGEMA_signal_6103), .Q (new_AGEMA_signal_6104) ) ;
    buf_clk new_AGEMA_reg_buffer_2645 ( .C (clk), .D (new_AGEMA_signal_6109), .Q (new_AGEMA_signal_6110) ) ;
    buf_clk new_AGEMA_reg_buffer_2651 ( .C (clk), .D (new_AGEMA_signal_6115), .Q (new_AGEMA_signal_6116) ) ;
    buf_clk new_AGEMA_reg_buffer_2657 ( .C (clk), .D (new_AGEMA_signal_6121), .Q (new_AGEMA_signal_6122) ) ;
    buf_clk new_AGEMA_reg_buffer_2663 ( .C (clk), .D (new_AGEMA_signal_6127), .Q (new_AGEMA_signal_6128) ) ;
    buf_clk new_AGEMA_reg_buffer_2669 ( .C (clk), .D (new_AGEMA_signal_6133), .Q (new_AGEMA_signal_6134) ) ;
    buf_clk new_AGEMA_reg_buffer_2675 ( .C (clk), .D (new_AGEMA_signal_6139), .Q (new_AGEMA_signal_6140) ) ;
    buf_clk new_AGEMA_reg_buffer_2681 ( .C (clk), .D (new_AGEMA_signal_6145), .Q (new_AGEMA_signal_6146) ) ;
    buf_clk new_AGEMA_reg_buffer_2687 ( .C (clk), .D (new_AGEMA_signal_6151), .Q (new_AGEMA_signal_6152) ) ;
    buf_clk new_AGEMA_reg_buffer_2693 ( .C (clk), .D (new_AGEMA_signal_6157), .Q (new_AGEMA_signal_6158) ) ;
    buf_clk new_AGEMA_reg_buffer_2699 ( .C (clk), .D (new_AGEMA_signal_6163), .Q (new_AGEMA_signal_6164) ) ;
    buf_clk new_AGEMA_reg_buffer_2705 ( .C (clk), .D (new_AGEMA_signal_6169), .Q (new_AGEMA_signal_6170) ) ;
    buf_clk new_AGEMA_reg_buffer_2711 ( .C (clk), .D (new_AGEMA_signal_6175), .Q (new_AGEMA_signal_6176) ) ;
    buf_clk new_AGEMA_reg_buffer_2717 ( .C (clk), .D (new_AGEMA_signal_6181), .Q (new_AGEMA_signal_6182) ) ;
    buf_clk new_AGEMA_reg_buffer_2723 ( .C (clk), .D (new_AGEMA_signal_6187), .Q (new_AGEMA_signal_6188) ) ;
    buf_clk new_AGEMA_reg_buffer_2729 ( .C (clk), .D (new_AGEMA_signal_6193), .Q (new_AGEMA_signal_6194) ) ;
    buf_clk new_AGEMA_reg_buffer_2735 ( .C (clk), .D (new_AGEMA_signal_6199), .Q (new_AGEMA_signal_6200) ) ;
    buf_clk new_AGEMA_reg_buffer_2741 ( .C (clk), .D (new_AGEMA_signal_6205), .Q (new_AGEMA_signal_6206) ) ;
    buf_clk new_AGEMA_reg_buffer_2747 ( .C (clk), .D (new_AGEMA_signal_6211), .Q (new_AGEMA_signal_6212) ) ;
    buf_clk new_AGEMA_reg_buffer_2753 ( .C (clk), .D (new_AGEMA_signal_6217), .Q (new_AGEMA_signal_6218) ) ;
    buf_clk new_AGEMA_reg_buffer_2759 ( .C (clk), .D (new_AGEMA_signal_6223), .Q (new_AGEMA_signal_6224) ) ;
    buf_clk new_AGEMA_reg_buffer_2765 ( .C (clk), .D (new_AGEMA_signal_6229), .Q (new_AGEMA_signal_6230) ) ;
    buf_clk new_AGEMA_reg_buffer_2771 ( .C (clk), .D (new_AGEMA_signal_6235), .Q (new_AGEMA_signal_6236) ) ;
    buf_clk new_AGEMA_reg_buffer_2777 ( .C (clk), .D (new_AGEMA_signal_6241), .Q (new_AGEMA_signal_6242) ) ;
    buf_clk new_AGEMA_reg_buffer_2783 ( .C (clk), .D (new_AGEMA_signal_6247), .Q (new_AGEMA_signal_6248) ) ;
    buf_clk new_AGEMA_reg_buffer_2789 ( .C (clk), .D (new_AGEMA_signal_6253), .Q (new_AGEMA_signal_6254) ) ;
    buf_clk new_AGEMA_reg_buffer_2795 ( .C (clk), .D (new_AGEMA_signal_6259), .Q (new_AGEMA_signal_6260) ) ;
    buf_clk new_AGEMA_reg_buffer_2801 ( .C (clk), .D (new_AGEMA_signal_6265), .Q (new_AGEMA_signal_6266) ) ;
    buf_clk new_AGEMA_reg_buffer_2807 ( .C (clk), .D (new_AGEMA_signal_6271), .Q (new_AGEMA_signal_6272) ) ;
    buf_clk new_AGEMA_reg_buffer_2813 ( .C (clk), .D (new_AGEMA_signal_6277), .Q (new_AGEMA_signal_6278) ) ;
    buf_clk new_AGEMA_reg_buffer_2819 ( .C (clk), .D (new_AGEMA_signal_6283), .Q (new_AGEMA_signal_6284) ) ;
    buf_clk new_AGEMA_reg_buffer_2825 ( .C (clk), .D (new_AGEMA_signal_6289), .Q (new_AGEMA_signal_6290) ) ;
    buf_clk new_AGEMA_reg_buffer_2831 ( .C (clk), .D (new_AGEMA_signal_6295), .Q (new_AGEMA_signal_6296) ) ;
    buf_clk new_AGEMA_reg_buffer_2837 ( .C (clk), .D (new_AGEMA_signal_6301), .Q (new_AGEMA_signal_6302) ) ;
    buf_clk new_AGEMA_reg_buffer_2843 ( .C (clk), .D (new_AGEMA_signal_6307), .Q (new_AGEMA_signal_6308) ) ;
    buf_clk new_AGEMA_reg_buffer_2849 ( .C (clk), .D (new_AGEMA_signal_6313), .Q (new_AGEMA_signal_6314) ) ;
    buf_clk new_AGEMA_reg_buffer_2855 ( .C (clk), .D (new_AGEMA_signal_6319), .Q (new_AGEMA_signal_6320) ) ;
    buf_clk new_AGEMA_reg_buffer_2861 ( .C (clk), .D (new_AGEMA_signal_6325), .Q (new_AGEMA_signal_6326) ) ;
    buf_clk new_AGEMA_reg_buffer_2867 ( .C (clk), .D (new_AGEMA_signal_6331), .Q (new_AGEMA_signal_6332) ) ;
    buf_clk new_AGEMA_reg_buffer_2873 ( .C (clk), .D (new_AGEMA_signal_6337), .Q (new_AGEMA_signal_6338) ) ;
    buf_clk new_AGEMA_reg_buffer_2879 ( .C (clk), .D (new_AGEMA_signal_6343), .Q (new_AGEMA_signal_6344) ) ;
    buf_clk new_AGEMA_reg_buffer_2885 ( .C (clk), .D (new_AGEMA_signal_6349), .Q (new_AGEMA_signal_6350) ) ;
    buf_clk new_AGEMA_reg_buffer_2891 ( .C (clk), .D (new_AGEMA_signal_6355), .Q (new_AGEMA_signal_6356) ) ;
    buf_clk new_AGEMA_reg_buffer_2897 ( .C (clk), .D (new_AGEMA_signal_6361), .Q (new_AGEMA_signal_6362) ) ;
    buf_clk new_AGEMA_reg_buffer_2903 ( .C (clk), .D (new_AGEMA_signal_6367), .Q (new_AGEMA_signal_6368) ) ;
    buf_clk new_AGEMA_reg_buffer_2909 ( .C (clk), .D (new_AGEMA_signal_6373), .Q (new_AGEMA_signal_6374) ) ;
    buf_clk new_AGEMA_reg_buffer_2915 ( .C (clk), .D (new_AGEMA_signal_6379), .Q (new_AGEMA_signal_6380) ) ;
    buf_clk new_AGEMA_reg_buffer_2921 ( .C (clk), .D (new_AGEMA_signal_6385), .Q (new_AGEMA_signal_6386) ) ;
    buf_clk new_AGEMA_reg_buffer_2927 ( .C (clk), .D (new_AGEMA_signal_6391), .Q (new_AGEMA_signal_6392) ) ;
    buf_clk new_AGEMA_reg_buffer_2933 ( .C (clk), .D (new_AGEMA_signal_6397), .Q (new_AGEMA_signal_6398) ) ;
    buf_clk new_AGEMA_reg_buffer_2939 ( .C (clk), .D (new_AGEMA_signal_6403), .Q (new_AGEMA_signal_6404) ) ;
    buf_clk new_AGEMA_reg_buffer_2945 ( .C (clk), .D (new_AGEMA_signal_6409), .Q (new_AGEMA_signal_6410) ) ;
    buf_clk new_AGEMA_reg_buffer_2951 ( .C (clk), .D (new_AGEMA_signal_6415), .Q (new_AGEMA_signal_6416) ) ;
    buf_clk new_AGEMA_reg_buffer_2957 ( .C (clk), .D (new_AGEMA_signal_6421), .Q (new_AGEMA_signal_6422) ) ;
    buf_clk new_AGEMA_reg_buffer_2963 ( .C (clk), .D (new_AGEMA_signal_6427), .Q (new_AGEMA_signal_6428) ) ;
    buf_clk new_AGEMA_reg_buffer_2969 ( .C (clk), .D (new_AGEMA_signal_6433), .Q (new_AGEMA_signal_6434) ) ;
    buf_clk new_AGEMA_reg_buffer_2975 ( .C (clk), .D (new_AGEMA_signal_6439), .Q (new_AGEMA_signal_6440) ) ;
    buf_clk new_AGEMA_reg_buffer_2981 ( .C (clk), .D (new_AGEMA_signal_6445), .Q (new_AGEMA_signal_6446) ) ;
    buf_clk new_AGEMA_reg_buffer_2987 ( .C (clk), .D (new_AGEMA_signal_6451), .Q (new_AGEMA_signal_6452) ) ;
    buf_clk new_AGEMA_reg_buffer_2993 ( .C (clk), .D (new_AGEMA_signal_6457), .Q (new_AGEMA_signal_6458) ) ;
    buf_clk new_AGEMA_reg_buffer_2999 ( .C (clk), .D (new_AGEMA_signal_6463), .Q (new_AGEMA_signal_6464) ) ;
    buf_clk new_AGEMA_reg_buffer_3005 ( .C (clk), .D (new_AGEMA_signal_6469), .Q (new_AGEMA_signal_6470) ) ;
    buf_clk new_AGEMA_reg_buffer_3011 ( .C (clk), .D (new_AGEMA_signal_6475), .Q (new_AGEMA_signal_6476) ) ;
    buf_clk new_AGEMA_reg_buffer_3017 ( .C (clk), .D (new_AGEMA_signal_6481), .Q (new_AGEMA_signal_6482) ) ;
    buf_clk new_AGEMA_reg_buffer_3023 ( .C (clk), .D (new_AGEMA_signal_6487), .Q (new_AGEMA_signal_6488) ) ;
    buf_clk new_AGEMA_reg_buffer_3029 ( .C (clk), .D (new_AGEMA_signal_6493), .Q (new_AGEMA_signal_6494) ) ;
    buf_clk new_AGEMA_reg_buffer_3035 ( .C (clk), .D (new_AGEMA_signal_6499), .Q (new_AGEMA_signal_6500) ) ;
    buf_clk new_AGEMA_reg_buffer_3041 ( .C (clk), .D (new_AGEMA_signal_6505), .Q (new_AGEMA_signal_6506) ) ;
    buf_clk new_AGEMA_reg_buffer_3047 ( .C (clk), .D (new_AGEMA_signal_6511), .Q (new_AGEMA_signal_6512) ) ;
    buf_clk new_AGEMA_reg_buffer_3053 ( .C (clk), .D (new_AGEMA_signal_6517), .Q (new_AGEMA_signal_6518) ) ;
    buf_clk new_AGEMA_reg_buffer_3059 ( .C (clk), .D (new_AGEMA_signal_6523), .Q (new_AGEMA_signal_6524) ) ;
    buf_clk new_AGEMA_reg_buffer_3065 ( .C (clk), .D (new_AGEMA_signal_6529), .Q (new_AGEMA_signal_6530) ) ;
    buf_clk new_AGEMA_reg_buffer_3071 ( .C (clk), .D (new_AGEMA_signal_6535), .Q (new_AGEMA_signal_6536) ) ;
    buf_clk new_AGEMA_reg_buffer_3077 ( .C (clk), .D (new_AGEMA_signal_6541), .Q (new_AGEMA_signal_6542) ) ;
    buf_clk new_AGEMA_reg_buffer_3083 ( .C (clk), .D (new_AGEMA_signal_6547), .Q (new_AGEMA_signal_6548) ) ;
    buf_clk new_AGEMA_reg_buffer_3089 ( .C (clk), .D (new_AGEMA_signal_6553), .Q (new_AGEMA_signal_6554) ) ;
    buf_clk new_AGEMA_reg_buffer_3095 ( .C (clk), .D (new_AGEMA_signal_6559), .Q (new_AGEMA_signal_6560) ) ;
    buf_clk new_AGEMA_reg_buffer_3101 ( .C (clk), .D (new_AGEMA_signal_6565), .Q (new_AGEMA_signal_6566) ) ;
    buf_clk new_AGEMA_reg_buffer_3107 ( .C (clk), .D (new_AGEMA_signal_6571), .Q (new_AGEMA_signal_6572) ) ;
    buf_clk new_AGEMA_reg_buffer_3113 ( .C (clk), .D (new_AGEMA_signal_6577), .Q (new_AGEMA_signal_6578) ) ;
    buf_clk new_AGEMA_reg_buffer_3119 ( .C (clk), .D (new_AGEMA_signal_6583), .Q (new_AGEMA_signal_6584) ) ;
    buf_clk new_AGEMA_reg_buffer_3125 ( .C (clk), .D (new_AGEMA_signal_6589), .Q (new_AGEMA_signal_6590) ) ;
    buf_clk new_AGEMA_reg_buffer_3131 ( .C (clk), .D (new_AGEMA_signal_6595), .Q (new_AGEMA_signal_6596) ) ;
    buf_clk new_AGEMA_reg_buffer_3137 ( .C (clk), .D (new_AGEMA_signal_6601), .Q (new_AGEMA_signal_6602) ) ;
    buf_clk new_AGEMA_reg_buffer_3143 ( .C (clk), .D (new_AGEMA_signal_6607), .Q (new_AGEMA_signal_6608) ) ;
    buf_clk new_AGEMA_reg_buffer_3149 ( .C (clk), .D (new_AGEMA_signal_6613), .Q (new_AGEMA_signal_6614) ) ;
    buf_clk new_AGEMA_reg_buffer_3155 ( .C (clk), .D (new_AGEMA_signal_6619), .Q (new_AGEMA_signal_6620) ) ;
    buf_clk new_AGEMA_reg_buffer_3161 ( .C (clk), .D (new_AGEMA_signal_6625), .Q (new_AGEMA_signal_6626) ) ;
    buf_clk new_AGEMA_reg_buffer_3167 ( .C (clk), .D (new_AGEMA_signal_6631), .Q (new_AGEMA_signal_6632) ) ;
    buf_clk new_AGEMA_reg_buffer_3173 ( .C (clk), .D (new_AGEMA_signal_6637), .Q (new_AGEMA_signal_6638) ) ;
    buf_clk new_AGEMA_reg_buffer_3179 ( .C (clk), .D (new_AGEMA_signal_6643), .Q (new_AGEMA_signal_6644) ) ;
    buf_clk new_AGEMA_reg_buffer_3185 ( .C (clk), .D (new_AGEMA_signal_6649), .Q (new_AGEMA_signal_6650) ) ;
    buf_clk new_AGEMA_reg_buffer_3191 ( .C (clk), .D (new_AGEMA_signal_6655), .Q (new_AGEMA_signal_6656) ) ;
    buf_clk new_AGEMA_reg_buffer_3197 ( .C (clk), .D (new_AGEMA_signal_6661), .Q (new_AGEMA_signal_6662) ) ;
    buf_clk new_AGEMA_reg_buffer_3203 ( .C (clk), .D (new_AGEMA_signal_6667), .Q (new_AGEMA_signal_6668) ) ;
    buf_clk new_AGEMA_reg_buffer_3209 ( .C (clk), .D (new_AGEMA_signal_6673), .Q (new_AGEMA_signal_6674) ) ;
    buf_clk new_AGEMA_reg_buffer_3215 ( .C (clk), .D (new_AGEMA_signal_6679), .Q (new_AGEMA_signal_6680) ) ;
    buf_clk new_AGEMA_reg_buffer_3221 ( .C (clk), .D (new_AGEMA_signal_6685), .Q (new_AGEMA_signal_6686) ) ;
    buf_clk new_AGEMA_reg_buffer_3227 ( .C (clk), .D (new_AGEMA_signal_6691), .Q (new_AGEMA_signal_6692) ) ;
    buf_clk new_AGEMA_reg_buffer_3233 ( .C (clk), .D (new_AGEMA_signal_6697), .Q (new_AGEMA_signal_6698) ) ;
    buf_clk new_AGEMA_reg_buffer_3239 ( .C (clk), .D (new_AGEMA_signal_6703), .Q (new_AGEMA_signal_6704) ) ;
    buf_clk new_AGEMA_reg_buffer_3245 ( .C (clk), .D (new_AGEMA_signal_6709), .Q (new_AGEMA_signal_6710) ) ;
    buf_clk new_AGEMA_reg_buffer_3251 ( .C (clk), .D (new_AGEMA_signal_6715), .Q (new_AGEMA_signal_6716) ) ;
    buf_clk new_AGEMA_reg_buffer_3257 ( .C (clk), .D (new_AGEMA_signal_6721), .Q (new_AGEMA_signal_6722) ) ;
    buf_clk new_AGEMA_reg_buffer_3263 ( .C (clk), .D (new_AGEMA_signal_6727), .Q (new_AGEMA_signal_6728) ) ;
    buf_clk new_AGEMA_reg_buffer_3269 ( .C (clk), .D (new_AGEMA_signal_6733), .Q (new_AGEMA_signal_6734) ) ;
    buf_clk new_AGEMA_reg_buffer_3275 ( .C (clk), .D (new_AGEMA_signal_6739), .Q (new_AGEMA_signal_6740) ) ;
    buf_clk new_AGEMA_reg_buffer_3281 ( .C (clk), .D (new_AGEMA_signal_6745), .Q (new_AGEMA_signal_6746) ) ;
    buf_clk new_AGEMA_reg_buffer_3287 ( .C (clk), .D (new_AGEMA_signal_6751), .Q (new_AGEMA_signal_6752) ) ;
    buf_clk new_AGEMA_reg_buffer_3293 ( .C (clk), .D (new_AGEMA_signal_6757), .Q (new_AGEMA_signal_6758) ) ;
    buf_clk new_AGEMA_reg_buffer_3299 ( .C (clk), .D (new_AGEMA_signal_6763), .Q (new_AGEMA_signal_6764) ) ;
    buf_clk new_AGEMA_reg_buffer_3305 ( .C (clk), .D (new_AGEMA_signal_6769), .Q (new_AGEMA_signal_6770) ) ;
    buf_clk new_AGEMA_reg_buffer_3311 ( .C (clk), .D (new_AGEMA_signal_6775), .Q (new_AGEMA_signal_6776) ) ;
    buf_clk new_AGEMA_reg_buffer_3317 ( .C (clk), .D (new_AGEMA_signal_6781), .Q (new_AGEMA_signal_6782) ) ;
    buf_clk new_AGEMA_reg_buffer_3323 ( .C (clk), .D (new_AGEMA_signal_6787), .Q (new_AGEMA_signal_6788) ) ;
    buf_clk new_AGEMA_reg_buffer_3329 ( .C (clk), .D (new_AGEMA_signal_6793), .Q (new_AGEMA_signal_6794) ) ;
    buf_clk new_AGEMA_reg_buffer_3335 ( .C (clk), .D (new_AGEMA_signal_6799), .Q (new_AGEMA_signal_6800) ) ;
    buf_clk new_AGEMA_reg_buffer_3341 ( .C (clk), .D (new_AGEMA_signal_6805), .Q (new_AGEMA_signal_6806) ) ;
    buf_clk new_AGEMA_reg_buffer_3347 ( .C (clk), .D (new_AGEMA_signal_6811), .Q (new_AGEMA_signal_6812) ) ;
    buf_clk new_AGEMA_reg_buffer_3353 ( .C (clk), .D (new_AGEMA_signal_6817), .Q (new_AGEMA_signal_6818) ) ;
    buf_clk new_AGEMA_reg_buffer_3359 ( .C (clk), .D (new_AGEMA_signal_6823), .Q (new_AGEMA_signal_6824) ) ;
    buf_clk new_AGEMA_reg_buffer_3365 ( .C (clk), .D (new_AGEMA_signal_6829), .Q (new_AGEMA_signal_6830) ) ;
    buf_clk new_AGEMA_reg_buffer_3371 ( .C (clk), .D (new_AGEMA_signal_6835), .Q (new_AGEMA_signal_6836) ) ;
    buf_clk new_AGEMA_reg_buffer_3377 ( .C (clk), .D (new_AGEMA_signal_6841), .Q (new_AGEMA_signal_6842) ) ;
    buf_clk new_AGEMA_reg_buffer_3383 ( .C (clk), .D (new_AGEMA_signal_6847), .Q (new_AGEMA_signal_6848) ) ;
    buf_clk new_AGEMA_reg_buffer_3389 ( .C (clk), .D (new_AGEMA_signal_6853), .Q (new_AGEMA_signal_6854) ) ;
    buf_clk new_AGEMA_reg_buffer_3395 ( .C (clk), .D (new_AGEMA_signal_6859), .Q (new_AGEMA_signal_6860) ) ;
    buf_clk new_AGEMA_reg_buffer_3401 ( .C (clk), .D (new_AGEMA_signal_6865), .Q (new_AGEMA_signal_6866) ) ;
    buf_clk new_AGEMA_reg_buffer_3407 ( .C (clk), .D (new_AGEMA_signal_6871), .Q (new_AGEMA_signal_6872) ) ;
    buf_clk new_AGEMA_reg_buffer_3413 ( .C (clk), .D (new_AGEMA_signal_6877), .Q (new_AGEMA_signal_6878) ) ;
    buf_clk new_AGEMA_reg_buffer_3419 ( .C (clk), .D (new_AGEMA_signal_6883), .Q (new_AGEMA_signal_6884) ) ;
    buf_clk new_AGEMA_reg_buffer_3425 ( .C (clk), .D (new_AGEMA_signal_6889), .Q (new_AGEMA_signal_6890) ) ;
    buf_clk new_AGEMA_reg_buffer_3431 ( .C (clk), .D (new_AGEMA_signal_6895), .Q (new_AGEMA_signal_6896) ) ;
    buf_clk new_AGEMA_reg_buffer_3437 ( .C (clk), .D (new_AGEMA_signal_6901), .Q (new_AGEMA_signal_6902) ) ;
    buf_clk new_AGEMA_reg_buffer_3443 ( .C (clk), .D (new_AGEMA_signal_6907), .Q (new_AGEMA_signal_6908) ) ;
    buf_clk new_AGEMA_reg_buffer_3449 ( .C (clk), .D (new_AGEMA_signal_6913), .Q (new_AGEMA_signal_6914) ) ;
    buf_clk new_AGEMA_reg_buffer_3455 ( .C (clk), .D (new_AGEMA_signal_6919), .Q (new_AGEMA_signal_6920) ) ;
    buf_clk new_AGEMA_reg_buffer_3461 ( .C (clk), .D (new_AGEMA_signal_6925), .Q (new_AGEMA_signal_6926) ) ;
    buf_clk new_AGEMA_reg_buffer_3467 ( .C (clk), .D (new_AGEMA_signal_6931), .Q (new_AGEMA_signal_6932) ) ;
    buf_clk new_AGEMA_reg_buffer_3473 ( .C (clk), .D (new_AGEMA_signal_6937), .Q (new_AGEMA_signal_6938) ) ;
    buf_clk new_AGEMA_reg_buffer_3479 ( .C (clk), .D (new_AGEMA_signal_6943), .Q (new_AGEMA_signal_6944) ) ;
    buf_clk new_AGEMA_reg_buffer_3485 ( .C (clk), .D (new_AGEMA_signal_6949), .Q (new_AGEMA_signal_6950) ) ;
    buf_clk new_AGEMA_reg_buffer_3491 ( .C (clk), .D (new_AGEMA_signal_6955), .Q (new_AGEMA_signal_6956) ) ;
    buf_clk new_AGEMA_reg_buffer_3497 ( .C (clk), .D (new_AGEMA_signal_6961), .Q (new_AGEMA_signal_6962) ) ;
    buf_clk new_AGEMA_reg_buffer_3503 ( .C (clk), .D (new_AGEMA_signal_6967), .Q (new_AGEMA_signal_6968) ) ;
    buf_clk new_AGEMA_reg_buffer_3509 ( .C (clk), .D (new_AGEMA_signal_6973), .Q (new_AGEMA_signal_6974) ) ;
    buf_clk new_AGEMA_reg_buffer_3515 ( .C (clk), .D (new_AGEMA_signal_6979), .Q (new_AGEMA_signal_6980) ) ;
    buf_clk new_AGEMA_reg_buffer_3521 ( .C (clk), .D (new_AGEMA_signal_6985), .Q (new_AGEMA_signal_6986) ) ;
    buf_clk new_AGEMA_reg_buffer_3527 ( .C (clk), .D (new_AGEMA_signal_6991), .Q (new_AGEMA_signal_6992) ) ;
    buf_clk new_AGEMA_reg_buffer_3533 ( .C (clk), .D (new_AGEMA_signal_6997), .Q (new_AGEMA_signal_6998) ) ;
    buf_clk new_AGEMA_reg_buffer_3539 ( .C (clk), .D (new_AGEMA_signal_7003), .Q (new_AGEMA_signal_7004) ) ;
    buf_clk new_AGEMA_reg_buffer_3545 ( .C (clk), .D (new_AGEMA_signal_7009), .Q (new_AGEMA_signal_7010) ) ;
    buf_clk new_AGEMA_reg_buffer_3551 ( .C (clk), .D (new_AGEMA_signal_7015), .Q (new_AGEMA_signal_7016) ) ;
    buf_clk new_AGEMA_reg_buffer_3557 ( .C (clk), .D (new_AGEMA_signal_7021), .Q (new_AGEMA_signal_7022) ) ;
    buf_clk new_AGEMA_reg_buffer_3563 ( .C (clk), .D (new_AGEMA_signal_7027), .Q (new_AGEMA_signal_7028) ) ;
    buf_clk new_AGEMA_reg_buffer_3569 ( .C (clk), .D (new_AGEMA_signal_7033), .Q (new_AGEMA_signal_7034) ) ;
    buf_clk new_AGEMA_reg_buffer_3573 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_0_n15), .Q (new_AGEMA_signal_7038) ) ;
    buf_clk new_AGEMA_reg_buffer_3575 ( .C (clk), .D (new_AGEMA_signal_2380), .Q (new_AGEMA_signal_7040) ) ;
    buf_clk new_AGEMA_reg_buffer_3577 ( .C (clk), .D (new_AGEMA_signal_2381), .Q (new_AGEMA_signal_7042) ) ;
    buf_clk new_AGEMA_reg_buffer_3579 ( .C (clk), .D (new_AGEMA_signal_4921), .Q (new_AGEMA_signal_7044) ) ;
    buf_clk new_AGEMA_reg_buffer_3581 ( .C (clk), .D (new_AGEMA_signal_4923), .Q (new_AGEMA_signal_7046) ) ;
    buf_clk new_AGEMA_reg_buffer_3583 ( .C (clk), .D (new_AGEMA_signal_4925), .Q (new_AGEMA_signal_7048) ) ;
    buf_clk new_AGEMA_reg_buffer_3585 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_0_n6), .Q (new_AGEMA_signal_7050) ) ;
    buf_clk new_AGEMA_reg_buffer_3587 ( .C (clk), .D (new_AGEMA_signal_2384), .Q (new_AGEMA_signal_7052) ) ;
    buf_clk new_AGEMA_reg_buffer_3589 ( .C (clk), .D (new_AGEMA_signal_2385), .Q (new_AGEMA_signal_7054) ) ;
    buf_clk new_AGEMA_reg_buffer_3591 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_1_n15), .Q (new_AGEMA_signal_7056) ) ;
    buf_clk new_AGEMA_reg_buffer_3593 ( .C (clk), .D (new_AGEMA_signal_2392), .Q (new_AGEMA_signal_7058) ) ;
    buf_clk new_AGEMA_reg_buffer_3595 ( .C (clk), .D (new_AGEMA_signal_2393), .Q (new_AGEMA_signal_7060) ) ;
    buf_clk new_AGEMA_reg_buffer_3597 ( .C (clk), .D (new_AGEMA_signal_4945), .Q (new_AGEMA_signal_7062) ) ;
    buf_clk new_AGEMA_reg_buffer_3599 ( .C (clk), .D (new_AGEMA_signal_4947), .Q (new_AGEMA_signal_7064) ) ;
    buf_clk new_AGEMA_reg_buffer_3601 ( .C (clk), .D (new_AGEMA_signal_4949), .Q (new_AGEMA_signal_7066) ) ;
    buf_clk new_AGEMA_reg_buffer_3603 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_1_n6), .Q (new_AGEMA_signal_7068) ) ;
    buf_clk new_AGEMA_reg_buffer_3605 ( .C (clk), .D (new_AGEMA_signal_2396), .Q (new_AGEMA_signal_7070) ) ;
    buf_clk new_AGEMA_reg_buffer_3607 ( .C (clk), .D (new_AGEMA_signal_2397), .Q (new_AGEMA_signal_7072) ) ;
    buf_clk new_AGEMA_reg_buffer_3609 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_2_n15), .Q (new_AGEMA_signal_7074) ) ;
    buf_clk new_AGEMA_reg_buffer_3611 ( .C (clk), .D (new_AGEMA_signal_2404), .Q (new_AGEMA_signal_7076) ) ;
    buf_clk new_AGEMA_reg_buffer_3613 ( .C (clk), .D (new_AGEMA_signal_2405), .Q (new_AGEMA_signal_7078) ) ;
    buf_clk new_AGEMA_reg_buffer_3615 ( .C (clk), .D (new_AGEMA_signal_4969), .Q (new_AGEMA_signal_7080) ) ;
    buf_clk new_AGEMA_reg_buffer_3617 ( .C (clk), .D (new_AGEMA_signal_4971), .Q (new_AGEMA_signal_7082) ) ;
    buf_clk new_AGEMA_reg_buffer_3619 ( .C (clk), .D (new_AGEMA_signal_4973), .Q (new_AGEMA_signal_7084) ) ;
    buf_clk new_AGEMA_reg_buffer_3621 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_2_n6), .Q (new_AGEMA_signal_7086) ) ;
    buf_clk new_AGEMA_reg_buffer_3623 ( .C (clk), .D (new_AGEMA_signal_2408), .Q (new_AGEMA_signal_7088) ) ;
    buf_clk new_AGEMA_reg_buffer_3625 ( .C (clk), .D (new_AGEMA_signal_2409), .Q (new_AGEMA_signal_7090) ) ;
    buf_clk new_AGEMA_reg_buffer_3627 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_3_n15), .Q (new_AGEMA_signal_7092) ) ;
    buf_clk new_AGEMA_reg_buffer_3629 ( .C (clk), .D (new_AGEMA_signal_2416), .Q (new_AGEMA_signal_7094) ) ;
    buf_clk new_AGEMA_reg_buffer_3631 ( .C (clk), .D (new_AGEMA_signal_2417), .Q (new_AGEMA_signal_7096) ) ;
    buf_clk new_AGEMA_reg_buffer_3633 ( .C (clk), .D (new_AGEMA_signal_4993), .Q (new_AGEMA_signal_7098) ) ;
    buf_clk new_AGEMA_reg_buffer_3635 ( .C (clk), .D (new_AGEMA_signal_4995), .Q (new_AGEMA_signal_7100) ) ;
    buf_clk new_AGEMA_reg_buffer_3637 ( .C (clk), .D (new_AGEMA_signal_4997), .Q (new_AGEMA_signal_7102) ) ;
    buf_clk new_AGEMA_reg_buffer_3639 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_3_n6), .Q (new_AGEMA_signal_7104) ) ;
    buf_clk new_AGEMA_reg_buffer_3641 ( .C (clk), .D (new_AGEMA_signal_2420), .Q (new_AGEMA_signal_7106) ) ;
    buf_clk new_AGEMA_reg_buffer_3643 ( .C (clk), .D (new_AGEMA_signal_2421), .Q (new_AGEMA_signal_7108) ) ;
    buf_clk new_AGEMA_reg_buffer_3645 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_4_n15), .Q (new_AGEMA_signal_7110) ) ;
    buf_clk new_AGEMA_reg_buffer_3647 ( .C (clk), .D (new_AGEMA_signal_2428), .Q (new_AGEMA_signal_7112) ) ;
    buf_clk new_AGEMA_reg_buffer_3649 ( .C (clk), .D (new_AGEMA_signal_2429), .Q (new_AGEMA_signal_7114) ) ;
    buf_clk new_AGEMA_reg_buffer_3651 ( .C (clk), .D (new_AGEMA_signal_5017), .Q (new_AGEMA_signal_7116) ) ;
    buf_clk new_AGEMA_reg_buffer_3653 ( .C (clk), .D (new_AGEMA_signal_5019), .Q (new_AGEMA_signal_7118) ) ;
    buf_clk new_AGEMA_reg_buffer_3655 ( .C (clk), .D (new_AGEMA_signal_5021), .Q (new_AGEMA_signal_7120) ) ;
    buf_clk new_AGEMA_reg_buffer_3657 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_4_n6), .Q (new_AGEMA_signal_7122) ) ;
    buf_clk new_AGEMA_reg_buffer_3659 ( .C (clk), .D (new_AGEMA_signal_2432), .Q (new_AGEMA_signal_7124) ) ;
    buf_clk new_AGEMA_reg_buffer_3661 ( .C (clk), .D (new_AGEMA_signal_2433), .Q (new_AGEMA_signal_7126) ) ;
    buf_clk new_AGEMA_reg_buffer_3663 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_5_n15), .Q (new_AGEMA_signal_7128) ) ;
    buf_clk new_AGEMA_reg_buffer_3665 ( .C (clk), .D (new_AGEMA_signal_2440), .Q (new_AGEMA_signal_7130) ) ;
    buf_clk new_AGEMA_reg_buffer_3667 ( .C (clk), .D (new_AGEMA_signal_2441), .Q (new_AGEMA_signal_7132) ) ;
    buf_clk new_AGEMA_reg_buffer_3669 ( .C (clk), .D (new_AGEMA_signal_5041), .Q (new_AGEMA_signal_7134) ) ;
    buf_clk new_AGEMA_reg_buffer_3671 ( .C (clk), .D (new_AGEMA_signal_5043), .Q (new_AGEMA_signal_7136) ) ;
    buf_clk new_AGEMA_reg_buffer_3673 ( .C (clk), .D (new_AGEMA_signal_5045), .Q (new_AGEMA_signal_7138) ) ;
    buf_clk new_AGEMA_reg_buffer_3675 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_5_n6), .Q (new_AGEMA_signal_7140) ) ;
    buf_clk new_AGEMA_reg_buffer_3677 ( .C (clk), .D (new_AGEMA_signal_2444), .Q (new_AGEMA_signal_7142) ) ;
    buf_clk new_AGEMA_reg_buffer_3679 ( .C (clk), .D (new_AGEMA_signal_2445), .Q (new_AGEMA_signal_7144) ) ;
    buf_clk new_AGEMA_reg_buffer_3681 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_6_n15), .Q (new_AGEMA_signal_7146) ) ;
    buf_clk new_AGEMA_reg_buffer_3683 ( .C (clk), .D (new_AGEMA_signal_2452), .Q (new_AGEMA_signal_7148) ) ;
    buf_clk new_AGEMA_reg_buffer_3685 ( .C (clk), .D (new_AGEMA_signal_2453), .Q (new_AGEMA_signal_7150) ) ;
    buf_clk new_AGEMA_reg_buffer_3687 ( .C (clk), .D (new_AGEMA_signal_5065), .Q (new_AGEMA_signal_7152) ) ;
    buf_clk new_AGEMA_reg_buffer_3689 ( .C (clk), .D (new_AGEMA_signal_5067), .Q (new_AGEMA_signal_7154) ) ;
    buf_clk new_AGEMA_reg_buffer_3691 ( .C (clk), .D (new_AGEMA_signal_5069), .Q (new_AGEMA_signal_7156) ) ;
    buf_clk new_AGEMA_reg_buffer_3693 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_6_n6), .Q (new_AGEMA_signal_7158) ) ;
    buf_clk new_AGEMA_reg_buffer_3695 ( .C (clk), .D (new_AGEMA_signal_2456), .Q (new_AGEMA_signal_7160) ) ;
    buf_clk new_AGEMA_reg_buffer_3697 ( .C (clk), .D (new_AGEMA_signal_2457), .Q (new_AGEMA_signal_7162) ) ;
    buf_clk new_AGEMA_reg_buffer_3699 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_7_n15), .Q (new_AGEMA_signal_7164) ) ;
    buf_clk new_AGEMA_reg_buffer_3701 ( .C (clk), .D (new_AGEMA_signal_2464), .Q (new_AGEMA_signal_7166) ) ;
    buf_clk new_AGEMA_reg_buffer_3703 ( .C (clk), .D (new_AGEMA_signal_2465), .Q (new_AGEMA_signal_7168) ) ;
    buf_clk new_AGEMA_reg_buffer_3705 ( .C (clk), .D (new_AGEMA_signal_5089), .Q (new_AGEMA_signal_7170) ) ;
    buf_clk new_AGEMA_reg_buffer_3707 ( .C (clk), .D (new_AGEMA_signal_5091), .Q (new_AGEMA_signal_7172) ) ;
    buf_clk new_AGEMA_reg_buffer_3709 ( .C (clk), .D (new_AGEMA_signal_5093), .Q (new_AGEMA_signal_7174) ) ;
    buf_clk new_AGEMA_reg_buffer_3711 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_7_n6), .Q (new_AGEMA_signal_7176) ) ;
    buf_clk new_AGEMA_reg_buffer_3713 ( .C (clk), .D (new_AGEMA_signal_2468), .Q (new_AGEMA_signal_7178) ) ;
    buf_clk new_AGEMA_reg_buffer_3715 ( .C (clk), .D (new_AGEMA_signal_2469), .Q (new_AGEMA_signal_7180) ) ;
    buf_clk new_AGEMA_reg_buffer_3717 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_8_n15), .Q (new_AGEMA_signal_7182) ) ;
    buf_clk new_AGEMA_reg_buffer_3719 ( .C (clk), .D (new_AGEMA_signal_2476), .Q (new_AGEMA_signal_7184) ) ;
    buf_clk new_AGEMA_reg_buffer_3721 ( .C (clk), .D (new_AGEMA_signal_2477), .Q (new_AGEMA_signal_7186) ) ;
    buf_clk new_AGEMA_reg_buffer_3723 ( .C (clk), .D (new_AGEMA_signal_5113), .Q (new_AGEMA_signal_7188) ) ;
    buf_clk new_AGEMA_reg_buffer_3725 ( .C (clk), .D (new_AGEMA_signal_5115), .Q (new_AGEMA_signal_7190) ) ;
    buf_clk new_AGEMA_reg_buffer_3727 ( .C (clk), .D (new_AGEMA_signal_5117), .Q (new_AGEMA_signal_7192) ) ;
    buf_clk new_AGEMA_reg_buffer_3729 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_8_n6), .Q (new_AGEMA_signal_7194) ) ;
    buf_clk new_AGEMA_reg_buffer_3731 ( .C (clk), .D (new_AGEMA_signal_2480), .Q (new_AGEMA_signal_7196) ) ;
    buf_clk new_AGEMA_reg_buffer_3733 ( .C (clk), .D (new_AGEMA_signal_2481), .Q (new_AGEMA_signal_7198) ) ;
    buf_clk new_AGEMA_reg_buffer_3735 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_9_n15), .Q (new_AGEMA_signal_7200) ) ;
    buf_clk new_AGEMA_reg_buffer_3737 ( .C (clk), .D (new_AGEMA_signal_2488), .Q (new_AGEMA_signal_7202) ) ;
    buf_clk new_AGEMA_reg_buffer_3739 ( .C (clk), .D (new_AGEMA_signal_2489), .Q (new_AGEMA_signal_7204) ) ;
    buf_clk new_AGEMA_reg_buffer_3741 ( .C (clk), .D (new_AGEMA_signal_5137), .Q (new_AGEMA_signal_7206) ) ;
    buf_clk new_AGEMA_reg_buffer_3743 ( .C (clk), .D (new_AGEMA_signal_5139), .Q (new_AGEMA_signal_7208) ) ;
    buf_clk new_AGEMA_reg_buffer_3745 ( .C (clk), .D (new_AGEMA_signal_5141), .Q (new_AGEMA_signal_7210) ) ;
    buf_clk new_AGEMA_reg_buffer_3747 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_9_n6), .Q (new_AGEMA_signal_7212) ) ;
    buf_clk new_AGEMA_reg_buffer_3749 ( .C (clk), .D (new_AGEMA_signal_2492), .Q (new_AGEMA_signal_7214) ) ;
    buf_clk new_AGEMA_reg_buffer_3751 ( .C (clk), .D (new_AGEMA_signal_2493), .Q (new_AGEMA_signal_7216) ) ;
    buf_clk new_AGEMA_reg_buffer_3753 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_10_n15), .Q (new_AGEMA_signal_7218) ) ;
    buf_clk new_AGEMA_reg_buffer_3755 ( .C (clk), .D (new_AGEMA_signal_2500), .Q (new_AGEMA_signal_7220) ) ;
    buf_clk new_AGEMA_reg_buffer_3757 ( .C (clk), .D (new_AGEMA_signal_2501), .Q (new_AGEMA_signal_7222) ) ;
    buf_clk new_AGEMA_reg_buffer_3759 ( .C (clk), .D (new_AGEMA_signal_5161), .Q (new_AGEMA_signal_7224) ) ;
    buf_clk new_AGEMA_reg_buffer_3761 ( .C (clk), .D (new_AGEMA_signal_5163), .Q (new_AGEMA_signal_7226) ) ;
    buf_clk new_AGEMA_reg_buffer_3763 ( .C (clk), .D (new_AGEMA_signal_5165), .Q (new_AGEMA_signal_7228) ) ;
    buf_clk new_AGEMA_reg_buffer_3765 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_10_n6), .Q (new_AGEMA_signal_7230) ) ;
    buf_clk new_AGEMA_reg_buffer_3767 ( .C (clk), .D (new_AGEMA_signal_2504), .Q (new_AGEMA_signal_7232) ) ;
    buf_clk new_AGEMA_reg_buffer_3769 ( .C (clk), .D (new_AGEMA_signal_2505), .Q (new_AGEMA_signal_7234) ) ;
    buf_clk new_AGEMA_reg_buffer_3771 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_11_n15), .Q (new_AGEMA_signal_7236) ) ;
    buf_clk new_AGEMA_reg_buffer_3773 ( .C (clk), .D (new_AGEMA_signal_2512), .Q (new_AGEMA_signal_7238) ) ;
    buf_clk new_AGEMA_reg_buffer_3775 ( .C (clk), .D (new_AGEMA_signal_2513), .Q (new_AGEMA_signal_7240) ) ;
    buf_clk new_AGEMA_reg_buffer_3777 ( .C (clk), .D (new_AGEMA_signal_5185), .Q (new_AGEMA_signal_7242) ) ;
    buf_clk new_AGEMA_reg_buffer_3779 ( .C (clk), .D (new_AGEMA_signal_5187), .Q (new_AGEMA_signal_7244) ) ;
    buf_clk new_AGEMA_reg_buffer_3781 ( .C (clk), .D (new_AGEMA_signal_5189), .Q (new_AGEMA_signal_7246) ) ;
    buf_clk new_AGEMA_reg_buffer_3783 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_11_n6), .Q (new_AGEMA_signal_7248) ) ;
    buf_clk new_AGEMA_reg_buffer_3785 ( .C (clk), .D (new_AGEMA_signal_2516), .Q (new_AGEMA_signal_7250) ) ;
    buf_clk new_AGEMA_reg_buffer_3787 ( .C (clk), .D (new_AGEMA_signal_2517), .Q (new_AGEMA_signal_7252) ) ;
    buf_clk new_AGEMA_reg_buffer_3789 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_12_n15), .Q (new_AGEMA_signal_7254) ) ;
    buf_clk new_AGEMA_reg_buffer_3791 ( .C (clk), .D (new_AGEMA_signal_2524), .Q (new_AGEMA_signal_7256) ) ;
    buf_clk new_AGEMA_reg_buffer_3793 ( .C (clk), .D (new_AGEMA_signal_2525), .Q (new_AGEMA_signal_7258) ) ;
    buf_clk new_AGEMA_reg_buffer_3795 ( .C (clk), .D (new_AGEMA_signal_5209), .Q (new_AGEMA_signal_7260) ) ;
    buf_clk new_AGEMA_reg_buffer_3797 ( .C (clk), .D (new_AGEMA_signal_5211), .Q (new_AGEMA_signal_7262) ) ;
    buf_clk new_AGEMA_reg_buffer_3799 ( .C (clk), .D (new_AGEMA_signal_5213), .Q (new_AGEMA_signal_7264) ) ;
    buf_clk new_AGEMA_reg_buffer_3801 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_12_n6), .Q (new_AGEMA_signal_7266) ) ;
    buf_clk new_AGEMA_reg_buffer_3803 ( .C (clk), .D (new_AGEMA_signal_2528), .Q (new_AGEMA_signal_7268) ) ;
    buf_clk new_AGEMA_reg_buffer_3805 ( .C (clk), .D (new_AGEMA_signal_2529), .Q (new_AGEMA_signal_7270) ) ;
    buf_clk new_AGEMA_reg_buffer_3807 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_13_n15), .Q (new_AGEMA_signal_7272) ) ;
    buf_clk new_AGEMA_reg_buffer_3809 ( .C (clk), .D (new_AGEMA_signal_2536), .Q (new_AGEMA_signal_7274) ) ;
    buf_clk new_AGEMA_reg_buffer_3811 ( .C (clk), .D (new_AGEMA_signal_2537), .Q (new_AGEMA_signal_7276) ) ;
    buf_clk new_AGEMA_reg_buffer_3813 ( .C (clk), .D (new_AGEMA_signal_5233), .Q (new_AGEMA_signal_7278) ) ;
    buf_clk new_AGEMA_reg_buffer_3815 ( .C (clk), .D (new_AGEMA_signal_5235), .Q (new_AGEMA_signal_7280) ) ;
    buf_clk new_AGEMA_reg_buffer_3817 ( .C (clk), .D (new_AGEMA_signal_5237), .Q (new_AGEMA_signal_7282) ) ;
    buf_clk new_AGEMA_reg_buffer_3819 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_13_n6), .Q (new_AGEMA_signal_7284) ) ;
    buf_clk new_AGEMA_reg_buffer_3821 ( .C (clk), .D (new_AGEMA_signal_2540), .Q (new_AGEMA_signal_7286) ) ;
    buf_clk new_AGEMA_reg_buffer_3823 ( .C (clk), .D (new_AGEMA_signal_2541), .Q (new_AGEMA_signal_7288) ) ;
    buf_clk new_AGEMA_reg_buffer_3825 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_14_n15), .Q (new_AGEMA_signal_7290) ) ;
    buf_clk new_AGEMA_reg_buffer_3827 ( .C (clk), .D (new_AGEMA_signal_2548), .Q (new_AGEMA_signal_7292) ) ;
    buf_clk new_AGEMA_reg_buffer_3829 ( .C (clk), .D (new_AGEMA_signal_2549), .Q (new_AGEMA_signal_7294) ) ;
    buf_clk new_AGEMA_reg_buffer_3831 ( .C (clk), .D (new_AGEMA_signal_5257), .Q (new_AGEMA_signal_7296) ) ;
    buf_clk new_AGEMA_reg_buffer_3833 ( .C (clk), .D (new_AGEMA_signal_5259), .Q (new_AGEMA_signal_7298) ) ;
    buf_clk new_AGEMA_reg_buffer_3835 ( .C (clk), .D (new_AGEMA_signal_5261), .Q (new_AGEMA_signal_7300) ) ;
    buf_clk new_AGEMA_reg_buffer_3837 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_14_n6), .Q (new_AGEMA_signal_7302) ) ;
    buf_clk new_AGEMA_reg_buffer_3839 ( .C (clk), .D (new_AGEMA_signal_2552), .Q (new_AGEMA_signal_7304) ) ;
    buf_clk new_AGEMA_reg_buffer_3841 ( .C (clk), .D (new_AGEMA_signal_2553), .Q (new_AGEMA_signal_7306) ) ;
    buf_clk new_AGEMA_reg_buffer_3843 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_15_n15), .Q (new_AGEMA_signal_7308) ) ;
    buf_clk new_AGEMA_reg_buffer_3845 ( .C (clk), .D (new_AGEMA_signal_2560), .Q (new_AGEMA_signal_7310) ) ;
    buf_clk new_AGEMA_reg_buffer_3847 ( .C (clk), .D (new_AGEMA_signal_2561), .Q (new_AGEMA_signal_7312) ) ;
    buf_clk new_AGEMA_reg_buffer_3849 ( .C (clk), .D (new_AGEMA_signal_5281), .Q (new_AGEMA_signal_7314) ) ;
    buf_clk new_AGEMA_reg_buffer_3851 ( .C (clk), .D (new_AGEMA_signal_5283), .Q (new_AGEMA_signal_7316) ) ;
    buf_clk new_AGEMA_reg_buffer_3853 ( .C (clk), .D (new_AGEMA_signal_5285), .Q (new_AGEMA_signal_7318) ) ;
    buf_clk new_AGEMA_reg_buffer_3855 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_15_n6), .Q (new_AGEMA_signal_7320) ) ;
    buf_clk new_AGEMA_reg_buffer_3857 ( .C (clk), .D (new_AGEMA_signal_2564), .Q (new_AGEMA_signal_7322) ) ;
    buf_clk new_AGEMA_reg_buffer_3859 ( .C (clk), .D (new_AGEMA_signal_2565), .Q (new_AGEMA_signal_7324) ) ;
    buf_clk new_AGEMA_reg_buffer_3863 ( .C (clk), .D (new_AGEMA_signal_7327), .Q (new_AGEMA_signal_7328) ) ;
    buf_clk new_AGEMA_reg_buffer_3869 ( .C (clk), .D (new_AGEMA_signal_7333), .Q (new_AGEMA_signal_7334) ) ;
    buf_clk new_AGEMA_reg_buffer_3877 ( .C (clk), .D (new_AGEMA_signal_7341), .Q (new_AGEMA_signal_7342) ) ;
    buf_clk new_AGEMA_reg_buffer_3885 ( .C (clk), .D (new_AGEMA_signal_7349), .Q (new_AGEMA_signal_7350) ) ;
    buf_clk new_AGEMA_reg_buffer_3893 ( .C (clk), .D (new_AGEMA_signal_7357), .Q (new_AGEMA_signal_7358) ) ;
    buf_clk new_AGEMA_reg_buffer_3901 ( .C (clk), .D (new_AGEMA_signal_7365), .Q (new_AGEMA_signal_7366) ) ;
    buf_clk new_AGEMA_reg_buffer_3909 ( .C (clk), .D (new_AGEMA_signal_7373), .Q (new_AGEMA_signal_7374) ) ;
    buf_clk new_AGEMA_reg_buffer_3917 ( .C (clk), .D (new_AGEMA_signal_7381), .Q (new_AGEMA_signal_7382) ) ;
    buf_clk new_AGEMA_reg_buffer_3925 ( .C (clk), .D (new_AGEMA_signal_7389), .Q (new_AGEMA_signal_7390) ) ;
    buf_clk new_AGEMA_reg_buffer_3933 ( .C (clk), .D (new_AGEMA_signal_7397), .Q (new_AGEMA_signal_7398) ) ;
    buf_clk new_AGEMA_reg_buffer_3941 ( .C (clk), .D (new_AGEMA_signal_7405), .Q (new_AGEMA_signal_7406) ) ;
    buf_clk new_AGEMA_reg_buffer_3949 ( .C (clk), .D (new_AGEMA_signal_7413), .Q (new_AGEMA_signal_7414) ) ;
    buf_clk new_AGEMA_reg_buffer_3957 ( .C (clk), .D (new_AGEMA_signal_7421), .Q (new_AGEMA_signal_7422) ) ;
    buf_clk new_AGEMA_reg_buffer_3965 ( .C (clk), .D (new_AGEMA_signal_7429), .Q (new_AGEMA_signal_7430) ) ;
    buf_clk new_AGEMA_reg_buffer_3973 ( .C (clk), .D (new_AGEMA_signal_7437), .Q (new_AGEMA_signal_7438) ) ;
    buf_clk new_AGEMA_reg_buffer_3981 ( .C (clk), .D (new_AGEMA_signal_7445), .Q (new_AGEMA_signal_7446) ) ;
    buf_clk new_AGEMA_reg_buffer_3989 ( .C (clk), .D (new_AGEMA_signal_7453), .Q (new_AGEMA_signal_7454) ) ;
    buf_clk new_AGEMA_reg_buffer_3997 ( .C (clk), .D (new_AGEMA_signal_7461), .Q (new_AGEMA_signal_7462) ) ;
    buf_clk new_AGEMA_reg_buffer_4005 ( .C (clk), .D (new_AGEMA_signal_7469), .Q (new_AGEMA_signal_7470) ) ;
    buf_clk new_AGEMA_reg_buffer_4013 ( .C (clk), .D (new_AGEMA_signal_7477), .Q (new_AGEMA_signal_7478) ) ;
    buf_clk new_AGEMA_reg_buffer_4021 ( .C (clk), .D (new_AGEMA_signal_7485), .Q (new_AGEMA_signal_7486) ) ;
    buf_clk new_AGEMA_reg_buffer_4029 ( .C (clk), .D (new_AGEMA_signal_7493), .Q (new_AGEMA_signal_7494) ) ;
    buf_clk new_AGEMA_reg_buffer_4037 ( .C (clk), .D (new_AGEMA_signal_7501), .Q (new_AGEMA_signal_7502) ) ;
    buf_clk new_AGEMA_reg_buffer_4045 ( .C (clk), .D (new_AGEMA_signal_7509), .Q (new_AGEMA_signal_7510) ) ;
    buf_clk new_AGEMA_reg_buffer_4053 ( .C (clk), .D (new_AGEMA_signal_7517), .Q (new_AGEMA_signal_7518) ) ;
    buf_clk new_AGEMA_reg_buffer_4061 ( .C (clk), .D (new_AGEMA_signal_7525), .Q (new_AGEMA_signal_7526) ) ;
    buf_clk new_AGEMA_reg_buffer_4069 ( .C (clk), .D (new_AGEMA_signal_7533), .Q (new_AGEMA_signal_7534) ) ;
    buf_clk new_AGEMA_reg_buffer_4077 ( .C (clk), .D (new_AGEMA_signal_7541), .Q (new_AGEMA_signal_7542) ) ;
    buf_clk new_AGEMA_reg_buffer_4085 ( .C (clk), .D (new_AGEMA_signal_7549), .Q (new_AGEMA_signal_7550) ) ;
    buf_clk new_AGEMA_reg_buffer_4093 ( .C (clk), .D (new_AGEMA_signal_7557), .Q (new_AGEMA_signal_7558) ) ;
    buf_clk new_AGEMA_reg_buffer_4101 ( .C (clk), .D (new_AGEMA_signal_7565), .Q (new_AGEMA_signal_7566) ) ;
    buf_clk new_AGEMA_reg_buffer_4109 ( .C (clk), .D (new_AGEMA_signal_7573), .Q (new_AGEMA_signal_7574) ) ;
    buf_clk new_AGEMA_reg_buffer_4117 ( .C (clk), .D (new_AGEMA_signal_7581), .Q (new_AGEMA_signal_7582) ) ;
    buf_clk new_AGEMA_reg_buffer_4125 ( .C (clk), .D (new_AGEMA_signal_7589), .Q (new_AGEMA_signal_7590) ) ;
    buf_clk new_AGEMA_reg_buffer_4133 ( .C (clk), .D (new_AGEMA_signal_7597), .Q (new_AGEMA_signal_7598) ) ;
    buf_clk new_AGEMA_reg_buffer_4141 ( .C (clk), .D (new_AGEMA_signal_7605), .Q (new_AGEMA_signal_7606) ) ;
    buf_clk new_AGEMA_reg_buffer_4149 ( .C (clk), .D (new_AGEMA_signal_7613), .Q (new_AGEMA_signal_7614) ) ;
    buf_clk new_AGEMA_reg_buffer_4157 ( .C (clk), .D (new_AGEMA_signal_7621), .Q (new_AGEMA_signal_7622) ) ;
    buf_clk new_AGEMA_reg_buffer_4165 ( .C (clk), .D (new_AGEMA_signal_7629), .Q (new_AGEMA_signal_7630) ) ;
    buf_clk new_AGEMA_reg_buffer_4173 ( .C (clk), .D (new_AGEMA_signal_7637), .Q (new_AGEMA_signal_7638) ) ;
    buf_clk new_AGEMA_reg_buffer_4181 ( .C (clk), .D (new_AGEMA_signal_7645), .Q (new_AGEMA_signal_7646) ) ;
    buf_clk new_AGEMA_reg_buffer_4189 ( .C (clk), .D (new_AGEMA_signal_7653), .Q (new_AGEMA_signal_7654) ) ;
    buf_clk new_AGEMA_reg_buffer_4197 ( .C (clk), .D (new_AGEMA_signal_7661), .Q (new_AGEMA_signal_7662) ) ;
    buf_clk new_AGEMA_reg_buffer_4205 ( .C (clk), .D (new_AGEMA_signal_7669), .Q (new_AGEMA_signal_7670) ) ;
    buf_clk new_AGEMA_reg_buffer_4213 ( .C (clk), .D (new_AGEMA_signal_7677), .Q (new_AGEMA_signal_7678) ) ;
    buf_clk new_AGEMA_reg_buffer_4221 ( .C (clk), .D (new_AGEMA_signal_7685), .Q (new_AGEMA_signal_7686) ) ;
    buf_clk new_AGEMA_reg_buffer_4229 ( .C (clk), .D (new_AGEMA_signal_7693), .Q (new_AGEMA_signal_7694) ) ;
    buf_clk new_AGEMA_reg_buffer_4237 ( .C (clk), .D (new_AGEMA_signal_7701), .Q (new_AGEMA_signal_7702) ) ;
    buf_clk new_AGEMA_reg_buffer_4245 ( .C (clk), .D (new_AGEMA_signal_7709), .Q (new_AGEMA_signal_7710) ) ;
    buf_clk new_AGEMA_reg_buffer_4253 ( .C (clk), .D (new_AGEMA_signal_7717), .Q (new_AGEMA_signal_7718) ) ;
    buf_clk new_AGEMA_reg_buffer_4261 ( .C (clk), .D (new_AGEMA_signal_7725), .Q (new_AGEMA_signal_7726) ) ;
    buf_clk new_AGEMA_reg_buffer_4269 ( .C (clk), .D (new_AGEMA_signal_7733), .Q (new_AGEMA_signal_7734) ) ;
    buf_clk new_AGEMA_reg_buffer_4277 ( .C (clk), .D (new_AGEMA_signal_7741), .Q (new_AGEMA_signal_7742) ) ;
    buf_clk new_AGEMA_reg_buffer_4285 ( .C (clk), .D (new_AGEMA_signal_7749), .Q (new_AGEMA_signal_7750) ) ;
    buf_clk new_AGEMA_reg_buffer_4293 ( .C (clk), .D (new_AGEMA_signal_7757), .Q (new_AGEMA_signal_7758) ) ;
    buf_clk new_AGEMA_reg_buffer_4301 ( .C (clk), .D (new_AGEMA_signal_7765), .Q (new_AGEMA_signal_7766) ) ;
    buf_clk new_AGEMA_reg_buffer_4309 ( .C (clk), .D (new_AGEMA_signal_7773), .Q (new_AGEMA_signal_7774) ) ;
    buf_clk new_AGEMA_reg_buffer_4317 ( .C (clk), .D (new_AGEMA_signal_7781), .Q (new_AGEMA_signal_7782) ) ;
    buf_clk new_AGEMA_reg_buffer_4325 ( .C (clk), .D (new_AGEMA_signal_7789), .Q (new_AGEMA_signal_7790) ) ;
    buf_clk new_AGEMA_reg_buffer_4333 ( .C (clk), .D (new_AGEMA_signal_7797), .Q (new_AGEMA_signal_7798) ) ;
    buf_clk new_AGEMA_reg_buffer_4341 ( .C (clk), .D (new_AGEMA_signal_7805), .Q (new_AGEMA_signal_7806) ) ;
    buf_clk new_AGEMA_reg_buffer_4349 ( .C (clk), .D (new_AGEMA_signal_7813), .Q (new_AGEMA_signal_7814) ) ;
    buf_clk new_AGEMA_reg_buffer_4357 ( .C (clk), .D (new_AGEMA_signal_7821), .Q (new_AGEMA_signal_7822) ) ;
    buf_clk new_AGEMA_reg_buffer_4365 ( .C (clk), .D (new_AGEMA_signal_7829), .Q (new_AGEMA_signal_7830) ) ;
    buf_clk new_AGEMA_reg_buffer_4373 ( .C (clk), .D (new_AGEMA_signal_7837), .Q (new_AGEMA_signal_7838) ) ;
    buf_clk new_AGEMA_reg_buffer_4381 ( .C (clk), .D (new_AGEMA_signal_7845), .Q (new_AGEMA_signal_7846) ) ;
    buf_clk new_AGEMA_reg_buffer_4389 ( .C (clk), .D (new_AGEMA_signal_7853), .Q (new_AGEMA_signal_7854) ) ;
    buf_clk new_AGEMA_reg_buffer_4397 ( .C (clk), .D (new_AGEMA_signal_7861), .Q (new_AGEMA_signal_7862) ) ;
    buf_clk new_AGEMA_reg_buffer_4405 ( .C (clk), .D (new_AGEMA_signal_7869), .Q (new_AGEMA_signal_7870) ) ;
    buf_clk new_AGEMA_reg_buffer_4413 ( .C (clk), .D (new_AGEMA_signal_7877), .Q (new_AGEMA_signal_7878) ) ;
    buf_clk new_AGEMA_reg_buffer_4421 ( .C (clk), .D (new_AGEMA_signal_7885), .Q (new_AGEMA_signal_7886) ) ;
    buf_clk new_AGEMA_reg_buffer_4429 ( .C (clk), .D (new_AGEMA_signal_7893), .Q (new_AGEMA_signal_7894) ) ;
    buf_clk new_AGEMA_reg_buffer_4437 ( .C (clk), .D (new_AGEMA_signal_7901), .Q (new_AGEMA_signal_7902) ) ;
    buf_clk new_AGEMA_reg_buffer_4445 ( .C (clk), .D (new_AGEMA_signal_7909), .Q (new_AGEMA_signal_7910) ) ;
    buf_clk new_AGEMA_reg_buffer_4453 ( .C (clk), .D (new_AGEMA_signal_7917), .Q (new_AGEMA_signal_7918) ) ;
    buf_clk new_AGEMA_reg_buffer_4461 ( .C (clk), .D (new_AGEMA_signal_7925), .Q (new_AGEMA_signal_7926) ) ;
    buf_clk new_AGEMA_reg_buffer_4469 ( .C (clk), .D (new_AGEMA_signal_7933), .Q (new_AGEMA_signal_7934) ) ;
    buf_clk new_AGEMA_reg_buffer_4477 ( .C (clk), .D (new_AGEMA_signal_7941), .Q (new_AGEMA_signal_7942) ) ;
    buf_clk new_AGEMA_reg_buffer_4485 ( .C (clk), .D (new_AGEMA_signal_7949), .Q (new_AGEMA_signal_7950) ) ;
    buf_clk new_AGEMA_reg_buffer_4493 ( .C (clk), .D (new_AGEMA_signal_7957), .Q (new_AGEMA_signal_7958) ) ;
    buf_clk new_AGEMA_reg_buffer_4501 ( .C (clk), .D (new_AGEMA_signal_7965), .Q (new_AGEMA_signal_7966) ) ;
    buf_clk new_AGEMA_reg_buffer_4509 ( .C (clk), .D (new_AGEMA_signal_7973), .Q (new_AGEMA_signal_7974) ) ;
    buf_clk new_AGEMA_reg_buffer_4517 ( .C (clk), .D (new_AGEMA_signal_7981), .Q (new_AGEMA_signal_7982) ) ;
    buf_clk new_AGEMA_reg_buffer_4525 ( .C (clk), .D (new_AGEMA_signal_7989), .Q (new_AGEMA_signal_7990) ) ;
    buf_clk new_AGEMA_reg_buffer_4533 ( .C (clk), .D (new_AGEMA_signal_7997), .Q (new_AGEMA_signal_7998) ) ;
    buf_clk new_AGEMA_reg_buffer_4541 ( .C (clk), .D (new_AGEMA_signal_8005), .Q (new_AGEMA_signal_8006) ) ;
    buf_clk new_AGEMA_reg_buffer_4549 ( .C (clk), .D (new_AGEMA_signal_8013), .Q (new_AGEMA_signal_8014) ) ;
    buf_clk new_AGEMA_reg_buffer_4557 ( .C (clk), .D (new_AGEMA_signal_8021), .Q (new_AGEMA_signal_8022) ) ;
    buf_clk new_AGEMA_reg_buffer_4565 ( .C (clk), .D (new_AGEMA_signal_8029), .Q (new_AGEMA_signal_8030) ) ;
    buf_clk new_AGEMA_reg_buffer_4573 ( .C (clk), .D (new_AGEMA_signal_8037), .Q (new_AGEMA_signal_8038) ) ;
    buf_clk new_AGEMA_reg_buffer_4581 ( .C (clk), .D (new_AGEMA_signal_8045), .Q (new_AGEMA_signal_8046) ) ;
    buf_clk new_AGEMA_reg_buffer_4589 ( .C (clk), .D (new_AGEMA_signal_8053), .Q (new_AGEMA_signal_8054) ) ;
    buf_clk new_AGEMA_reg_buffer_4597 ( .C (clk), .D (new_AGEMA_signal_8061), .Q (new_AGEMA_signal_8062) ) ;
    buf_clk new_AGEMA_reg_buffer_4605 ( .C (clk), .D (new_AGEMA_signal_8069), .Q (new_AGEMA_signal_8070) ) ;
    buf_clk new_AGEMA_reg_buffer_4613 ( .C (clk), .D (new_AGEMA_signal_8077), .Q (new_AGEMA_signal_8078) ) ;
    buf_clk new_AGEMA_reg_buffer_4621 ( .C (clk), .D (new_AGEMA_signal_8085), .Q (new_AGEMA_signal_8086) ) ;
    buf_clk new_AGEMA_reg_buffer_4629 ( .C (clk), .D (new_AGEMA_signal_8093), .Q (new_AGEMA_signal_8094) ) ;
    buf_clk new_AGEMA_reg_buffer_4637 ( .C (clk), .D (new_AGEMA_signal_8101), .Q (new_AGEMA_signal_8102) ) ;
    buf_clk new_AGEMA_reg_buffer_4645 ( .C (clk), .D (new_AGEMA_signal_8109), .Q (new_AGEMA_signal_8110) ) ;
    buf_clk new_AGEMA_reg_buffer_4653 ( .C (clk), .D (new_AGEMA_signal_8117), .Q (new_AGEMA_signal_8118) ) ;
    buf_clk new_AGEMA_reg_buffer_4661 ( .C (clk), .D (new_AGEMA_signal_8125), .Q (new_AGEMA_signal_8126) ) ;
    buf_clk new_AGEMA_reg_buffer_4669 ( .C (clk), .D (new_AGEMA_signal_8133), .Q (new_AGEMA_signal_8134) ) ;
    buf_clk new_AGEMA_reg_buffer_4677 ( .C (clk), .D (new_AGEMA_signal_8141), .Q (new_AGEMA_signal_8142) ) ;
    buf_clk new_AGEMA_reg_buffer_4685 ( .C (clk), .D (new_AGEMA_signal_8149), .Q (new_AGEMA_signal_8150) ) ;
    buf_clk new_AGEMA_reg_buffer_4693 ( .C (clk), .D (new_AGEMA_signal_8157), .Q (new_AGEMA_signal_8158) ) ;
    buf_clk new_AGEMA_reg_buffer_4701 ( .C (clk), .D (new_AGEMA_signal_8165), .Q (new_AGEMA_signal_8166) ) ;
    buf_clk new_AGEMA_reg_buffer_4709 ( .C (clk), .D (new_AGEMA_signal_8173), .Q (new_AGEMA_signal_8174) ) ;
    buf_clk new_AGEMA_reg_buffer_4717 ( .C (clk), .D (new_AGEMA_signal_8181), .Q (new_AGEMA_signal_8182) ) ;
    buf_clk new_AGEMA_reg_buffer_4725 ( .C (clk), .D (new_AGEMA_signal_8189), .Q (new_AGEMA_signal_8190) ) ;
    buf_clk new_AGEMA_reg_buffer_4733 ( .C (clk), .D (new_AGEMA_signal_8197), .Q (new_AGEMA_signal_8198) ) ;
    buf_clk new_AGEMA_reg_buffer_4741 ( .C (clk), .D (new_AGEMA_signal_8205), .Q (new_AGEMA_signal_8206) ) ;
    buf_clk new_AGEMA_reg_buffer_4749 ( .C (clk), .D (new_AGEMA_signal_8213), .Q (new_AGEMA_signal_8214) ) ;
    buf_clk new_AGEMA_reg_buffer_4757 ( .C (clk), .D (new_AGEMA_signal_8221), .Q (new_AGEMA_signal_8222) ) ;
    buf_clk new_AGEMA_reg_buffer_4765 ( .C (clk), .D (new_AGEMA_signal_8229), .Q (new_AGEMA_signal_8230) ) ;
    buf_clk new_AGEMA_reg_buffer_4773 ( .C (clk), .D (new_AGEMA_signal_8237), .Q (new_AGEMA_signal_8238) ) ;
    buf_clk new_AGEMA_reg_buffer_4781 ( .C (clk), .D (new_AGEMA_signal_8245), .Q (new_AGEMA_signal_8246) ) ;
    buf_clk new_AGEMA_reg_buffer_4789 ( .C (clk), .D (new_AGEMA_signal_8253), .Q (new_AGEMA_signal_8254) ) ;
    buf_clk new_AGEMA_reg_buffer_4797 ( .C (clk), .D (new_AGEMA_signal_8261), .Q (new_AGEMA_signal_8262) ) ;
    buf_clk new_AGEMA_reg_buffer_4805 ( .C (clk), .D (new_AGEMA_signal_8269), .Q (new_AGEMA_signal_8270) ) ;
    buf_clk new_AGEMA_reg_buffer_4813 ( .C (clk), .D (new_AGEMA_signal_8277), .Q (new_AGEMA_signal_8278) ) ;
    buf_clk new_AGEMA_reg_buffer_4821 ( .C (clk), .D (new_AGEMA_signal_8285), .Q (new_AGEMA_signal_8286) ) ;
    buf_clk new_AGEMA_reg_buffer_4829 ( .C (clk), .D (new_AGEMA_signal_8293), .Q (new_AGEMA_signal_8294) ) ;
    buf_clk new_AGEMA_reg_buffer_4837 ( .C (clk), .D (new_AGEMA_signal_8301), .Q (new_AGEMA_signal_8302) ) ;
    buf_clk new_AGEMA_reg_buffer_4845 ( .C (clk), .D (new_AGEMA_signal_8309), .Q (new_AGEMA_signal_8310) ) ;
    buf_clk new_AGEMA_reg_buffer_4853 ( .C (clk), .D (new_AGEMA_signal_8317), .Q (new_AGEMA_signal_8318) ) ;
    buf_clk new_AGEMA_reg_buffer_4861 ( .C (clk), .D (new_AGEMA_signal_8325), .Q (new_AGEMA_signal_8326) ) ;
    buf_clk new_AGEMA_reg_buffer_4869 ( .C (clk), .D (new_AGEMA_signal_8333), .Q (new_AGEMA_signal_8334) ) ;
    buf_clk new_AGEMA_reg_buffer_4877 ( .C (clk), .D (new_AGEMA_signal_8341), .Q (new_AGEMA_signal_8342) ) ;
    buf_clk new_AGEMA_reg_buffer_4885 ( .C (clk), .D (new_AGEMA_signal_8349), .Q (new_AGEMA_signal_8350) ) ;
    buf_clk new_AGEMA_reg_buffer_4893 ( .C (clk), .D (new_AGEMA_signal_8357), .Q (new_AGEMA_signal_8358) ) ;
    buf_clk new_AGEMA_reg_buffer_4901 ( .C (clk), .D (new_AGEMA_signal_8365), .Q (new_AGEMA_signal_8366) ) ;
    buf_clk new_AGEMA_reg_buffer_4909 ( .C (clk), .D (new_AGEMA_signal_8373), .Q (new_AGEMA_signal_8374) ) ;
    buf_clk new_AGEMA_reg_buffer_4917 ( .C (clk), .D (new_AGEMA_signal_8381), .Q (new_AGEMA_signal_8382) ) ;
    buf_clk new_AGEMA_reg_buffer_4925 ( .C (clk), .D (new_AGEMA_signal_8389), .Q (new_AGEMA_signal_8390) ) ;
    buf_clk new_AGEMA_reg_buffer_4933 ( .C (clk), .D (new_AGEMA_signal_8397), .Q (new_AGEMA_signal_8398) ) ;
    buf_clk new_AGEMA_reg_buffer_4941 ( .C (clk), .D (new_AGEMA_signal_8405), .Q (new_AGEMA_signal_8406) ) ;
    buf_clk new_AGEMA_reg_buffer_4949 ( .C (clk), .D (new_AGEMA_signal_8413), .Q (new_AGEMA_signal_8414) ) ;
    buf_clk new_AGEMA_reg_buffer_4957 ( .C (clk), .D (new_AGEMA_signal_8421), .Q (new_AGEMA_signal_8422) ) ;
    buf_clk new_AGEMA_reg_buffer_4965 ( .C (clk), .D (new_AGEMA_signal_8429), .Q (new_AGEMA_signal_8430) ) ;
    buf_clk new_AGEMA_reg_buffer_4973 ( .C (clk), .D (new_AGEMA_signal_8437), .Q (new_AGEMA_signal_8438) ) ;
    buf_clk new_AGEMA_reg_buffer_4981 ( .C (clk), .D (new_AGEMA_signal_8445), .Q (new_AGEMA_signal_8446) ) ;
    buf_clk new_AGEMA_reg_buffer_4989 ( .C (clk), .D (new_AGEMA_signal_8453), .Q (new_AGEMA_signal_8454) ) ;
    buf_clk new_AGEMA_reg_buffer_4997 ( .C (clk), .D (new_AGEMA_signal_8461), .Q (new_AGEMA_signal_8462) ) ;
    buf_clk new_AGEMA_reg_buffer_5005 ( .C (clk), .D (new_AGEMA_signal_8469), .Q (new_AGEMA_signal_8470) ) ;
    buf_clk new_AGEMA_reg_buffer_5013 ( .C (clk), .D (new_AGEMA_signal_8477), .Q (new_AGEMA_signal_8478) ) ;
    buf_clk new_AGEMA_reg_buffer_5021 ( .C (clk), .D (new_AGEMA_signal_8485), .Q (new_AGEMA_signal_8486) ) ;
    buf_clk new_AGEMA_reg_buffer_5029 ( .C (clk), .D (new_AGEMA_signal_8493), .Q (new_AGEMA_signal_8494) ) ;
    buf_clk new_AGEMA_reg_buffer_5037 ( .C (clk), .D (new_AGEMA_signal_8501), .Q (new_AGEMA_signal_8502) ) ;
    buf_clk new_AGEMA_reg_buffer_5045 ( .C (clk), .D (new_AGEMA_signal_8509), .Q (new_AGEMA_signal_8510) ) ;
    buf_clk new_AGEMA_reg_buffer_5053 ( .C (clk), .D (new_AGEMA_signal_8517), .Q (new_AGEMA_signal_8518) ) ;
    buf_clk new_AGEMA_reg_buffer_5061 ( .C (clk), .D (new_AGEMA_signal_8525), .Q (new_AGEMA_signal_8526) ) ;
    buf_clk new_AGEMA_reg_buffer_5069 ( .C (clk), .D (new_AGEMA_signal_8533), .Q (new_AGEMA_signal_8534) ) ;
    buf_clk new_AGEMA_reg_buffer_5077 ( .C (clk), .D (new_AGEMA_signal_8541), .Q (new_AGEMA_signal_8542) ) ;
    buf_clk new_AGEMA_reg_buffer_5085 ( .C (clk), .D (new_AGEMA_signal_8549), .Q (new_AGEMA_signal_8550) ) ;
    buf_clk new_AGEMA_reg_buffer_5093 ( .C (clk), .D (new_AGEMA_signal_8557), .Q (new_AGEMA_signal_8558) ) ;
    buf_clk new_AGEMA_reg_buffer_5101 ( .C (clk), .D (new_AGEMA_signal_8565), .Q (new_AGEMA_signal_8566) ) ;
    buf_clk new_AGEMA_reg_buffer_5109 ( .C (clk), .D (new_AGEMA_signal_8573), .Q (new_AGEMA_signal_8574) ) ;
    buf_clk new_AGEMA_reg_buffer_5117 ( .C (clk), .D (new_AGEMA_signal_8581), .Q (new_AGEMA_signal_8582) ) ;
    buf_clk new_AGEMA_reg_buffer_5125 ( .C (clk), .D (new_AGEMA_signal_8589), .Q (new_AGEMA_signal_8590) ) ;
    buf_clk new_AGEMA_reg_buffer_5133 ( .C (clk), .D (new_AGEMA_signal_8597), .Q (new_AGEMA_signal_8598) ) ;
    buf_clk new_AGEMA_reg_buffer_5141 ( .C (clk), .D (new_AGEMA_signal_8605), .Q (new_AGEMA_signal_8606) ) ;
    buf_clk new_AGEMA_reg_buffer_5149 ( .C (clk), .D (new_AGEMA_signal_8613), .Q (new_AGEMA_signal_8614) ) ;
    buf_clk new_AGEMA_reg_buffer_5157 ( .C (clk), .D (new_AGEMA_signal_8621), .Q (new_AGEMA_signal_8622) ) ;
    buf_clk new_AGEMA_reg_buffer_5165 ( .C (clk), .D (new_AGEMA_signal_8629), .Q (new_AGEMA_signal_8630) ) ;
    buf_clk new_AGEMA_reg_buffer_5173 ( .C (clk), .D (new_AGEMA_signal_8637), .Q (new_AGEMA_signal_8638) ) ;
    buf_clk new_AGEMA_reg_buffer_5181 ( .C (clk), .D (new_AGEMA_signal_8645), .Q (new_AGEMA_signal_8646) ) ;
    buf_clk new_AGEMA_reg_buffer_5189 ( .C (clk), .D (new_AGEMA_signal_8653), .Q (new_AGEMA_signal_8654) ) ;
    buf_clk new_AGEMA_reg_buffer_5197 ( .C (clk), .D (new_AGEMA_signal_8661), .Q (new_AGEMA_signal_8662) ) ;
    buf_clk new_AGEMA_reg_buffer_5205 ( .C (clk), .D (new_AGEMA_signal_8669), .Q (new_AGEMA_signal_8670) ) ;
    buf_clk new_AGEMA_reg_buffer_5213 ( .C (clk), .D (new_AGEMA_signal_8677), .Q (new_AGEMA_signal_8678) ) ;
    buf_clk new_AGEMA_reg_buffer_5221 ( .C (clk), .D (new_AGEMA_signal_8685), .Q (new_AGEMA_signal_8686) ) ;
    buf_clk new_AGEMA_reg_buffer_5229 ( .C (clk), .D (new_AGEMA_signal_8693), .Q (new_AGEMA_signal_8694) ) ;
    buf_clk new_AGEMA_reg_buffer_5237 ( .C (clk), .D (new_AGEMA_signal_8701), .Q (new_AGEMA_signal_8702) ) ;
    buf_clk new_AGEMA_reg_buffer_5245 ( .C (clk), .D (new_AGEMA_signal_8709), .Q (new_AGEMA_signal_8710) ) ;
    buf_clk new_AGEMA_reg_buffer_5253 ( .C (clk), .D (new_AGEMA_signal_8717), .Q (new_AGEMA_signal_8718) ) ;
    buf_clk new_AGEMA_reg_buffer_5261 ( .C (clk), .D (new_AGEMA_signal_8725), .Q (new_AGEMA_signal_8726) ) ;
    buf_clk new_AGEMA_reg_buffer_5269 ( .C (clk), .D (new_AGEMA_signal_8733), .Q (new_AGEMA_signal_8734) ) ;
    buf_clk new_AGEMA_reg_buffer_5277 ( .C (clk), .D (new_AGEMA_signal_8741), .Q (new_AGEMA_signal_8742) ) ;
    buf_clk new_AGEMA_reg_buffer_5285 ( .C (clk), .D (new_AGEMA_signal_8749), .Q (new_AGEMA_signal_8750) ) ;
    buf_clk new_AGEMA_reg_buffer_5293 ( .C (clk), .D (new_AGEMA_signal_8757), .Q (new_AGEMA_signal_8758) ) ;
    buf_clk new_AGEMA_reg_buffer_5301 ( .C (clk), .D (new_AGEMA_signal_8765), .Q (new_AGEMA_signal_8766) ) ;
    buf_clk new_AGEMA_reg_buffer_5309 ( .C (clk), .D (new_AGEMA_signal_8773), .Q (new_AGEMA_signal_8774) ) ;
    buf_clk new_AGEMA_reg_buffer_5317 ( .C (clk), .D (new_AGEMA_signal_8781), .Q (new_AGEMA_signal_8782) ) ;
    buf_clk new_AGEMA_reg_buffer_5325 ( .C (clk), .D (new_AGEMA_signal_8789), .Q (new_AGEMA_signal_8790) ) ;
    buf_clk new_AGEMA_reg_buffer_5333 ( .C (clk), .D (new_AGEMA_signal_8797), .Q (new_AGEMA_signal_8798) ) ;
    buf_clk new_AGEMA_reg_buffer_5341 ( .C (clk), .D (new_AGEMA_signal_8805), .Q (new_AGEMA_signal_8806) ) ;
    buf_clk new_AGEMA_reg_buffer_5349 ( .C (clk), .D (new_AGEMA_signal_8813), .Q (new_AGEMA_signal_8814) ) ;
    buf_clk new_AGEMA_reg_buffer_5357 ( .C (clk), .D (new_AGEMA_signal_8821), .Q (new_AGEMA_signal_8822) ) ;
    buf_clk new_AGEMA_reg_buffer_5365 ( .C (clk), .D (new_AGEMA_signal_8829), .Q (new_AGEMA_signal_8830) ) ;
    buf_clk new_AGEMA_reg_buffer_5373 ( .C (clk), .D (new_AGEMA_signal_8837), .Q (new_AGEMA_signal_8838) ) ;
    buf_clk new_AGEMA_reg_buffer_5381 ( .C (clk), .D (new_AGEMA_signal_8845), .Q (new_AGEMA_signal_8846) ) ;
    buf_clk new_AGEMA_reg_buffer_5389 ( .C (clk), .D (new_AGEMA_signal_8853), .Q (new_AGEMA_signal_8854) ) ;
    buf_clk new_AGEMA_reg_buffer_5397 ( .C (clk), .D (new_AGEMA_signal_8861), .Q (new_AGEMA_signal_8862) ) ;
    buf_clk new_AGEMA_reg_buffer_5407 ( .C (clk), .D (new_AGEMA_signal_8871), .Q (new_AGEMA_signal_8872) ) ;
    buf_clk new_AGEMA_reg_buffer_5415 ( .C (clk), .D (new_AGEMA_signal_8879), .Q (new_AGEMA_signal_8880) ) ;
    buf_clk new_AGEMA_reg_buffer_5423 ( .C (clk), .D (new_AGEMA_signal_8887), .Q (new_AGEMA_signal_8888) ) ;
    buf_clk new_AGEMA_reg_buffer_5431 ( .C (clk), .D (new_AGEMA_signal_8895), .Q (new_AGEMA_signal_8896) ) ;
    buf_clk new_AGEMA_reg_buffer_5439 ( .C (clk), .D (new_AGEMA_signal_8903), .Q (new_AGEMA_signal_8904) ) ;
    buf_clk new_AGEMA_reg_buffer_5447 ( .C (clk), .D (new_AGEMA_signal_8911), .Q (new_AGEMA_signal_8912) ) ;
    buf_clk new_AGEMA_reg_buffer_5455 ( .C (clk), .D (new_AGEMA_signal_8919), .Q (new_AGEMA_signal_8920) ) ;
    buf_clk new_AGEMA_reg_buffer_5463 ( .C (clk), .D (new_AGEMA_signal_8927), .Q (new_AGEMA_signal_8928) ) ;
    buf_clk new_AGEMA_reg_buffer_5471 ( .C (clk), .D (new_AGEMA_signal_8935), .Q (new_AGEMA_signal_8936) ) ;
    buf_clk new_AGEMA_reg_buffer_5479 ( .C (clk), .D (new_AGEMA_signal_8943), .Q (new_AGEMA_signal_8944) ) ;
    buf_clk new_AGEMA_reg_buffer_5487 ( .C (clk), .D (new_AGEMA_signal_8951), .Q (new_AGEMA_signal_8952) ) ;
    buf_clk new_AGEMA_reg_buffer_5495 ( .C (clk), .D (new_AGEMA_signal_8959), .Q (new_AGEMA_signal_8960) ) ;
    buf_clk new_AGEMA_reg_buffer_5503 ( .C (clk), .D (new_AGEMA_signal_8967), .Q (new_AGEMA_signal_8968) ) ;
    buf_clk new_AGEMA_reg_buffer_5511 ( .C (clk), .D (new_AGEMA_signal_8975), .Q (new_AGEMA_signal_8976) ) ;
    buf_clk new_AGEMA_reg_buffer_5519 ( .C (clk), .D (new_AGEMA_signal_8983), .Q (new_AGEMA_signal_8984) ) ;
    buf_clk new_AGEMA_reg_buffer_5527 ( .C (clk), .D (new_AGEMA_signal_8991), .Q (new_AGEMA_signal_8992) ) ;
    buf_clk new_AGEMA_reg_buffer_5535 ( .C (clk), .D (new_AGEMA_signal_8999), .Q (new_AGEMA_signal_9000) ) ;
    buf_clk new_AGEMA_reg_buffer_5543 ( .C (clk), .D (new_AGEMA_signal_9007), .Q (new_AGEMA_signal_9008) ) ;
    buf_clk new_AGEMA_reg_buffer_5551 ( .C (clk), .D (new_AGEMA_signal_9015), .Q (new_AGEMA_signal_9016) ) ;
    buf_clk new_AGEMA_reg_buffer_5559 ( .C (clk), .D (new_AGEMA_signal_9023), .Q (new_AGEMA_signal_9024) ) ;
    buf_clk new_AGEMA_reg_buffer_5567 ( .C (clk), .D (new_AGEMA_signal_9031), .Q (new_AGEMA_signal_9032) ) ;
    buf_clk new_AGEMA_reg_buffer_5575 ( .C (clk), .D (new_AGEMA_signal_9039), .Q (new_AGEMA_signal_9040) ) ;
    buf_clk new_AGEMA_reg_buffer_5583 ( .C (clk), .D (new_AGEMA_signal_9047), .Q (new_AGEMA_signal_9048) ) ;
    buf_clk new_AGEMA_reg_buffer_5591 ( .C (clk), .D (new_AGEMA_signal_9055), .Q (new_AGEMA_signal_9056) ) ;
    buf_clk new_AGEMA_reg_buffer_5599 ( .C (clk), .D (new_AGEMA_signal_9063), .Q (new_AGEMA_signal_9064) ) ;
    buf_clk new_AGEMA_reg_buffer_5607 ( .C (clk), .D (new_AGEMA_signal_9071), .Q (new_AGEMA_signal_9072) ) ;
    buf_clk new_AGEMA_reg_buffer_5615 ( .C (clk), .D (new_AGEMA_signal_9079), .Q (new_AGEMA_signal_9080) ) ;
    buf_clk new_AGEMA_reg_buffer_5623 ( .C (clk), .D (new_AGEMA_signal_9087), .Q (new_AGEMA_signal_9088) ) ;
    buf_clk new_AGEMA_reg_buffer_5631 ( .C (clk), .D (new_AGEMA_signal_9095), .Q (new_AGEMA_signal_9096) ) ;
    buf_clk new_AGEMA_reg_buffer_5639 ( .C (clk), .D (new_AGEMA_signal_9103), .Q (new_AGEMA_signal_9104) ) ;
    buf_clk new_AGEMA_reg_buffer_5647 ( .C (clk), .D (new_AGEMA_signal_9111), .Q (new_AGEMA_signal_9112) ) ;
    buf_clk new_AGEMA_reg_buffer_5655 ( .C (clk), .D (new_AGEMA_signal_9119), .Q (new_AGEMA_signal_9120) ) ;
    buf_clk new_AGEMA_reg_buffer_5663 ( .C (clk), .D (new_AGEMA_signal_9127), .Q (new_AGEMA_signal_9128) ) ;
    buf_clk new_AGEMA_reg_buffer_5671 ( .C (clk), .D (new_AGEMA_signal_9135), .Q (new_AGEMA_signal_9136) ) ;
    buf_clk new_AGEMA_reg_buffer_5679 ( .C (clk), .D (new_AGEMA_signal_9143), .Q (new_AGEMA_signal_9144) ) ;
    buf_clk new_AGEMA_reg_buffer_5687 ( .C (clk), .D (new_AGEMA_signal_9151), .Q (new_AGEMA_signal_9152) ) ;
    buf_clk new_AGEMA_reg_buffer_5695 ( .C (clk), .D (new_AGEMA_signal_9159), .Q (new_AGEMA_signal_9160) ) ;
    buf_clk new_AGEMA_reg_buffer_5703 ( .C (clk), .D (new_AGEMA_signal_9167), .Q (new_AGEMA_signal_9168) ) ;
    buf_clk new_AGEMA_reg_buffer_5711 ( .C (clk), .D (new_AGEMA_signal_9175), .Q (new_AGEMA_signal_9176) ) ;
    buf_clk new_AGEMA_reg_buffer_5719 ( .C (clk), .D (new_AGEMA_signal_9183), .Q (new_AGEMA_signal_9184) ) ;
    buf_clk new_AGEMA_reg_buffer_5727 ( .C (clk), .D (new_AGEMA_signal_9191), .Q (new_AGEMA_signal_9192) ) ;
    buf_clk new_AGEMA_reg_buffer_5735 ( .C (clk), .D (new_AGEMA_signal_9199), .Q (new_AGEMA_signal_9200) ) ;
    buf_clk new_AGEMA_reg_buffer_5743 ( .C (clk), .D (new_AGEMA_signal_9207), .Q (new_AGEMA_signal_9208) ) ;
    buf_clk new_AGEMA_reg_buffer_5751 ( .C (clk), .D (new_AGEMA_signal_9215), .Q (new_AGEMA_signal_9216) ) ;
    buf_clk new_AGEMA_reg_buffer_5759 ( .C (clk), .D (new_AGEMA_signal_9223), .Q (new_AGEMA_signal_9224) ) ;
    buf_clk new_AGEMA_reg_buffer_5767 ( .C (clk), .D (new_AGEMA_signal_9231), .Q (new_AGEMA_signal_9232) ) ;
    buf_clk new_AGEMA_reg_buffer_5775 ( .C (clk), .D (new_AGEMA_signal_9239), .Q (new_AGEMA_signal_9240) ) ;
    buf_clk new_AGEMA_reg_buffer_5783 ( .C (clk), .D (new_AGEMA_signal_9247), .Q (new_AGEMA_signal_9248) ) ;
    buf_clk new_AGEMA_reg_buffer_5791 ( .C (clk), .D (new_AGEMA_signal_9255), .Q (new_AGEMA_signal_9256) ) ;
    buf_clk new_AGEMA_reg_buffer_5799 ( .C (clk), .D (new_AGEMA_signal_9263), .Q (new_AGEMA_signal_9264) ) ;
    buf_clk new_AGEMA_reg_buffer_5807 ( .C (clk), .D (new_AGEMA_signal_9271), .Q (new_AGEMA_signal_9272) ) ;
    buf_clk new_AGEMA_reg_buffer_5815 ( .C (clk), .D (new_AGEMA_signal_9279), .Q (new_AGEMA_signal_9280) ) ;
    buf_clk new_AGEMA_reg_buffer_5823 ( .C (clk), .D (new_AGEMA_signal_9287), .Q (new_AGEMA_signal_9288) ) ;
    buf_clk new_AGEMA_reg_buffer_5831 ( .C (clk), .D (new_AGEMA_signal_9295), .Q (new_AGEMA_signal_9296) ) ;
    buf_clk new_AGEMA_reg_buffer_5839 ( .C (clk), .D (new_AGEMA_signal_9303), .Q (new_AGEMA_signal_9304) ) ;
    buf_clk new_AGEMA_reg_buffer_5847 ( .C (clk), .D (new_AGEMA_signal_9311), .Q (new_AGEMA_signal_9312) ) ;
    buf_clk new_AGEMA_reg_buffer_5855 ( .C (clk), .D (new_AGEMA_signal_9319), .Q (new_AGEMA_signal_9320) ) ;
    buf_clk new_AGEMA_reg_buffer_5863 ( .C (clk), .D (new_AGEMA_signal_9327), .Q (new_AGEMA_signal_9328) ) ;
    buf_clk new_AGEMA_reg_buffer_5871 ( .C (clk), .D (new_AGEMA_signal_9335), .Q (new_AGEMA_signal_9336) ) ;
    buf_clk new_AGEMA_reg_buffer_5879 ( .C (clk), .D (new_AGEMA_signal_9343), .Q (new_AGEMA_signal_9344) ) ;
    buf_clk new_AGEMA_reg_buffer_5887 ( .C (clk), .D (new_AGEMA_signal_9351), .Q (new_AGEMA_signal_9352) ) ;
    buf_clk new_AGEMA_reg_buffer_5895 ( .C (clk), .D (new_AGEMA_signal_9359), .Q (new_AGEMA_signal_9360) ) ;
    buf_clk new_AGEMA_reg_buffer_5903 ( .C (clk), .D (new_AGEMA_signal_9367), .Q (new_AGEMA_signal_9368) ) ;
    buf_clk new_AGEMA_reg_buffer_5911 ( .C (clk), .D (new_AGEMA_signal_9375), .Q (new_AGEMA_signal_9376) ) ;
    buf_clk new_AGEMA_reg_buffer_5919 ( .C (clk), .D (new_AGEMA_signal_9383), .Q (new_AGEMA_signal_9384) ) ;
    buf_clk new_AGEMA_reg_buffer_5927 ( .C (clk), .D (new_AGEMA_signal_9391), .Q (new_AGEMA_signal_9392) ) ;
    buf_clk new_AGEMA_reg_buffer_5935 ( .C (clk), .D (new_AGEMA_signal_9399), .Q (new_AGEMA_signal_9400) ) ;
    buf_clk new_AGEMA_reg_buffer_5943 ( .C (clk), .D (new_AGEMA_signal_9407), .Q (new_AGEMA_signal_9408) ) ;
    buf_clk new_AGEMA_reg_buffer_5951 ( .C (clk), .D (new_AGEMA_signal_9415), .Q (new_AGEMA_signal_9416) ) ;
    buf_clk new_AGEMA_reg_buffer_5959 ( .C (clk), .D (new_AGEMA_signal_9423), .Q (new_AGEMA_signal_9424) ) ;
    buf_clk new_AGEMA_reg_buffer_5967 ( .C (clk), .D (new_AGEMA_signal_9431), .Q (new_AGEMA_signal_9432) ) ;
    buf_clk new_AGEMA_reg_buffer_5975 ( .C (clk), .D (new_AGEMA_signal_9439), .Q (new_AGEMA_signal_9440) ) ;
    buf_clk new_AGEMA_reg_buffer_5983 ( .C (clk), .D (new_AGEMA_signal_9447), .Q (new_AGEMA_signal_9448) ) ;
    buf_clk new_AGEMA_reg_buffer_5991 ( .C (clk), .D (new_AGEMA_signal_9455), .Q (new_AGEMA_signal_9456) ) ;
    buf_clk new_AGEMA_reg_buffer_5999 ( .C (clk), .D (new_AGEMA_signal_9463), .Q (new_AGEMA_signal_9464) ) ;
    buf_clk new_AGEMA_reg_buffer_6007 ( .C (clk), .D (new_AGEMA_signal_9471), .Q (new_AGEMA_signal_9472) ) ;
    buf_clk new_AGEMA_reg_buffer_6015 ( .C (clk), .D (new_AGEMA_signal_9479), .Q (new_AGEMA_signal_9480) ) ;
    buf_clk new_AGEMA_reg_buffer_6023 ( .C (clk), .D (new_AGEMA_signal_9487), .Q (new_AGEMA_signal_9488) ) ;
    buf_clk new_AGEMA_reg_buffer_6031 ( .C (clk), .D (new_AGEMA_signal_9495), .Q (new_AGEMA_signal_9496) ) ;
    buf_clk new_AGEMA_reg_buffer_6039 ( .C (clk), .D (new_AGEMA_signal_9503), .Q (new_AGEMA_signal_9504) ) ;
    buf_clk new_AGEMA_reg_buffer_6047 ( .C (clk), .D (new_AGEMA_signal_9511), .Q (new_AGEMA_signal_9512) ) ;
    buf_clk new_AGEMA_reg_buffer_6055 ( .C (clk), .D (new_AGEMA_signal_9519), .Q (new_AGEMA_signal_9520) ) ;
    buf_clk new_AGEMA_reg_buffer_6063 ( .C (clk), .D (new_AGEMA_signal_9527), .Q (new_AGEMA_signal_9528) ) ;
    buf_clk new_AGEMA_reg_buffer_6071 ( .C (clk), .D (new_AGEMA_signal_9535), .Q (new_AGEMA_signal_9536) ) ;
    buf_clk new_AGEMA_reg_buffer_6079 ( .C (clk), .D (new_AGEMA_signal_9543), .Q (new_AGEMA_signal_9544) ) ;
    buf_clk new_AGEMA_reg_buffer_6087 ( .C (clk), .D (new_AGEMA_signal_9551), .Q (new_AGEMA_signal_9552) ) ;
    buf_clk new_AGEMA_reg_buffer_6095 ( .C (clk), .D (new_AGEMA_signal_9559), .Q (new_AGEMA_signal_9560) ) ;
    buf_clk new_AGEMA_reg_buffer_6103 ( .C (clk), .D (new_AGEMA_signal_9567), .Q (new_AGEMA_signal_9568) ) ;
    buf_clk new_AGEMA_reg_buffer_6111 ( .C (clk), .D (new_AGEMA_signal_9575), .Q (new_AGEMA_signal_9576) ) ;
    buf_clk new_AGEMA_reg_buffer_6119 ( .C (clk), .D (new_AGEMA_signal_9583), .Q (new_AGEMA_signal_9584) ) ;
    buf_clk new_AGEMA_reg_buffer_6127 ( .C (clk), .D (new_AGEMA_signal_9591), .Q (new_AGEMA_signal_9592) ) ;
    buf_clk new_AGEMA_reg_buffer_6135 ( .C (clk), .D (new_AGEMA_signal_9599), .Q (new_AGEMA_signal_9600) ) ;
    buf_clk new_AGEMA_reg_buffer_6143 ( .C (clk), .D (new_AGEMA_signal_9607), .Q (new_AGEMA_signal_9608) ) ;
    buf_clk new_AGEMA_reg_buffer_6151 ( .C (clk), .D (new_AGEMA_signal_9615), .Q (new_AGEMA_signal_9616) ) ;
    buf_clk new_AGEMA_reg_buffer_6159 ( .C (clk), .D (new_AGEMA_signal_9623), .Q (new_AGEMA_signal_9624) ) ;
    buf_clk new_AGEMA_reg_buffer_6167 ( .C (clk), .D (new_AGEMA_signal_9631), .Q (new_AGEMA_signal_9632) ) ;
    buf_clk new_AGEMA_reg_buffer_6179 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_0_n13), .Q (new_AGEMA_signal_9644) ) ;
    buf_clk new_AGEMA_reg_buffer_6183 ( .C (clk), .D (new_AGEMA_signal_2388), .Q (new_AGEMA_signal_9648) ) ;
    buf_clk new_AGEMA_reg_buffer_6187 ( .C (clk), .D (new_AGEMA_signal_2389), .Q (new_AGEMA_signal_9652) ) ;
    buf_clk new_AGEMA_reg_buffer_6197 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_1_n13), .Q (new_AGEMA_signal_9662) ) ;
    buf_clk new_AGEMA_reg_buffer_6201 ( .C (clk), .D (new_AGEMA_signal_2400), .Q (new_AGEMA_signal_9666) ) ;
    buf_clk new_AGEMA_reg_buffer_6205 ( .C (clk), .D (new_AGEMA_signal_2401), .Q (new_AGEMA_signal_9670) ) ;
    buf_clk new_AGEMA_reg_buffer_6215 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_2_n13), .Q (new_AGEMA_signal_9680) ) ;
    buf_clk new_AGEMA_reg_buffer_6219 ( .C (clk), .D (new_AGEMA_signal_2412), .Q (new_AGEMA_signal_9684) ) ;
    buf_clk new_AGEMA_reg_buffer_6223 ( .C (clk), .D (new_AGEMA_signal_2413), .Q (new_AGEMA_signal_9688) ) ;
    buf_clk new_AGEMA_reg_buffer_6233 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_3_n13), .Q (new_AGEMA_signal_9698) ) ;
    buf_clk new_AGEMA_reg_buffer_6237 ( .C (clk), .D (new_AGEMA_signal_2424), .Q (new_AGEMA_signal_9702) ) ;
    buf_clk new_AGEMA_reg_buffer_6241 ( .C (clk), .D (new_AGEMA_signal_2425), .Q (new_AGEMA_signal_9706) ) ;
    buf_clk new_AGEMA_reg_buffer_6251 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_4_n13), .Q (new_AGEMA_signal_9716) ) ;
    buf_clk new_AGEMA_reg_buffer_6255 ( .C (clk), .D (new_AGEMA_signal_2436), .Q (new_AGEMA_signal_9720) ) ;
    buf_clk new_AGEMA_reg_buffer_6259 ( .C (clk), .D (new_AGEMA_signal_2437), .Q (new_AGEMA_signal_9724) ) ;
    buf_clk new_AGEMA_reg_buffer_6269 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_5_n13), .Q (new_AGEMA_signal_9734) ) ;
    buf_clk new_AGEMA_reg_buffer_6273 ( .C (clk), .D (new_AGEMA_signal_2448), .Q (new_AGEMA_signal_9738) ) ;
    buf_clk new_AGEMA_reg_buffer_6277 ( .C (clk), .D (new_AGEMA_signal_2449), .Q (new_AGEMA_signal_9742) ) ;
    buf_clk new_AGEMA_reg_buffer_6287 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_6_n13), .Q (new_AGEMA_signal_9752) ) ;
    buf_clk new_AGEMA_reg_buffer_6291 ( .C (clk), .D (new_AGEMA_signal_2460), .Q (new_AGEMA_signal_9756) ) ;
    buf_clk new_AGEMA_reg_buffer_6295 ( .C (clk), .D (new_AGEMA_signal_2461), .Q (new_AGEMA_signal_9760) ) ;
    buf_clk new_AGEMA_reg_buffer_6305 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_7_n13), .Q (new_AGEMA_signal_9770) ) ;
    buf_clk new_AGEMA_reg_buffer_6309 ( .C (clk), .D (new_AGEMA_signal_2472), .Q (new_AGEMA_signal_9774) ) ;
    buf_clk new_AGEMA_reg_buffer_6313 ( .C (clk), .D (new_AGEMA_signal_2473), .Q (new_AGEMA_signal_9778) ) ;
    buf_clk new_AGEMA_reg_buffer_6323 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_8_n13), .Q (new_AGEMA_signal_9788) ) ;
    buf_clk new_AGEMA_reg_buffer_6327 ( .C (clk), .D (new_AGEMA_signal_2484), .Q (new_AGEMA_signal_9792) ) ;
    buf_clk new_AGEMA_reg_buffer_6331 ( .C (clk), .D (new_AGEMA_signal_2485), .Q (new_AGEMA_signal_9796) ) ;
    buf_clk new_AGEMA_reg_buffer_6341 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_9_n13), .Q (new_AGEMA_signal_9806) ) ;
    buf_clk new_AGEMA_reg_buffer_6345 ( .C (clk), .D (new_AGEMA_signal_2496), .Q (new_AGEMA_signal_9810) ) ;
    buf_clk new_AGEMA_reg_buffer_6349 ( .C (clk), .D (new_AGEMA_signal_2497), .Q (new_AGEMA_signal_9814) ) ;
    buf_clk new_AGEMA_reg_buffer_6359 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_10_n13), .Q (new_AGEMA_signal_9824) ) ;
    buf_clk new_AGEMA_reg_buffer_6363 ( .C (clk), .D (new_AGEMA_signal_2508), .Q (new_AGEMA_signal_9828) ) ;
    buf_clk new_AGEMA_reg_buffer_6367 ( .C (clk), .D (new_AGEMA_signal_2509), .Q (new_AGEMA_signal_9832) ) ;
    buf_clk new_AGEMA_reg_buffer_6377 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_11_n13), .Q (new_AGEMA_signal_9842) ) ;
    buf_clk new_AGEMA_reg_buffer_6381 ( .C (clk), .D (new_AGEMA_signal_2520), .Q (new_AGEMA_signal_9846) ) ;
    buf_clk new_AGEMA_reg_buffer_6385 ( .C (clk), .D (new_AGEMA_signal_2521), .Q (new_AGEMA_signal_9850) ) ;
    buf_clk new_AGEMA_reg_buffer_6395 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_12_n13), .Q (new_AGEMA_signal_9860) ) ;
    buf_clk new_AGEMA_reg_buffer_6399 ( .C (clk), .D (new_AGEMA_signal_2532), .Q (new_AGEMA_signal_9864) ) ;
    buf_clk new_AGEMA_reg_buffer_6403 ( .C (clk), .D (new_AGEMA_signal_2533), .Q (new_AGEMA_signal_9868) ) ;
    buf_clk new_AGEMA_reg_buffer_6413 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_13_n13), .Q (new_AGEMA_signal_9878) ) ;
    buf_clk new_AGEMA_reg_buffer_6417 ( .C (clk), .D (new_AGEMA_signal_2544), .Q (new_AGEMA_signal_9882) ) ;
    buf_clk new_AGEMA_reg_buffer_6421 ( .C (clk), .D (new_AGEMA_signal_2545), .Q (new_AGEMA_signal_9886) ) ;
    buf_clk new_AGEMA_reg_buffer_6431 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_14_n13), .Q (new_AGEMA_signal_9896) ) ;
    buf_clk new_AGEMA_reg_buffer_6435 ( .C (clk), .D (new_AGEMA_signal_2556), .Q (new_AGEMA_signal_9900) ) ;
    buf_clk new_AGEMA_reg_buffer_6439 ( .C (clk), .D (new_AGEMA_signal_2557), .Q (new_AGEMA_signal_9904) ) ;
    buf_clk new_AGEMA_reg_buffer_6449 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_15_n13), .Q (new_AGEMA_signal_9914) ) ;
    buf_clk new_AGEMA_reg_buffer_6453 ( .C (clk), .D (new_AGEMA_signal_2568), .Q (new_AGEMA_signal_9918) ) ;
    buf_clk new_AGEMA_reg_buffer_6457 ( .C (clk), .D (new_AGEMA_signal_2569), .Q (new_AGEMA_signal_9922) ) ;
    buf_clk new_AGEMA_reg_buffer_6465 ( .C (clk), .D (new_AGEMA_signal_9929), .Q (new_AGEMA_signal_9930) ) ;
    buf_clk new_AGEMA_reg_buffer_6473 ( .C (clk), .D (new_AGEMA_signal_9937), .Q (new_AGEMA_signal_9938) ) ;
    buf_clk new_AGEMA_reg_buffer_6481 ( .C (clk), .D (new_AGEMA_signal_9945), .Q (new_AGEMA_signal_9946) ) ;
    buf_clk new_AGEMA_reg_buffer_6489 ( .C (clk), .D (new_AGEMA_signal_9953), .Q (new_AGEMA_signal_9954) ) ;

    /* cells in depth 4 */
    or_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U18 ( .a ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, Midori_rounds_sub_sBox_PRINCE_0_n13}), .b ({new_AGEMA_signal_4925, new_AGEMA_signal_4923, new_AGEMA_signal_4921}), .clk (clk), .r ({Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, Midori_rounds_sub_sBox_PRINCE_0_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U15 ( .a ({new_AGEMA_signal_1871, new_AGEMA_signal_1870, Midori_rounds_sub_sBox_PRINCE_0_n10}), .b ({new_AGEMA_signal_4931, new_AGEMA_signal_4929, new_AGEMA_signal_4927}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291]}), .c ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, Midori_rounds_sub_sBox_PRINCE_0_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U11 ( .a ({new_AGEMA_signal_4937, new_AGEMA_signal_4935, new_AGEMA_signal_4933}), .b ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, Midori_rounds_sub_sBox_PRINCE_0_n4}), .clk (clk), .r ({Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, Midori_rounds_sub_sBox_PRINCE_0_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U6 ( .a ({new_AGEMA_signal_4943, new_AGEMA_signal_4941, new_AGEMA_signal_4939}), .b ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, Midori_rounds_sub_sBox_PRINCE_0_n1}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297]}), .c ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, Midori_rounds_sub_sBox_PRINCE_0_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U18 ( .a ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, Midori_rounds_sub_sBox_PRINCE_1_n13}), .b ({new_AGEMA_signal_4949, new_AGEMA_signal_4947, new_AGEMA_signal_4945}), .clk (clk), .r ({Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, Midori_rounds_sub_sBox_PRINCE_1_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U15 ( .a ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, Midori_rounds_sub_sBox_PRINCE_1_n10}), .b ({new_AGEMA_signal_4955, new_AGEMA_signal_4953, new_AGEMA_signal_4951}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303]}), .c ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, Midori_rounds_sub_sBox_PRINCE_1_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U11 ( .a ({new_AGEMA_signal_4961, new_AGEMA_signal_4959, new_AGEMA_signal_4957}), .b ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, Midori_rounds_sub_sBox_PRINCE_1_n4}), .clk (clk), .r ({Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, Midori_rounds_sub_sBox_PRINCE_1_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U6 ( .a ({new_AGEMA_signal_4967, new_AGEMA_signal_4965, new_AGEMA_signal_4963}), .b ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, Midori_rounds_sub_sBox_PRINCE_1_n1}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309]}), .c ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, Midori_rounds_sub_sBox_PRINCE_1_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U18 ( .a ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, Midori_rounds_sub_sBox_PRINCE_2_n13}), .b ({new_AGEMA_signal_4973, new_AGEMA_signal_4971, new_AGEMA_signal_4969}), .clk (clk), .r ({Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, Midori_rounds_sub_sBox_PRINCE_2_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U15 ( .a ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, Midori_rounds_sub_sBox_PRINCE_2_n10}), .b ({new_AGEMA_signal_4979, new_AGEMA_signal_4977, new_AGEMA_signal_4975}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315]}), .c ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, Midori_rounds_sub_sBox_PRINCE_2_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U11 ( .a ({new_AGEMA_signal_4985, new_AGEMA_signal_4983, new_AGEMA_signal_4981}), .b ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, Midori_rounds_sub_sBox_PRINCE_2_n4}), .clk (clk), .r ({Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, Midori_rounds_sub_sBox_PRINCE_2_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U6 ( .a ({new_AGEMA_signal_4991, new_AGEMA_signal_4989, new_AGEMA_signal_4987}), .b ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, Midori_rounds_sub_sBox_PRINCE_2_n1}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321]}), .c ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, Midori_rounds_sub_sBox_PRINCE_2_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U18 ( .a ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, Midori_rounds_sub_sBox_PRINCE_3_n13}), .b ({new_AGEMA_signal_4997, new_AGEMA_signal_4995, new_AGEMA_signal_4993}), .clk (clk), .r ({Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, Midori_rounds_sub_sBox_PRINCE_3_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U15 ( .a ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, Midori_rounds_sub_sBox_PRINCE_3_n10}), .b ({new_AGEMA_signal_5003, new_AGEMA_signal_5001, new_AGEMA_signal_4999}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327]}), .c ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, Midori_rounds_sub_sBox_PRINCE_3_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U11 ( .a ({new_AGEMA_signal_5009, new_AGEMA_signal_5007, new_AGEMA_signal_5005}), .b ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, Midori_rounds_sub_sBox_PRINCE_3_n4}), .clk (clk), .r ({Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, Midori_rounds_sub_sBox_PRINCE_3_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U6 ( .a ({new_AGEMA_signal_5015, new_AGEMA_signal_5013, new_AGEMA_signal_5011}), .b ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, Midori_rounds_sub_sBox_PRINCE_3_n1}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333]}), .c ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, Midori_rounds_sub_sBox_PRINCE_3_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U18 ( .a ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, Midori_rounds_sub_sBox_PRINCE_4_n13}), .b ({new_AGEMA_signal_5021, new_AGEMA_signal_5019, new_AGEMA_signal_5017}), .clk (clk), .r ({Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, Midori_rounds_sub_sBox_PRINCE_4_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U15 ( .a ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, Midori_rounds_sub_sBox_PRINCE_4_n10}), .b ({new_AGEMA_signal_5027, new_AGEMA_signal_5025, new_AGEMA_signal_5023}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339]}), .c ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, Midori_rounds_sub_sBox_PRINCE_4_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U11 ( .a ({new_AGEMA_signal_5033, new_AGEMA_signal_5031, new_AGEMA_signal_5029}), .b ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, Midori_rounds_sub_sBox_PRINCE_4_n4}), .clk (clk), .r ({Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, Midori_rounds_sub_sBox_PRINCE_4_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U6 ( .a ({new_AGEMA_signal_5039, new_AGEMA_signal_5037, new_AGEMA_signal_5035}), .b ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, Midori_rounds_sub_sBox_PRINCE_4_n1}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345]}), .c ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, Midori_rounds_sub_sBox_PRINCE_4_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U18 ( .a ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, Midori_rounds_sub_sBox_PRINCE_5_n13}), .b ({new_AGEMA_signal_5045, new_AGEMA_signal_5043, new_AGEMA_signal_5041}), .clk (clk), .r ({Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, Midori_rounds_sub_sBox_PRINCE_5_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U15 ( .a ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, Midori_rounds_sub_sBox_PRINCE_5_n10}), .b ({new_AGEMA_signal_5051, new_AGEMA_signal_5049, new_AGEMA_signal_5047}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351]}), .c ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, Midori_rounds_sub_sBox_PRINCE_5_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U11 ( .a ({new_AGEMA_signal_5057, new_AGEMA_signal_5055, new_AGEMA_signal_5053}), .b ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, Midori_rounds_sub_sBox_PRINCE_5_n4}), .clk (clk), .r ({Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, Midori_rounds_sub_sBox_PRINCE_5_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U6 ( .a ({new_AGEMA_signal_5063, new_AGEMA_signal_5061, new_AGEMA_signal_5059}), .b ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, Midori_rounds_sub_sBox_PRINCE_5_n1}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357]}), .c ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, Midori_rounds_sub_sBox_PRINCE_5_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U18 ( .a ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, Midori_rounds_sub_sBox_PRINCE_6_n13}), .b ({new_AGEMA_signal_5069, new_AGEMA_signal_5067, new_AGEMA_signal_5065}), .clk (clk), .r ({Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, Midori_rounds_sub_sBox_PRINCE_6_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U15 ( .a ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, Midori_rounds_sub_sBox_PRINCE_6_n10}), .b ({new_AGEMA_signal_5075, new_AGEMA_signal_5073, new_AGEMA_signal_5071}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363]}), .c ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, Midori_rounds_sub_sBox_PRINCE_6_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U11 ( .a ({new_AGEMA_signal_5081, new_AGEMA_signal_5079, new_AGEMA_signal_5077}), .b ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, Midori_rounds_sub_sBox_PRINCE_6_n4}), .clk (clk), .r ({Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, Midori_rounds_sub_sBox_PRINCE_6_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U6 ( .a ({new_AGEMA_signal_5087, new_AGEMA_signal_5085, new_AGEMA_signal_5083}), .b ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, Midori_rounds_sub_sBox_PRINCE_6_n1}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369]}), .c ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, Midori_rounds_sub_sBox_PRINCE_6_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U18 ( .a ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, Midori_rounds_sub_sBox_PRINCE_7_n13}), .b ({new_AGEMA_signal_5093, new_AGEMA_signal_5091, new_AGEMA_signal_5089}), .clk (clk), .r ({Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, Midori_rounds_sub_sBox_PRINCE_7_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U15 ( .a ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, Midori_rounds_sub_sBox_PRINCE_7_n10}), .b ({new_AGEMA_signal_5099, new_AGEMA_signal_5097, new_AGEMA_signal_5095}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375]}), .c ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, Midori_rounds_sub_sBox_PRINCE_7_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U11 ( .a ({new_AGEMA_signal_5105, new_AGEMA_signal_5103, new_AGEMA_signal_5101}), .b ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, Midori_rounds_sub_sBox_PRINCE_7_n4}), .clk (clk), .r ({Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, Midori_rounds_sub_sBox_PRINCE_7_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U6 ( .a ({new_AGEMA_signal_5111, new_AGEMA_signal_5109, new_AGEMA_signal_5107}), .b ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, Midori_rounds_sub_sBox_PRINCE_7_n1}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381]}), .c ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, Midori_rounds_sub_sBox_PRINCE_7_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U18 ( .a ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, Midori_rounds_sub_sBox_PRINCE_8_n13}), .b ({new_AGEMA_signal_5117, new_AGEMA_signal_5115, new_AGEMA_signal_5113}), .clk (clk), .r ({Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, Midori_rounds_sub_sBox_PRINCE_8_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U15 ( .a ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, Midori_rounds_sub_sBox_PRINCE_8_n10}), .b ({new_AGEMA_signal_5123, new_AGEMA_signal_5121, new_AGEMA_signal_5119}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387]}), .c ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, Midori_rounds_sub_sBox_PRINCE_8_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U11 ( .a ({new_AGEMA_signal_5129, new_AGEMA_signal_5127, new_AGEMA_signal_5125}), .b ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, Midori_rounds_sub_sBox_PRINCE_8_n4}), .clk (clk), .r ({Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, Midori_rounds_sub_sBox_PRINCE_8_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U6 ( .a ({new_AGEMA_signal_5135, new_AGEMA_signal_5133, new_AGEMA_signal_5131}), .b ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, Midori_rounds_sub_sBox_PRINCE_8_n1}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393]}), .c ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, Midori_rounds_sub_sBox_PRINCE_8_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U18 ( .a ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, Midori_rounds_sub_sBox_PRINCE_9_n13}), .b ({new_AGEMA_signal_5141, new_AGEMA_signal_5139, new_AGEMA_signal_5137}), .clk (clk), .r ({Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, Midori_rounds_sub_sBox_PRINCE_9_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U15 ( .a ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, Midori_rounds_sub_sBox_PRINCE_9_n10}), .b ({new_AGEMA_signal_5147, new_AGEMA_signal_5145, new_AGEMA_signal_5143}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399]}), .c ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, Midori_rounds_sub_sBox_PRINCE_9_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U11 ( .a ({new_AGEMA_signal_5153, new_AGEMA_signal_5151, new_AGEMA_signal_5149}), .b ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, Midori_rounds_sub_sBox_PRINCE_9_n4}), .clk (clk), .r ({Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, Midori_rounds_sub_sBox_PRINCE_9_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U6 ( .a ({new_AGEMA_signal_5159, new_AGEMA_signal_5157, new_AGEMA_signal_5155}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, Midori_rounds_sub_sBox_PRINCE_9_n1}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405]}), .c ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, Midori_rounds_sub_sBox_PRINCE_9_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U18 ( .a ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, Midori_rounds_sub_sBox_PRINCE_10_n13}), .b ({new_AGEMA_signal_5165, new_AGEMA_signal_5163, new_AGEMA_signal_5161}), .clk (clk), .r ({Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, Midori_rounds_sub_sBox_PRINCE_10_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U15 ( .a ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, Midori_rounds_sub_sBox_PRINCE_10_n10}), .b ({new_AGEMA_signal_5171, new_AGEMA_signal_5169, new_AGEMA_signal_5167}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411]}), .c ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, Midori_rounds_sub_sBox_PRINCE_10_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U11 ( .a ({new_AGEMA_signal_5177, new_AGEMA_signal_5175, new_AGEMA_signal_5173}), .b ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, Midori_rounds_sub_sBox_PRINCE_10_n4}), .clk (clk), .r ({Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, Midori_rounds_sub_sBox_PRINCE_10_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U6 ( .a ({new_AGEMA_signal_5183, new_AGEMA_signal_5181, new_AGEMA_signal_5179}), .b ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, Midori_rounds_sub_sBox_PRINCE_10_n1}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417]}), .c ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, Midori_rounds_sub_sBox_PRINCE_10_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U18 ( .a ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, Midori_rounds_sub_sBox_PRINCE_11_n13}), .b ({new_AGEMA_signal_5189, new_AGEMA_signal_5187, new_AGEMA_signal_5185}), .clk (clk), .r ({Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, Midori_rounds_sub_sBox_PRINCE_11_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U15 ( .a ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, Midori_rounds_sub_sBox_PRINCE_11_n10}), .b ({new_AGEMA_signal_5195, new_AGEMA_signal_5193, new_AGEMA_signal_5191}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423]}), .c ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, Midori_rounds_sub_sBox_PRINCE_11_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U11 ( .a ({new_AGEMA_signal_5201, new_AGEMA_signal_5199, new_AGEMA_signal_5197}), .b ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, Midori_rounds_sub_sBox_PRINCE_11_n4}), .clk (clk), .r ({Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, Midori_rounds_sub_sBox_PRINCE_11_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U6 ( .a ({new_AGEMA_signal_5207, new_AGEMA_signal_5205, new_AGEMA_signal_5203}), .b ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, Midori_rounds_sub_sBox_PRINCE_11_n1}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429]}), .c ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, Midori_rounds_sub_sBox_PRINCE_11_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U18 ( .a ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, Midori_rounds_sub_sBox_PRINCE_12_n13}), .b ({new_AGEMA_signal_5213, new_AGEMA_signal_5211, new_AGEMA_signal_5209}), .clk (clk), .r ({Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, Midori_rounds_sub_sBox_PRINCE_12_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U15 ( .a ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, Midori_rounds_sub_sBox_PRINCE_12_n10}), .b ({new_AGEMA_signal_5219, new_AGEMA_signal_5217, new_AGEMA_signal_5215}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435]}), .c ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, Midori_rounds_sub_sBox_PRINCE_12_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U11 ( .a ({new_AGEMA_signal_5225, new_AGEMA_signal_5223, new_AGEMA_signal_5221}), .b ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, Midori_rounds_sub_sBox_PRINCE_12_n4}), .clk (clk), .r ({Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, Midori_rounds_sub_sBox_PRINCE_12_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U6 ( .a ({new_AGEMA_signal_5231, new_AGEMA_signal_5229, new_AGEMA_signal_5227}), .b ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, Midori_rounds_sub_sBox_PRINCE_12_n1}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441]}), .c ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, Midori_rounds_sub_sBox_PRINCE_12_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U18 ( .a ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, Midori_rounds_sub_sBox_PRINCE_13_n13}), .b ({new_AGEMA_signal_5237, new_AGEMA_signal_5235, new_AGEMA_signal_5233}), .clk (clk), .r ({Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, Midori_rounds_sub_sBox_PRINCE_13_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U15 ( .a ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, Midori_rounds_sub_sBox_PRINCE_13_n10}), .b ({new_AGEMA_signal_5243, new_AGEMA_signal_5241, new_AGEMA_signal_5239}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447]}), .c ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, Midori_rounds_sub_sBox_PRINCE_13_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U11 ( .a ({new_AGEMA_signal_5249, new_AGEMA_signal_5247, new_AGEMA_signal_5245}), .b ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, Midori_rounds_sub_sBox_PRINCE_13_n4}), .clk (clk), .r ({Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, Midori_rounds_sub_sBox_PRINCE_13_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U6 ( .a ({new_AGEMA_signal_5255, new_AGEMA_signal_5253, new_AGEMA_signal_5251}), .b ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, Midori_rounds_sub_sBox_PRINCE_13_n1}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453]}), .c ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, Midori_rounds_sub_sBox_PRINCE_13_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U18 ( .a ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, Midori_rounds_sub_sBox_PRINCE_14_n13}), .b ({new_AGEMA_signal_5261, new_AGEMA_signal_5259, new_AGEMA_signal_5257}), .clk (clk), .r ({Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_2815, new_AGEMA_signal_2814, Midori_rounds_sub_sBox_PRINCE_14_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U15 ( .a ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, Midori_rounds_sub_sBox_PRINCE_14_n10}), .b ({new_AGEMA_signal_5267, new_AGEMA_signal_5265, new_AGEMA_signal_5263}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459]}), .c ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, Midori_rounds_sub_sBox_PRINCE_14_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U11 ( .a ({new_AGEMA_signal_5273, new_AGEMA_signal_5271, new_AGEMA_signal_5269}), .b ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, Midori_rounds_sub_sBox_PRINCE_14_n4}), .clk (clk), .r ({Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, Midori_rounds_sub_sBox_PRINCE_14_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U6 ( .a ({new_AGEMA_signal_5279, new_AGEMA_signal_5277, new_AGEMA_signal_5275}), .b ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, Midori_rounds_sub_sBox_PRINCE_14_n1}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465]}), .c ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, Midori_rounds_sub_sBox_PRINCE_14_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U18 ( .a ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, Midori_rounds_sub_sBox_PRINCE_15_n13}), .b ({new_AGEMA_signal_5285, new_AGEMA_signal_5283, new_AGEMA_signal_5281}), .clk (clk), .r ({Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, Midori_rounds_sub_sBox_PRINCE_15_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U15 ( .a ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, Midori_rounds_sub_sBox_PRINCE_15_n10}), .b ({new_AGEMA_signal_5291, new_AGEMA_signal_5289, new_AGEMA_signal_5287}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471]}), .c ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, Midori_rounds_sub_sBox_PRINCE_15_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U11 ( .a ({new_AGEMA_signal_5297, new_AGEMA_signal_5295, new_AGEMA_signal_5293}), .b ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, Midori_rounds_sub_sBox_PRINCE_15_n4}), .clk (clk), .r ({Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, Midori_rounds_sub_sBox_PRINCE_15_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U6 ( .a ({new_AGEMA_signal_5303, new_AGEMA_signal_5301, new_AGEMA_signal_5299}), .b ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, Midori_rounds_sub_sBox_PRINCE_15_n1}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477]}), .c ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, Midori_rounds_sub_sBox_PRINCE_15_n2}) ) ;
    buf_clk new_AGEMA_reg_buffer_1322 ( .C (clk), .D (new_AGEMA_signal_4787), .Q (new_AGEMA_signal_4788) ) ;
    buf_clk new_AGEMA_reg_buffer_1842 ( .C (clk), .D (new_AGEMA_signal_5306), .Q (new_AGEMA_signal_5307) ) ;
    buf_clk new_AGEMA_reg_buffer_1848 ( .C (clk), .D (new_AGEMA_signal_5312), .Q (new_AGEMA_signal_5313) ) ;
    buf_clk new_AGEMA_reg_buffer_1854 ( .C (clk), .D (new_AGEMA_signal_5318), .Q (new_AGEMA_signal_5319) ) ;
    buf_clk new_AGEMA_reg_buffer_1860 ( .C (clk), .D (new_AGEMA_signal_5324), .Q (new_AGEMA_signal_5325) ) ;
    buf_clk new_AGEMA_reg_buffer_1866 ( .C (clk), .D (new_AGEMA_signal_5330), .Q (new_AGEMA_signal_5331) ) ;
    buf_clk new_AGEMA_reg_buffer_1872 ( .C (clk), .D (new_AGEMA_signal_5336), .Q (new_AGEMA_signal_5337) ) ;
    buf_clk new_AGEMA_reg_buffer_1878 ( .C (clk), .D (new_AGEMA_signal_5342), .Q (new_AGEMA_signal_5343) ) ;
    buf_clk new_AGEMA_reg_buffer_1884 ( .C (clk), .D (new_AGEMA_signal_5348), .Q (new_AGEMA_signal_5349) ) ;
    buf_clk new_AGEMA_reg_buffer_1890 ( .C (clk), .D (new_AGEMA_signal_5354), .Q (new_AGEMA_signal_5355) ) ;
    buf_clk new_AGEMA_reg_buffer_1896 ( .C (clk), .D (new_AGEMA_signal_5360), .Q (new_AGEMA_signal_5361) ) ;
    buf_clk new_AGEMA_reg_buffer_1902 ( .C (clk), .D (new_AGEMA_signal_5366), .Q (new_AGEMA_signal_5367) ) ;
    buf_clk new_AGEMA_reg_buffer_1908 ( .C (clk), .D (new_AGEMA_signal_5372), .Q (new_AGEMA_signal_5373) ) ;
    buf_clk new_AGEMA_reg_buffer_1914 ( .C (clk), .D (new_AGEMA_signal_5378), .Q (new_AGEMA_signal_5379) ) ;
    buf_clk new_AGEMA_reg_buffer_1920 ( .C (clk), .D (new_AGEMA_signal_5384), .Q (new_AGEMA_signal_5385) ) ;
    buf_clk new_AGEMA_reg_buffer_1926 ( .C (clk), .D (new_AGEMA_signal_5390), .Q (new_AGEMA_signal_5391) ) ;
    buf_clk new_AGEMA_reg_buffer_1932 ( .C (clk), .D (new_AGEMA_signal_5396), .Q (new_AGEMA_signal_5397) ) ;
    buf_clk new_AGEMA_reg_buffer_1938 ( .C (clk), .D (new_AGEMA_signal_5402), .Q (new_AGEMA_signal_5403) ) ;
    buf_clk new_AGEMA_reg_buffer_1944 ( .C (clk), .D (new_AGEMA_signal_5408), .Q (new_AGEMA_signal_5409) ) ;
    buf_clk new_AGEMA_reg_buffer_1950 ( .C (clk), .D (new_AGEMA_signal_5414), .Q (new_AGEMA_signal_5415) ) ;
    buf_clk new_AGEMA_reg_buffer_1956 ( .C (clk), .D (new_AGEMA_signal_5420), .Q (new_AGEMA_signal_5421) ) ;
    buf_clk new_AGEMA_reg_buffer_1962 ( .C (clk), .D (new_AGEMA_signal_5426), .Q (new_AGEMA_signal_5427) ) ;
    buf_clk new_AGEMA_reg_buffer_1968 ( .C (clk), .D (new_AGEMA_signal_5432), .Q (new_AGEMA_signal_5433) ) ;
    buf_clk new_AGEMA_reg_buffer_1974 ( .C (clk), .D (new_AGEMA_signal_5438), .Q (new_AGEMA_signal_5439) ) ;
    buf_clk new_AGEMA_reg_buffer_1980 ( .C (clk), .D (new_AGEMA_signal_5444), .Q (new_AGEMA_signal_5445) ) ;
    buf_clk new_AGEMA_reg_buffer_1986 ( .C (clk), .D (new_AGEMA_signal_5450), .Q (new_AGEMA_signal_5451) ) ;
    buf_clk new_AGEMA_reg_buffer_1992 ( .C (clk), .D (new_AGEMA_signal_5456), .Q (new_AGEMA_signal_5457) ) ;
    buf_clk new_AGEMA_reg_buffer_1998 ( .C (clk), .D (new_AGEMA_signal_5462), .Q (new_AGEMA_signal_5463) ) ;
    buf_clk new_AGEMA_reg_buffer_2004 ( .C (clk), .D (new_AGEMA_signal_5468), .Q (new_AGEMA_signal_5469) ) ;
    buf_clk new_AGEMA_reg_buffer_2010 ( .C (clk), .D (new_AGEMA_signal_5474), .Q (new_AGEMA_signal_5475) ) ;
    buf_clk new_AGEMA_reg_buffer_2016 ( .C (clk), .D (new_AGEMA_signal_5480), .Q (new_AGEMA_signal_5481) ) ;
    buf_clk new_AGEMA_reg_buffer_2022 ( .C (clk), .D (new_AGEMA_signal_5486), .Q (new_AGEMA_signal_5487) ) ;
    buf_clk new_AGEMA_reg_buffer_2028 ( .C (clk), .D (new_AGEMA_signal_5492), .Q (new_AGEMA_signal_5493) ) ;
    buf_clk new_AGEMA_reg_buffer_2034 ( .C (clk), .D (new_AGEMA_signal_5498), .Q (new_AGEMA_signal_5499) ) ;
    buf_clk new_AGEMA_reg_buffer_2040 ( .C (clk), .D (new_AGEMA_signal_5504), .Q (new_AGEMA_signal_5505) ) ;
    buf_clk new_AGEMA_reg_buffer_2046 ( .C (clk), .D (new_AGEMA_signal_5510), .Q (new_AGEMA_signal_5511) ) ;
    buf_clk new_AGEMA_reg_buffer_2052 ( .C (clk), .D (new_AGEMA_signal_5516), .Q (new_AGEMA_signal_5517) ) ;
    buf_clk new_AGEMA_reg_buffer_2058 ( .C (clk), .D (new_AGEMA_signal_5522), .Q (new_AGEMA_signal_5523) ) ;
    buf_clk new_AGEMA_reg_buffer_2064 ( .C (clk), .D (new_AGEMA_signal_5528), .Q (new_AGEMA_signal_5529) ) ;
    buf_clk new_AGEMA_reg_buffer_2070 ( .C (clk), .D (new_AGEMA_signal_5534), .Q (new_AGEMA_signal_5535) ) ;
    buf_clk new_AGEMA_reg_buffer_2076 ( .C (clk), .D (new_AGEMA_signal_5540), .Q (new_AGEMA_signal_5541) ) ;
    buf_clk new_AGEMA_reg_buffer_2082 ( .C (clk), .D (new_AGEMA_signal_5546), .Q (new_AGEMA_signal_5547) ) ;
    buf_clk new_AGEMA_reg_buffer_2088 ( .C (clk), .D (new_AGEMA_signal_5552), .Q (new_AGEMA_signal_5553) ) ;
    buf_clk new_AGEMA_reg_buffer_2094 ( .C (clk), .D (new_AGEMA_signal_5558), .Q (new_AGEMA_signal_5559) ) ;
    buf_clk new_AGEMA_reg_buffer_2100 ( .C (clk), .D (new_AGEMA_signal_5564), .Q (new_AGEMA_signal_5565) ) ;
    buf_clk new_AGEMA_reg_buffer_2106 ( .C (clk), .D (new_AGEMA_signal_5570), .Q (new_AGEMA_signal_5571) ) ;
    buf_clk new_AGEMA_reg_buffer_2112 ( .C (clk), .D (new_AGEMA_signal_5576), .Q (new_AGEMA_signal_5577) ) ;
    buf_clk new_AGEMA_reg_buffer_2118 ( .C (clk), .D (new_AGEMA_signal_5582), .Q (new_AGEMA_signal_5583) ) ;
    buf_clk new_AGEMA_reg_buffer_2124 ( .C (clk), .D (new_AGEMA_signal_5588), .Q (new_AGEMA_signal_5589) ) ;
    buf_clk new_AGEMA_reg_buffer_2130 ( .C (clk), .D (new_AGEMA_signal_5594), .Q (new_AGEMA_signal_5595) ) ;
    buf_clk new_AGEMA_reg_buffer_2136 ( .C (clk), .D (new_AGEMA_signal_5600), .Q (new_AGEMA_signal_5601) ) ;
    buf_clk new_AGEMA_reg_buffer_2142 ( .C (clk), .D (new_AGEMA_signal_5606), .Q (new_AGEMA_signal_5607) ) ;
    buf_clk new_AGEMA_reg_buffer_2148 ( .C (clk), .D (new_AGEMA_signal_5612), .Q (new_AGEMA_signal_5613) ) ;
    buf_clk new_AGEMA_reg_buffer_2154 ( .C (clk), .D (new_AGEMA_signal_5618), .Q (new_AGEMA_signal_5619) ) ;
    buf_clk new_AGEMA_reg_buffer_2160 ( .C (clk), .D (new_AGEMA_signal_5624), .Q (new_AGEMA_signal_5625) ) ;
    buf_clk new_AGEMA_reg_buffer_2166 ( .C (clk), .D (new_AGEMA_signal_5630), .Q (new_AGEMA_signal_5631) ) ;
    buf_clk new_AGEMA_reg_buffer_2172 ( .C (clk), .D (new_AGEMA_signal_5636), .Q (new_AGEMA_signal_5637) ) ;
    buf_clk new_AGEMA_reg_buffer_2178 ( .C (clk), .D (new_AGEMA_signal_5642), .Q (new_AGEMA_signal_5643) ) ;
    buf_clk new_AGEMA_reg_buffer_2184 ( .C (clk), .D (new_AGEMA_signal_5648), .Q (new_AGEMA_signal_5649) ) ;
    buf_clk new_AGEMA_reg_buffer_2190 ( .C (clk), .D (new_AGEMA_signal_5654), .Q (new_AGEMA_signal_5655) ) ;
    buf_clk new_AGEMA_reg_buffer_2196 ( .C (clk), .D (new_AGEMA_signal_5660), .Q (new_AGEMA_signal_5661) ) ;
    buf_clk new_AGEMA_reg_buffer_2202 ( .C (clk), .D (new_AGEMA_signal_5666), .Q (new_AGEMA_signal_5667) ) ;
    buf_clk new_AGEMA_reg_buffer_2208 ( .C (clk), .D (new_AGEMA_signal_5672), .Q (new_AGEMA_signal_5673) ) ;
    buf_clk new_AGEMA_reg_buffer_2214 ( .C (clk), .D (new_AGEMA_signal_5678), .Q (new_AGEMA_signal_5679) ) ;
    buf_clk new_AGEMA_reg_buffer_2220 ( .C (clk), .D (new_AGEMA_signal_5684), .Q (new_AGEMA_signal_5685) ) ;
    buf_clk new_AGEMA_reg_buffer_2226 ( .C (clk), .D (new_AGEMA_signal_5690), .Q (new_AGEMA_signal_5691) ) ;
    buf_clk new_AGEMA_reg_buffer_2232 ( .C (clk), .D (new_AGEMA_signal_5696), .Q (new_AGEMA_signal_5697) ) ;
    buf_clk new_AGEMA_reg_buffer_2238 ( .C (clk), .D (new_AGEMA_signal_5702), .Q (new_AGEMA_signal_5703) ) ;
    buf_clk new_AGEMA_reg_buffer_2244 ( .C (clk), .D (new_AGEMA_signal_5708), .Q (new_AGEMA_signal_5709) ) ;
    buf_clk new_AGEMA_reg_buffer_2250 ( .C (clk), .D (new_AGEMA_signal_5714), .Q (new_AGEMA_signal_5715) ) ;
    buf_clk new_AGEMA_reg_buffer_2256 ( .C (clk), .D (new_AGEMA_signal_5720), .Q (new_AGEMA_signal_5721) ) ;
    buf_clk new_AGEMA_reg_buffer_2262 ( .C (clk), .D (new_AGEMA_signal_5726), .Q (new_AGEMA_signal_5727) ) ;
    buf_clk new_AGEMA_reg_buffer_2268 ( .C (clk), .D (new_AGEMA_signal_5732), .Q (new_AGEMA_signal_5733) ) ;
    buf_clk new_AGEMA_reg_buffer_2274 ( .C (clk), .D (new_AGEMA_signal_5738), .Q (new_AGEMA_signal_5739) ) ;
    buf_clk new_AGEMA_reg_buffer_2280 ( .C (clk), .D (new_AGEMA_signal_5744), .Q (new_AGEMA_signal_5745) ) ;
    buf_clk new_AGEMA_reg_buffer_2286 ( .C (clk), .D (new_AGEMA_signal_5750), .Q (new_AGEMA_signal_5751) ) ;
    buf_clk new_AGEMA_reg_buffer_2292 ( .C (clk), .D (new_AGEMA_signal_5756), .Q (new_AGEMA_signal_5757) ) ;
    buf_clk new_AGEMA_reg_buffer_2298 ( .C (clk), .D (new_AGEMA_signal_5762), .Q (new_AGEMA_signal_5763) ) ;
    buf_clk new_AGEMA_reg_buffer_2304 ( .C (clk), .D (new_AGEMA_signal_5768), .Q (new_AGEMA_signal_5769) ) ;
    buf_clk new_AGEMA_reg_buffer_2310 ( .C (clk), .D (new_AGEMA_signal_5774), .Q (new_AGEMA_signal_5775) ) ;
    buf_clk new_AGEMA_reg_buffer_2316 ( .C (clk), .D (new_AGEMA_signal_5780), .Q (new_AGEMA_signal_5781) ) ;
    buf_clk new_AGEMA_reg_buffer_2322 ( .C (clk), .D (new_AGEMA_signal_5786), .Q (new_AGEMA_signal_5787) ) ;
    buf_clk new_AGEMA_reg_buffer_2328 ( .C (clk), .D (new_AGEMA_signal_5792), .Q (new_AGEMA_signal_5793) ) ;
    buf_clk new_AGEMA_reg_buffer_2334 ( .C (clk), .D (new_AGEMA_signal_5798), .Q (new_AGEMA_signal_5799) ) ;
    buf_clk new_AGEMA_reg_buffer_2340 ( .C (clk), .D (new_AGEMA_signal_5804), .Q (new_AGEMA_signal_5805) ) ;
    buf_clk new_AGEMA_reg_buffer_2346 ( .C (clk), .D (new_AGEMA_signal_5810), .Q (new_AGEMA_signal_5811) ) ;
    buf_clk new_AGEMA_reg_buffer_2352 ( .C (clk), .D (new_AGEMA_signal_5816), .Q (new_AGEMA_signal_5817) ) ;
    buf_clk new_AGEMA_reg_buffer_2358 ( .C (clk), .D (new_AGEMA_signal_5822), .Q (new_AGEMA_signal_5823) ) ;
    buf_clk new_AGEMA_reg_buffer_2364 ( .C (clk), .D (new_AGEMA_signal_5828), .Q (new_AGEMA_signal_5829) ) ;
    buf_clk new_AGEMA_reg_buffer_2370 ( .C (clk), .D (new_AGEMA_signal_5834), .Q (new_AGEMA_signal_5835) ) ;
    buf_clk new_AGEMA_reg_buffer_2376 ( .C (clk), .D (new_AGEMA_signal_5840), .Q (new_AGEMA_signal_5841) ) ;
    buf_clk new_AGEMA_reg_buffer_2382 ( .C (clk), .D (new_AGEMA_signal_5846), .Q (new_AGEMA_signal_5847) ) ;
    buf_clk new_AGEMA_reg_buffer_2388 ( .C (clk), .D (new_AGEMA_signal_5852), .Q (new_AGEMA_signal_5853) ) ;
    buf_clk new_AGEMA_reg_buffer_2394 ( .C (clk), .D (new_AGEMA_signal_5858), .Q (new_AGEMA_signal_5859) ) ;
    buf_clk new_AGEMA_reg_buffer_2400 ( .C (clk), .D (new_AGEMA_signal_5864), .Q (new_AGEMA_signal_5865) ) ;
    buf_clk new_AGEMA_reg_buffer_2406 ( .C (clk), .D (new_AGEMA_signal_5870), .Q (new_AGEMA_signal_5871) ) ;
    buf_clk new_AGEMA_reg_buffer_2412 ( .C (clk), .D (new_AGEMA_signal_5876), .Q (new_AGEMA_signal_5877) ) ;
    buf_clk new_AGEMA_reg_buffer_2418 ( .C (clk), .D (new_AGEMA_signal_5882), .Q (new_AGEMA_signal_5883) ) ;
    buf_clk new_AGEMA_reg_buffer_2424 ( .C (clk), .D (new_AGEMA_signal_5888), .Q (new_AGEMA_signal_5889) ) ;
    buf_clk new_AGEMA_reg_buffer_2430 ( .C (clk), .D (new_AGEMA_signal_5894), .Q (new_AGEMA_signal_5895) ) ;
    buf_clk new_AGEMA_reg_buffer_2436 ( .C (clk), .D (new_AGEMA_signal_5900), .Q (new_AGEMA_signal_5901) ) ;
    buf_clk new_AGEMA_reg_buffer_2442 ( .C (clk), .D (new_AGEMA_signal_5906), .Q (new_AGEMA_signal_5907) ) ;
    buf_clk new_AGEMA_reg_buffer_2448 ( .C (clk), .D (new_AGEMA_signal_5912), .Q (new_AGEMA_signal_5913) ) ;
    buf_clk new_AGEMA_reg_buffer_2454 ( .C (clk), .D (new_AGEMA_signal_5918), .Q (new_AGEMA_signal_5919) ) ;
    buf_clk new_AGEMA_reg_buffer_2460 ( .C (clk), .D (new_AGEMA_signal_5924), .Q (new_AGEMA_signal_5925) ) ;
    buf_clk new_AGEMA_reg_buffer_2466 ( .C (clk), .D (new_AGEMA_signal_5930), .Q (new_AGEMA_signal_5931) ) ;
    buf_clk new_AGEMA_reg_buffer_2472 ( .C (clk), .D (new_AGEMA_signal_5936), .Q (new_AGEMA_signal_5937) ) ;
    buf_clk new_AGEMA_reg_buffer_2478 ( .C (clk), .D (new_AGEMA_signal_5942), .Q (new_AGEMA_signal_5943) ) ;
    buf_clk new_AGEMA_reg_buffer_2484 ( .C (clk), .D (new_AGEMA_signal_5948), .Q (new_AGEMA_signal_5949) ) ;
    buf_clk new_AGEMA_reg_buffer_2490 ( .C (clk), .D (new_AGEMA_signal_5954), .Q (new_AGEMA_signal_5955) ) ;
    buf_clk new_AGEMA_reg_buffer_2496 ( .C (clk), .D (new_AGEMA_signal_5960), .Q (new_AGEMA_signal_5961) ) ;
    buf_clk new_AGEMA_reg_buffer_2502 ( .C (clk), .D (new_AGEMA_signal_5966), .Q (new_AGEMA_signal_5967) ) ;
    buf_clk new_AGEMA_reg_buffer_2508 ( .C (clk), .D (new_AGEMA_signal_5972), .Q (new_AGEMA_signal_5973) ) ;
    buf_clk new_AGEMA_reg_buffer_2514 ( .C (clk), .D (new_AGEMA_signal_5978), .Q (new_AGEMA_signal_5979) ) ;
    buf_clk new_AGEMA_reg_buffer_2520 ( .C (clk), .D (new_AGEMA_signal_5984), .Q (new_AGEMA_signal_5985) ) ;
    buf_clk new_AGEMA_reg_buffer_2526 ( .C (clk), .D (new_AGEMA_signal_5990), .Q (new_AGEMA_signal_5991) ) ;
    buf_clk new_AGEMA_reg_buffer_2532 ( .C (clk), .D (new_AGEMA_signal_5996), .Q (new_AGEMA_signal_5997) ) ;
    buf_clk new_AGEMA_reg_buffer_2538 ( .C (clk), .D (new_AGEMA_signal_6002), .Q (new_AGEMA_signal_6003) ) ;
    buf_clk new_AGEMA_reg_buffer_2544 ( .C (clk), .D (new_AGEMA_signal_6008), .Q (new_AGEMA_signal_6009) ) ;
    buf_clk new_AGEMA_reg_buffer_2550 ( .C (clk), .D (new_AGEMA_signal_6014), .Q (new_AGEMA_signal_6015) ) ;
    buf_clk new_AGEMA_reg_buffer_2556 ( .C (clk), .D (new_AGEMA_signal_6020), .Q (new_AGEMA_signal_6021) ) ;
    buf_clk new_AGEMA_reg_buffer_2562 ( .C (clk), .D (new_AGEMA_signal_6026), .Q (new_AGEMA_signal_6027) ) ;
    buf_clk new_AGEMA_reg_buffer_2568 ( .C (clk), .D (new_AGEMA_signal_6032), .Q (new_AGEMA_signal_6033) ) ;
    buf_clk new_AGEMA_reg_buffer_2574 ( .C (clk), .D (new_AGEMA_signal_6038), .Q (new_AGEMA_signal_6039) ) ;
    buf_clk new_AGEMA_reg_buffer_2580 ( .C (clk), .D (new_AGEMA_signal_6044), .Q (new_AGEMA_signal_6045) ) ;
    buf_clk new_AGEMA_reg_buffer_2586 ( .C (clk), .D (new_AGEMA_signal_6050), .Q (new_AGEMA_signal_6051) ) ;
    buf_clk new_AGEMA_reg_buffer_2592 ( .C (clk), .D (new_AGEMA_signal_6056), .Q (new_AGEMA_signal_6057) ) ;
    buf_clk new_AGEMA_reg_buffer_2598 ( .C (clk), .D (new_AGEMA_signal_6062), .Q (new_AGEMA_signal_6063) ) ;
    buf_clk new_AGEMA_reg_buffer_2604 ( .C (clk), .D (new_AGEMA_signal_6068), .Q (new_AGEMA_signal_6069) ) ;
    buf_clk new_AGEMA_reg_buffer_2610 ( .C (clk), .D (new_AGEMA_signal_6074), .Q (new_AGEMA_signal_6075) ) ;
    buf_clk new_AGEMA_reg_buffer_2616 ( .C (clk), .D (new_AGEMA_signal_6080), .Q (new_AGEMA_signal_6081) ) ;
    buf_clk new_AGEMA_reg_buffer_2622 ( .C (clk), .D (new_AGEMA_signal_6086), .Q (new_AGEMA_signal_6087) ) ;
    buf_clk new_AGEMA_reg_buffer_2628 ( .C (clk), .D (new_AGEMA_signal_6092), .Q (new_AGEMA_signal_6093) ) ;
    buf_clk new_AGEMA_reg_buffer_2634 ( .C (clk), .D (new_AGEMA_signal_6098), .Q (new_AGEMA_signal_6099) ) ;
    buf_clk new_AGEMA_reg_buffer_2640 ( .C (clk), .D (new_AGEMA_signal_6104), .Q (new_AGEMA_signal_6105) ) ;
    buf_clk new_AGEMA_reg_buffer_2646 ( .C (clk), .D (new_AGEMA_signal_6110), .Q (new_AGEMA_signal_6111) ) ;
    buf_clk new_AGEMA_reg_buffer_2652 ( .C (clk), .D (new_AGEMA_signal_6116), .Q (new_AGEMA_signal_6117) ) ;
    buf_clk new_AGEMA_reg_buffer_2658 ( .C (clk), .D (new_AGEMA_signal_6122), .Q (new_AGEMA_signal_6123) ) ;
    buf_clk new_AGEMA_reg_buffer_2664 ( .C (clk), .D (new_AGEMA_signal_6128), .Q (new_AGEMA_signal_6129) ) ;
    buf_clk new_AGEMA_reg_buffer_2670 ( .C (clk), .D (new_AGEMA_signal_6134), .Q (new_AGEMA_signal_6135) ) ;
    buf_clk new_AGEMA_reg_buffer_2676 ( .C (clk), .D (new_AGEMA_signal_6140), .Q (new_AGEMA_signal_6141) ) ;
    buf_clk new_AGEMA_reg_buffer_2682 ( .C (clk), .D (new_AGEMA_signal_6146), .Q (new_AGEMA_signal_6147) ) ;
    buf_clk new_AGEMA_reg_buffer_2688 ( .C (clk), .D (new_AGEMA_signal_6152), .Q (new_AGEMA_signal_6153) ) ;
    buf_clk new_AGEMA_reg_buffer_2694 ( .C (clk), .D (new_AGEMA_signal_6158), .Q (new_AGEMA_signal_6159) ) ;
    buf_clk new_AGEMA_reg_buffer_2700 ( .C (clk), .D (new_AGEMA_signal_6164), .Q (new_AGEMA_signal_6165) ) ;
    buf_clk new_AGEMA_reg_buffer_2706 ( .C (clk), .D (new_AGEMA_signal_6170), .Q (new_AGEMA_signal_6171) ) ;
    buf_clk new_AGEMA_reg_buffer_2712 ( .C (clk), .D (new_AGEMA_signal_6176), .Q (new_AGEMA_signal_6177) ) ;
    buf_clk new_AGEMA_reg_buffer_2718 ( .C (clk), .D (new_AGEMA_signal_6182), .Q (new_AGEMA_signal_6183) ) ;
    buf_clk new_AGEMA_reg_buffer_2724 ( .C (clk), .D (new_AGEMA_signal_6188), .Q (new_AGEMA_signal_6189) ) ;
    buf_clk new_AGEMA_reg_buffer_2730 ( .C (clk), .D (new_AGEMA_signal_6194), .Q (new_AGEMA_signal_6195) ) ;
    buf_clk new_AGEMA_reg_buffer_2736 ( .C (clk), .D (new_AGEMA_signal_6200), .Q (new_AGEMA_signal_6201) ) ;
    buf_clk new_AGEMA_reg_buffer_2742 ( .C (clk), .D (new_AGEMA_signal_6206), .Q (new_AGEMA_signal_6207) ) ;
    buf_clk new_AGEMA_reg_buffer_2748 ( .C (clk), .D (new_AGEMA_signal_6212), .Q (new_AGEMA_signal_6213) ) ;
    buf_clk new_AGEMA_reg_buffer_2754 ( .C (clk), .D (new_AGEMA_signal_6218), .Q (new_AGEMA_signal_6219) ) ;
    buf_clk new_AGEMA_reg_buffer_2760 ( .C (clk), .D (new_AGEMA_signal_6224), .Q (new_AGEMA_signal_6225) ) ;
    buf_clk new_AGEMA_reg_buffer_2766 ( .C (clk), .D (new_AGEMA_signal_6230), .Q (new_AGEMA_signal_6231) ) ;
    buf_clk new_AGEMA_reg_buffer_2772 ( .C (clk), .D (new_AGEMA_signal_6236), .Q (new_AGEMA_signal_6237) ) ;
    buf_clk new_AGEMA_reg_buffer_2778 ( .C (clk), .D (new_AGEMA_signal_6242), .Q (new_AGEMA_signal_6243) ) ;
    buf_clk new_AGEMA_reg_buffer_2784 ( .C (clk), .D (new_AGEMA_signal_6248), .Q (new_AGEMA_signal_6249) ) ;
    buf_clk new_AGEMA_reg_buffer_2790 ( .C (clk), .D (new_AGEMA_signal_6254), .Q (new_AGEMA_signal_6255) ) ;
    buf_clk new_AGEMA_reg_buffer_2796 ( .C (clk), .D (new_AGEMA_signal_6260), .Q (new_AGEMA_signal_6261) ) ;
    buf_clk new_AGEMA_reg_buffer_2802 ( .C (clk), .D (new_AGEMA_signal_6266), .Q (new_AGEMA_signal_6267) ) ;
    buf_clk new_AGEMA_reg_buffer_2808 ( .C (clk), .D (new_AGEMA_signal_6272), .Q (new_AGEMA_signal_6273) ) ;
    buf_clk new_AGEMA_reg_buffer_2814 ( .C (clk), .D (new_AGEMA_signal_6278), .Q (new_AGEMA_signal_6279) ) ;
    buf_clk new_AGEMA_reg_buffer_2820 ( .C (clk), .D (new_AGEMA_signal_6284), .Q (new_AGEMA_signal_6285) ) ;
    buf_clk new_AGEMA_reg_buffer_2826 ( .C (clk), .D (new_AGEMA_signal_6290), .Q (new_AGEMA_signal_6291) ) ;
    buf_clk new_AGEMA_reg_buffer_2832 ( .C (clk), .D (new_AGEMA_signal_6296), .Q (new_AGEMA_signal_6297) ) ;
    buf_clk new_AGEMA_reg_buffer_2838 ( .C (clk), .D (new_AGEMA_signal_6302), .Q (new_AGEMA_signal_6303) ) ;
    buf_clk new_AGEMA_reg_buffer_2844 ( .C (clk), .D (new_AGEMA_signal_6308), .Q (new_AGEMA_signal_6309) ) ;
    buf_clk new_AGEMA_reg_buffer_2850 ( .C (clk), .D (new_AGEMA_signal_6314), .Q (new_AGEMA_signal_6315) ) ;
    buf_clk new_AGEMA_reg_buffer_2856 ( .C (clk), .D (new_AGEMA_signal_6320), .Q (new_AGEMA_signal_6321) ) ;
    buf_clk new_AGEMA_reg_buffer_2862 ( .C (clk), .D (new_AGEMA_signal_6326), .Q (new_AGEMA_signal_6327) ) ;
    buf_clk new_AGEMA_reg_buffer_2868 ( .C (clk), .D (new_AGEMA_signal_6332), .Q (new_AGEMA_signal_6333) ) ;
    buf_clk new_AGEMA_reg_buffer_2874 ( .C (clk), .D (new_AGEMA_signal_6338), .Q (new_AGEMA_signal_6339) ) ;
    buf_clk new_AGEMA_reg_buffer_2880 ( .C (clk), .D (new_AGEMA_signal_6344), .Q (new_AGEMA_signal_6345) ) ;
    buf_clk new_AGEMA_reg_buffer_2886 ( .C (clk), .D (new_AGEMA_signal_6350), .Q (new_AGEMA_signal_6351) ) ;
    buf_clk new_AGEMA_reg_buffer_2892 ( .C (clk), .D (new_AGEMA_signal_6356), .Q (new_AGEMA_signal_6357) ) ;
    buf_clk new_AGEMA_reg_buffer_2898 ( .C (clk), .D (new_AGEMA_signal_6362), .Q (new_AGEMA_signal_6363) ) ;
    buf_clk new_AGEMA_reg_buffer_2904 ( .C (clk), .D (new_AGEMA_signal_6368), .Q (new_AGEMA_signal_6369) ) ;
    buf_clk new_AGEMA_reg_buffer_2910 ( .C (clk), .D (new_AGEMA_signal_6374), .Q (new_AGEMA_signal_6375) ) ;
    buf_clk new_AGEMA_reg_buffer_2916 ( .C (clk), .D (new_AGEMA_signal_6380), .Q (new_AGEMA_signal_6381) ) ;
    buf_clk new_AGEMA_reg_buffer_2922 ( .C (clk), .D (new_AGEMA_signal_6386), .Q (new_AGEMA_signal_6387) ) ;
    buf_clk new_AGEMA_reg_buffer_2928 ( .C (clk), .D (new_AGEMA_signal_6392), .Q (new_AGEMA_signal_6393) ) ;
    buf_clk new_AGEMA_reg_buffer_2934 ( .C (clk), .D (new_AGEMA_signal_6398), .Q (new_AGEMA_signal_6399) ) ;
    buf_clk new_AGEMA_reg_buffer_2940 ( .C (clk), .D (new_AGEMA_signal_6404), .Q (new_AGEMA_signal_6405) ) ;
    buf_clk new_AGEMA_reg_buffer_2946 ( .C (clk), .D (new_AGEMA_signal_6410), .Q (new_AGEMA_signal_6411) ) ;
    buf_clk new_AGEMA_reg_buffer_2952 ( .C (clk), .D (new_AGEMA_signal_6416), .Q (new_AGEMA_signal_6417) ) ;
    buf_clk new_AGEMA_reg_buffer_2958 ( .C (clk), .D (new_AGEMA_signal_6422), .Q (new_AGEMA_signal_6423) ) ;
    buf_clk new_AGEMA_reg_buffer_2964 ( .C (clk), .D (new_AGEMA_signal_6428), .Q (new_AGEMA_signal_6429) ) ;
    buf_clk new_AGEMA_reg_buffer_2970 ( .C (clk), .D (new_AGEMA_signal_6434), .Q (new_AGEMA_signal_6435) ) ;
    buf_clk new_AGEMA_reg_buffer_2976 ( .C (clk), .D (new_AGEMA_signal_6440), .Q (new_AGEMA_signal_6441) ) ;
    buf_clk new_AGEMA_reg_buffer_2982 ( .C (clk), .D (new_AGEMA_signal_6446), .Q (new_AGEMA_signal_6447) ) ;
    buf_clk new_AGEMA_reg_buffer_2988 ( .C (clk), .D (new_AGEMA_signal_6452), .Q (new_AGEMA_signal_6453) ) ;
    buf_clk new_AGEMA_reg_buffer_2994 ( .C (clk), .D (new_AGEMA_signal_6458), .Q (new_AGEMA_signal_6459) ) ;
    buf_clk new_AGEMA_reg_buffer_3000 ( .C (clk), .D (new_AGEMA_signal_6464), .Q (new_AGEMA_signal_6465) ) ;
    buf_clk new_AGEMA_reg_buffer_3006 ( .C (clk), .D (new_AGEMA_signal_6470), .Q (new_AGEMA_signal_6471) ) ;
    buf_clk new_AGEMA_reg_buffer_3012 ( .C (clk), .D (new_AGEMA_signal_6476), .Q (new_AGEMA_signal_6477) ) ;
    buf_clk new_AGEMA_reg_buffer_3018 ( .C (clk), .D (new_AGEMA_signal_6482), .Q (new_AGEMA_signal_6483) ) ;
    buf_clk new_AGEMA_reg_buffer_3024 ( .C (clk), .D (new_AGEMA_signal_6488), .Q (new_AGEMA_signal_6489) ) ;
    buf_clk new_AGEMA_reg_buffer_3030 ( .C (clk), .D (new_AGEMA_signal_6494), .Q (new_AGEMA_signal_6495) ) ;
    buf_clk new_AGEMA_reg_buffer_3036 ( .C (clk), .D (new_AGEMA_signal_6500), .Q (new_AGEMA_signal_6501) ) ;
    buf_clk new_AGEMA_reg_buffer_3042 ( .C (clk), .D (new_AGEMA_signal_6506), .Q (new_AGEMA_signal_6507) ) ;
    buf_clk new_AGEMA_reg_buffer_3048 ( .C (clk), .D (new_AGEMA_signal_6512), .Q (new_AGEMA_signal_6513) ) ;
    buf_clk new_AGEMA_reg_buffer_3054 ( .C (clk), .D (new_AGEMA_signal_6518), .Q (new_AGEMA_signal_6519) ) ;
    buf_clk new_AGEMA_reg_buffer_3060 ( .C (clk), .D (new_AGEMA_signal_6524), .Q (new_AGEMA_signal_6525) ) ;
    buf_clk new_AGEMA_reg_buffer_3066 ( .C (clk), .D (new_AGEMA_signal_6530), .Q (new_AGEMA_signal_6531) ) ;
    buf_clk new_AGEMA_reg_buffer_3072 ( .C (clk), .D (new_AGEMA_signal_6536), .Q (new_AGEMA_signal_6537) ) ;
    buf_clk new_AGEMA_reg_buffer_3078 ( .C (clk), .D (new_AGEMA_signal_6542), .Q (new_AGEMA_signal_6543) ) ;
    buf_clk new_AGEMA_reg_buffer_3084 ( .C (clk), .D (new_AGEMA_signal_6548), .Q (new_AGEMA_signal_6549) ) ;
    buf_clk new_AGEMA_reg_buffer_3090 ( .C (clk), .D (new_AGEMA_signal_6554), .Q (new_AGEMA_signal_6555) ) ;
    buf_clk new_AGEMA_reg_buffer_3096 ( .C (clk), .D (new_AGEMA_signal_6560), .Q (new_AGEMA_signal_6561) ) ;
    buf_clk new_AGEMA_reg_buffer_3102 ( .C (clk), .D (new_AGEMA_signal_6566), .Q (new_AGEMA_signal_6567) ) ;
    buf_clk new_AGEMA_reg_buffer_3108 ( .C (clk), .D (new_AGEMA_signal_6572), .Q (new_AGEMA_signal_6573) ) ;
    buf_clk new_AGEMA_reg_buffer_3114 ( .C (clk), .D (new_AGEMA_signal_6578), .Q (new_AGEMA_signal_6579) ) ;
    buf_clk new_AGEMA_reg_buffer_3120 ( .C (clk), .D (new_AGEMA_signal_6584), .Q (new_AGEMA_signal_6585) ) ;
    buf_clk new_AGEMA_reg_buffer_3126 ( .C (clk), .D (new_AGEMA_signal_6590), .Q (new_AGEMA_signal_6591) ) ;
    buf_clk new_AGEMA_reg_buffer_3132 ( .C (clk), .D (new_AGEMA_signal_6596), .Q (new_AGEMA_signal_6597) ) ;
    buf_clk new_AGEMA_reg_buffer_3138 ( .C (clk), .D (new_AGEMA_signal_6602), .Q (new_AGEMA_signal_6603) ) ;
    buf_clk new_AGEMA_reg_buffer_3144 ( .C (clk), .D (new_AGEMA_signal_6608), .Q (new_AGEMA_signal_6609) ) ;
    buf_clk new_AGEMA_reg_buffer_3150 ( .C (clk), .D (new_AGEMA_signal_6614), .Q (new_AGEMA_signal_6615) ) ;
    buf_clk new_AGEMA_reg_buffer_3156 ( .C (clk), .D (new_AGEMA_signal_6620), .Q (new_AGEMA_signal_6621) ) ;
    buf_clk new_AGEMA_reg_buffer_3162 ( .C (clk), .D (new_AGEMA_signal_6626), .Q (new_AGEMA_signal_6627) ) ;
    buf_clk new_AGEMA_reg_buffer_3168 ( .C (clk), .D (new_AGEMA_signal_6632), .Q (new_AGEMA_signal_6633) ) ;
    buf_clk new_AGEMA_reg_buffer_3174 ( .C (clk), .D (new_AGEMA_signal_6638), .Q (new_AGEMA_signal_6639) ) ;
    buf_clk new_AGEMA_reg_buffer_3180 ( .C (clk), .D (new_AGEMA_signal_6644), .Q (new_AGEMA_signal_6645) ) ;
    buf_clk new_AGEMA_reg_buffer_3186 ( .C (clk), .D (new_AGEMA_signal_6650), .Q (new_AGEMA_signal_6651) ) ;
    buf_clk new_AGEMA_reg_buffer_3192 ( .C (clk), .D (new_AGEMA_signal_6656), .Q (new_AGEMA_signal_6657) ) ;
    buf_clk new_AGEMA_reg_buffer_3198 ( .C (clk), .D (new_AGEMA_signal_6662), .Q (new_AGEMA_signal_6663) ) ;
    buf_clk new_AGEMA_reg_buffer_3204 ( .C (clk), .D (new_AGEMA_signal_6668), .Q (new_AGEMA_signal_6669) ) ;
    buf_clk new_AGEMA_reg_buffer_3210 ( .C (clk), .D (new_AGEMA_signal_6674), .Q (new_AGEMA_signal_6675) ) ;
    buf_clk new_AGEMA_reg_buffer_3216 ( .C (clk), .D (new_AGEMA_signal_6680), .Q (new_AGEMA_signal_6681) ) ;
    buf_clk new_AGEMA_reg_buffer_3222 ( .C (clk), .D (new_AGEMA_signal_6686), .Q (new_AGEMA_signal_6687) ) ;
    buf_clk new_AGEMA_reg_buffer_3228 ( .C (clk), .D (new_AGEMA_signal_6692), .Q (new_AGEMA_signal_6693) ) ;
    buf_clk new_AGEMA_reg_buffer_3234 ( .C (clk), .D (new_AGEMA_signal_6698), .Q (new_AGEMA_signal_6699) ) ;
    buf_clk new_AGEMA_reg_buffer_3240 ( .C (clk), .D (new_AGEMA_signal_6704), .Q (new_AGEMA_signal_6705) ) ;
    buf_clk new_AGEMA_reg_buffer_3246 ( .C (clk), .D (new_AGEMA_signal_6710), .Q (new_AGEMA_signal_6711) ) ;
    buf_clk new_AGEMA_reg_buffer_3252 ( .C (clk), .D (new_AGEMA_signal_6716), .Q (new_AGEMA_signal_6717) ) ;
    buf_clk new_AGEMA_reg_buffer_3258 ( .C (clk), .D (new_AGEMA_signal_6722), .Q (new_AGEMA_signal_6723) ) ;
    buf_clk new_AGEMA_reg_buffer_3264 ( .C (clk), .D (new_AGEMA_signal_6728), .Q (new_AGEMA_signal_6729) ) ;
    buf_clk new_AGEMA_reg_buffer_3270 ( .C (clk), .D (new_AGEMA_signal_6734), .Q (new_AGEMA_signal_6735) ) ;
    buf_clk new_AGEMA_reg_buffer_3276 ( .C (clk), .D (new_AGEMA_signal_6740), .Q (new_AGEMA_signal_6741) ) ;
    buf_clk new_AGEMA_reg_buffer_3282 ( .C (clk), .D (new_AGEMA_signal_6746), .Q (new_AGEMA_signal_6747) ) ;
    buf_clk new_AGEMA_reg_buffer_3288 ( .C (clk), .D (new_AGEMA_signal_6752), .Q (new_AGEMA_signal_6753) ) ;
    buf_clk new_AGEMA_reg_buffer_3294 ( .C (clk), .D (new_AGEMA_signal_6758), .Q (new_AGEMA_signal_6759) ) ;
    buf_clk new_AGEMA_reg_buffer_3300 ( .C (clk), .D (new_AGEMA_signal_6764), .Q (new_AGEMA_signal_6765) ) ;
    buf_clk new_AGEMA_reg_buffer_3306 ( .C (clk), .D (new_AGEMA_signal_6770), .Q (new_AGEMA_signal_6771) ) ;
    buf_clk new_AGEMA_reg_buffer_3312 ( .C (clk), .D (new_AGEMA_signal_6776), .Q (new_AGEMA_signal_6777) ) ;
    buf_clk new_AGEMA_reg_buffer_3318 ( .C (clk), .D (new_AGEMA_signal_6782), .Q (new_AGEMA_signal_6783) ) ;
    buf_clk new_AGEMA_reg_buffer_3324 ( .C (clk), .D (new_AGEMA_signal_6788), .Q (new_AGEMA_signal_6789) ) ;
    buf_clk new_AGEMA_reg_buffer_3330 ( .C (clk), .D (new_AGEMA_signal_6794), .Q (new_AGEMA_signal_6795) ) ;
    buf_clk new_AGEMA_reg_buffer_3336 ( .C (clk), .D (new_AGEMA_signal_6800), .Q (new_AGEMA_signal_6801) ) ;
    buf_clk new_AGEMA_reg_buffer_3342 ( .C (clk), .D (new_AGEMA_signal_6806), .Q (new_AGEMA_signal_6807) ) ;
    buf_clk new_AGEMA_reg_buffer_3348 ( .C (clk), .D (new_AGEMA_signal_6812), .Q (new_AGEMA_signal_6813) ) ;
    buf_clk new_AGEMA_reg_buffer_3354 ( .C (clk), .D (new_AGEMA_signal_6818), .Q (new_AGEMA_signal_6819) ) ;
    buf_clk new_AGEMA_reg_buffer_3360 ( .C (clk), .D (new_AGEMA_signal_6824), .Q (new_AGEMA_signal_6825) ) ;
    buf_clk new_AGEMA_reg_buffer_3366 ( .C (clk), .D (new_AGEMA_signal_6830), .Q (new_AGEMA_signal_6831) ) ;
    buf_clk new_AGEMA_reg_buffer_3372 ( .C (clk), .D (new_AGEMA_signal_6836), .Q (new_AGEMA_signal_6837) ) ;
    buf_clk new_AGEMA_reg_buffer_3378 ( .C (clk), .D (new_AGEMA_signal_6842), .Q (new_AGEMA_signal_6843) ) ;
    buf_clk new_AGEMA_reg_buffer_3384 ( .C (clk), .D (new_AGEMA_signal_6848), .Q (new_AGEMA_signal_6849) ) ;
    buf_clk new_AGEMA_reg_buffer_3390 ( .C (clk), .D (new_AGEMA_signal_6854), .Q (new_AGEMA_signal_6855) ) ;
    buf_clk new_AGEMA_reg_buffer_3396 ( .C (clk), .D (new_AGEMA_signal_6860), .Q (new_AGEMA_signal_6861) ) ;
    buf_clk new_AGEMA_reg_buffer_3402 ( .C (clk), .D (new_AGEMA_signal_6866), .Q (new_AGEMA_signal_6867) ) ;
    buf_clk new_AGEMA_reg_buffer_3408 ( .C (clk), .D (new_AGEMA_signal_6872), .Q (new_AGEMA_signal_6873) ) ;
    buf_clk new_AGEMA_reg_buffer_3414 ( .C (clk), .D (new_AGEMA_signal_6878), .Q (new_AGEMA_signal_6879) ) ;
    buf_clk new_AGEMA_reg_buffer_3420 ( .C (clk), .D (new_AGEMA_signal_6884), .Q (new_AGEMA_signal_6885) ) ;
    buf_clk new_AGEMA_reg_buffer_3426 ( .C (clk), .D (new_AGEMA_signal_6890), .Q (new_AGEMA_signal_6891) ) ;
    buf_clk new_AGEMA_reg_buffer_3432 ( .C (clk), .D (new_AGEMA_signal_6896), .Q (new_AGEMA_signal_6897) ) ;
    buf_clk new_AGEMA_reg_buffer_3438 ( .C (clk), .D (new_AGEMA_signal_6902), .Q (new_AGEMA_signal_6903) ) ;
    buf_clk new_AGEMA_reg_buffer_3444 ( .C (clk), .D (new_AGEMA_signal_6908), .Q (new_AGEMA_signal_6909) ) ;
    buf_clk new_AGEMA_reg_buffer_3450 ( .C (clk), .D (new_AGEMA_signal_6914), .Q (new_AGEMA_signal_6915) ) ;
    buf_clk new_AGEMA_reg_buffer_3456 ( .C (clk), .D (new_AGEMA_signal_6920), .Q (new_AGEMA_signal_6921) ) ;
    buf_clk new_AGEMA_reg_buffer_3462 ( .C (clk), .D (new_AGEMA_signal_6926), .Q (new_AGEMA_signal_6927) ) ;
    buf_clk new_AGEMA_reg_buffer_3468 ( .C (clk), .D (new_AGEMA_signal_6932), .Q (new_AGEMA_signal_6933) ) ;
    buf_clk new_AGEMA_reg_buffer_3474 ( .C (clk), .D (new_AGEMA_signal_6938), .Q (new_AGEMA_signal_6939) ) ;
    buf_clk new_AGEMA_reg_buffer_3480 ( .C (clk), .D (new_AGEMA_signal_6944), .Q (new_AGEMA_signal_6945) ) ;
    buf_clk new_AGEMA_reg_buffer_3486 ( .C (clk), .D (new_AGEMA_signal_6950), .Q (new_AGEMA_signal_6951) ) ;
    buf_clk new_AGEMA_reg_buffer_3492 ( .C (clk), .D (new_AGEMA_signal_6956), .Q (new_AGEMA_signal_6957) ) ;
    buf_clk new_AGEMA_reg_buffer_3498 ( .C (clk), .D (new_AGEMA_signal_6962), .Q (new_AGEMA_signal_6963) ) ;
    buf_clk new_AGEMA_reg_buffer_3504 ( .C (clk), .D (new_AGEMA_signal_6968), .Q (new_AGEMA_signal_6969) ) ;
    buf_clk new_AGEMA_reg_buffer_3510 ( .C (clk), .D (new_AGEMA_signal_6974), .Q (new_AGEMA_signal_6975) ) ;
    buf_clk new_AGEMA_reg_buffer_3516 ( .C (clk), .D (new_AGEMA_signal_6980), .Q (new_AGEMA_signal_6981) ) ;
    buf_clk new_AGEMA_reg_buffer_3522 ( .C (clk), .D (new_AGEMA_signal_6986), .Q (new_AGEMA_signal_6987) ) ;
    buf_clk new_AGEMA_reg_buffer_3528 ( .C (clk), .D (new_AGEMA_signal_6992), .Q (new_AGEMA_signal_6993) ) ;
    buf_clk new_AGEMA_reg_buffer_3534 ( .C (clk), .D (new_AGEMA_signal_6998), .Q (new_AGEMA_signal_6999) ) ;
    buf_clk new_AGEMA_reg_buffer_3540 ( .C (clk), .D (new_AGEMA_signal_7004), .Q (new_AGEMA_signal_7005) ) ;
    buf_clk new_AGEMA_reg_buffer_3546 ( .C (clk), .D (new_AGEMA_signal_7010), .Q (new_AGEMA_signal_7011) ) ;
    buf_clk new_AGEMA_reg_buffer_3552 ( .C (clk), .D (new_AGEMA_signal_7016), .Q (new_AGEMA_signal_7017) ) ;
    buf_clk new_AGEMA_reg_buffer_3558 ( .C (clk), .D (new_AGEMA_signal_7022), .Q (new_AGEMA_signal_7023) ) ;
    buf_clk new_AGEMA_reg_buffer_3564 ( .C (clk), .D (new_AGEMA_signal_7028), .Q (new_AGEMA_signal_7029) ) ;
    buf_clk new_AGEMA_reg_buffer_3570 ( .C (clk), .D (new_AGEMA_signal_7034), .Q (new_AGEMA_signal_7035) ) ;
    buf_clk new_AGEMA_reg_buffer_3574 ( .C (clk), .D (new_AGEMA_signal_7038), .Q (new_AGEMA_signal_7039) ) ;
    buf_clk new_AGEMA_reg_buffer_3576 ( .C (clk), .D (new_AGEMA_signal_7040), .Q (new_AGEMA_signal_7041) ) ;
    buf_clk new_AGEMA_reg_buffer_3578 ( .C (clk), .D (new_AGEMA_signal_7042), .Q (new_AGEMA_signal_7043) ) ;
    buf_clk new_AGEMA_reg_buffer_3580 ( .C (clk), .D (new_AGEMA_signal_7044), .Q (new_AGEMA_signal_7045) ) ;
    buf_clk new_AGEMA_reg_buffer_3582 ( .C (clk), .D (new_AGEMA_signal_7046), .Q (new_AGEMA_signal_7047) ) ;
    buf_clk new_AGEMA_reg_buffer_3584 ( .C (clk), .D (new_AGEMA_signal_7048), .Q (new_AGEMA_signal_7049) ) ;
    buf_clk new_AGEMA_reg_buffer_3586 ( .C (clk), .D (new_AGEMA_signal_7050), .Q (new_AGEMA_signal_7051) ) ;
    buf_clk new_AGEMA_reg_buffer_3588 ( .C (clk), .D (new_AGEMA_signal_7052), .Q (new_AGEMA_signal_7053) ) ;
    buf_clk new_AGEMA_reg_buffer_3590 ( .C (clk), .D (new_AGEMA_signal_7054), .Q (new_AGEMA_signal_7055) ) ;
    buf_clk new_AGEMA_reg_buffer_3592 ( .C (clk), .D (new_AGEMA_signal_7056), .Q (new_AGEMA_signal_7057) ) ;
    buf_clk new_AGEMA_reg_buffer_3594 ( .C (clk), .D (new_AGEMA_signal_7058), .Q (new_AGEMA_signal_7059) ) ;
    buf_clk new_AGEMA_reg_buffer_3596 ( .C (clk), .D (new_AGEMA_signal_7060), .Q (new_AGEMA_signal_7061) ) ;
    buf_clk new_AGEMA_reg_buffer_3598 ( .C (clk), .D (new_AGEMA_signal_7062), .Q (new_AGEMA_signal_7063) ) ;
    buf_clk new_AGEMA_reg_buffer_3600 ( .C (clk), .D (new_AGEMA_signal_7064), .Q (new_AGEMA_signal_7065) ) ;
    buf_clk new_AGEMA_reg_buffer_3602 ( .C (clk), .D (new_AGEMA_signal_7066), .Q (new_AGEMA_signal_7067) ) ;
    buf_clk new_AGEMA_reg_buffer_3604 ( .C (clk), .D (new_AGEMA_signal_7068), .Q (new_AGEMA_signal_7069) ) ;
    buf_clk new_AGEMA_reg_buffer_3606 ( .C (clk), .D (new_AGEMA_signal_7070), .Q (new_AGEMA_signal_7071) ) ;
    buf_clk new_AGEMA_reg_buffer_3608 ( .C (clk), .D (new_AGEMA_signal_7072), .Q (new_AGEMA_signal_7073) ) ;
    buf_clk new_AGEMA_reg_buffer_3610 ( .C (clk), .D (new_AGEMA_signal_7074), .Q (new_AGEMA_signal_7075) ) ;
    buf_clk new_AGEMA_reg_buffer_3612 ( .C (clk), .D (new_AGEMA_signal_7076), .Q (new_AGEMA_signal_7077) ) ;
    buf_clk new_AGEMA_reg_buffer_3614 ( .C (clk), .D (new_AGEMA_signal_7078), .Q (new_AGEMA_signal_7079) ) ;
    buf_clk new_AGEMA_reg_buffer_3616 ( .C (clk), .D (new_AGEMA_signal_7080), .Q (new_AGEMA_signal_7081) ) ;
    buf_clk new_AGEMA_reg_buffer_3618 ( .C (clk), .D (new_AGEMA_signal_7082), .Q (new_AGEMA_signal_7083) ) ;
    buf_clk new_AGEMA_reg_buffer_3620 ( .C (clk), .D (new_AGEMA_signal_7084), .Q (new_AGEMA_signal_7085) ) ;
    buf_clk new_AGEMA_reg_buffer_3622 ( .C (clk), .D (new_AGEMA_signal_7086), .Q (new_AGEMA_signal_7087) ) ;
    buf_clk new_AGEMA_reg_buffer_3624 ( .C (clk), .D (new_AGEMA_signal_7088), .Q (new_AGEMA_signal_7089) ) ;
    buf_clk new_AGEMA_reg_buffer_3626 ( .C (clk), .D (new_AGEMA_signal_7090), .Q (new_AGEMA_signal_7091) ) ;
    buf_clk new_AGEMA_reg_buffer_3628 ( .C (clk), .D (new_AGEMA_signal_7092), .Q (new_AGEMA_signal_7093) ) ;
    buf_clk new_AGEMA_reg_buffer_3630 ( .C (clk), .D (new_AGEMA_signal_7094), .Q (new_AGEMA_signal_7095) ) ;
    buf_clk new_AGEMA_reg_buffer_3632 ( .C (clk), .D (new_AGEMA_signal_7096), .Q (new_AGEMA_signal_7097) ) ;
    buf_clk new_AGEMA_reg_buffer_3634 ( .C (clk), .D (new_AGEMA_signal_7098), .Q (new_AGEMA_signal_7099) ) ;
    buf_clk new_AGEMA_reg_buffer_3636 ( .C (clk), .D (new_AGEMA_signal_7100), .Q (new_AGEMA_signal_7101) ) ;
    buf_clk new_AGEMA_reg_buffer_3638 ( .C (clk), .D (new_AGEMA_signal_7102), .Q (new_AGEMA_signal_7103) ) ;
    buf_clk new_AGEMA_reg_buffer_3640 ( .C (clk), .D (new_AGEMA_signal_7104), .Q (new_AGEMA_signal_7105) ) ;
    buf_clk new_AGEMA_reg_buffer_3642 ( .C (clk), .D (new_AGEMA_signal_7106), .Q (new_AGEMA_signal_7107) ) ;
    buf_clk new_AGEMA_reg_buffer_3644 ( .C (clk), .D (new_AGEMA_signal_7108), .Q (new_AGEMA_signal_7109) ) ;
    buf_clk new_AGEMA_reg_buffer_3646 ( .C (clk), .D (new_AGEMA_signal_7110), .Q (new_AGEMA_signal_7111) ) ;
    buf_clk new_AGEMA_reg_buffer_3648 ( .C (clk), .D (new_AGEMA_signal_7112), .Q (new_AGEMA_signal_7113) ) ;
    buf_clk new_AGEMA_reg_buffer_3650 ( .C (clk), .D (new_AGEMA_signal_7114), .Q (new_AGEMA_signal_7115) ) ;
    buf_clk new_AGEMA_reg_buffer_3652 ( .C (clk), .D (new_AGEMA_signal_7116), .Q (new_AGEMA_signal_7117) ) ;
    buf_clk new_AGEMA_reg_buffer_3654 ( .C (clk), .D (new_AGEMA_signal_7118), .Q (new_AGEMA_signal_7119) ) ;
    buf_clk new_AGEMA_reg_buffer_3656 ( .C (clk), .D (new_AGEMA_signal_7120), .Q (new_AGEMA_signal_7121) ) ;
    buf_clk new_AGEMA_reg_buffer_3658 ( .C (clk), .D (new_AGEMA_signal_7122), .Q (new_AGEMA_signal_7123) ) ;
    buf_clk new_AGEMA_reg_buffer_3660 ( .C (clk), .D (new_AGEMA_signal_7124), .Q (new_AGEMA_signal_7125) ) ;
    buf_clk new_AGEMA_reg_buffer_3662 ( .C (clk), .D (new_AGEMA_signal_7126), .Q (new_AGEMA_signal_7127) ) ;
    buf_clk new_AGEMA_reg_buffer_3664 ( .C (clk), .D (new_AGEMA_signal_7128), .Q (new_AGEMA_signal_7129) ) ;
    buf_clk new_AGEMA_reg_buffer_3666 ( .C (clk), .D (new_AGEMA_signal_7130), .Q (new_AGEMA_signal_7131) ) ;
    buf_clk new_AGEMA_reg_buffer_3668 ( .C (clk), .D (new_AGEMA_signal_7132), .Q (new_AGEMA_signal_7133) ) ;
    buf_clk new_AGEMA_reg_buffer_3670 ( .C (clk), .D (new_AGEMA_signal_7134), .Q (new_AGEMA_signal_7135) ) ;
    buf_clk new_AGEMA_reg_buffer_3672 ( .C (clk), .D (new_AGEMA_signal_7136), .Q (new_AGEMA_signal_7137) ) ;
    buf_clk new_AGEMA_reg_buffer_3674 ( .C (clk), .D (new_AGEMA_signal_7138), .Q (new_AGEMA_signal_7139) ) ;
    buf_clk new_AGEMA_reg_buffer_3676 ( .C (clk), .D (new_AGEMA_signal_7140), .Q (new_AGEMA_signal_7141) ) ;
    buf_clk new_AGEMA_reg_buffer_3678 ( .C (clk), .D (new_AGEMA_signal_7142), .Q (new_AGEMA_signal_7143) ) ;
    buf_clk new_AGEMA_reg_buffer_3680 ( .C (clk), .D (new_AGEMA_signal_7144), .Q (new_AGEMA_signal_7145) ) ;
    buf_clk new_AGEMA_reg_buffer_3682 ( .C (clk), .D (new_AGEMA_signal_7146), .Q (new_AGEMA_signal_7147) ) ;
    buf_clk new_AGEMA_reg_buffer_3684 ( .C (clk), .D (new_AGEMA_signal_7148), .Q (new_AGEMA_signal_7149) ) ;
    buf_clk new_AGEMA_reg_buffer_3686 ( .C (clk), .D (new_AGEMA_signal_7150), .Q (new_AGEMA_signal_7151) ) ;
    buf_clk new_AGEMA_reg_buffer_3688 ( .C (clk), .D (new_AGEMA_signal_7152), .Q (new_AGEMA_signal_7153) ) ;
    buf_clk new_AGEMA_reg_buffer_3690 ( .C (clk), .D (new_AGEMA_signal_7154), .Q (new_AGEMA_signal_7155) ) ;
    buf_clk new_AGEMA_reg_buffer_3692 ( .C (clk), .D (new_AGEMA_signal_7156), .Q (new_AGEMA_signal_7157) ) ;
    buf_clk new_AGEMA_reg_buffer_3694 ( .C (clk), .D (new_AGEMA_signal_7158), .Q (new_AGEMA_signal_7159) ) ;
    buf_clk new_AGEMA_reg_buffer_3696 ( .C (clk), .D (new_AGEMA_signal_7160), .Q (new_AGEMA_signal_7161) ) ;
    buf_clk new_AGEMA_reg_buffer_3698 ( .C (clk), .D (new_AGEMA_signal_7162), .Q (new_AGEMA_signal_7163) ) ;
    buf_clk new_AGEMA_reg_buffer_3700 ( .C (clk), .D (new_AGEMA_signal_7164), .Q (new_AGEMA_signal_7165) ) ;
    buf_clk new_AGEMA_reg_buffer_3702 ( .C (clk), .D (new_AGEMA_signal_7166), .Q (new_AGEMA_signal_7167) ) ;
    buf_clk new_AGEMA_reg_buffer_3704 ( .C (clk), .D (new_AGEMA_signal_7168), .Q (new_AGEMA_signal_7169) ) ;
    buf_clk new_AGEMA_reg_buffer_3706 ( .C (clk), .D (new_AGEMA_signal_7170), .Q (new_AGEMA_signal_7171) ) ;
    buf_clk new_AGEMA_reg_buffer_3708 ( .C (clk), .D (new_AGEMA_signal_7172), .Q (new_AGEMA_signal_7173) ) ;
    buf_clk new_AGEMA_reg_buffer_3710 ( .C (clk), .D (new_AGEMA_signal_7174), .Q (new_AGEMA_signal_7175) ) ;
    buf_clk new_AGEMA_reg_buffer_3712 ( .C (clk), .D (new_AGEMA_signal_7176), .Q (new_AGEMA_signal_7177) ) ;
    buf_clk new_AGEMA_reg_buffer_3714 ( .C (clk), .D (new_AGEMA_signal_7178), .Q (new_AGEMA_signal_7179) ) ;
    buf_clk new_AGEMA_reg_buffer_3716 ( .C (clk), .D (new_AGEMA_signal_7180), .Q (new_AGEMA_signal_7181) ) ;
    buf_clk new_AGEMA_reg_buffer_3718 ( .C (clk), .D (new_AGEMA_signal_7182), .Q (new_AGEMA_signal_7183) ) ;
    buf_clk new_AGEMA_reg_buffer_3720 ( .C (clk), .D (new_AGEMA_signal_7184), .Q (new_AGEMA_signal_7185) ) ;
    buf_clk new_AGEMA_reg_buffer_3722 ( .C (clk), .D (new_AGEMA_signal_7186), .Q (new_AGEMA_signal_7187) ) ;
    buf_clk new_AGEMA_reg_buffer_3724 ( .C (clk), .D (new_AGEMA_signal_7188), .Q (new_AGEMA_signal_7189) ) ;
    buf_clk new_AGEMA_reg_buffer_3726 ( .C (clk), .D (new_AGEMA_signal_7190), .Q (new_AGEMA_signal_7191) ) ;
    buf_clk new_AGEMA_reg_buffer_3728 ( .C (clk), .D (new_AGEMA_signal_7192), .Q (new_AGEMA_signal_7193) ) ;
    buf_clk new_AGEMA_reg_buffer_3730 ( .C (clk), .D (new_AGEMA_signal_7194), .Q (new_AGEMA_signal_7195) ) ;
    buf_clk new_AGEMA_reg_buffer_3732 ( .C (clk), .D (new_AGEMA_signal_7196), .Q (new_AGEMA_signal_7197) ) ;
    buf_clk new_AGEMA_reg_buffer_3734 ( .C (clk), .D (new_AGEMA_signal_7198), .Q (new_AGEMA_signal_7199) ) ;
    buf_clk new_AGEMA_reg_buffer_3736 ( .C (clk), .D (new_AGEMA_signal_7200), .Q (new_AGEMA_signal_7201) ) ;
    buf_clk new_AGEMA_reg_buffer_3738 ( .C (clk), .D (new_AGEMA_signal_7202), .Q (new_AGEMA_signal_7203) ) ;
    buf_clk new_AGEMA_reg_buffer_3740 ( .C (clk), .D (new_AGEMA_signal_7204), .Q (new_AGEMA_signal_7205) ) ;
    buf_clk new_AGEMA_reg_buffer_3742 ( .C (clk), .D (new_AGEMA_signal_7206), .Q (new_AGEMA_signal_7207) ) ;
    buf_clk new_AGEMA_reg_buffer_3744 ( .C (clk), .D (new_AGEMA_signal_7208), .Q (new_AGEMA_signal_7209) ) ;
    buf_clk new_AGEMA_reg_buffer_3746 ( .C (clk), .D (new_AGEMA_signal_7210), .Q (new_AGEMA_signal_7211) ) ;
    buf_clk new_AGEMA_reg_buffer_3748 ( .C (clk), .D (new_AGEMA_signal_7212), .Q (new_AGEMA_signal_7213) ) ;
    buf_clk new_AGEMA_reg_buffer_3750 ( .C (clk), .D (new_AGEMA_signal_7214), .Q (new_AGEMA_signal_7215) ) ;
    buf_clk new_AGEMA_reg_buffer_3752 ( .C (clk), .D (new_AGEMA_signal_7216), .Q (new_AGEMA_signal_7217) ) ;
    buf_clk new_AGEMA_reg_buffer_3754 ( .C (clk), .D (new_AGEMA_signal_7218), .Q (new_AGEMA_signal_7219) ) ;
    buf_clk new_AGEMA_reg_buffer_3756 ( .C (clk), .D (new_AGEMA_signal_7220), .Q (new_AGEMA_signal_7221) ) ;
    buf_clk new_AGEMA_reg_buffer_3758 ( .C (clk), .D (new_AGEMA_signal_7222), .Q (new_AGEMA_signal_7223) ) ;
    buf_clk new_AGEMA_reg_buffer_3760 ( .C (clk), .D (new_AGEMA_signal_7224), .Q (new_AGEMA_signal_7225) ) ;
    buf_clk new_AGEMA_reg_buffer_3762 ( .C (clk), .D (new_AGEMA_signal_7226), .Q (new_AGEMA_signal_7227) ) ;
    buf_clk new_AGEMA_reg_buffer_3764 ( .C (clk), .D (new_AGEMA_signal_7228), .Q (new_AGEMA_signal_7229) ) ;
    buf_clk new_AGEMA_reg_buffer_3766 ( .C (clk), .D (new_AGEMA_signal_7230), .Q (new_AGEMA_signal_7231) ) ;
    buf_clk new_AGEMA_reg_buffer_3768 ( .C (clk), .D (new_AGEMA_signal_7232), .Q (new_AGEMA_signal_7233) ) ;
    buf_clk new_AGEMA_reg_buffer_3770 ( .C (clk), .D (new_AGEMA_signal_7234), .Q (new_AGEMA_signal_7235) ) ;
    buf_clk new_AGEMA_reg_buffer_3772 ( .C (clk), .D (new_AGEMA_signal_7236), .Q (new_AGEMA_signal_7237) ) ;
    buf_clk new_AGEMA_reg_buffer_3774 ( .C (clk), .D (new_AGEMA_signal_7238), .Q (new_AGEMA_signal_7239) ) ;
    buf_clk new_AGEMA_reg_buffer_3776 ( .C (clk), .D (new_AGEMA_signal_7240), .Q (new_AGEMA_signal_7241) ) ;
    buf_clk new_AGEMA_reg_buffer_3778 ( .C (clk), .D (new_AGEMA_signal_7242), .Q (new_AGEMA_signal_7243) ) ;
    buf_clk new_AGEMA_reg_buffer_3780 ( .C (clk), .D (new_AGEMA_signal_7244), .Q (new_AGEMA_signal_7245) ) ;
    buf_clk new_AGEMA_reg_buffer_3782 ( .C (clk), .D (new_AGEMA_signal_7246), .Q (new_AGEMA_signal_7247) ) ;
    buf_clk new_AGEMA_reg_buffer_3784 ( .C (clk), .D (new_AGEMA_signal_7248), .Q (new_AGEMA_signal_7249) ) ;
    buf_clk new_AGEMA_reg_buffer_3786 ( .C (clk), .D (new_AGEMA_signal_7250), .Q (new_AGEMA_signal_7251) ) ;
    buf_clk new_AGEMA_reg_buffer_3788 ( .C (clk), .D (new_AGEMA_signal_7252), .Q (new_AGEMA_signal_7253) ) ;
    buf_clk new_AGEMA_reg_buffer_3790 ( .C (clk), .D (new_AGEMA_signal_7254), .Q (new_AGEMA_signal_7255) ) ;
    buf_clk new_AGEMA_reg_buffer_3792 ( .C (clk), .D (new_AGEMA_signal_7256), .Q (new_AGEMA_signal_7257) ) ;
    buf_clk new_AGEMA_reg_buffer_3794 ( .C (clk), .D (new_AGEMA_signal_7258), .Q (new_AGEMA_signal_7259) ) ;
    buf_clk new_AGEMA_reg_buffer_3796 ( .C (clk), .D (new_AGEMA_signal_7260), .Q (new_AGEMA_signal_7261) ) ;
    buf_clk new_AGEMA_reg_buffer_3798 ( .C (clk), .D (new_AGEMA_signal_7262), .Q (new_AGEMA_signal_7263) ) ;
    buf_clk new_AGEMA_reg_buffer_3800 ( .C (clk), .D (new_AGEMA_signal_7264), .Q (new_AGEMA_signal_7265) ) ;
    buf_clk new_AGEMA_reg_buffer_3802 ( .C (clk), .D (new_AGEMA_signal_7266), .Q (new_AGEMA_signal_7267) ) ;
    buf_clk new_AGEMA_reg_buffer_3804 ( .C (clk), .D (new_AGEMA_signal_7268), .Q (new_AGEMA_signal_7269) ) ;
    buf_clk new_AGEMA_reg_buffer_3806 ( .C (clk), .D (new_AGEMA_signal_7270), .Q (new_AGEMA_signal_7271) ) ;
    buf_clk new_AGEMA_reg_buffer_3808 ( .C (clk), .D (new_AGEMA_signal_7272), .Q (new_AGEMA_signal_7273) ) ;
    buf_clk new_AGEMA_reg_buffer_3810 ( .C (clk), .D (new_AGEMA_signal_7274), .Q (new_AGEMA_signal_7275) ) ;
    buf_clk new_AGEMA_reg_buffer_3812 ( .C (clk), .D (new_AGEMA_signal_7276), .Q (new_AGEMA_signal_7277) ) ;
    buf_clk new_AGEMA_reg_buffer_3814 ( .C (clk), .D (new_AGEMA_signal_7278), .Q (new_AGEMA_signal_7279) ) ;
    buf_clk new_AGEMA_reg_buffer_3816 ( .C (clk), .D (new_AGEMA_signal_7280), .Q (new_AGEMA_signal_7281) ) ;
    buf_clk new_AGEMA_reg_buffer_3818 ( .C (clk), .D (new_AGEMA_signal_7282), .Q (new_AGEMA_signal_7283) ) ;
    buf_clk new_AGEMA_reg_buffer_3820 ( .C (clk), .D (new_AGEMA_signal_7284), .Q (new_AGEMA_signal_7285) ) ;
    buf_clk new_AGEMA_reg_buffer_3822 ( .C (clk), .D (new_AGEMA_signal_7286), .Q (new_AGEMA_signal_7287) ) ;
    buf_clk new_AGEMA_reg_buffer_3824 ( .C (clk), .D (new_AGEMA_signal_7288), .Q (new_AGEMA_signal_7289) ) ;
    buf_clk new_AGEMA_reg_buffer_3826 ( .C (clk), .D (new_AGEMA_signal_7290), .Q (new_AGEMA_signal_7291) ) ;
    buf_clk new_AGEMA_reg_buffer_3828 ( .C (clk), .D (new_AGEMA_signal_7292), .Q (new_AGEMA_signal_7293) ) ;
    buf_clk new_AGEMA_reg_buffer_3830 ( .C (clk), .D (new_AGEMA_signal_7294), .Q (new_AGEMA_signal_7295) ) ;
    buf_clk new_AGEMA_reg_buffer_3832 ( .C (clk), .D (new_AGEMA_signal_7296), .Q (new_AGEMA_signal_7297) ) ;
    buf_clk new_AGEMA_reg_buffer_3834 ( .C (clk), .D (new_AGEMA_signal_7298), .Q (new_AGEMA_signal_7299) ) ;
    buf_clk new_AGEMA_reg_buffer_3836 ( .C (clk), .D (new_AGEMA_signal_7300), .Q (new_AGEMA_signal_7301) ) ;
    buf_clk new_AGEMA_reg_buffer_3838 ( .C (clk), .D (new_AGEMA_signal_7302), .Q (new_AGEMA_signal_7303) ) ;
    buf_clk new_AGEMA_reg_buffer_3840 ( .C (clk), .D (new_AGEMA_signal_7304), .Q (new_AGEMA_signal_7305) ) ;
    buf_clk new_AGEMA_reg_buffer_3842 ( .C (clk), .D (new_AGEMA_signal_7306), .Q (new_AGEMA_signal_7307) ) ;
    buf_clk new_AGEMA_reg_buffer_3844 ( .C (clk), .D (new_AGEMA_signal_7308), .Q (new_AGEMA_signal_7309) ) ;
    buf_clk new_AGEMA_reg_buffer_3846 ( .C (clk), .D (new_AGEMA_signal_7310), .Q (new_AGEMA_signal_7311) ) ;
    buf_clk new_AGEMA_reg_buffer_3848 ( .C (clk), .D (new_AGEMA_signal_7312), .Q (new_AGEMA_signal_7313) ) ;
    buf_clk new_AGEMA_reg_buffer_3850 ( .C (clk), .D (new_AGEMA_signal_7314), .Q (new_AGEMA_signal_7315) ) ;
    buf_clk new_AGEMA_reg_buffer_3852 ( .C (clk), .D (new_AGEMA_signal_7316), .Q (new_AGEMA_signal_7317) ) ;
    buf_clk new_AGEMA_reg_buffer_3854 ( .C (clk), .D (new_AGEMA_signal_7318), .Q (new_AGEMA_signal_7319) ) ;
    buf_clk new_AGEMA_reg_buffer_3856 ( .C (clk), .D (new_AGEMA_signal_7320), .Q (new_AGEMA_signal_7321) ) ;
    buf_clk new_AGEMA_reg_buffer_3858 ( .C (clk), .D (new_AGEMA_signal_7322), .Q (new_AGEMA_signal_7323) ) ;
    buf_clk new_AGEMA_reg_buffer_3860 ( .C (clk), .D (new_AGEMA_signal_7324), .Q (new_AGEMA_signal_7325) ) ;
    buf_clk new_AGEMA_reg_buffer_3864 ( .C (clk), .D (new_AGEMA_signal_7328), .Q (new_AGEMA_signal_7329) ) ;
    buf_clk new_AGEMA_reg_buffer_3870 ( .C (clk), .D (new_AGEMA_signal_7334), .Q (new_AGEMA_signal_7335) ) ;
    buf_clk new_AGEMA_reg_buffer_3878 ( .C (clk), .D (new_AGEMA_signal_7342), .Q (new_AGEMA_signal_7343) ) ;
    buf_clk new_AGEMA_reg_buffer_3886 ( .C (clk), .D (new_AGEMA_signal_7350), .Q (new_AGEMA_signal_7351) ) ;
    buf_clk new_AGEMA_reg_buffer_3894 ( .C (clk), .D (new_AGEMA_signal_7358), .Q (new_AGEMA_signal_7359) ) ;
    buf_clk new_AGEMA_reg_buffer_3902 ( .C (clk), .D (new_AGEMA_signal_7366), .Q (new_AGEMA_signal_7367) ) ;
    buf_clk new_AGEMA_reg_buffer_3910 ( .C (clk), .D (new_AGEMA_signal_7374), .Q (new_AGEMA_signal_7375) ) ;
    buf_clk new_AGEMA_reg_buffer_3918 ( .C (clk), .D (new_AGEMA_signal_7382), .Q (new_AGEMA_signal_7383) ) ;
    buf_clk new_AGEMA_reg_buffer_3926 ( .C (clk), .D (new_AGEMA_signal_7390), .Q (new_AGEMA_signal_7391) ) ;
    buf_clk new_AGEMA_reg_buffer_3934 ( .C (clk), .D (new_AGEMA_signal_7398), .Q (new_AGEMA_signal_7399) ) ;
    buf_clk new_AGEMA_reg_buffer_3942 ( .C (clk), .D (new_AGEMA_signal_7406), .Q (new_AGEMA_signal_7407) ) ;
    buf_clk new_AGEMA_reg_buffer_3950 ( .C (clk), .D (new_AGEMA_signal_7414), .Q (new_AGEMA_signal_7415) ) ;
    buf_clk new_AGEMA_reg_buffer_3958 ( .C (clk), .D (new_AGEMA_signal_7422), .Q (new_AGEMA_signal_7423) ) ;
    buf_clk new_AGEMA_reg_buffer_3966 ( .C (clk), .D (new_AGEMA_signal_7430), .Q (new_AGEMA_signal_7431) ) ;
    buf_clk new_AGEMA_reg_buffer_3974 ( .C (clk), .D (new_AGEMA_signal_7438), .Q (new_AGEMA_signal_7439) ) ;
    buf_clk new_AGEMA_reg_buffer_3982 ( .C (clk), .D (new_AGEMA_signal_7446), .Q (new_AGEMA_signal_7447) ) ;
    buf_clk new_AGEMA_reg_buffer_3990 ( .C (clk), .D (new_AGEMA_signal_7454), .Q (new_AGEMA_signal_7455) ) ;
    buf_clk new_AGEMA_reg_buffer_3998 ( .C (clk), .D (new_AGEMA_signal_7462), .Q (new_AGEMA_signal_7463) ) ;
    buf_clk new_AGEMA_reg_buffer_4006 ( .C (clk), .D (new_AGEMA_signal_7470), .Q (new_AGEMA_signal_7471) ) ;
    buf_clk new_AGEMA_reg_buffer_4014 ( .C (clk), .D (new_AGEMA_signal_7478), .Q (new_AGEMA_signal_7479) ) ;
    buf_clk new_AGEMA_reg_buffer_4022 ( .C (clk), .D (new_AGEMA_signal_7486), .Q (new_AGEMA_signal_7487) ) ;
    buf_clk new_AGEMA_reg_buffer_4030 ( .C (clk), .D (new_AGEMA_signal_7494), .Q (new_AGEMA_signal_7495) ) ;
    buf_clk new_AGEMA_reg_buffer_4038 ( .C (clk), .D (new_AGEMA_signal_7502), .Q (new_AGEMA_signal_7503) ) ;
    buf_clk new_AGEMA_reg_buffer_4046 ( .C (clk), .D (new_AGEMA_signal_7510), .Q (new_AGEMA_signal_7511) ) ;
    buf_clk new_AGEMA_reg_buffer_4054 ( .C (clk), .D (new_AGEMA_signal_7518), .Q (new_AGEMA_signal_7519) ) ;
    buf_clk new_AGEMA_reg_buffer_4062 ( .C (clk), .D (new_AGEMA_signal_7526), .Q (new_AGEMA_signal_7527) ) ;
    buf_clk new_AGEMA_reg_buffer_4070 ( .C (clk), .D (new_AGEMA_signal_7534), .Q (new_AGEMA_signal_7535) ) ;
    buf_clk new_AGEMA_reg_buffer_4078 ( .C (clk), .D (new_AGEMA_signal_7542), .Q (new_AGEMA_signal_7543) ) ;
    buf_clk new_AGEMA_reg_buffer_4086 ( .C (clk), .D (new_AGEMA_signal_7550), .Q (new_AGEMA_signal_7551) ) ;
    buf_clk new_AGEMA_reg_buffer_4094 ( .C (clk), .D (new_AGEMA_signal_7558), .Q (new_AGEMA_signal_7559) ) ;
    buf_clk new_AGEMA_reg_buffer_4102 ( .C (clk), .D (new_AGEMA_signal_7566), .Q (new_AGEMA_signal_7567) ) ;
    buf_clk new_AGEMA_reg_buffer_4110 ( .C (clk), .D (new_AGEMA_signal_7574), .Q (new_AGEMA_signal_7575) ) ;
    buf_clk new_AGEMA_reg_buffer_4118 ( .C (clk), .D (new_AGEMA_signal_7582), .Q (new_AGEMA_signal_7583) ) ;
    buf_clk new_AGEMA_reg_buffer_4126 ( .C (clk), .D (new_AGEMA_signal_7590), .Q (new_AGEMA_signal_7591) ) ;
    buf_clk new_AGEMA_reg_buffer_4134 ( .C (clk), .D (new_AGEMA_signal_7598), .Q (new_AGEMA_signal_7599) ) ;
    buf_clk new_AGEMA_reg_buffer_4142 ( .C (clk), .D (new_AGEMA_signal_7606), .Q (new_AGEMA_signal_7607) ) ;
    buf_clk new_AGEMA_reg_buffer_4150 ( .C (clk), .D (new_AGEMA_signal_7614), .Q (new_AGEMA_signal_7615) ) ;
    buf_clk new_AGEMA_reg_buffer_4158 ( .C (clk), .D (new_AGEMA_signal_7622), .Q (new_AGEMA_signal_7623) ) ;
    buf_clk new_AGEMA_reg_buffer_4166 ( .C (clk), .D (new_AGEMA_signal_7630), .Q (new_AGEMA_signal_7631) ) ;
    buf_clk new_AGEMA_reg_buffer_4174 ( .C (clk), .D (new_AGEMA_signal_7638), .Q (new_AGEMA_signal_7639) ) ;
    buf_clk new_AGEMA_reg_buffer_4182 ( .C (clk), .D (new_AGEMA_signal_7646), .Q (new_AGEMA_signal_7647) ) ;
    buf_clk new_AGEMA_reg_buffer_4190 ( .C (clk), .D (new_AGEMA_signal_7654), .Q (new_AGEMA_signal_7655) ) ;
    buf_clk new_AGEMA_reg_buffer_4198 ( .C (clk), .D (new_AGEMA_signal_7662), .Q (new_AGEMA_signal_7663) ) ;
    buf_clk new_AGEMA_reg_buffer_4206 ( .C (clk), .D (new_AGEMA_signal_7670), .Q (new_AGEMA_signal_7671) ) ;
    buf_clk new_AGEMA_reg_buffer_4214 ( .C (clk), .D (new_AGEMA_signal_7678), .Q (new_AGEMA_signal_7679) ) ;
    buf_clk new_AGEMA_reg_buffer_4222 ( .C (clk), .D (new_AGEMA_signal_7686), .Q (new_AGEMA_signal_7687) ) ;
    buf_clk new_AGEMA_reg_buffer_4230 ( .C (clk), .D (new_AGEMA_signal_7694), .Q (new_AGEMA_signal_7695) ) ;
    buf_clk new_AGEMA_reg_buffer_4238 ( .C (clk), .D (new_AGEMA_signal_7702), .Q (new_AGEMA_signal_7703) ) ;
    buf_clk new_AGEMA_reg_buffer_4246 ( .C (clk), .D (new_AGEMA_signal_7710), .Q (new_AGEMA_signal_7711) ) ;
    buf_clk new_AGEMA_reg_buffer_4254 ( .C (clk), .D (new_AGEMA_signal_7718), .Q (new_AGEMA_signal_7719) ) ;
    buf_clk new_AGEMA_reg_buffer_4262 ( .C (clk), .D (new_AGEMA_signal_7726), .Q (new_AGEMA_signal_7727) ) ;
    buf_clk new_AGEMA_reg_buffer_4270 ( .C (clk), .D (new_AGEMA_signal_7734), .Q (new_AGEMA_signal_7735) ) ;
    buf_clk new_AGEMA_reg_buffer_4278 ( .C (clk), .D (new_AGEMA_signal_7742), .Q (new_AGEMA_signal_7743) ) ;
    buf_clk new_AGEMA_reg_buffer_4286 ( .C (clk), .D (new_AGEMA_signal_7750), .Q (new_AGEMA_signal_7751) ) ;
    buf_clk new_AGEMA_reg_buffer_4294 ( .C (clk), .D (new_AGEMA_signal_7758), .Q (new_AGEMA_signal_7759) ) ;
    buf_clk new_AGEMA_reg_buffer_4302 ( .C (clk), .D (new_AGEMA_signal_7766), .Q (new_AGEMA_signal_7767) ) ;
    buf_clk new_AGEMA_reg_buffer_4310 ( .C (clk), .D (new_AGEMA_signal_7774), .Q (new_AGEMA_signal_7775) ) ;
    buf_clk new_AGEMA_reg_buffer_4318 ( .C (clk), .D (new_AGEMA_signal_7782), .Q (new_AGEMA_signal_7783) ) ;
    buf_clk new_AGEMA_reg_buffer_4326 ( .C (clk), .D (new_AGEMA_signal_7790), .Q (new_AGEMA_signal_7791) ) ;
    buf_clk new_AGEMA_reg_buffer_4334 ( .C (clk), .D (new_AGEMA_signal_7798), .Q (new_AGEMA_signal_7799) ) ;
    buf_clk new_AGEMA_reg_buffer_4342 ( .C (clk), .D (new_AGEMA_signal_7806), .Q (new_AGEMA_signal_7807) ) ;
    buf_clk new_AGEMA_reg_buffer_4350 ( .C (clk), .D (new_AGEMA_signal_7814), .Q (new_AGEMA_signal_7815) ) ;
    buf_clk new_AGEMA_reg_buffer_4358 ( .C (clk), .D (new_AGEMA_signal_7822), .Q (new_AGEMA_signal_7823) ) ;
    buf_clk new_AGEMA_reg_buffer_4366 ( .C (clk), .D (new_AGEMA_signal_7830), .Q (new_AGEMA_signal_7831) ) ;
    buf_clk new_AGEMA_reg_buffer_4374 ( .C (clk), .D (new_AGEMA_signal_7838), .Q (new_AGEMA_signal_7839) ) ;
    buf_clk new_AGEMA_reg_buffer_4382 ( .C (clk), .D (new_AGEMA_signal_7846), .Q (new_AGEMA_signal_7847) ) ;
    buf_clk new_AGEMA_reg_buffer_4390 ( .C (clk), .D (new_AGEMA_signal_7854), .Q (new_AGEMA_signal_7855) ) ;
    buf_clk new_AGEMA_reg_buffer_4398 ( .C (clk), .D (new_AGEMA_signal_7862), .Q (new_AGEMA_signal_7863) ) ;
    buf_clk new_AGEMA_reg_buffer_4406 ( .C (clk), .D (new_AGEMA_signal_7870), .Q (new_AGEMA_signal_7871) ) ;
    buf_clk new_AGEMA_reg_buffer_4414 ( .C (clk), .D (new_AGEMA_signal_7878), .Q (new_AGEMA_signal_7879) ) ;
    buf_clk new_AGEMA_reg_buffer_4422 ( .C (clk), .D (new_AGEMA_signal_7886), .Q (new_AGEMA_signal_7887) ) ;
    buf_clk new_AGEMA_reg_buffer_4430 ( .C (clk), .D (new_AGEMA_signal_7894), .Q (new_AGEMA_signal_7895) ) ;
    buf_clk new_AGEMA_reg_buffer_4438 ( .C (clk), .D (new_AGEMA_signal_7902), .Q (new_AGEMA_signal_7903) ) ;
    buf_clk new_AGEMA_reg_buffer_4446 ( .C (clk), .D (new_AGEMA_signal_7910), .Q (new_AGEMA_signal_7911) ) ;
    buf_clk new_AGEMA_reg_buffer_4454 ( .C (clk), .D (new_AGEMA_signal_7918), .Q (new_AGEMA_signal_7919) ) ;
    buf_clk new_AGEMA_reg_buffer_4462 ( .C (clk), .D (new_AGEMA_signal_7926), .Q (new_AGEMA_signal_7927) ) ;
    buf_clk new_AGEMA_reg_buffer_4470 ( .C (clk), .D (new_AGEMA_signal_7934), .Q (new_AGEMA_signal_7935) ) ;
    buf_clk new_AGEMA_reg_buffer_4478 ( .C (clk), .D (new_AGEMA_signal_7942), .Q (new_AGEMA_signal_7943) ) ;
    buf_clk new_AGEMA_reg_buffer_4486 ( .C (clk), .D (new_AGEMA_signal_7950), .Q (new_AGEMA_signal_7951) ) ;
    buf_clk new_AGEMA_reg_buffer_4494 ( .C (clk), .D (new_AGEMA_signal_7958), .Q (new_AGEMA_signal_7959) ) ;
    buf_clk new_AGEMA_reg_buffer_4502 ( .C (clk), .D (new_AGEMA_signal_7966), .Q (new_AGEMA_signal_7967) ) ;
    buf_clk new_AGEMA_reg_buffer_4510 ( .C (clk), .D (new_AGEMA_signal_7974), .Q (new_AGEMA_signal_7975) ) ;
    buf_clk new_AGEMA_reg_buffer_4518 ( .C (clk), .D (new_AGEMA_signal_7982), .Q (new_AGEMA_signal_7983) ) ;
    buf_clk new_AGEMA_reg_buffer_4526 ( .C (clk), .D (new_AGEMA_signal_7990), .Q (new_AGEMA_signal_7991) ) ;
    buf_clk new_AGEMA_reg_buffer_4534 ( .C (clk), .D (new_AGEMA_signal_7998), .Q (new_AGEMA_signal_7999) ) ;
    buf_clk new_AGEMA_reg_buffer_4542 ( .C (clk), .D (new_AGEMA_signal_8006), .Q (new_AGEMA_signal_8007) ) ;
    buf_clk new_AGEMA_reg_buffer_4550 ( .C (clk), .D (new_AGEMA_signal_8014), .Q (new_AGEMA_signal_8015) ) ;
    buf_clk new_AGEMA_reg_buffer_4558 ( .C (clk), .D (new_AGEMA_signal_8022), .Q (new_AGEMA_signal_8023) ) ;
    buf_clk new_AGEMA_reg_buffer_4566 ( .C (clk), .D (new_AGEMA_signal_8030), .Q (new_AGEMA_signal_8031) ) ;
    buf_clk new_AGEMA_reg_buffer_4574 ( .C (clk), .D (new_AGEMA_signal_8038), .Q (new_AGEMA_signal_8039) ) ;
    buf_clk new_AGEMA_reg_buffer_4582 ( .C (clk), .D (new_AGEMA_signal_8046), .Q (new_AGEMA_signal_8047) ) ;
    buf_clk new_AGEMA_reg_buffer_4590 ( .C (clk), .D (new_AGEMA_signal_8054), .Q (new_AGEMA_signal_8055) ) ;
    buf_clk new_AGEMA_reg_buffer_4598 ( .C (clk), .D (new_AGEMA_signal_8062), .Q (new_AGEMA_signal_8063) ) ;
    buf_clk new_AGEMA_reg_buffer_4606 ( .C (clk), .D (new_AGEMA_signal_8070), .Q (new_AGEMA_signal_8071) ) ;
    buf_clk new_AGEMA_reg_buffer_4614 ( .C (clk), .D (new_AGEMA_signal_8078), .Q (new_AGEMA_signal_8079) ) ;
    buf_clk new_AGEMA_reg_buffer_4622 ( .C (clk), .D (new_AGEMA_signal_8086), .Q (new_AGEMA_signal_8087) ) ;
    buf_clk new_AGEMA_reg_buffer_4630 ( .C (clk), .D (new_AGEMA_signal_8094), .Q (new_AGEMA_signal_8095) ) ;
    buf_clk new_AGEMA_reg_buffer_4638 ( .C (clk), .D (new_AGEMA_signal_8102), .Q (new_AGEMA_signal_8103) ) ;
    buf_clk new_AGEMA_reg_buffer_4646 ( .C (clk), .D (new_AGEMA_signal_8110), .Q (new_AGEMA_signal_8111) ) ;
    buf_clk new_AGEMA_reg_buffer_4654 ( .C (clk), .D (new_AGEMA_signal_8118), .Q (new_AGEMA_signal_8119) ) ;
    buf_clk new_AGEMA_reg_buffer_4662 ( .C (clk), .D (new_AGEMA_signal_8126), .Q (new_AGEMA_signal_8127) ) ;
    buf_clk new_AGEMA_reg_buffer_4670 ( .C (clk), .D (new_AGEMA_signal_8134), .Q (new_AGEMA_signal_8135) ) ;
    buf_clk new_AGEMA_reg_buffer_4678 ( .C (clk), .D (new_AGEMA_signal_8142), .Q (new_AGEMA_signal_8143) ) ;
    buf_clk new_AGEMA_reg_buffer_4686 ( .C (clk), .D (new_AGEMA_signal_8150), .Q (new_AGEMA_signal_8151) ) ;
    buf_clk new_AGEMA_reg_buffer_4694 ( .C (clk), .D (new_AGEMA_signal_8158), .Q (new_AGEMA_signal_8159) ) ;
    buf_clk new_AGEMA_reg_buffer_4702 ( .C (clk), .D (new_AGEMA_signal_8166), .Q (new_AGEMA_signal_8167) ) ;
    buf_clk new_AGEMA_reg_buffer_4710 ( .C (clk), .D (new_AGEMA_signal_8174), .Q (new_AGEMA_signal_8175) ) ;
    buf_clk new_AGEMA_reg_buffer_4718 ( .C (clk), .D (new_AGEMA_signal_8182), .Q (new_AGEMA_signal_8183) ) ;
    buf_clk new_AGEMA_reg_buffer_4726 ( .C (clk), .D (new_AGEMA_signal_8190), .Q (new_AGEMA_signal_8191) ) ;
    buf_clk new_AGEMA_reg_buffer_4734 ( .C (clk), .D (new_AGEMA_signal_8198), .Q (new_AGEMA_signal_8199) ) ;
    buf_clk new_AGEMA_reg_buffer_4742 ( .C (clk), .D (new_AGEMA_signal_8206), .Q (new_AGEMA_signal_8207) ) ;
    buf_clk new_AGEMA_reg_buffer_4750 ( .C (clk), .D (new_AGEMA_signal_8214), .Q (new_AGEMA_signal_8215) ) ;
    buf_clk new_AGEMA_reg_buffer_4758 ( .C (clk), .D (new_AGEMA_signal_8222), .Q (new_AGEMA_signal_8223) ) ;
    buf_clk new_AGEMA_reg_buffer_4766 ( .C (clk), .D (new_AGEMA_signal_8230), .Q (new_AGEMA_signal_8231) ) ;
    buf_clk new_AGEMA_reg_buffer_4774 ( .C (clk), .D (new_AGEMA_signal_8238), .Q (new_AGEMA_signal_8239) ) ;
    buf_clk new_AGEMA_reg_buffer_4782 ( .C (clk), .D (new_AGEMA_signal_8246), .Q (new_AGEMA_signal_8247) ) ;
    buf_clk new_AGEMA_reg_buffer_4790 ( .C (clk), .D (new_AGEMA_signal_8254), .Q (new_AGEMA_signal_8255) ) ;
    buf_clk new_AGEMA_reg_buffer_4798 ( .C (clk), .D (new_AGEMA_signal_8262), .Q (new_AGEMA_signal_8263) ) ;
    buf_clk new_AGEMA_reg_buffer_4806 ( .C (clk), .D (new_AGEMA_signal_8270), .Q (new_AGEMA_signal_8271) ) ;
    buf_clk new_AGEMA_reg_buffer_4814 ( .C (clk), .D (new_AGEMA_signal_8278), .Q (new_AGEMA_signal_8279) ) ;
    buf_clk new_AGEMA_reg_buffer_4822 ( .C (clk), .D (new_AGEMA_signal_8286), .Q (new_AGEMA_signal_8287) ) ;
    buf_clk new_AGEMA_reg_buffer_4830 ( .C (clk), .D (new_AGEMA_signal_8294), .Q (new_AGEMA_signal_8295) ) ;
    buf_clk new_AGEMA_reg_buffer_4838 ( .C (clk), .D (new_AGEMA_signal_8302), .Q (new_AGEMA_signal_8303) ) ;
    buf_clk new_AGEMA_reg_buffer_4846 ( .C (clk), .D (new_AGEMA_signal_8310), .Q (new_AGEMA_signal_8311) ) ;
    buf_clk new_AGEMA_reg_buffer_4854 ( .C (clk), .D (new_AGEMA_signal_8318), .Q (new_AGEMA_signal_8319) ) ;
    buf_clk new_AGEMA_reg_buffer_4862 ( .C (clk), .D (new_AGEMA_signal_8326), .Q (new_AGEMA_signal_8327) ) ;
    buf_clk new_AGEMA_reg_buffer_4870 ( .C (clk), .D (new_AGEMA_signal_8334), .Q (new_AGEMA_signal_8335) ) ;
    buf_clk new_AGEMA_reg_buffer_4878 ( .C (clk), .D (new_AGEMA_signal_8342), .Q (new_AGEMA_signal_8343) ) ;
    buf_clk new_AGEMA_reg_buffer_4886 ( .C (clk), .D (new_AGEMA_signal_8350), .Q (new_AGEMA_signal_8351) ) ;
    buf_clk new_AGEMA_reg_buffer_4894 ( .C (clk), .D (new_AGEMA_signal_8358), .Q (new_AGEMA_signal_8359) ) ;
    buf_clk new_AGEMA_reg_buffer_4902 ( .C (clk), .D (new_AGEMA_signal_8366), .Q (new_AGEMA_signal_8367) ) ;
    buf_clk new_AGEMA_reg_buffer_4910 ( .C (clk), .D (new_AGEMA_signal_8374), .Q (new_AGEMA_signal_8375) ) ;
    buf_clk new_AGEMA_reg_buffer_4918 ( .C (clk), .D (new_AGEMA_signal_8382), .Q (new_AGEMA_signal_8383) ) ;
    buf_clk new_AGEMA_reg_buffer_4926 ( .C (clk), .D (new_AGEMA_signal_8390), .Q (new_AGEMA_signal_8391) ) ;
    buf_clk new_AGEMA_reg_buffer_4934 ( .C (clk), .D (new_AGEMA_signal_8398), .Q (new_AGEMA_signal_8399) ) ;
    buf_clk new_AGEMA_reg_buffer_4942 ( .C (clk), .D (new_AGEMA_signal_8406), .Q (new_AGEMA_signal_8407) ) ;
    buf_clk new_AGEMA_reg_buffer_4950 ( .C (clk), .D (new_AGEMA_signal_8414), .Q (new_AGEMA_signal_8415) ) ;
    buf_clk new_AGEMA_reg_buffer_4958 ( .C (clk), .D (new_AGEMA_signal_8422), .Q (new_AGEMA_signal_8423) ) ;
    buf_clk new_AGEMA_reg_buffer_4966 ( .C (clk), .D (new_AGEMA_signal_8430), .Q (new_AGEMA_signal_8431) ) ;
    buf_clk new_AGEMA_reg_buffer_4974 ( .C (clk), .D (new_AGEMA_signal_8438), .Q (new_AGEMA_signal_8439) ) ;
    buf_clk new_AGEMA_reg_buffer_4982 ( .C (clk), .D (new_AGEMA_signal_8446), .Q (new_AGEMA_signal_8447) ) ;
    buf_clk new_AGEMA_reg_buffer_4990 ( .C (clk), .D (new_AGEMA_signal_8454), .Q (new_AGEMA_signal_8455) ) ;
    buf_clk new_AGEMA_reg_buffer_4998 ( .C (clk), .D (new_AGEMA_signal_8462), .Q (new_AGEMA_signal_8463) ) ;
    buf_clk new_AGEMA_reg_buffer_5006 ( .C (clk), .D (new_AGEMA_signal_8470), .Q (new_AGEMA_signal_8471) ) ;
    buf_clk new_AGEMA_reg_buffer_5014 ( .C (clk), .D (new_AGEMA_signal_8478), .Q (new_AGEMA_signal_8479) ) ;
    buf_clk new_AGEMA_reg_buffer_5022 ( .C (clk), .D (new_AGEMA_signal_8486), .Q (new_AGEMA_signal_8487) ) ;
    buf_clk new_AGEMA_reg_buffer_5030 ( .C (clk), .D (new_AGEMA_signal_8494), .Q (new_AGEMA_signal_8495) ) ;
    buf_clk new_AGEMA_reg_buffer_5038 ( .C (clk), .D (new_AGEMA_signal_8502), .Q (new_AGEMA_signal_8503) ) ;
    buf_clk new_AGEMA_reg_buffer_5046 ( .C (clk), .D (new_AGEMA_signal_8510), .Q (new_AGEMA_signal_8511) ) ;
    buf_clk new_AGEMA_reg_buffer_5054 ( .C (clk), .D (new_AGEMA_signal_8518), .Q (new_AGEMA_signal_8519) ) ;
    buf_clk new_AGEMA_reg_buffer_5062 ( .C (clk), .D (new_AGEMA_signal_8526), .Q (new_AGEMA_signal_8527) ) ;
    buf_clk new_AGEMA_reg_buffer_5070 ( .C (clk), .D (new_AGEMA_signal_8534), .Q (new_AGEMA_signal_8535) ) ;
    buf_clk new_AGEMA_reg_buffer_5078 ( .C (clk), .D (new_AGEMA_signal_8542), .Q (new_AGEMA_signal_8543) ) ;
    buf_clk new_AGEMA_reg_buffer_5086 ( .C (clk), .D (new_AGEMA_signal_8550), .Q (new_AGEMA_signal_8551) ) ;
    buf_clk new_AGEMA_reg_buffer_5094 ( .C (clk), .D (new_AGEMA_signal_8558), .Q (new_AGEMA_signal_8559) ) ;
    buf_clk new_AGEMA_reg_buffer_5102 ( .C (clk), .D (new_AGEMA_signal_8566), .Q (new_AGEMA_signal_8567) ) ;
    buf_clk new_AGEMA_reg_buffer_5110 ( .C (clk), .D (new_AGEMA_signal_8574), .Q (new_AGEMA_signal_8575) ) ;
    buf_clk new_AGEMA_reg_buffer_5118 ( .C (clk), .D (new_AGEMA_signal_8582), .Q (new_AGEMA_signal_8583) ) ;
    buf_clk new_AGEMA_reg_buffer_5126 ( .C (clk), .D (new_AGEMA_signal_8590), .Q (new_AGEMA_signal_8591) ) ;
    buf_clk new_AGEMA_reg_buffer_5134 ( .C (clk), .D (new_AGEMA_signal_8598), .Q (new_AGEMA_signal_8599) ) ;
    buf_clk new_AGEMA_reg_buffer_5142 ( .C (clk), .D (new_AGEMA_signal_8606), .Q (new_AGEMA_signal_8607) ) ;
    buf_clk new_AGEMA_reg_buffer_5150 ( .C (clk), .D (new_AGEMA_signal_8614), .Q (new_AGEMA_signal_8615) ) ;
    buf_clk new_AGEMA_reg_buffer_5158 ( .C (clk), .D (new_AGEMA_signal_8622), .Q (new_AGEMA_signal_8623) ) ;
    buf_clk new_AGEMA_reg_buffer_5166 ( .C (clk), .D (new_AGEMA_signal_8630), .Q (new_AGEMA_signal_8631) ) ;
    buf_clk new_AGEMA_reg_buffer_5174 ( .C (clk), .D (new_AGEMA_signal_8638), .Q (new_AGEMA_signal_8639) ) ;
    buf_clk new_AGEMA_reg_buffer_5182 ( .C (clk), .D (new_AGEMA_signal_8646), .Q (new_AGEMA_signal_8647) ) ;
    buf_clk new_AGEMA_reg_buffer_5190 ( .C (clk), .D (new_AGEMA_signal_8654), .Q (new_AGEMA_signal_8655) ) ;
    buf_clk new_AGEMA_reg_buffer_5198 ( .C (clk), .D (new_AGEMA_signal_8662), .Q (new_AGEMA_signal_8663) ) ;
    buf_clk new_AGEMA_reg_buffer_5206 ( .C (clk), .D (new_AGEMA_signal_8670), .Q (new_AGEMA_signal_8671) ) ;
    buf_clk new_AGEMA_reg_buffer_5214 ( .C (clk), .D (new_AGEMA_signal_8678), .Q (new_AGEMA_signal_8679) ) ;
    buf_clk new_AGEMA_reg_buffer_5222 ( .C (clk), .D (new_AGEMA_signal_8686), .Q (new_AGEMA_signal_8687) ) ;
    buf_clk new_AGEMA_reg_buffer_5230 ( .C (clk), .D (new_AGEMA_signal_8694), .Q (new_AGEMA_signal_8695) ) ;
    buf_clk new_AGEMA_reg_buffer_5238 ( .C (clk), .D (new_AGEMA_signal_8702), .Q (new_AGEMA_signal_8703) ) ;
    buf_clk new_AGEMA_reg_buffer_5246 ( .C (clk), .D (new_AGEMA_signal_8710), .Q (new_AGEMA_signal_8711) ) ;
    buf_clk new_AGEMA_reg_buffer_5254 ( .C (clk), .D (new_AGEMA_signal_8718), .Q (new_AGEMA_signal_8719) ) ;
    buf_clk new_AGEMA_reg_buffer_5262 ( .C (clk), .D (new_AGEMA_signal_8726), .Q (new_AGEMA_signal_8727) ) ;
    buf_clk new_AGEMA_reg_buffer_5270 ( .C (clk), .D (new_AGEMA_signal_8734), .Q (new_AGEMA_signal_8735) ) ;
    buf_clk new_AGEMA_reg_buffer_5278 ( .C (clk), .D (new_AGEMA_signal_8742), .Q (new_AGEMA_signal_8743) ) ;
    buf_clk new_AGEMA_reg_buffer_5286 ( .C (clk), .D (new_AGEMA_signal_8750), .Q (new_AGEMA_signal_8751) ) ;
    buf_clk new_AGEMA_reg_buffer_5294 ( .C (clk), .D (new_AGEMA_signal_8758), .Q (new_AGEMA_signal_8759) ) ;
    buf_clk new_AGEMA_reg_buffer_5302 ( .C (clk), .D (new_AGEMA_signal_8766), .Q (new_AGEMA_signal_8767) ) ;
    buf_clk new_AGEMA_reg_buffer_5310 ( .C (clk), .D (new_AGEMA_signal_8774), .Q (new_AGEMA_signal_8775) ) ;
    buf_clk new_AGEMA_reg_buffer_5318 ( .C (clk), .D (new_AGEMA_signal_8782), .Q (new_AGEMA_signal_8783) ) ;
    buf_clk new_AGEMA_reg_buffer_5326 ( .C (clk), .D (new_AGEMA_signal_8790), .Q (new_AGEMA_signal_8791) ) ;
    buf_clk new_AGEMA_reg_buffer_5334 ( .C (clk), .D (new_AGEMA_signal_8798), .Q (new_AGEMA_signal_8799) ) ;
    buf_clk new_AGEMA_reg_buffer_5342 ( .C (clk), .D (new_AGEMA_signal_8806), .Q (new_AGEMA_signal_8807) ) ;
    buf_clk new_AGEMA_reg_buffer_5350 ( .C (clk), .D (new_AGEMA_signal_8814), .Q (new_AGEMA_signal_8815) ) ;
    buf_clk new_AGEMA_reg_buffer_5358 ( .C (clk), .D (new_AGEMA_signal_8822), .Q (new_AGEMA_signal_8823) ) ;
    buf_clk new_AGEMA_reg_buffer_5366 ( .C (clk), .D (new_AGEMA_signal_8830), .Q (new_AGEMA_signal_8831) ) ;
    buf_clk new_AGEMA_reg_buffer_5374 ( .C (clk), .D (new_AGEMA_signal_8838), .Q (new_AGEMA_signal_8839) ) ;
    buf_clk new_AGEMA_reg_buffer_5382 ( .C (clk), .D (new_AGEMA_signal_8846), .Q (new_AGEMA_signal_8847) ) ;
    buf_clk new_AGEMA_reg_buffer_5390 ( .C (clk), .D (new_AGEMA_signal_8854), .Q (new_AGEMA_signal_8855) ) ;
    buf_clk new_AGEMA_reg_buffer_5398 ( .C (clk), .D (new_AGEMA_signal_8862), .Q (new_AGEMA_signal_8863) ) ;
    buf_clk new_AGEMA_reg_buffer_5408 ( .C (clk), .D (new_AGEMA_signal_8872), .Q (new_AGEMA_signal_8873) ) ;
    buf_clk new_AGEMA_reg_buffer_5416 ( .C (clk), .D (new_AGEMA_signal_8880), .Q (new_AGEMA_signal_8881) ) ;
    buf_clk new_AGEMA_reg_buffer_5424 ( .C (clk), .D (new_AGEMA_signal_8888), .Q (new_AGEMA_signal_8889) ) ;
    buf_clk new_AGEMA_reg_buffer_5432 ( .C (clk), .D (new_AGEMA_signal_8896), .Q (new_AGEMA_signal_8897) ) ;
    buf_clk new_AGEMA_reg_buffer_5440 ( .C (clk), .D (new_AGEMA_signal_8904), .Q (new_AGEMA_signal_8905) ) ;
    buf_clk new_AGEMA_reg_buffer_5448 ( .C (clk), .D (new_AGEMA_signal_8912), .Q (new_AGEMA_signal_8913) ) ;
    buf_clk new_AGEMA_reg_buffer_5456 ( .C (clk), .D (new_AGEMA_signal_8920), .Q (new_AGEMA_signal_8921) ) ;
    buf_clk new_AGEMA_reg_buffer_5464 ( .C (clk), .D (new_AGEMA_signal_8928), .Q (new_AGEMA_signal_8929) ) ;
    buf_clk new_AGEMA_reg_buffer_5472 ( .C (clk), .D (new_AGEMA_signal_8936), .Q (new_AGEMA_signal_8937) ) ;
    buf_clk new_AGEMA_reg_buffer_5480 ( .C (clk), .D (new_AGEMA_signal_8944), .Q (new_AGEMA_signal_8945) ) ;
    buf_clk new_AGEMA_reg_buffer_5488 ( .C (clk), .D (new_AGEMA_signal_8952), .Q (new_AGEMA_signal_8953) ) ;
    buf_clk new_AGEMA_reg_buffer_5496 ( .C (clk), .D (new_AGEMA_signal_8960), .Q (new_AGEMA_signal_8961) ) ;
    buf_clk new_AGEMA_reg_buffer_5504 ( .C (clk), .D (new_AGEMA_signal_8968), .Q (new_AGEMA_signal_8969) ) ;
    buf_clk new_AGEMA_reg_buffer_5512 ( .C (clk), .D (new_AGEMA_signal_8976), .Q (new_AGEMA_signal_8977) ) ;
    buf_clk new_AGEMA_reg_buffer_5520 ( .C (clk), .D (new_AGEMA_signal_8984), .Q (new_AGEMA_signal_8985) ) ;
    buf_clk new_AGEMA_reg_buffer_5528 ( .C (clk), .D (new_AGEMA_signal_8992), .Q (new_AGEMA_signal_8993) ) ;
    buf_clk new_AGEMA_reg_buffer_5536 ( .C (clk), .D (new_AGEMA_signal_9000), .Q (new_AGEMA_signal_9001) ) ;
    buf_clk new_AGEMA_reg_buffer_5544 ( .C (clk), .D (new_AGEMA_signal_9008), .Q (new_AGEMA_signal_9009) ) ;
    buf_clk new_AGEMA_reg_buffer_5552 ( .C (clk), .D (new_AGEMA_signal_9016), .Q (new_AGEMA_signal_9017) ) ;
    buf_clk new_AGEMA_reg_buffer_5560 ( .C (clk), .D (new_AGEMA_signal_9024), .Q (new_AGEMA_signal_9025) ) ;
    buf_clk new_AGEMA_reg_buffer_5568 ( .C (clk), .D (new_AGEMA_signal_9032), .Q (new_AGEMA_signal_9033) ) ;
    buf_clk new_AGEMA_reg_buffer_5576 ( .C (clk), .D (new_AGEMA_signal_9040), .Q (new_AGEMA_signal_9041) ) ;
    buf_clk new_AGEMA_reg_buffer_5584 ( .C (clk), .D (new_AGEMA_signal_9048), .Q (new_AGEMA_signal_9049) ) ;
    buf_clk new_AGEMA_reg_buffer_5592 ( .C (clk), .D (new_AGEMA_signal_9056), .Q (new_AGEMA_signal_9057) ) ;
    buf_clk new_AGEMA_reg_buffer_5600 ( .C (clk), .D (new_AGEMA_signal_9064), .Q (new_AGEMA_signal_9065) ) ;
    buf_clk new_AGEMA_reg_buffer_5608 ( .C (clk), .D (new_AGEMA_signal_9072), .Q (new_AGEMA_signal_9073) ) ;
    buf_clk new_AGEMA_reg_buffer_5616 ( .C (clk), .D (new_AGEMA_signal_9080), .Q (new_AGEMA_signal_9081) ) ;
    buf_clk new_AGEMA_reg_buffer_5624 ( .C (clk), .D (new_AGEMA_signal_9088), .Q (new_AGEMA_signal_9089) ) ;
    buf_clk new_AGEMA_reg_buffer_5632 ( .C (clk), .D (new_AGEMA_signal_9096), .Q (new_AGEMA_signal_9097) ) ;
    buf_clk new_AGEMA_reg_buffer_5640 ( .C (clk), .D (new_AGEMA_signal_9104), .Q (new_AGEMA_signal_9105) ) ;
    buf_clk new_AGEMA_reg_buffer_5648 ( .C (clk), .D (new_AGEMA_signal_9112), .Q (new_AGEMA_signal_9113) ) ;
    buf_clk new_AGEMA_reg_buffer_5656 ( .C (clk), .D (new_AGEMA_signal_9120), .Q (new_AGEMA_signal_9121) ) ;
    buf_clk new_AGEMA_reg_buffer_5664 ( .C (clk), .D (new_AGEMA_signal_9128), .Q (new_AGEMA_signal_9129) ) ;
    buf_clk new_AGEMA_reg_buffer_5672 ( .C (clk), .D (new_AGEMA_signal_9136), .Q (new_AGEMA_signal_9137) ) ;
    buf_clk new_AGEMA_reg_buffer_5680 ( .C (clk), .D (new_AGEMA_signal_9144), .Q (new_AGEMA_signal_9145) ) ;
    buf_clk new_AGEMA_reg_buffer_5688 ( .C (clk), .D (new_AGEMA_signal_9152), .Q (new_AGEMA_signal_9153) ) ;
    buf_clk new_AGEMA_reg_buffer_5696 ( .C (clk), .D (new_AGEMA_signal_9160), .Q (new_AGEMA_signal_9161) ) ;
    buf_clk new_AGEMA_reg_buffer_5704 ( .C (clk), .D (new_AGEMA_signal_9168), .Q (new_AGEMA_signal_9169) ) ;
    buf_clk new_AGEMA_reg_buffer_5712 ( .C (clk), .D (new_AGEMA_signal_9176), .Q (new_AGEMA_signal_9177) ) ;
    buf_clk new_AGEMA_reg_buffer_5720 ( .C (clk), .D (new_AGEMA_signal_9184), .Q (new_AGEMA_signal_9185) ) ;
    buf_clk new_AGEMA_reg_buffer_5728 ( .C (clk), .D (new_AGEMA_signal_9192), .Q (new_AGEMA_signal_9193) ) ;
    buf_clk new_AGEMA_reg_buffer_5736 ( .C (clk), .D (new_AGEMA_signal_9200), .Q (new_AGEMA_signal_9201) ) ;
    buf_clk new_AGEMA_reg_buffer_5744 ( .C (clk), .D (new_AGEMA_signal_9208), .Q (new_AGEMA_signal_9209) ) ;
    buf_clk new_AGEMA_reg_buffer_5752 ( .C (clk), .D (new_AGEMA_signal_9216), .Q (new_AGEMA_signal_9217) ) ;
    buf_clk new_AGEMA_reg_buffer_5760 ( .C (clk), .D (new_AGEMA_signal_9224), .Q (new_AGEMA_signal_9225) ) ;
    buf_clk new_AGEMA_reg_buffer_5768 ( .C (clk), .D (new_AGEMA_signal_9232), .Q (new_AGEMA_signal_9233) ) ;
    buf_clk new_AGEMA_reg_buffer_5776 ( .C (clk), .D (new_AGEMA_signal_9240), .Q (new_AGEMA_signal_9241) ) ;
    buf_clk new_AGEMA_reg_buffer_5784 ( .C (clk), .D (new_AGEMA_signal_9248), .Q (new_AGEMA_signal_9249) ) ;
    buf_clk new_AGEMA_reg_buffer_5792 ( .C (clk), .D (new_AGEMA_signal_9256), .Q (new_AGEMA_signal_9257) ) ;
    buf_clk new_AGEMA_reg_buffer_5800 ( .C (clk), .D (new_AGEMA_signal_9264), .Q (new_AGEMA_signal_9265) ) ;
    buf_clk new_AGEMA_reg_buffer_5808 ( .C (clk), .D (new_AGEMA_signal_9272), .Q (new_AGEMA_signal_9273) ) ;
    buf_clk new_AGEMA_reg_buffer_5816 ( .C (clk), .D (new_AGEMA_signal_9280), .Q (new_AGEMA_signal_9281) ) ;
    buf_clk new_AGEMA_reg_buffer_5824 ( .C (clk), .D (new_AGEMA_signal_9288), .Q (new_AGEMA_signal_9289) ) ;
    buf_clk new_AGEMA_reg_buffer_5832 ( .C (clk), .D (new_AGEMA_signal_9296), .Q (new_AGEMA_signal_9297) ) ;
    buf_clk new_AGEMA_reg_buffer_5840 ( .C (clk), .D (new_AGEMA_signal_9304), .Q (new_AGEMA_signal_9305) ) ;
    buf_clk new_AGEMA_reg_buffer_5848 ( .C (clk), .D (new_AGEMA_signal_9312), .Q (new_AGEMA_signal_9313) ) ;
    buf_clk new_AGEMA_reg_buffer_5856 ( .C (clk), .D (new_AGEMA_signal_9320), .Q (new_AGEMA_signal_9321) ) ;
    buf_clk new_AGEMA_reg_buffer_5864 ( .C (clk), .D (new_AGEMA_signal_9328), .Q (new_AGEMA_signal_9329) ) ;
    buf_clk new_AGEMA_reg_buffer_5872 ( .C (clk), .D (new_AGEMA_signal_9336), .Q (new_AGEMA_signal_9337) ) ;
    buf_clk new_AGEMA_reg_buffer_5880 ( .C (clk), .D (new_AGEMA_signal_9344), .Q (new_AGEMA_signal_9345) ) ;
    buf_clk new_AGEMA_reg_buffer_5888 ( .C (clk), .D (new_AGEMA_signal_9352), .Q (new_AGEMA_signal_9353) ) ;
    buf_clk new_AGEMA_reg_buffer_5896 ( .C (clk), .D (new_AGEMA_signal_9360), .Q (new_AGEMA_signal_9361) ) ;
    buf_clk new_AGEMA_reg_buffer_5904 ( .C (clk), .D (new_AGEMA_signal_9368), .Q (new_AGEMA_signal_9369) ) ;
    buf_clk new_AGEMA_reg_buffer_5912 ( .C (clk), .D (new_AGEMA_signal_9376), .Q (new_AGEMA_signal_9377) ) ;
    buf_clk new_AGEMA_reg_buffer_5920 ( .C (clk), .D (new_AGEMA_signal_9384), .Q (new_AGEMA_signal_9385) ) ;
    buf_clk new_AGEMA_reg_buffer_5928 ( .C (clk), .D (new_AGEMA_signal_9392), .Q (new_AGEMA_signal_9393) ) ;
    buf_clk new_AGEMA_reg_buffer_5936 ( .C (clk), .D (new_AGEMA_signal_9400), .Q (new_AGEMA_signal_9401) ) ;
    buf_clk new_AGEMA_reg_buffer_5944 ( .C (clk), .D (new_AGEMA_signal_9408), .Q (new_AGEMA_signal_9409) ) ;
    buf_clk new_AGEMA_reg_buffer_5952 ( .C (clk), .D (new_AGEMA_signal_9416), .Q (new_AGEMA_signal_9417) ) ;
    buf_clk new_AGEMA_reg_buffer_5960 ( .C (clk), .D (new_AGEMA_signal_9424), .Q (new_AGEMA_signal_9425) ) ;
    buf_clk new_AGEMA_reg_buffer_5968 ( .C (clk), .D (new_AGEMA_signal_9432), .Q (new_AGEMA_signal_9433) ) ;
    buf_clk new_AGEMA_reg_buffer_5976 ( .C (clk), .D (new_AGEMA_signal_9440), .Q (new_AGEMA_signal_9441) ) ;
    buf_clk new_AGEMA_reg_buffer_5984 ( .C (clk), .D (new_AGEMA_signal_9448), .Q (new_AGEMA_signal_9449) ) ;
    buf_clk new_AGEMA_reg_buffer_5992 ( .C (clk), .D (new_AGEMA_signal_9456), .Q (new_AGEMA_signal_9457) ) ;
    buf_clk new_AGEMA_reg_buffer_6000 ( .C (clk), .D (new_AGEMA_signal_9464), .Q (new_AGEMA_signal_9465) ) ;
    buf_clk new_AGEMA_reg_buffer_6008 ( .C (clk), .D (new_AGEMA_signal_9472), .Q (new_AGEMA_signal_9473) ) ;
    buf_clk new_AGEMA_reg_buffer_6016 ( .C (clk), .D (new_AGEMA_signal_9480), .Q (new_AGEMA_signal_9481) ) ;
    buf_clk new_AGEMA_reg_buffer_6024 ( .C (clk), .D (new_AGEMA_signal_9488), .Q (new_AGEMA_signal_9489) ) ;
    buf_clk new_AGEMA_reg_buffer_6032 ( .C (clk), .D (new_AGEMA_signal_9496), .Q (new_AGEMA_signal_9497) ) ;
    buf_clk new_AGEMA_reg_buffer_6040 ( .C (clk), .D (new_AGEMA_signal_9504), .Q (new_AGEMA_signal_9505) ) ;
    buf_clk new_AGEMA_reg_buffer_6048 ( .C (clk), .D (new_AGEMA_signal_9512), .Q (new_AGEMA_signal_9513) ) ;
    buf_clk new_AGEMA_reg_buffer_6056 ( .C (clk), .D (new_AGEMA_signal_9520), .Q (new_AGEMA_signal_9521) ) ;
    buf_clk new_AGEMA_reg_buffer_6064 ( .C (clk), .D (new_AGEMA_signal_9528), .Q (new_AGEMA_signal_9529) ) ;
    buf_clk new_AGEMA_reg_buffer_6072 ( .C (clk), .D (new_AGEMA_signal_9536), .Q (new_AGEMA_signal_9537) ) ;
    buf_clk new_AGEMA_reg_buffer_6080 ( .C (clk), .D (new_AGEMA_signal_9544), .Q (new_AGEMA_signal_9545) ) ;
    buf_clk new_AGEMA_reg_buffer_6088 ( .C (clk), .D (new_AGEMA_signal_9552), .Q (new_AGEMA_signal_9553) ) ;
    buf_clk new_AGEMA_reg_buffer_6096 ( .C (clk), .D (new_AGEMA_signal_9560), .Q (new_AGEMA_signal_9561) ) ;
    buf_clk new_AGEMA_reg_buffer_6104 ( .C (clk), .D (new_AGEMA_signal_9568), .Q (new_AGEMA_signal_9569) ) ;
    buf_clk new_AGEMA_reg_buffer_6112 ( .C (clk), .D (new_AGEMA_signal_9576), .Q (new_AGEMA_signal_9577) ) ;
    buf_clk new_AGEMA_reg_buffer_6120 ( .C (clk), .D (new_AGEMA_signal_9584), .Q (new_AGEMA_signal_9585) ) ;
    buf_clk new_AGEMA_reg_buffer_6128 ( .C (clk), .D (new_AGEMA_signal_9592), .Q (new_AGEMA_signal_9593) ) ;
    buf_clk new_AGEMA_reg_buffer_6136 ( .C (clk), .D (new_AGEMA_signal_9600), .Q (new_AGEMA_signal_9601) ) ;
    buf_clk new_AGEMA_reg_buffer_6144 ( .C (clk), .D (new_AGEMA_signal_9608), .Q (new_AGEMA_signal_9609) ) ;
    buf_clk new_AGEMA_reg_buffer_6152 ( .C (clk), .D (new_AGEMA_signal_9616), .Q (new_AGEMA_signal_9617) ) ;
    buf_clk new_AGEMA_reg_buffer_6160 ( .C (clk), .D (new_AGEMA_signal_9624), .Q (new_AGEMA_signal_9625) ) ;
    buf_clk new_AGEMA_reg_buffer_6168 ( .C (clk), .D (new_AGEMA_signal_9632), .Q (new_AGEMA_signal_9633) ) ;
    buf_clk new_AGEMA_reg_buffer_6180 ( .C (clk), .D (new_AGEMA_signal_9644), .Q (new_AGEMA_signal_9645) ) ;
    buf_clk new_AGEMA_reg_buffer_6184 ( .C (clk), .D (new_AGEMA_signal_9648), .Q (new_AGEMA_signal_9649) ) ;
    buf_clk new_AGEMA_reg_buffer_6188 ( .C (clk), .D (new_AGEMA_signal_9652), .Q (new_AGEMA_signal_9653) ) ;
    buf_clk new_AGEMA_reg_buffer_6198 ( .C (clk), .D (new_AGEMA_signal_9662), .Q (new_AGEMA_signal_9663) ) ;
    buf_clk new_AGEMA_reg_buffer_6202 ( .C (clk), .D (new_AGEMA_signal_9666), .Q (new_AGEMA_signal_9667) ) ;
    buf_clk new_AGEMA_reg_buffer_6206 ( .C (clk), .D (new_AGEMA_signal_9670), .Q (new_AGEMA_signal_9671) ) ;
    buf_clk new_AGEMA_reg_buffer_6216 ( .C (clk), .D (new_AGEMA_signal_9680), .Q (new_AGEMA_signal_9681) ) ;
    buf_clk new_AGEMA_reg_buffer_6220 ( .C (clk), .D (new_AGEMA_signal_9684), .Q (new_AGEMA_signal_9685) ) ;
    buf_clk new_AGEMA_reg_buffer_6224 ( .C (clk), .D (new_AGEMA_signal_9688), .Q (new_AGEMA_signal_9689) ) ;
    buf_clk new_AGEMA_reg_buffer_6234 ( .C (clk), .D (new_AGEMA_signal_9698), .Q (new_AGEMA_signal_9699) ) ;
    buf_clk new_AGEMA_reg_buffer_6238 ( .C (clk), .D (new_AGEMA_signal_9702), .Q (new_AGEMA_signal_9703) ) ;
    buf_clk new_AGEMA_reg_buffer_6242 ( .C (clk), .D (new_AGEMA_signal_9706), .Q (new_AGEMA_signal_9707) ) ;
    buf_clk new_AGEMA_reg_buffer_6252 ( .C (clk), .D (new_AGEMA_signal_9716), .Q (new_AGEMA_signal_9717) ) ;
    buf_clk new_AGEMA_reg_buffer_6256 ( .C (clk), .D (new_AGEMA_signal_9720), .Q (new_AGEMA_signal_9721) ) ;
    buf_clk new_AGEMA_reg_buffer_6260 ( .C (clk), .D (new_AGEMA_signal_9724), .Q (new_AGEMA_signal_9725) ) ;
    buf_clk new_AGEMA_reg_buffer_6270 ( .C (clk), .D (new_AGEMA_signal_9734), .Q (new_AGEMA_signal_9735) ) ;
    buf_clk new_AGEMA_reg_buffer_6274 ( .C (clk), .D (new_AGEMA_signal_9738), .Q (new_AGEMA_signal_9739) ) ;
    buf_clk new_AGEMA_reg_buffer_6278 ( .C (clk), .D (new_AGEMA_signal_9742), .Q (new_AGEMA_signal_9743) ) ;
    buf_clk new_AGEMA_reg_buffer_6288 ( .C (clk), .D (new_AGEMA_signal_9752), .Q (new_AGEMA_signal_9753) ) ;
    buf_clk new_AGEMA_reg_buffer_6292 ( .C (clk), .D (new_AGEMA_signal_9756), .Q (new_AGEMA_signal_9757) ) ;
    buf_clk new_AGEMA_reg_buffer_6296 ( .C (clk), .D (new_AGEMA_signal_9760), .Q (new_AGEMA_signal_9761) ) ;
    buf_clk new_AGEMA_reg_buffer_6306 ( .C (clk), .D (new_AGEMA_signal_9770), .Q (new_AGEMA_signal_9771) ) ;
    buf_clk new_AGEMA_reg_buffer_6310 ( .C (clk), .D (new_AGEMA_signal_9774), .Q (new_AGEMA_signal_9775) ) ;
    buf_clk new_AGEMA_reg_buffer_6314 ( .C (clk), .D (new_AGEMA_signal_9778), .Q (new_AGEMA_signal_9779) ) ;
    buf_clk new_AGEMA_reg_buffer_6324 ( .C (clk), .D (new_AGEMA_signal_9788), .Q (new_AGEMA_signal_9789) ) ;
    buf_clk new_AGEMA_reg_buffer_6328 ( .C (clk), .D (new_AGEMA_signal_9792), .Q (new_AGEMA_signal_9793) ) ;
    buf_clk new_AGEMA_reg_buffer_6332 ( .C (clk), .D (new_AGEMA_signal_9796), .Q (new_AGEMA_signal_9797) ) ;
    buf_clk new_AGEMA_reg_buffer_6342 ( .C (clk), .D (new_AGEMA_signal_9806), .Q (new_AGEMA_signal_9807) ) ;
    buf_clk new_AGEMA_reg_buffer_6346 ( .C (clk), .D (new_AGEMA_signal_9810), .Q (new_AGEMA_signal_9811) ) ;
    buf_clk new_AGEMA_reg_buffer_6350 ( .C (clk), .D (new_AGEMA_signal_9814), .Q (new_AGEMA_signal_9815) ) ;
    buf_clk new_AGEMA_reg_buffer_6360 ( .C (clk), .D (new_AGEMA_signal_9824), .Q (new_AGEMA_signal_9825) ) ;
    buf_clk new_AGEMA_reg_buffer_6364 ( .C (clk), .D (new_AGEMA_signal_9828), .Q (new_AGEMA_signal_9829) ) ;
    buf_clk new_AGEMA_reg_buffer_6368 ( .C (clk), .D (new_AGEMA_signal_9832), .Q (new_AGEMA_signal_9833) ) ;
    buf_clk new_AGEMA_reg_buffer_6378 ( .C (clk), .D (new_AGEMA_signal_9842), .Q (new_AGEMA_signal_9843) ) ;
    buf_clk new_AGEMA_reg_buffer_6382 ( .C (clk), .D (new_AGEMA_signal_9846), .Q (new_AGEMA_signal_9847) ) ;
    buf_clk new_AGEMA_reg_buffer_6386 ( .C (clk), .D (new_AGEMA_signal_9850), .Q (new_AGEMA_signal_9851) ) ;
    buf_clk new_AGEMA_reg_buffer_6396 ( .C (clk), .D (new_AGEMA_signal_9860), .Q (new_AGEMA_signal_9861) ) ;
    buf_clk new_AGEMA_reg_buffer_6400 ( .C (clk), .D (new_AGEMA_signal_9864), .Q (new_AGEMA_signal_9865) ) ;
    buf_clk new_AGEMA_reg_buffer_6404 ( .C (clk), .D (new_AGEMA_signal_9868), .Q (new_AGEMA_signal_9869) ) ;
    buf_clk new_AGEMA_reg_buffer_6414 ( .C (clk), .D (new_AGEMA_signal_9878), .Q (new_AGEMA_signal_9879) ) ;
    buf_clk new_AGEMA_reg_buffer_6418 ( .C (clk), .D (new_AGEMA_signal_9882), .Q (new_AGEMA_signal_9883) ) ;
    buf_clk new_AGEMA_reg_buffer_6422 ( .C (clk), .D (new_AGEMA_signal_9886), .Q (new_AGEMA_signal_9887) ) ;
    buf_clk new_AGEMA_reg_buffer_6432 ( .C (clk), .D (new_AGEMA_signal_9896), .Q (new_AGEMA_signal_9897) ) ;
    buf_clk new_AGEMA_reg_buffer_6436 ( .C (clk), .D (new_AGEMA_signal_9900), .Q (new_AGEMA_signal_9901) ) ;
    buf_clk new_AGEMA_reg_buffer_6440 ( .C (clk), .D (new_AGEMA_signal_9904), .Q (new_AGEMA_signal_9905) ) ;
    buf_clk new_AGEMA_reg_buffer_6450 ( .C (clk), .D (new_AGEMA_signal_9914), .Q (new_AGEMA_signal_9915) ) ;
    buf_clk new_AGEMA_reg_buffer_6454 ( .C (clk), .D (new_AGEMA_signal_9918), .Q (new_AGEMA_signal_9919) ) ;
    buf_clk new_AGEMA_reg_buffer_6458 ( .C (clk), .D (new_AGEMA_signal_9922), .Q (new_AGEMA_signal_9923) ) ;
    buf_clk new_AGEMA_reg_buffer_6466 ( .C (clk), .D (new_AGEMA_signal_9930), .Q (new_AGEMA_signal_9931) ) ;
    buf_clk new_AGEMA_reg_buffer_6474 ( .C (clk), .D (new_AGEMA_signal_9938), .Q (new_AGEMA_signal_9939) ) ;
    buf_clk new_AGEMA_reg_buffer_6482 ( .C (clk), .D (new_AGEMA_signal_9946), .Q (new_AGEMA_signal_9947) ) ;
    buf_clk new_AGEMA_reg_buffer_6490 ( .C (clk), .D (new_AGEMA_signal_9954), .Q (new_AGEMA_signal_9955) ) ;

    /* cells in depth 5 */
    buf_clk new_AGEMA_reg_buffer_1323 ( .C (clk), .D (new_AGEMA_signal_4788), .Q (new_AGEMA_signal_4789) ) ;
    buf_clk new_AGEMA_reg_buffer_1843 ( .C (clk), .D (new_AGEMA_signal_5307), .Q (new_AGEMA_signal_5308) ) ;
    buf_clk new_AGEMA_reg_buffer_1849 ( .C (clk), .D (new_AGEMA_signal_5313), .Q (new_AGEMA_signal_5314) ) ;
    buf_clk new_AGEMA_reg_buffer_1855 ( .C (clk), .D (new_AGEMA_signal_5319), .Q (new_AGEMA_signal_5320) ) ;
    buf_clk new_AGEMA_reg_buffer_1861 ( .C (clk), .D (new_AGEMA_signal_5325), .Q (new_AGEMA_signal_5326) ) ;
    buf_clk new_AGEMA_reg_buffer_1867 ( .C (clk), .D (new_AGEMA_signal_5331), .Q (new_AGEMA_signal_5332) ) ;
    buf_clk new_AGEMA_reg_buffer_1873 ( .C (clk), .D (new_AGEMA_signal_5337), .Q (new_AGEMA_signal_5338) ) ;
    buf_clk new_AGEMA_reg_buffer_1879 ( .C (clk), .D (new_AGEMA_signal_5343), .Q (new_AGEMA_signal_5344) ) ;
    buf_clk new_AGEMA_reg_buffer_1885 ( .C (clk), .D (new_AGEMA_signal_5349), .Q (new_AGEMA_signal_5350) ) ;
    buf_clk new_AGEMA_reg_buffer_1891 ( .C (clk), .D (new_AGEMA_signal_5355), .Q (new_AGEMA_signal_5356) ) ;
    buf_clk new_AGEMA_reg_buffer_1897 ( .C (clk), .D (new_AGEMA_signal_5361), .Q (new_AGEMA_signal_5362) ) ;
    buf_clk new_AGEMA_reg_buffer_1903 ( .C (clk), .D (new_AGEMA_signal_5367), .Q (new_AGEMA_signal_5368) ) ;
    buf_clk new_AGEMA_reg_buffer_1909 ( .C (clk), .D (new_AGEMA_signal_5373), .Q (new_AGEMA_signal_5374) ) ;
    buf_clk new_AGEMA_reg_buffer_1915 ( .C (clk), .D (new_AGEMA_signal_5379), .Q (new_AGEMA_signal_5380) ) ;
    buf_clk new_AGEMA_reg_buffer_1921 ( .C (clk), .D (new_AGEMA_signal_5385), .Q (new_AGEMA_signal_5386) ) ;
    buf_clk new_AGEMA_reg_buffer_1927 ( .C (clk), .D (new_AGEMA_signal_5391), .Q (new_AGEMA_signal_5392) ) ;
    buf_clk new_AGEMA_reg_buffer_1933 ( .C (clk), .D (new_AGEMA_signal_5397), .Q (new_AGEMA_signal_5398) ) ;
    buf_clk new_AGEMA_reg_buffer_1939 ( .C (clk), .D (new_AGEMA_signal_5403), .Q (new_AGEMA_signal_5404) ) ;
    buf_clk new_AGEMA_reg_buffer_1945 ( .C (clk), .D (new_AGEMA_signal_5409), .Q (new_AGEMA_signal_5410) ) ;
    buf_clk new_AGEMA_reg_buffer_1951 ( .C (clk), .D (new_AGEMA_signal_5415), .Q (new_AGEMA_signal_5416) ) ;
    buf_clk new_AGEMA_reg_buffer_1957 ( .C (clk), .D (new_AGEMA_signal_5421), .Q (new_AGEMA_signal_5422) ) ;
    buf_clk new_AGEMA_reg_buffer_1963 ( .C (clk), .D (new_AGEMA_signal_5427), .Q (new_AGEMA_signal_5428) ) ;
    buf_clk new_AGEMA_reg_buffer_1969 ( .C (clk), .D (new_AGEMA_signal_5433), .Q (new_AGEMA_signal_5434) ) ;
    buf_clk new_AGEMA_reg_buffer_1975 ( .C (clk), .D (new_AGEMA_signal_5439), .Q (new_AGEMA_signal_5440) ) ;
    buf_clk new_AGEMA_reg_buffer_1981 ( .C (clk), .D (new_AGEMA_signal_5445), .Q (new_AGEMA_signal_5446) ) ;
    buf_clk new_AGEMA_reg_buffer_1987 ( .C (clk), .D (new_AGEMA_signal_5451), .Q (new_AGEMA_signal_5452) ) ;
    buf_clk new_AGEMA_reg_buffer_1993 ( .C (clk), .D (new_AGEMA_signal_5457), .Q (new_AGEMA_signal_5458) ) ;
    buf_clk new_AGEMA_reg_buffer_1999 ( .C (clk), .D (new_AGEMA_signal_5463), .Q (new_AGEMA_signal_5464) ) ;
    buf_clk new_AGEMA_reg_buffer_2005 ( .C (clk), .D (new_AGEMA_signal_5469), .Q (new_AGEMA_signal_5470) ) ;
    buf_clk new_AGEMA_reg_buffer_2011 ( .C (clk), .D (new_AGEMA_signal_5475), .Q (new_AGEMA_signal_5476) ) ;
    buf_clk new_AGEMA_reg_buffer_2017 ( .C (clk), .D (new_AGEMA_signal_5481), .Q (new_AGEMA_signal_5482) ) ;
    buf_clk new_AGEMA_reg_buffer_2023 ( .C (clk), .D (new_AGEMA_signal_5487), .Q (new_AGEMA_signal_5488) ) ;
    buf_clk new_AGEMA_reg_buffer_2029 ( .C (clk), .D (new_AGEMA_signal_5493), .Q (new_AGEMA_signal_5494) ) ;
    buf_clk new_AGEMA_reg_buffer_2035 ( .C (clk), .D (new_AGEMA_signal_5499), .Q (new_AGEMA_signal_5500) ) ;
    buf_clk new_AGEMA_reg_buffer_2041 ( .C (clk), .D (new_AGEMA_signal_5505), .Q (new_AGEMA_signal_5506) ) ;
    buf_clk new_AGEMA_reg_buffer_2047 ( .C (clk), .D (new_AGEMA_signal_5511), .Q (new_AGEMA_signal_5512) ) ;
    buf_clk new_AGEMA_reg_buffer_2053 ( .C (clk), .D (new_AGEMA_signal_5517), .Q (new_AGEMA_signal_5518) ) ;
    buf_clk new_AGEMA_reg_buffer_2059 ( .C (clk), .D (new_AGEMA_signal_5523), .Q (new_AGEMA_signal_5524) ) ;
    buf_clk new_AGEMA_reg_buffer_2065 ( .C (clk), .D (new_AGEMA_signal_5529), .Q (new_AGEMA_signal_5530) ) ;
    buf_clk new_AGEMA_reg_buffer_2071 ( .C (clk), .D (new_AGEMA_signal_5535), .Q (new_AGEMA_signal_5536) ) ;
    buf_clk new_AGEMA_reg_buffer_2077 ( .C (clk), .D (new_AGEMA_signal_5541), .Q (new_AGEMA_signal_5542) ) ;
    buf_clk new_AGEMA_reg_buffer_2083 ( .C (clk), .D (new_AGEMA_signal_5547), .Q (new_AGEMA_signal_5548) ) ;
    buf_clk new_AGEMA_reg_buffer_2089 ( .C (clk), .D (new_AGEMA_signal_5553), .Q (new_AGEMA_signal_5554) ) ;
    buf_clk new_AGEMA_reg_buffer_2095 ( .C (clk), .D (new_AGEMA_signal_5559), .Q (new_AGEMA_signal_5560) ) ;
    buf_clk new_AGEMA_reg_buffer_2101 ( .C (clk), .D (new_AGEMA_signal_5565), .Q (new_AGEMA_signal_5566) ) ;
    buf_clk new_AGEMA_reg_buffer_2107 ( .C (clk), .D (new_AGEMA_signal_5571), .Q (new_AGEMA_signal_5572) ) ;
    buf_clk new_AGEMA_reg_buffer_2113 ( .C (clk), .D (new_AGEMA_signal_5577), .Q (new_AGEMA_signal_5578) ) ;
    buf_clk new_AGEMA_reg_buffer_2119 ( .C (clk), .D (new_AGEMA_signal_5583), .Q (new_AGEMA_signal_5584) ) ;
    buf_clk new_AGEMA_reg_buffer_2125 ( .C (clk), .D (new_AGEMA_signal_5589), .Q (new_AGEMA_signal_5590) ) ;
    buf_clk new_AGEMA_reg_buffer_2131 ( .C (clk), .D (new_AGEMA_signal_5595), .Q (new_AGEMA_signal_5596) ) ;
    buf_clk new_AGEMA_reg_buffer_2137 ( .C (clk), .D (new_AGEMA_signal_5601), .Q (new_AGEMA_signal_5602) ) ;
    buf_clk new_AGEMA_reg_buffer_2143 ( .C (clk), .D (new_AGEMA_signal_5607), .Q (new_AGEMA_signal_5608) ) ;
    buf_clk new_AGEMA_reg_buffer_2149 ( .C (clk), .D (new_AGEMA_signal_5613), .Q (new_AGEMA_signal_5614) ) ;
    buf_clk new_AGEMA_reg_buffer_2155 ( .C (clk), .D (new_AGEMA_signal_5619), .Q (new_AGEMA_signal_5620) ) ;
    buf_clk new_AGEMA_reg_buffer_2161 ( .C (clk), .D (new_AGEMA_signal_5625), .Q (new_AGEMA_signal_5626) ) ;
    buf_clk new_AGEMA_reg_buffer_2167 ( .C (clk), .D (new_AGEMA_signal_5631), .Q (new_AGEMA_signal_5632) ) ;
    buf_clk new_AGEMA_reg_buffer_2173 ( .C (clk), .D (new_AGEMA_signal_5637), .Q (new_AGEMA_signal_5638) ) ;
    buf_clk new_AGEMA_reg_buffer_2179 ( .C (clk), .D (new_AGEMA_signal_5643), .Q (new_AGEMA_signal_5644) ) ;
    buf_clk new_AGEMA_reg_buffer_2185 ( .C (clk), .D (new_AGEMA_signal_5649), .Q (new_AGEMA_signal_5650) ) ;
    buf_clk new_AGEMA_reg_buffer_2191 ( .C (clk), .D (new_AGEMA_signal_5655), .Q (new_AGEMA_signal_5656) ) ;
    buf_clk new_AGEMA_reg_buffer_2197 ( .C (clk), .D (new_AGEMA_signal_5661), .Q (new_AGEMA_signal_5662) ) ;
    buf_clk new_AGEMA_reg_buffer_2203 ( .C (clk), .D (new_AGEMA_signal_5667), .Q (new_AGEMA_signal_5668) ) ;
    buf_clk new_AGEMA_reg_buffer_2209 ( .C (clk), .D (new_AGEMA_signal_5673), .Q (new_AGEMA_signal_5674) ) ;
    buf_clk new_AGEMA_reg_buffer_2215 ( .C (clk), .D (new_AGEMA_signal_5679), .Q (new_AGEMA_signal_5680) ) ;
    buf_clk new_AGEMA_reg_buffer_2221 ( .C (clk), .D (new_AGEMA_signal_5685), .Q (new_AGEMA_signal_5686) ) ;
    buf_clk new_AGEMA_reg_buffer_2227 ( .C (clk), .D (new_AGEMA_signal_5691), .Q (new_AGEMA_signal_5692) ) ;
    buf_clk new_AGEMA_reg_buffer_2233 ( .C (clk), .D (new_AGEMA_signal_5697), .Q (new_AGEMA_signal_5698) ) ;
    buf_clk new_AGEMA_reg_buffer_2239 ( .C (clk), .D (new_AGEMA_signal_5703), .Q (new_AGEMA_signal_5704) ) ;
    buf_clk new_AGEMA_reg_buffer_2245 ( .C (clk), .D (new_AGEMA_signal_5709), .Q (new_AGEMA_signal_5710) ) ;
    buf_clk new_AGEMA_reg_buffer_2251 ( .C (clk), .D (new_AGEMA_signal_5715), .Q (new_AGEMA_signal_5716) ) ;
    buf_clk new_AGEMA_reg_buffer_2257 ( .C (clk), .D (new_AGEMA_signal_5721), .Q (new_AGEMA_signal_5722) ) ;
    buf_clk new_AGEMA_reg_buffer_2263 ( .C (clk), .D (new_AGEMA_signal_5727), .Q (new_AGEMA_signal_5728) ) ;
    buf_clk new_AGEMA_reg_buffer_2269 ( .C (clk), .D (new_AGEMA_signal_5733), .Q (new_AGEMA_signal_5734) ) ;
    buf_clk new_AGEMA_reg_buffer_2275 ( .C (clk), .D (new_AGEMA_signal_5739), .Q (new_AGEMA_signal_5740) ) ;
    buf_clk new_AGEMA_reg_buffer_2281 ( .C (clk), .D (new_AGEMA_signal_5745), .Q (new_AGEMA_signal_5746) ) ;
    buf_clk new_AGEMA_reg_buffer_2287 ( .C (clk), .D (new_AGEMA_signal_5751), .Q (new_AGEMA_signal_5752) ) ;
    buf_clk new_AGEMA_reg_buffer_2293 ( .C (clk), .D (new_AGEMA_signal_5757), .Q (new_AGEMA_signal_5758) ) ;
    buf_clk new_AGEMA_reg_buffer_2299 ( .C (clk), .D (new_AGEMA_signal_5763), .Q (new_AGEMA_signal_5764) ) ;
    buf_clk new_AGEMA_reg_buffer_2305 ( .C (clk), .D (new_AGEMA_signal_5769), .Q (new_AGEMA_signal_5770) ) ;
    buf_clk new_AGEMA_reg_buffer_2311 ( .C (clk), .D (new_AGEMA_signal_5775), .Q (new_AGEMA_signal_5776) ) ;
    buf_clk new_AGEMA_reg_buffer_2317 ( .C (clk), .D (new_AGEMA_signal_5781), .Q (new_AGEMA_signal_5782) ) ;
    buf_clk new_AGEMA_reg_buffer_2323 ( .C (clk), .D (new_AGEMA_signal_5787), .Q (new_AGEMA_signal_5788) ) ;
    buf_clk new_AGEMA_reg_buffer_2329 ( .C (clk), .D (new_AGEMA_signal_5793), .Q (new_AGEMA_signal_5794) ) ;
    buf_clk new_AGEMA_reg_buffer_2335 ( .C (clk), .D (new_AGEMA_signal_5799), .Q (new_AGEMA_signal_5800) ) ;
    buf_clk new_AGEMA_reg_buffer_2341 ( .C (clk), .D (new_AGEMA_signal_5805), .Q (new_AGEMA_signal_5806) ) ;
    buf_clk new_AGEMA_reg_buffer_2347 ( .C (clk), .D (new_AGEMA_signal_5811), .Q (new_AGEMA_signal_5812) ) ;
    buf_clk new_AGEMA_reg_buffer_2353 ( .C (clk), .D (new_AGEMA_signal_5817), .Q (new_AGEMA_signal_5818) ) ;
    buf_clk new_AGEMA_reg_buffer_2359 ( .C (clk), .D (new_AGEMA_signal_5823), .Q (new_AGEMA_signal_5824) ) ;
    buf_clk new_AGEMA_reg_buffer_2365 ( .C (clk), .D (new_AGEMA_signal_5829), .Q (new_AGEMA_signal_5830) ) ;
    buf_clk new_AGEMA_reg_buffer_2371 ( .C (clk), .D (new_AGEMA_signal_5835), .Q (new_AGEMA_signal_5836) ) ;
    buf_clk new_AGEMA_reg_buffer_2377 ( .C (clk), .D (new_AGEMA_signal_5841), .Q (new_AGEMA_signal_5842) ) ;
    buf_clk new_AGEMA_reg_buffer_2383 ( .C (clk), .D (new_AGEMA_signal_5847), .Q (new_AGEMA_signal_5848) ) ;
    buf_clk new_AGEMA_reg_buffer_2389 ( .C (clk), .D (new_AGEMA_signal_5853), .Q (new_AGEMA_signal_5854) ) ;
    buf_clk new_AGEMA_reg_buffer_2395 ( .C (clk), .D (new_AGEMA_signal_5859), .Q (new_AGEMA_signal_5860) ) ;
    buf_clk new_AGEMA_reg_buffer_2401 ( .C (clk), .D (new_AGEMA_signal_5865), .Q (new_AGEMA_signal_5866) ) ;
    buf_clk new_AGEMA_reg_buffer_2407 ( .C (clk), .D (new_AGEMA_signal_5871), .Q (new_AGEMA_signal_5872) ) ;
    buf_clk new_AGEMA_reg_buffer_2413 ( .C (clk), .D (new_AGEMA_signal_5877), .Q (new_AGEMA_signal_5878) ) ;
    buf_clk new_AGEMA_reg_buffer_2419 ( .C (clk), .D (new_AGEMA_signal_5883), .Q (new_AGEMA_signal_5884) ) ;
    buf_clk new_AGEMA_reg_buffer_2425 ( .C (clk), .D (new_AGEMA_signal_5889), .Q (new_AGEMA_signal_5890) ) ;
    buf_clk new_AGEMA_reg_buffer_2431 ( .C (clk), .D (new_AGEMA_signal_5895), .Q (new_AGEMA_signal_5896) ) ;
    buf_clk new_AGEMA_reg_buffer_2437 ( .C (clk), .D (new_AGEMA_signal_5901), .Q (new_AGEMA_signal_5902) ) ;
    buf_clk new_AGEMA_reg_buffer_2443 ( .C (clk), .D (new_AGEMA_signal_5907), .Q (new_AGEMA_signal_5908) ) ;
    buf_clk new_AGEMA_reg_buffer_2449 ( .C (clk), .D (new_AGEMA_signal_5913), .Q (new_AGEMA_signal_5914) ) ;
    buf_clk new_AGEMA_reg_buffer_2455 ( .C (clk), .D (new_AGEMA_signal_5919), .Q (new_AGEMA_signal_5920) ) ;
    buf_clk new_AGEMA_reg_buffer_2461 ( .C (clk), .D (new_AGEMA_signal_5925), .Q (new_AGEMA_signal_5926) ) ;
    buf_clk new_AGEMA_reg_buffer_2467 ( .C (clk), .D (new_AGEMA_signal_5931), .Q (new_AGEMA_signal_5932) ) ;
    buf_clk new_AGEMA_reg_buffer_2473 ( .C (clk), .D (new_AGEMA_signal_5937), .Q (new_AGEMA_signal_5938) ) ;
    buf_clk new_AGEMA_reg_buffer_2479 ( .C (clk), .D (new_AGEMA_signal_5943), .Q (new_AGEMA_signal_5944) ) ;
    buf_clk new_AGEMA_reg_buffer_2485 ( .C (clk), .D (new_AGEMA_signal_5949), .Q (new_AGEMA_signal_5950) ) ;
    buf_clk new_AGEMA_reg_buffer_2491 ( .C (clk), .D (new_AGEMA_signal_5955), .Q (new_AGEMA_signal_5956) ) ;
    buf_clk new_AGEMA_reg_buffer_2497 ( .C (clk), .D (new_AGEMA_signal_5961), .Q (new_AGEMA_signal_5962) ) ;
    buf_clk new_AGEMA_reg_buffer_2503 ( .C (clk), .D (new_AGEMA_signal_5967), .Q (new_AGEMA_signal_5968) ) ;
    buf_clk new_AGEMA_reg_buffer_2509 ( .C (clk), .D (new_AGEMA_signal_5973), .Q (new_AGEMA_signal_5974) ) ;
    buf_clk new_AGEMA_reg_buffer_2515 ( .C (clk), .D (new_AGEMA_signal_5979), .Q (new_AGEMA_signal_5980) ) ;
    buf_clk new_AGEMA_reg_buffer_2521 ( .C (clk), .D (new_AGEMA_signal_5985), .Q (new_AGEMA_signal_5986) ) ;
    buf_clk new_AGEMA_reg_buffer_2527 ( .C (clk), .D (new_AGEMA_signal_5991), .Q (new_AGEMA_signal_5992) ) ;
    buf_clk new_AGEMA_reg_buffer_2533 ( .C (clk), .D (new_AGEMA_signal_5997), .Q (new_AGEMA_signal_5998) ) ;
    buf_clk new_AGEMA_reg_buffer_2539 ( .C (clk), .D (new_AGEMA_signal_6003), .Q (new_AGEMA_signal_6004) ) ;
    buf_clk new_AGEMA_reg_buffer_2545 ( .C (clk), .D (new_AGEMA_signal_6009), .Q (new_AGEMA_signal_6010) ) ;
    buf_clk new_AGEMA_reg_buffer_2551 ( .C (clk), .D (new_AGEMA_signal_6015), .Q (new_AGEMA_signal_6016) ) ;
    buf_clk new_AGEMA_reg_buffer_2557 ( .C (clk), .D (new_AGEMA_signal_6021), .Q (new_AGEMA_signal_6022) ) ;
    buf_clk new_AGEMA_reg_buffer_2563 ( .C (clk), .D (new_AGEMA_signal_6027), .Q (new_AGEMA_signal_6028) ) ;
    buf_clk new_AGEMA_reg_buffer_2569 ( .C (clk), .D (new_AGEMA_signal_6033), .Q (new_AGEMA_signal_6034) ) ;
    buf_clk new_AGEMA_reg_buffer_2575 ( .C (clk), .D (new_AGEMA_signal_6039), .Q (new_AGEMA_signal_6040) ) ;
    buf_clk new_AGEMA_reg_buffer_2581 ( .C (clk), .D (new_AGEMA_signal_6045), .Q (new_AGEMA_signal_6046) ) ;
    buf_clk new_AGEMA_reg_buffer_2587 ( .C (clk), .D (new_AGEMA_signal_6051), .Q (new_AGEMA_signal_6052) ) ;
    buf_clk new_AGEMA_reg_buffer_2593 ( .C (clk), .D (new_AGEMA_signal_6057), .Q (new_AGEMA_signal_6058) ) ;
    buf_clk new_AGEMA_reg_buffer_2599 ( .C (clk), .D (new_AGEMA_signal_6063), .Q (new_AGEMA_signal_6064) ) ;
    buf_clk new_AGEMA_reg_buffer_2605 ( .C (clk), .D (new_AGEMA_signal_6069), .Q (new_AGEMA_signal_6070) ) ;
    buf_clk new_AGEMA_reg_buffer_2611 ( .C (clk), .D (new_AGEMA_signal_6075), .Q (new_AGEMA_signal_6076) ) ;
    buf_clk new_AGEMA_reg_buffer_2617 ( .C (clk), .D (new_AGEMA_signal_6081), .Q (new_AGEMA_signal_6082) ) ;
    buf_clk new_AGEMA_reg_buffer_2623 ( .C (clk), .D (new_AGEMA_signal_6087), .Q (new_AGEMA_signal_6088) ) ;
    buf_clk new_AGEMA_reg_buffer_2629 ( .C (clk), .D (new_AGEMA_signal_6093), .Q (new_AGEMA_signal_6094) ) ;
    buf_clk new_AGEMA_reg_buffer_2635 ( .C (clk), .D (new_AGEMA_signal_6099), .Q (new_AGEMA_signal_6100) ) ;
    buf_clk new_AGEMA_reg_buffer_2641 ( .C (clk), .D (new_AGEMA_signal_6105), .Q (new_AGEMA_signal_6106) ) ;
    buf_clk new_AGEMA_reg_buffer_2647 ( .C (clk), .D (new_AGEMA_signal_6111), .Q (new_AGEMA_signal_6112) ) ;
    buf_clk new_AGEMA_reg_buffer_2653 ( .C (clk), .D (new_AGEMA_signal_6117), .Q (new_AGEMA_signal_6118) ) ;
    buf_clk new_AGEMA_reg_buffer_2659 ( .C (clk), .D (new_AGEMA_signal_6123), .Q (new_AGEMA_signal_6124) ) ;
    buf_clk new_AGEMA_reg_buffer_2665 ( .C (clk), .D (new_AGEMA_signal_6129), .Q (new_AGEMA_signal_6130) ) ;
    buf_clk new_AGEMA_reg_buffer_2671 ( .C (clk), .D (new_AGEMA_signal_6135), .Q (new_AGEMA_signal_6136) ) ;
    buf_clk new_AGEMA_reg_buffer_2677 ( .C (clk), .D (new_AGEMA_signal_6141), .Q (new_AGEMA_signal_6142) ) ;
    buf_clk new_AGEMA_reg_buffer_2683 ( .C (clk), .D (new_AGEMA_signal_6147), .Q (new_AGEMA_signal_6148) ) ;
    buf_clk new_AGEMA_reg_buffer_2689 ( .C (clk), .D (new_AGEMA_signal_6153), .Q (new_AGEMA_signal_6154) ) ;
    buf_clk new_AGEMA_reg_buffer_2695 ( .C (clk), .D (new_AGEMA_signal_6159), .Q (new_AGEMA_signal_6160) ) ;
    buf_clk new_AGEMA_reg_buffer_2701 ( .C (clk), .D (new_AGEMA_signal_6165), .Q (new_AGEMA_signal_6166) ) ;
    buf_clk new_AGEMA_reg_buffer_2707 ( .C (clk), .D (new_AGEMA_signal_6171), .Q (new_AGEMA_signal_6172) ) ;
    buf_clk new_AGEMA_reg_buffer_2713 ( .C (clk), .D (new_AGEMA_signal_6177), .Q (new_AGEMA_signal_6178) ) ;
    buf_clk new_AGEMA_reg_buffer_2719 ( .C (clk), .D (new_AGEMA_signal_6183), .Q (new_AGEMA_signal_6184) ) ;
    buf_clk new_AGEMA_reg_buffer_2725 ( .C (clk), .D (new_AGEMA_signal_6189), .Q (new_AGEMA_signal_6190) ) ;
    buf_clk new_AGEMA_reg_buffer_2731 ( .C (clk), .D (new_AGEMA_signal_6195), .Q (new_AGEMA_signal_6196) ) ;
    buf_clk new_AGEMA_reg_buffer_2737 ( .C (clk), .D (new_AGEMA_signal_6201), .Q (new_AGEMA_signal_6202) ) ;
    buf_clk new_AGEMA_reg_buffer_2743 ( .C (clk), .D (new_AGEMA_signal_6207), .Q (new_AGEMA_signal_6208) ) ;
    buf_clk new_AGEMA_reg_buffer_2749 ( .C (clk), .D (new_AGEMA_signal_6213), .Q (new_AGEMA_signal_6214) ) ;
    buf_clk new_AGEMA_reg_buffer_2755 ( .C (clk), .D (new_AGEMA_signal_6219), .Q (new_AGEMA_signal_6220) ) ;
    buf_clk new_AGEMA_reg_buffer_2761 ( .C (clk), .D (new_AGEMA_signal_6225), .Q (new_AGEMA_signal_6226) ) ;
    buf_clk new_AGEMA_reg_buffer_2767 ( .C (clk), .D (new_AGEMA_signal_6231), .Q (new_AGEMA_signal_6232) ) ;
    buf_clk new_AGEMA_reg_buffer_2773 ( .C (clk), .D (new_AGEMA_signal_6237), .Q (new_AGEMA_signal_6238) ) ;
    buf_clk new_AGEMA_reg_buffer_2779 ( .C (clk), .D (new_AGEMA_signal_6243), .Q (new_AGEMA_signal_6244) ) ;
    buf_clk new_AGEMA_reg_buffer_2785 ( .C (clk), .D (new_AGEMA_signal_6249), .Q (new_AGEMA_signal_6250) ) ;
    buf_clk new_AGEMA_reg_buffer_2791 ( .C (clk), .D (new_AGEMA_signal_6255), .Q (new_AGEMA_signal_6256) ) ;
    buf_clk new_AGEMA_reg_buffer_2797 ( .C (clk), .D (new_AGEMA_signal_6261), .Q (new_AGEMA_signal_6262) ) ;
    buf_clk new_AGEMA_reg_buffer_2803 ( .C (clk), .D (new_AGEMA_signal_6267), .Q (new_AGEMA_signal_6268) ) ;
    buf_clk new_AGEMA_reg_buffer_2809 ( .C (clk), .D (new_AGEMA_signal_6273), .Q (new_AGEMA_signal_6274) ) ;
    buf_clk new_AGEMA_reg_buffer_2815 ( .C (clk), .D (new_AGEMA_signal_6279), .Q (new_AGEMA_signal_6280) ) ;
    buf_clk new_AGEMA_reg_buffer_2821 ( .C (clk), .D (new_AGEMA_signal_6285), .Q (new_AGEMA_signal_6286) ) ;
    buf_clk new_AGEMA_reg_buffer_2827 ( .C (clk), .D (new_AGEMA_signal_6291), .Q (new_AGEMA_signal_6292) ) ;
    buf_clk new_AGEMA_reg_buffer_2833 ( .C (clk), .D (new_AGEMA_signal_6297), .Q (new_AGEMA_signal_6298) ) ;
    buf_clk new_AGEMA_reg_buffer_2839 ( .C (clk), .D (new_AGEMA_signal_6303), .Q (new_AGEMA_signal_6304) ) ;
    buf_clk new_AGEMA_reg_buffer_2845 ( .C (clk), .D (new_AGEMA_signal_6309), .Q (new_AGEMA_signal_6310) ) ;
    buf_clk new_AGEMA_reg_buffer_2851 ( .C (clk), .D (new_AGEMA_signal_6315), .Q (new_AGEMA_signal_6316) ) ;
    buf_clk new_AGEMA_reg_buffer_2857 ( .C (clk), .D (new_AGEMA_signal_6321), .Q (new_AGEMA_signal_6322) ) ;
    buf_clk new_AGEMA_reg_buffer_2863 ( .C (clk), .D (new_AGEMA_signal_6327), .Q (new_AGEMA_signal_6328) ) ;
    buf_clk new_AGEMA_reg_buffer_2869 ( .C (clk), .D (new_AGEMA_signal_6333), .Q (new_AGEMA_signal_6334) ) ;
    buf_clk new_AGEMA_reg_buffer_2875 ( .C (clk), .D (new_AGEMA_signal_6339), .Q (new_AGEMA_signal_6340) ) ;
    buf_clk new_AGEMA_reg_buffer_2881 ( .C (clk), .D (new_AGEMA_signal_6345), .Q (new_AGEMA_signal_6346) ) ;
    buf_clk new_AGEMA_reg_buffer_2887 ( .C (clk), .D (new_AGEMA_signal_6351), .Q (new_AGEMA_signal_6352) ) ;
    buf_clk new_AGEMA_reg_buffer_2893 ( .C (clk), .D (new_AGEMA_signal_6357), .Q (new_AGEMA_signal_6358) ) ;
    buf_clk new_AGEMA_reg_buffer_2899 ( .C (clk), .D (new_AGEMA_signal_6363), .Q (new_AGEMA_signal_6364) ) ;
    buf_clk new_AGEMA_reg_buffer_2905 ( .C (clk), .D (new_AGEMA_signal_6369), .Q (new_AGEMA_signal_6370) ) ;
    buf_clk new_AGEMA_reg_buffer_2911 ( .C (clk), .D (new_AGEMA_signal_6375), .Q (new_AGEMA_signal_6376) ) ;
    buf_clk new_AGEMA_reg_buffer_2917 ( .C (clk), .D (new_AGEMA_signal_6381), .Q (new_AGEMA_signal_6382) ) ;
    buf_clk new_AGEMA_reg_buffer_2923 ( .C (clk), .D (new_AGEMA_signal_6387), .Q (new_AGEMA_signal_6388) ) ;
    buf_clk new_AGEMA_reg_buffer_2929 ( .C (clk), .D (new_AGEMA_signal_6393), .Q (new_AGEMA_signal_6394) ) ;
    buf_clk new_AGEMA_reg_buffer_2935 ( .C (clk), .D (new_AGEMA_signal_6399), .Q (new_AGEMA_signal_6400) ) ;
    buf_clk new_AGEMA_reg_buffer_2941 ( .C (clk), .D (new_AGEMA_signal_6405), .Q (new_AGEMA_signal_6406) ) ;
    buf_clk new_AGEMA_reg_buffer_2947 ( .C (clk), .D (new_AGEMA_signal_6411), .Q (new_AGEMA_signal_6412) ) ;
    buf_clk new_AGEMA_reg_buffer_2953 ( .C (clk), .D (new_AGEMA_signal_6417), .Q (new_AGEMA_signal_6418) ) ;
    buf_clk new_AGEMA_reg_buffer_2959 ( .C (clk), .D (new_AGEMA_signal_6423), .Q (new_AGEMA_signal_6424) ) ;
    buf_clk new_AGEMA_reg_buffer_2965 ( .C (clk), .D (new_AGEMA_signal_6429), .Q (new_AGEMA_signal_6430) ) ;
    buf_clk new_AGEMA_reg_buffer_2971 ( .C (clk), .D (new_AGEMA_signal_6435), .Q (new_AGEMA_signal_6436) ) ;
    buf_clk new_AGEMA_reg_buffer_2977 ( .C (clk), .D (new_AGEMA_signal_6441), .Q (new_AGEMA_signal_6442) ) ;
    buf_clk new_AGEMA_reg_buffer_2983 ( .C (clk), .D (new_AGEMA_signal_6447), .Q (new_AGEMA_signal_6448) ) ;
    buf_clk new_AGEMA_reg_buffer_2989 ( .C (clk), .D (new_AGEMA_signal_6453), .Q (new_AGEMA_signal_6454) ) ;
    buf_clk new_AGEMA_reg_buffer_2995 ( .C (clk), .D (new_AGEMA_signal_6459), .Q (new_AGEMA_signal_6460) ) ;
    buf_clk new_AGEMA_reg_buffer_3001 ( .C (clk), .D (new_AGEMA_signal_6465), .Q (new_AGEMA_signal_6466) ) ;
    buf_clk new_AGEMA_reg_buffer_3007 ( .C (clk), .D (new_AGEMA_signal_6471), .Q (new_AGEMA_signal_6472) ) ;
    buf_clk new_AGEMA_reg_buffer_3013 ( .C (clk), .D (new_AGEMA_signal_6477), .Q (new_AGEMA_signal_6478) ) ;
    buf_clk new_AGEMA_reg_buffer_3019 ( .C (clk), .D (new_AGEMA_signal_6483), .Q (new_AGEMA_signal_6484) ) ;
    buf_clk new_AGEMA_reg_buffer_3025 ( .C (clk), .D (new_AGEMA_signal_6489), .Q (new_AGEMA_signal_6490) ) ;
    buf_clk new_AGEMA_reg_buffer_3031 ( .C (clk), .D (new_AGEMA_signal_6495), .Q (new_AGEMA_signal_6496) ) ;
    buf_clk new_AGEMA_reg_buffer_3037 ( .C (clk), .D (new_AGEMA_signal_6501), .Q (new_AGEMA_signal_6502) ) ;
    buf_clk new_AGEMA_reg_buffer_3043 ( .C (clk), .D (new_AGEMA_signal_6507), .Q (new_AGEMA_signal_6508) ) ;
    buf_clk new_AGEMA_reg_buffer_3049 ( .C (clk), .D (new_AGEMA_signal_6513), .Q (new_AGEMA_signal_6514) ) ;
    buf_clk new_AGEMA_reg_buffer_3055 ( .C (clk), .D (new_AGEMA_signal_6519), .Q (new_AGEMA_signal_6520) ) ;
    buf_clk new_AGEMA_reg_buffer_3061 ( .C (clk), .D (new_AGEMA_signal_6525), .Q (new_AGEMA_signal_6526) ) ;
    buf_clk new_AGEMA_reg_buffer_3067 ( .C (clk), .D (new_AGEMA_signal_6531), .Q (new_AGEMA_signal_6532) ) ;
    buf_clk new_AGEMA_reg_buffer_3073 ( .C (clk), .D (new_AGEMA_signal_6537), .Q (new_AGEMA_signal_6538) ) ;
    buf_clk new_AGEMA_reg_buffer_3079 ( .C (clk), .D (new_AGEMA_signal_6543), .Q (new_AGEMA_signal_6544) ) ;
    buf_clk new_AGEMA_reg_buffer_3085 ( .C (clk), .D (new_AGEMA_signal_6549), .Q (new_AGEMA_signal_6550) ) ;
    buf_clk new_AGEMA_reg_buffer_3091 ( .C (clk), .D (new_AGEMA_signal_6555), .Q (new_AGEMA_signal_6556) ) ;
    buf_clk new_AGEMA_reg_buffer_3097 ( .C (clk), .D (new_AGEMA_signal_6561), .Q (new_AGEMA_signal_6562) ) ;
    buf_clk new_AGEMA_reg_buffer_3103 ( .C (clk), .D (new_AGEMA_signal_6567), .Q (new_AGEMA_signal_6568) ) ;
    buf_clk new_AGEMA_reg_buffer_3109 ( .C (clk), .D (new_AGEMA_signal_6573), .Q (new_AGEMA_signal_6574) ) ;
    buf_clk new_AGEMA_reg_buffer_3115 ( .C (clk), .D (new_AGEMA_signal_6579), .Q (new_AGEMA_signal_6580) ) ;
    buf_clk new_AGEMA_reg_buffer_3121 ( .C (clk), .D (new_AGEMA_signal_6585), .Q (new_AGEMA_signal_6586) ) ;
    buf_clk new_AGEMA_reg_buffer_3127 ( .C (clk), .D (new_AGEMA_signal_6591), .Q (new_AGEMA_signal_6592) ) ;
    buf_clk new_AGEMA_reg_buffer_3133 ( .C (clk), .D (new_AGEMA_signal_6597), .Q (new_AGEMA_signal_6598) ) ;
    buf_clk new_AGEMA_reg_buffer_3139 ( .C (clk), .D (new_AGEMA_signal_6603), .Q (new_AGEMA_signal_6604) ) ;
    buf_clk new_AGEMA_reg_buffer_3145 ( .C (clk), .D (new_AGEMA_signal_6609), .Q (new_AGEMA_signal_6610) ) ;
    buf_clk new_AGEMA_reg_buffer_3151 ( .C (clk), .D (new_AGEMA_signal_6615), .Q (new_AGEMA_signal_6616) ) ;
    buf_clk new_AGEMA_reg_buffer_3157 ( .C (clk), .D (new_AGEMA_signal_6621), .Q (new_AGEMA_signal_6622) ) ;
    buf_clk new_AGEMA_reg_buffer_3163 ( .C (clk), .D (new_AGEMA_signal_6627), .Q (new_AGEMA_signal_6628) ) ;
    buf_clk new_AGEMA_reg_buffer_3169 ( .C (clk), .D (new_AGEMA_signal_6633), .Q (new_AGEMA_signal_6634) ) ;
    buf_clk new_AGEMA_reg_buffer_3175 ( .C (clk), .D (new_AGEMA_signal_6639), .Q (new_AGEMA_signal_6640) ) ;
    buf_clk new_AGEMA_reg_buffer_3181 ( .C (clk), .D (new_AGEMA_signal_6645), .Q (new_AGEMA_signal_6646) ) ;
    buf_clk new_AGEMA_reg_buffer_3187 ( .C (clk), .D (new_AGEMA_signal_6651), .Q (new_AGEMA_signal_6652) ) ;
    buf_clk new_AGEMA_reg_buffer_3193 ( .C (clk), .D (new_AGEMA_signal_6657), .Q (new_AGEMA_signal_6658) ) ;
    buf_clk new_AGEMA_reg_buffer_3199 ( .C (clk), .D (new_AGEMA_signal_6663), .Q (new_AGEMA_signal_6664) ) ;
    buf_clk new_AGEMA_reg_buffer_3205 ( .C (clk), .D (new_AGEMA_signal_6669), .Q (new_AGEMA_signal_6670) ) ;
    buf_clk new_AGEMA_reg_buffer_3211 ( .C (clk), .D (new_AGEMA_signal_6675), .Q (new_AGEMA_signal_6676) ) ;
    buf_clk new_AGEMA_reg_buffer_3217 ( .C (clk), .D (new_AGEMA_signal_6681), .Q (new_AGEMA_signal_6682) ) ;
    buf_clk new_AGEMA_reg_buffer_3223 ( .C (clk), .D (new_AGEMA_signal_6687), .Q (new_AGEMA_signal_6688) ) ;
    buf_clk new_AGEMA_reg_buffer_3229 ( .C (clk), .D (new_AGEMA_signal_6693), .Q (new_AGEMA_signal_6694) ) ;
    buf_clk new_AGEMA_reg_buffer_3235 ( .C (clk), .D (new_AGEMA_signal_6699), .Q (new_AGEMA_signal_6700) ) ;
    buf_clk new_AGEMA_reg_buffer_3241 ( .C (clk), .D (new_AGEMA_signal_6705), .Q (new_AGEMA_signal_6706) ) ;
    buf_clk new_AGEMA_reg_buffer_3247 ( .C (clk), .D (new_AGEMA_signal_6711), .Q (new_AGEMA_signal_6712) ) ;
    buf_clk new_AGEMA_reg_buffer_3253 ( .C (clk), .D (new_AGEMA_signal_6717), .Q (new_AGEMA_signal_6718) ) ;
    buf_clk new_AGEMA_reg_buffer_3259 ( .C (clk), .D (new_AGEMA_signal_6723), .Q (new_AGEMA_signal_6724) ) ;
    buf_clk new_AGEMA_reg_buffer_3265 ( .C (clk), .D (new_AGEMA_signal_6729), .Q (new_AGEMA_signal_6730) ) ;
    buf_clk new_AGEMA_reg_buffer_3271 ( .C (clk), .D (new_AGEMA_signal_6735), .Q (new_AGEMA_signal_6736) ) ;
    buf_clk new_AGEMA_reg_buffer_3277 ( .C (clk), .D (new_AGEMA_signal_6741), .Q (new_AGEMA_signal_6742) ) ;
    buf_clk new_AGEMA_reg_buffer_3283 ( .C (clk), .D (new_AGEMA_signal_6747), .Q (new_AGEMA_signal_6748) ) ;
    buf_clk new_AGEMA_reg_buffer_3289 ( .C (clk), .D (new_AGEMA_signal_6753), .Q (new_AGEMA_signal_6754) ) ;
    buf_clk new_AGEMA_reg_buffer_3295 ( .C (clk), .D (new_AGEMA_signal_6759), .Q (new_AGEMA_signal_6760) ) ;
    buf_clk new_AGEMA_reg_buffer_3301 ( .C (clk), .D (new_AGEMA_signal_6765), .Q (new_AGEMA_signal_6766) ) ;
    buf_clk new_AGEMA_reg_buffer_3307 ( .C (clk), .D (new_AGEMA_signal_6771), .Q (new_AGEMA_signal_6772) ) ;
    buf_clk new_AGEMA_reg_buffer_3313 ( .C (clk), .D (new_AGEMA_signal_6777), .Q (new_AGEMA_signal_6778) ) ;
    buf_clk new_AGEMA_reg_buffer_3319 ( .C (clk), .D (new_AGEMA_signal_6783), .Q (new_AGEMA_signal_6784) ) ;
    buf_clk new_AGEMA_reg_buffer_3325 ( .C (clk), .D (new_AGEMA_signal_6789), .Q (new_AGEMA_signal_6790) ) ;
    buf_clk new_AGEMA_reg_buffer_3331 ( .C (clk), .D (new_AGEMA_signal_6795), .Q (new_AGEMA_signal_6796) ) ;
    buf_clk new_AGEMA_reg_buffer_3337 ( .C (clk), .D (new_AGEMA_signal_6801), .Q (new_AGEMA_signal_6802) ) ;
    buf_clk new_AGEMA_reg_buffer_3343 ( .C (clk), .D (new_AGEMA_signal_6807), .Q (new_AGEMA_signal_6808) ) ;
    buf_clk new_AGEMA_reg_buffer_3349 ( .C (clk), .D (new_AGEMA_signal_6813), .Q (new_AGEMA_signal_6814) ) ;
    buf_clk new_AGEMA_reg_buffer_3355 ( .C (clk), .D (new_AGEMA_signal_6819), .Q (new_AGEMA_signal_6820) ) ;
    buf_clk new_AGEMA_reg_buffer_3361 ( .C (clk), .D (new_AGEMA_signal_6825), .Q (new_AGEMA_signal_6826) ) ;
    buf_clk new_AGEMA_reg_buffer_3367 ( .C (clk), .D (new_AGEMA_signal_6831), .Q (new_AGEMA_signal_6832) ) ;
    buf_clk new_AGEMA_reg_buffer_3373 ( .C (clk), .D (new_AGEMA_signal_6837), .Q (new_AGEMA_signal_6838) ) ;
    buf_clk new_AGEMA_reg_buffer_3379 ( .C (clk), .D (new_AGEMA_signal_6843), .Q (new_AGEMA_signal_6844) ) ;
    buf_clk new_AGEMA_reg_buffer_3385 ( .C (clk), .D (new_AGEMA_signal_6849), .Q (new_AGEMA_signal_6850) ) ;
    buf_clk new_AGEMA_reg_buffer_3391 ( .C (clk), .D (new_AGEMA_signal_6855), .Q (new_AGEMA_signal_6856) ) ;
    buf_clk new_AGEMA_reg_buffer_3397 ( .C (clk), .D (new_AGEMA_signal_6861), .Q (new_AGEMA_signal_6862) ) ;
    buf_clk new_AGEMA_reg_buffer_3403 ( .C (clk), .D (new_AGEMA_signal_6867), .Q (new_AGEMA_signal_6868) ) ;
    buf_clk new_AGEMA_reg_buffer_3409 ( .C (clk), .D (new_AGEMA_signal_6873), .Q (new_AGEMA_signal_6874) ) ;
    buf_clk new_AGEMA_reg_buffer_3415 ( .C (clk), .D (new_AGEMA_signal_6879), .Q (new_AGEMA_signal_6880) ) ;
    buf_clk new_AGEMA_reg_buffer_3421 ( .C (clk), .D (new_AGEMA_signal_6885), .Q (new_AGEMA_signal_6886) ) ;
    buf_clk new_AGEMA_reg_buffer_3427 ( .C (clk), .D (new_AGEMA_signal_6891), .Q (new_AGEMA_signal_6892) ) ;
    buf_clk new_AGEMA_reg_buffer_3433 ( .C (clk), .D (new_AGEMA_signal_6897), .Q (new_AGEMA_signal_6898) ) ;
    buf_clk new_AGEMA_reg_buffer_3439 ( .C (clk), .D (new_AGEMA_signal_6903), .Q (new_AGEMA_signal_6904) ) ;
    buf_clk new_AGEMA_reg_buffer_3445 ( .C (clk), .D (new_AGEMA_signal_6909), .Q (new_AGEMA_signal_6910) ) ;
    buf_clk new_AGEMA_reg_buffer_3451 ( .C (clk), .D (new_AGEMA_signal_6915), .Q (new_AGEMA_signal_6916) ) ;
    buf_clk new_AGEMA_reg_buffer_3457 ( .C (clk), .D (new_AGEMA_signal_6921), .Q (new_AGEMA_signal_6922) ) ;
    buf_clk new_AGEMA_reg_buffer_3463 ( .C (clk), .D (new_AGEMA_signal_6927), .Q (new_AGEMA_signal_6928) ) ;
    buf_clk new_AGEMA_reg_buffer_3469 ( .C (clk), .D (new_AGEMA_signal_6933), .Q (new_AGEMA_signal_6934) ) ;
    buf_clk new_AGEMA_reg_buffer_3475 ( .C (clk), .D (new_AGEMA_signal_6939), .Q (new_AGEMA_signal_6940) ) ;
    buf_clk new_AGEMA_reg_buffer_3481 ( .C (clk), .D (new_AGEMA_signal_6945), .Q (new_AGEMA_signal_6946) ) ;
    buf_clk new_AGEMA_reg_buffer_3487 ( .C (clk), .D (new_AGEMA_signal_6951), .Q (new_AGEMA_signal_6952) ) ;
    buf_clk new_AGEMA_reg_buffer_3493 ( .C (clk), .D (new_AGEMA_signal_6957), .Q (new_AGEMA_signal_6958) ) ;
    buf_clk new_AGEMA_reg_buffer_3499 ( .C (clk), .D (new_AGEMA_signal_6963), .Q (new_AGEMA_signal_6964) ) ;
    buf_clk new_AGEMA_reg_buffer_3505 ( .C (clk), .D (new_AGEMA_signal_6969), .Q (new_AGEMA_signal_6970) ) ;
    buf_clk new_AGEMA_reg_buffer_3511 ( .C (clk), .D (new_AGEMA_signal_6975), .Q (new_AGEMA_signal_6976) ) ;
    buf_clk new_AGEMA_reg_buffer_3517 ( .C (clk), .D (new_AGEMA_signal_6981), .Q (new_AGEMA_signal_6982) ) ;
    buf_clk new_AGEMA_reg_buffer_3523 ( .C (clk), .D (new_AGEMA_signal_6987), .Q (new_AGEMA_signal_6988) ) ;
    buf_clk new_AGEMA_reg_buffer_3529 ( .C (clk), .D (new_AGEMA_signal_6993), .Q (new_AGEMA_signal_6994) ) ;
    buf_clk new_AGEMA_reg_buffer_3535 ( .C (clk), .D (new_AGEMA_signal_6999), .Q (new_AGEMA_signal_7000) ) ;
    buf_clk new_AGEMA_reg_buffer_3541 ( .C (clk), .D (new_AGEMA_signal_7005), .Q (new_AGEMA_signal_7006) ) ;
    buf_clk new_AGEMA_reg_buffer_3547 ( .C (clk), .D (new_AGEMA_signal_7011), .Q (new_AGEMA_signal_7012) ) ;
    buf_clk new_AGEMA_reg_buffer_3553 ( .C (clk), .D (new_AGEMA_signal_7017), .Q (new_AGEMA_signal_7018) ) ;
    buf_clk new_AGEMA_reg_buffer_3559 ( .C (clk), .D (new_AGEMA_signal_7023), .Q (new_AGEMA_signal_7024) ) ;
    buf_clk new_AGEMA_reg_buffer_3565 ( .C (clk), .D (new_AGEMA_signal_7029), .Q (new_AGEMA_signal_7030) ) ;
    buf_clk new_AGEMA_reg_buffer_3571 ( .C (clk), .D (new_AGEMA_signal_7035), .Q (new_AGEMA_signal_7036) ) ;
    buf_clk new_AGEMA_reg_buffer_3865 ( .C (clk), .D (new_AGEMA_signal_7329), .Q (new_AGEMA_signal_7330) ) ;
    buf_clk new_AGEMA_reg_buffer_3871 ( .C (clk), .D (new_AGEMA_signal_7335), .Q (new_AGEMA_signal_7336) ) ;
    buf_clk new_AGEMA_reg_buffer_3879 ( .C (clk), .D (new_AGEMA_signal_7343), .Q (new_AGEMA_signal_7344) ) ;
    buf_clk new_AGEMA_reg_buffer_3887 ( .C (clk), .D (new_AGEMA_signal_7351), .Q (new_AGEMA_signal_7352) ) ;
    buf_clk new_AGEMA_reg_buffer_3895 ( .C (clk), .D (new_AGEMA_signal_7359), .Q (new_AGEMA_signal_7360) ) ;
    buf_clk new_AGEMA_reg_buffer_3903 ( .C (clk), .D (new_AGEMA_signal_7367), .Q (new_AGEMA_signal_7368) ) ;
    buf_clk new_AGEMA_reg_buffer_3911 ( .C (clk), .D (new_AGEMA_signal_7375), .Q (new_AGEMA_signal_7376) ) ;
    buf_clk new_AGEMA_reg_buffer_3919 ( .C (clk), .D (new_AGEMA_signal_7383), .Q (new_AGEMA_signal_7384) ) ;
    buf_clk new_AGEMA_reg_buffer_3927 ( .C (clk), .D (new_AGEMA_signal_7391), .Q (new_AGEMA_signal_7392) ) ;
    buf_clk new_AGEMA_reg_buffer_3935 ( .C (clk), .D (new_AGEMA_signal_7399), .Q (new_AGEMA_signal_7400) ) ;
    buf_clk new_AGEMA_reg_buffer_3943 ( .C (clk), .D (new_AGEMA_signal_7407), .Q (new_AGEMA_signal_7408) ) ;
    buf_clk new_AGEMA_reg_buffer_3951 ( .C (clk), .D (new_AGEMA_signal_7415), .Q (new_AGEMA_signal_7416) ) ;
    buf_clk new_AGEMA_reg_buffer_3959 ( .C (clk), .D (new_AGEMA_signal_7423), .Q (new_AGEMA_signal_7424) ) ;
    buf_clk new_AGEMA_reg_buffer_3967 ( .C (clk), .D (new_AGEMA_signal_7431), .Q (new_AGEMA_signal_7432) ) ;
    buf_clk new_AGEMA_reg_buffer_3975 ( .C (clk), .D (new_AGEMA_signal_7439), .Q (new_AGEMA_signal_7440) ) ;
    buf_clk new_AGEMA_reg_buffer_3983 ( .C (clk), .D (new_AGEMA_signal_7447), .Q (new_AGEMA_signal_7448) ) ;
    buf_clk new_AGEMA_reg_buffer_3991 ( .C (clk), .D (new_AGEMA_signal_7455), .Q (new_AGEMA_signal_7456) ) ;
    buf_clk new_AGEMA_reg_buffer_3999 ( .C (clk), .D (new_AGEMA_signal_7463), .Q (new_AGEMA_signal_7464) ) ;
    buf_clk new_AGEMA_reg_buffer_4007 ( .C (clk), .D (new_AGEMA_signal_7471), .Q (new_AGEMA_signal_7472) ) ;
    buf_clk new_AGEMA_reg_buffer_4015 ( .C (clk), .D (new_AGEMA_signal_7479), .Q (new_AGEMA_signal_7480) ) ;
    buf_clk new_AGEMA_reg_buffer_4023 ( .C (clk), .D (new_AGEMA_signal_7487), .Q (new_AGEMA_signal_7488) ) ;
    buf_clk new_AGEMA_reg_buffer_4031 ( .C (clk), .D (new_AGEMA_signal_7495), .Q (new_AGEMA_signal_7496) ) ;
    buf_clk new_AGEMA_reg_buffer_4039 ( .C (clk), .D (new_AGEMA_signal_7503), .Q (new_AGEMA_signal_7504) ) ;
    buf_clk new_AGEMA_reg_buffer_4047 ( .C (clk), .D (new_AGEMA_signal_7511), .Q (new_AGEMA_signal_7512) ) ;
    buf_clk new_AGEMA_reg_buffer_4055 ( .C (clk), .D (new_AGEMA_signal_7519), .Q (new_AGEMA_signal_7520) ) ;
    buf_clk new_AGEMA_reg_buffer_4063 ( .C (clk), .D (new_AGEMA_signal_7527), .Q (new_AGEMA_signal_7528) ) ;
    buf_clk new_AGEMA_reg_buffer_4071 ( .C (clk), .D (new_AGEMA_signal_7535), .Q (new_AGEMA_signal_7536) ) ;
    buf_clk new_AGEMA_reg_buffer_4079 ( .C (clk), .D (new_AGEMA_signal_7543), .Q (new_AGEMA_signal_7544) ) ;
    buf_clk new_AGEMA_reg_buffer_4087 ( .C (clk), .D (new_AGEMA_signal_7551), .Q (new_AGEMA_signal_7552) ) ;
    buf_clk new_AGEMA_reg_buffer_4095 ( .C (clk), .D (new_AGEMA_signal_7559), .Q (new_AGEMA_signal_7560) ) ;
    buf_clk new_AGEMA_reg_buffer_4103 ( .C (clk), .D (new_AGEMA_signal_7567), .Q (new_AGEMA_signal_7568) ) ;
    buf_clk new_AGEMA_reg_buffer_4111 ( .C (clk), .D (new_AGEMA_signal_7575), .Q (new_AGEMA_signal_7576) ) ;
    buf_clk new_AGEMA_reg_buffer_4119 ( .C (clk), .D (new_AGEMA_signal_7583), .Q (new_AGEMA_signal_7584) ) ;
    buf_clk new_AGEMA_reg_buffer_4127 ( .C (clk), .D (new_AGEMA_signal_7591), .Q (new_AGEMA_signal_7592) ) ;
    buf_clk new_AGEMA_reg_buffer_4135 ( .C (clk), .D (new_AGEMA_signal_7599), .Q (new_AGEMA_signal_7600) ) ;
    buf_clk new_AGEMA_reg_buffer_4143 ( .C (clk), .D (new_AGEMA_signal_7607), .Q (new_AGEMA_signal_7608) ) ;
    buf_clk new_AGEMA_reg_buffer_4151 ( .C (clk), .D (new_AGEMA_signal_7615), .Q (new_AGEMA_signal_7616) ) ;
    buf_clk new_AGEMA_reg_buffer_4159 ( .C (clk), .D (new_AGEMA_signal_7623), .Q (new_AGEMA_signal_7624) ) ;
    buf_clk new_AGEMA_reg_buffer_4167 ( .C (clk), .D (new_AGEMA_signal_7631), .Q (new_AGEMA_signal_7632) ) ;
    buf_clk new_AGEMA_reg_buffer_4175 ( .C (clk), .D (new_AGEMA_signal_7639), .Q (new_AGEMA_signal_7640) ) ;
    buf_clk new_AGEMA_reg_buffer_4183 ( .C (clk), .D (new_AGEMA_signal_7647), .Q (new_AGEMA_signal_7648) ) ;
    buf_clk new_AGEMA_reg_buffer_4191 ( .C (clk), .D (new_AGEMA_signal_7655), .Q (new_AGEMA_signal_7656) ) ;
    buf_clk new_AGEMA_reg_buffer_4199 ( .C (clk), .D (new_AGEMA_signal_7663), .Q (new_AGEMA_signal_7664) ) ;
    buf_clk new_AGEMA_reg_buffer_4207 ( .C (clk), .D (new_AGEMA_signal_7671), .Q (new_AGEMA_signal_7672) ) ;
    buf_clk new_AGEMA_reg_buffer_4215 ( .C (clk), .D (new_AGEMA_signal_7679), .Q (new_AGEMA_signal_7680) ) ;
    buf_clk new_AGEMA_reg_buffer_4223 ( .C (clk), .D (new_AGEMA_signal_7687), .Q (new_AGEMA_signal_7688) ) ;
    buf_clk new_AGEMA_reg_buffer_4231 ( .C (clk), .D (new_AGEMA_signal_7695), .Q (new_AGEMA_signal_7696) ) ;
    buf_clk new_AGEMA_reg_buffer_4239 ( .C (clk), .D (new_AGEMA_signal_7703), .Q (new_AGEMA_signal_7704) ) ;
    buf_clk new_AGEMA_reg_buffer_4247 ( .C (clk), .D (new_AGEMA_signal_7711), .Q (new_AGEMA_signal_7712) ) ;
    buf_clk new_AGEMA_reg_buffer_4255 ( .C (clk), .D (new_AGEMA_signal_7719), .Q (new_AGEMA_signal_7720) ) ;
    buf_clk new_AGEMA_reg_buffer_4263 ( .C (clk), .D (new_AGEMA_signal_7727), .Q (new_AGEMA_signal_7728) ) ;
    buf_clk new_AGEMA_reg_buffer_4271 ( .C (clk), .D (new_AGEMA_signal_7735), .Q (new_AGEMA_signal_7736) ) ;
    buf_clk new_AGEMA_reg_buffer_4279 ( .C (clk), .D (new_AGEMA_signal_7743), .Q (new_AGEMA_signal_7744) ) ;
    buf_clk new_AGEMA_reg_buffer_4287 ( .C (clk), .D (new_AGEMA_signal_7751), .Q (new_AGEMA_signal_7752) ) ;
    buf_clk new_AGEMA_reg_buffer_4295 ( .C (clk), .D (new_AGEMA_signal_7759), .Q (new_AGEMA_signal_7760) ) ;
    buf_clk new_AGEMA_reg_buffer_4303 ( .C (clk), .D (new_AGEMA_signal_7767), .Q (new_AGEMA_signal_7768) ) ;
    buf_clk new_AGEMA_reg_buffer_4311 ( .C (clk), .D (new_AGEMA_signal_7775), .Q (new_AGEMA_signal_7776) ) ;
    buf_clk new_AGEMA_reg_buffer_4319 ( .C (clk), .D (new_AGEMA_signal_7783), .Q (new_AGEMA_signal_7784) ) ;
    buf_clk new_AGEMA_reg_buffer_4327 ( .C (clk), .D (new_AGEMA_signal_7791), .Q (new_AGEMA_signal_7792) ) ;
    buf_clk new_AGEMA_reg_buffer_4335 ( .C (clk), .D (new_AGEMA_signal_7799), .Q (new_AGEMA_signal_7800) ) ;
    buf_clk new_AGEMA_reg_buffer_4343 ( .C (clk), .D (new_AGEMA_signal_7807), .Q (new_AGEMA_signal_7808) ) ;
    buf_clk new_AGEMA_reg_buffer_4351 ( .C (clk), .D (new_AGEMA_signal_7815), .Q (new_AGEMA_signal_7816) ) ;
    buf_clk new_AGEMA_reg_buffer_4359 ( .C (clk), .D (new_AGEMA_signal_7823), .Q (new_AGEMA_signal_7824) ) ;
    buf_clk new_AGEMA_reg_buffer_4367 ( .C (clk), .D (new_AGEMA_signal_7831), .Q (new_AGEMA_signal_7832) ) ;
    buf_clk new_AGEMA_reg_buffer_4375 ( .C (clk), .D (new_AGEMA_signal_7839), .Q (new_AGEMA_signal_7840) ) ;
    buf_clk new_AGEMA_reg_buffer_4383 ( .C (clk), .D (new_AGEMA_signal_7847), .Q (new_AGEMA_signal_7848) ) ;
    buf_clk new_AGEMA_reg_buffer_4391 ( .C (clk), .D (new_AGEMA_signal_7855), .Q (new_AGEMA_signal_7856) ) ;
    buf_clk new_AGEMA_reg_buffer_4399 ( .C (clk), .D (new_AGEMA_signal_7863), .Q (new_AGEMA_signal_7864) ) ;
    buf_clk new_AGEMA_reg_buffer_4407 ( .C (clk), .D (new_AGEMA_signal_7871), .Q (new_AGEMA_signal_7872) ) ;
    buf_clk new_AGEMA_reg_buffer_4415 ( .C (clk), .D (new_AGEMA_signal_7879), .Q (new_AGEMA_signal_7880) ) ;
    buf_clk new_AGEMA_reg_buffer_4423 ( .C (clk), .D (new_AGEMA_signal_7887), .Q (new_AGEMA_signal_7888) ) ;
    buf_clk new_AGEMA_reg_buffer_4431 ( .C (clk), .D (new_AGEMA_signal_7895), .Q (new_AGEMA_signal_7896) ) ;
    buf_clk new_AGEMA_reg_buffer_4439 ( .C (clk), .D (new_AGEMA_signal_7903), .Q (new_AGEMA_signal_7904) ) ;
    buf_clk new_AGEMA_reg_buffer_4447 ( .C (clk), .D (new_AGEMA_signal_7911), .Q (new_AGEMA_signal_7912) ) ;
    buf_clk new_AGEMA_reg_buffer_4455 ( .C (clk), .D (new_AGEMA_signal_7919), .Q (new_AGEMA_signal_7920) ) ;
    buf_clk new_AGEMA_reg_buffer_4463 ( .C (clk), .D (new_AGEMA_signal_7927), .Q (new_AGEMA_signal_7928) ) ;
    buf_clk new_AGEMA_reg_buffer_4471 ( .C (clk), .D (new_AGEMA_signal_7935), .Q (new_AGEMA_signal_7936) ) ;
    buf_clk new_AGEMA_reg_buffer_4479 ( .C (clk), .D (new_AGEMA_signal_7943), .Q (new_AGEMA_signal_7944) ) ;
    buf_clk new_AGEMA_reg_buffer_4487 ( .C (clk), .D (new_AGEMA_signal_7951), .Q (new_AGEMA_signal_7952) ) ;
    buf_clk new_AGEMA_reg_buffer_4495 ( .C (clk), .D (new_AGEMA_signal_7959), .Q (new_AGEMA_signal_7960) ) ;
    buf_clk new_AGEMA_reg_buffer_4503 ( .C (clk), .D (new_AGEMA_signal_7967), .Q (new_AGEMA_signal_7968) ) ;
    buf_clk new_AGEMA_reg_buffer_4511 ( .C (clk), .D (new_AGEMA_signal_7975), .Q (new_AGEMA_signal_7976) ) ;
    buf_clk new_AGEMA_reg_buffer_4519 ( .C (clk), .D (new_AGEMA_signal_7983), .Q (new_AGEMA_signal_7984) ) ;
    buf_clk new_AGEMA_reg_buffer_4527 ( .C (clk), .D (new_AGEMA_signal_7991), .Q (new_AGEMA_signal_7992) ) ;
    buf_clk new_AGEMA_reg_buffer_4535 ( .C (clk), .D (new_AGEMA_signal_7999), .Q (new_AGEMA_signal_8000) ) ;
    buf_clk new_AGEMA_reg_buffer_4543 ( .C (clk), .D (new_AGEMA_signal_8007), .Q (new_AGEMA_signal_8008) ) ;
    buf_clk new_AGEMA_reg_buffer_4551 ( .C (clk), .D (new_AGEMA_signal_8015), .Q (new_AGEMA_signal_8016) ) ;
    buf_clk new_AGEMA_reg_buffer_4559 ( .C (clk), .D (new_AGEMA_signal_8023), .Q (new_AGEMA_signal_8024) ) ;
    buf_clk new_AGEMA_reg_buffer_4567 ( .C (clk), .D (new_AGEMA_signal_8031), .Q (new_AGEMA_signal_8032) ) ;
    buf_clk new_AGEMA_reg_buffer_4575 ( .C (clk), .D (new_AGEMA_signal_8039), .Q (new_AGEMA_signal_8040) ) ;
    buf_clk new_AGEMA_reg_buffer_4583 ( .C (clk), .D (new_AGEMA_signal_8047), .Q (new_AGEMA_signal_8048) ) ;
    buf_clk new_AGEMA_reg_buffer_4591 ( .C (clk), .D (new_AGEMA_signal_8055), .Q (new_AGEMA_signal_8056) ) ;
    buf_clk new_AGEMA_reg_buffer_4599 ( .C (clk), .D (new_AGEMA_signal_8063), .Q (new_AGEMA_signal_8064) ) ;
    buf_clk new_AGEMA_reg_buffer_4607 ( .C (clk), .D (new_AGEMA_signal_8071), .Q (new_AGEMA_signal_8072) ) ;
    buf_clk new_AGEMA_reg_buffer_4615 ( .C (clk), .D (new_AGEMA_signal_8079), .Q (new_AGEMA_signal_8080) ) ;
    buf_clk new_AGEMA_reg_buffer_4623 ( .C (clk), .D (new_AGEMA_signal_8087), .Q (new_AGEMA_signal_8088) ) ;
    buf_clk new_AGEMA_reg_buffer_4631 ( .C (clk), .D (new_AGEMA_signal_8095), .Q (new_AGEMA_signal_8096) ) ;
    buf_clk new_AGEMA_reg_buffer_4639 ( .C (clk), .D (new_AGEMA_signal_8103), .Q (new_AGEMA_signal_8104) ) ;
    buf_clk new_AGEMA_reg_buffer_4647 ( .C (clk), .D (new_AGEMA_signal_8111), .Q (new_AGEMA_signal_8112) ) ;
    buf_clk new_AGEMA_reg_buffer_4655 ( .C (clk), .D (new_AGEMA_signal_8119), .Q (new_AGEMA_signal_8120) ) ;
    buf_clk new_AGEMA_reg_buffer_4663 ( .C (clk), .D (new_AGEMA_signal_8127), .Q (new_AGEMA_signal_8128) ) ;
    buf_clk new_AGEMA_reg_buffer_4671 ( .C (clk), .D (new_AGEMA_signal_8135), .Q (new_AGEMA_signal_8136) ) ;
    buf_clk new_AGEMA_reg_buffer_4679 ( .C (clk), .D (new_AGEMA_signal_8143), .Q (new_AGEMA_signal_8144) ) ;
    buf_clk new_AGEMA_reg_buffer_4687 ( .C (clk), .D (new_AGEMA_signal_8151), .Q (new_AGEMA_signal_8152) ) ;
    buf_clk new_AGEMA_reg_buffer_4695 ( .C (clk), .D (new_AGEMA_signal_8159), .Q (new_AGEMA_signal_8160) ) ;
    buf_clk new_AGEMA_reg_buffer_4703 ( .C (clk), .D (new_AGEMA_signal_8167), .Q (new_AGEMA_signal_8168) ) ;
    buf_clk new_AGEMA_reg_buffer_4711 ( .C (clk), .D (new_AGEMA_signal_8175), .Q (new_AGEMA_signal_8176) ) ;
    buf_clk new_AGEMA_reg_buffer_4719 ( .C (clk), .D (new_AGEMA_signal_8183), .Q (new_AGEMA_signal_8184) ) ;
    buf_clk new_AGEMA_reg_buffer_4727 ( .C (clk), .D (new_AGEMA_signal_8191), .Q (new_AGEMA_signal_8192) ) ;
    buf_clk new_AGEMA_reg_buffer_4735 ( .C (clk), .D (new_AGEMA_signal_8199), .Q (new_AGEMA_signal_8200) ) ;
    buf_clk new_AGEMA_reg_buffer_4743 ( .C (clk), .D (new_AGEMA_signal_8207), .Q (new_AGEMA_signal_8208) ) ;
    buf_clk new_AGEMA_reg_buffer_4751 ( .C (clk), .D (new_AGEMA_signal_8215), .Q (new_AGEMA_signal_8216) ) ;
    buf_clk new_AGEMA_reg_buffer_4759 ( .C (clk), .D (new_AGEMA_signal_8223), .Q (new_AGEMA_signal_8224) ) ;
    buf_clk new_AGEMA_reg_buffer_4767 ( .C (clk), .D (new_AGEMA_signal_8231), .Q (new_AGEMA_signal_8232) ) ;
    buf_clk new_AGEMA_reg_buffer_4775 ( .C (clk), .D (new_AGEMA_signal_8239), .Q (new_AGEMA_signal_8240) ) ;
    buf_clk new_AGEMA_reg_buffer_4783 ( .C (clk), .D (new_AGEMA_signal_8247), .Q (new_AGEMA_signal_8248) ) ;
    buf_clk new_AGEMA_reg_buffer_4791 ( .C (clk), .D (new_AGEMA_signal_8255), .Q (new_AGEMA_signal_8256) ) ;
    buf_clk new_AGEMA_reg_buffer_4799 ( .C (clk), .D (new_AGEMA_signal_8263), .Q (new_AGEMA_signal_8264) ) ;
    buf_clk new_AGEMA_reg_buffer_4807 ( .C (clk), .D (new_AGEMA_signal_8271), .Q (new_AGEMA_signal_8272) ) ;
    buf_clk new_AGEMA_reg_buffer_4815 ( .C (clk), .D (new_AGEMA_signal_8279), .Q (new_AGEMA_signal_8280) ) ;
    buf_clk new_AGEMA_reg_buffer_4823 ( .C (clk), .D (new_AGEMA_signal_8287), .Q (new_AGEMA_signal_8288) ) ;
    buf_clk new_AGEMA_reg_buffer_4831 ( .C (clk), .D (new_AGEMA_signal_8295), .Q (new_AGEMA_signal_8296) ) ;
    buf_clk new_AGEMA_reg_buffer_4839 ( .C (clk), .D (new_AGEMA_signal_8303), .Q (new_AGEMA_signal_8304) ) ;
    buf_clk new_AGEMA_reg_buffer_4847 ( .C (clk), .D (new_AGEMA_signal_8311), .Q (new_AGEMA_signal_8312) ) ;
    buf_clk new_AGEMA_reg_buffer_4855 ( .C (clk), .D (new_AGEMA_signal_8319), .Q (new_AGEMA_signal_8320) ) ;
    buf_clk new_AGEMA_reg_buffer_4863 ( .C (clk), .D (new_AGEMA_signal_8327), .Q (new_AGEMA_signal_8328) ) ;
    buf_clk new_AGEMA_reg_buffer_4871 ( .C (clk), .D (new_AGEMA_signal_8335), .Q (new_AGEMA_signal_8336) ) ;
    buf_clk new_AGEMA_reg_buffer_4879 ( .C (clk), .D (new_AGEMA_signal_8343), .Q (new_AGEMA_signal_8344) ) ;
    buf_clk new_AGEMA_reg_buffer_4887 ( .C (clk), .D (new_AGEMA_signal_8351), .Q (new_AGEMA_signal_8352) ) ;
    buf_clk new_AGEMA_reg_buffer_4895 ( .C (clk), .D (new_AGEMA_signal_8359), .Q (new_AGEMA_signal_8360) ) ;
    buf_clk new_AGEMA_reg_buffer_4903 ( .C (clk), .D (new_AGEMA_signal_8367), .Q (new_AGEMA_signal_8368) ) ;
    buf_clk new_AGEMA_reg_buffer_4911 ( .C (clk), .D (new_AGEMA_signal_8375), .Q (new_AGEMA_signal_8376) ) ;
    buf_clk new_AGEMA_reg_buffer_4919 ( .C (clk), .D (new_AGEMA_signal_8383), .Q (new_AGEMA_signal_8384) ) ;
    buf_clk new_AGEMA_reg_buffer_4927 ( .C (clk), .D (new_AGEMA_signal_8391), .Q (new_AGEMA_signal_8392) ) ;
    buf_clk new_AGEMA_reg_buffer_4935 ( .C (clk), .D (new_AGEMA_signal_8399), .Q (new_AGEMA_signal_8400) ) ;
    buf_clk new_AGEMA_reg_buffer_4943 ( .C (clk), .D (new_AGEMA_signal_8407), .Q (new_AGEMA_signal_8408) ) ;
    buf_clk new_AGEMA_reg_buffer_4951 ( .C (clk), .D (new_AGEMA_signal_8415), .Q (new_AGEMA_signal_8416) ) ;
    buf_clk new_AGEMA_reg_buffer_4959 ( .C (clk), .D (new_AGEMA_signal_8423), .Q (new_AGEMA_signal_8424) ) ;
    buf_clk new_AGEMA_reg_buffer_4967 ( .C (clk), .D (new_AGEMA_signal_8431), .Q (new_AGEMA_signal_8432) ) ;
    buf_clk new_AGEMA_reg_buffer_4975 ( .C (clk), .D (new_AGEMA_signal_8439), .Q (new_AGEMA_signal_8440) ) ;
    buf_clk new_AGEMA_reg_buffer_4983 ( .C (clk), .D (new_AGEMA_signal_8447), .Q (new_AGEMA_signal_8448) ) ;
    buf_clk new_AGEMA_reg_buffer_4991 ( .C (clk), .D (new_AGEMA_signal_8455), .Q (new_AGEMA_signal_8456) ) ;
    buf_clk new_AGEMA_reg_buffer_4999 ( .C (clk), .D (new_AGEMA_signal_8463), .Q (new_AGEMA_signal_8464) ) ;
    buf_clk new_AGEMA_reg_buffer_5007 ( .C (clk), .D (new_AGEMA_signal_8471), .Q (new_AGEMA_signal_8472) ) ;
    buf_clk new_AGEMA_reg_buffer_5015 ( .C (clk), .D (new_AGEMA_signal_8479), .Q (new_AGEMA_signal_8480) ) ;
    buf_clk new_AGEMA_reg_buffer_5023 ( .C (clk), .D (new_AGEMA_signal_8487), .Q (new_AGEMA_signal_8488) ) ;
    buf_clk new_AGEMA_reg_buffer_5031 ( .C (clk), .D (new_AGEMA_signal_8495), .Q (new_AGEMA_signal_8496) ) ;
    buf_clk new_AGEMA_reg_buffer_5039 ( .C (clk), .D (new_AGEMA_signal_8503), .Q (new_AGEMA_signal_8504) ) ;
    buf_clk new_AGEMA_reg_buffer_5047 ( .C (clk), .D (new_AGEMA_signal_8511), .Q (new_AGEMA_signal_8512) ) ;
    buf_clk new_AGEMA_reg_buffer_5055 ( .C (clk), .D (new_AGEMA_signal_8519), .Q (new_AGEMA_signal_8520) ) ;
    buf_clk new_AGEMA_reg_buffer_5063 ( .C (clk), .D (new_AGEMA_signal_8527), .Q (new_AGEMA_signal_8528) ) ;
    buf_clk new_AGEMA_reg_buffer_5071 ( .C (clk), .D (new_AGEMA_signal_8535), .Q (new_AGEMA_signal_8536) ) ;
    buf_clk new_AGEMA_reg_buffer_5079 ( .C (clk), .D (new_AGEMA_signal_8543), .Q (new_AGEMA_signal_8544) ) ;
    buf_clk new_AGEMA_reg_buffer_5087 ( .C (clk), .D (new_AGEMA_signal_8551), .Q (new_AGEMA_signal_8552) ) ;
    buf_clk new_AGEMA_reg_buffer_5095 ( .C (clk), .D (new_AGEMA_signal_8559), .Q (new_AGEMA_signal_8560) ) ;
    buf_clk new_AGEMA_reg_buffer_5103 ( .C (clk), .D (new_AGEMA_signal_8567), .Q (new_AGEMA_signal_8568) ) ;
    buf_clk new_AGEMA_reg_buffer_5111 ( .C (clk), .D (new_AGEMA_signal_8575), .Q (new_AGEMA_signal_8576) ) ;
    buf_clk new_AGEMA_reg_buffer_5119 ( .C (clk), .D (new_AGEMA_signal_8583), .Q (new_AGEMA_signal_8584) ) ;
    buf_clk new_AGEMA_reg_buffer_5127 ( .C (clk), .D (new_AGEMA_signal_8591), .Q (new_AGEMA_signal_8592) ) ;
    buf_clk new_AGEMA_reg_buffer_5135 ( .C (clk), .D (new_AGEMA_signal_8599), .Q (new_AGEMA_signal_8600) ) ;
    buf_clk new_AGEMA_reg_buffer_5143 ( .C (clk), .D (new_AGEMA_signal_8607), .Q (new_AGEMA_signal_8608) ) ;
    buf_clk new_AGEMA_reg_buffer_5151 ( .C (clk), .D (new_AGEMA_signal_8615), .Q (new_AGEMA_signal_8616) ) ;
    buf_clk new_AGEMA_reg_buffer_5159 ( .C (clk), .D (new_AGEMA_signal_8623), .Q (new_AGEMA_signal_8624) ) ;
    buf_clk new_AGEMA_reg_buffer_5167 ( .C (clk), .D (new_AGEMA_signal_8631), .Q (new_AGEMA_signal_8632) ) ;
    buf_clk new_AGEMA_reg_buffer_5175 ( .C (clk), .D (new_AGEMA_signal_8639), .Q (new_AGEMA_signal_8640) ) ;
    buf_clk new_AGEMA_reg_buffer_5183 ( .C (clk), .D (new_AGEMA_signal_8647), .Q (new_AGEMA_signal_8648) ) ;
    buf_clk new_AGEMA_reg_buffer_5191 ( .C (clk), .D (new_AGEMA_signal_8655), .Q (new_AGEMA_signal_8656) ) ;
    buf_clk new_AGEMA_reg_buffer_5199 ( .C (clk), .D (new_AGEMA_signal_8663), .Q (new_AGEMA_signal_8664) ) ;
    buf_clk new_AGEMA_reg_buffer_5207 ( .C (clk), .D (new_AGEMA_signal_8671), .Q (new_AGEMA_signal_8672) ) ;
    buf_clk new_AGEMA_reg_buffer_5215 ( .C (clk), .D (new_AGEMA_signal_8679), .Q (new_AGEMA_signal_8680) ) ;
    buf_clk new_AGEMA_reg_buffer_5223 ( .C (clk), .D (new_AGEMA_signal_8687), .Q (new_AGEMA_signal_8688) ) ;
    buf_clk new_AGEMA_reg_buffer_5231 ( .C (clk), .D (new_AGEMA_signal_8695), .Q (new_AGEMA_signal_8696) ) ;
    buf_clk new_AGEMA_reg_buffer_5239 ( .C (clk), .D (new_AGEMA_signal_8703), .Q (new_AGEMA_signal_8704) ) ;
    buf_clk new_AGEMA_reg_buffer_5247 ( .C (clk), .D (new_AGEMA_signal_8711), .Q (new_AGEMA_signal_8712) ) ;
    buf_clk new_AGEMA_reg_buffer_5255 ( .C (clk), .D (new_AGEMA_signal_8719), .Q (new_AGEMA_signal_8720) ) ;
    buf_clk new_AGEMA_reg_buffer_5263 ( .C (clk), .D (new_AGEMA_signal_8727), .Q (new_AGEMA_signal_8728) ) ;
    buf_clk new_AGEMA_reg_buffer_5271 ( .C (clk), .D (new_AGEMA_signal_8735), .Q (new_AGEMA_signal_8736) ) ;
    buf_clk new_AGEMA_reg_buffer_5279 ( .C (clk), .D (new_AGEMA_signal_8743), .Q (new_AGEMA_signal_8744) ) ;
    buf_clk new_AGEMA_reg_buffer_5287 ( .C (clk), .D (new_AGEMA_signal_8751), .Q (new_AGEMA_signal_8752) ) ;
    buf_clk new_AGEMA_reg_buffer_5295 ( .C (clk), .D (new_AGEMA_signal_8759), .Q (new_AGEMA_signal_8760) ) ;
    buf_clk new_AGEMA_reg_buffer_5303 ( .C (clk), .D (new_AGEMA_signal_8767), .Q (new_AGEMA_signal_8768) ) ;
    buf_clk new_AGEMA_reg_buffer_5311 ( .C (clk), .D (new_AGEMA_signal_8775), .Q (new_AGEMA_signal_8776) ) ;
    buf_clk new_AGEMA_reg_buffer_5319 ( .C (clk), .D (new_AGEMA_signal_8783), .Q (new_AGEMA_signal_8784) ) ;
    buf_clk new_AGEMA_reg_buffer_5327 ( .C (clk), .D (new_AGEMA_signal_8791), .Q (new_AGEMA_signal_8792) ) ;
    buf_clk new_AGEMA_reg_buffer_5335 ( .C (clk), .D (new_AGEMA_signal_8799), .Q (new_AGEMA_signal_8800) ) ;
    buf_clk new_AGEMA_reg_buffer_5343 ( .C (clk), .D (new_AGEMA_signal_8807), .Q (new_AGEMA_signal_8808) ) ;
    buf_clk new_AGEMA_reg_buffer_5351 ( .C (clk), .D (new_AGEMA_signal_8815), .Q (new_AGEMA_signal_8816) ) ;
    buf_clk new_AGEMA_reg_buffer_5359 ( .C (clk), .D (new_AGEMA_signal_8823), .Q (new_AGEMA_signal_8824) ) ;
    buf_clk new_AGEMA_reg_buffer_5367 ( .C (clk), .D (new_AGEMA_signal_8831), .Q (new_AGEMA_signal_8832) ) ;
    buf_clk new_AGEMA_reg_buffer_5375 ( .C (clk), .D (new_AGEMA_signal_8839), .Q (new_AGEMA_signal_8840) ) ;
    buf_clk new_AGEMA_reg_buffer_5383 ( .C (clk), .D (new_AGEMA_signal_8847), .Q (new_AGEMA_signal_8848) ) ;
    buf_clk new_AGEMA_reg_buffer_5391 ( .C (clk), .D (new_AGEMA_signal_8855), .Q (new_AGEMA_signal_8856) ) ;
    buf_clk new_AGEMA_reg_buffer_5399 ( .C (clk), .D (new_AGEMA_signal_8863), .Q (new_AGEMA_signal_8864) ) ;
    buf_clk new_AGEMA_reg_buffer_5409 ( .C (clk), .D (new_AGEMA_signal_8873), .Q (new_AGEMA_signal_8874) ) ;
    buf_clk new_AGEMA_reg_buffer_5417 ( .C (clk), .D (new_AGEMA_signal_8881), .Q (new_AGEMA_signal_8882) ) ;
    buf_clk new_AGEMA_reg_buffer_5425 ( .C (clk), .D (new_AGEMA_signal_8889), .Q (new_AGEMA_signal_8890) ) ;
    buf_clk new_AGEMA_reg_buffer_5433 ( .C (clk), .D (new_AGEMA_signal_8897), .Q (new_AGEMA_signal_8898) ) ;
    buf_clk new_AGEMA_reg_buffer_5441 ( .C (clk), .D (new_AGEMA_signal_8905), .Q (new_AGEMA_signal_8906) ) ;
    buf_clk new_AGEMA_reg_buffer_5449 ( .C (clk), .D (new_AGEMA_signal_8913), .Q (new_AGEMA_signal_8914) ) ;
    buf_clk new_AGEMA_reg_buffer_5457 ( .C (clk), .D (new_AGEMA_signal_8921), .Q (new_AGEMA_signal_8922) ) ;
    buf_clk new_AGEMA_reg_buffer_5465 ( .C (clk), .D (new_AGEMA_signal_8929), .Q (new_AGEMA_signal_8930) ) ;
    buf_clk new_AGEMA_reg_buffer_5473 ( .C (clk), .D (new_AGEMA_signal_8937), .Q (new_AGEMA_signal_8938) ) ;
    buf_clk new_AGEMA_reg_buffer_5481 ( .C (clk), .D (new_AGEMA_signal_8945), .Q (new_AGEMA_signal_8946) ) ;
    buf_clk new_AGEMA_reg_buffer_5489 ( .C (clk), .D (new_AGEMA_signal_8953), .Q (new_AGEMA_signal_8954) ) ;
    buf_clk new_AGEMA_reg_buffer_5497 ( .C (clk), .D (new_AGEMA_signal_8961), .Q (new_AGEMA_signal_8962) ) ;
    buf_clk new_AGEMA_reg_buffer_5505 ( .C (clk), .D (new_AGEMA_signal_8969), .Q (new_AGEMA_signal_8970) ) ;
    buf_clk new_AGEMA_reg_buffer_5513 ( .C (clk), .D (new_AGEMA_signal_8977), .Q (new_AGEMA_signal_8978) ) ;
    buf_clk new_AGEMA_reg_buffer_5521 ( .C (clk), .D (new_AGEMA_signal_8985), .Q (new_AGEMA_signal_8986) ) ;
    buf_clk new_AGEMA_reg_buffer_5529 ( .C (clk), .D (new_AGEMA_signal_8993), .Q (new_AGEMA_signal_8994) ) ;
    buf_clk new_AGEMA_reg_buffer_5537 ( .C (clk), .D (new_AGEMA_signal_9001), .Q (new_AGEMA_signal_9002) ) ;
    buf_clk new_AGEMA_reg_buffer_5545 ( .C (clk), .D (new_AGEMA_signal_9009), .Q (new_AGEMA_signal_9010) ) ;
    buf_clk new_AGEMA_reg_buffer_5553 ( .C (clk), .D (new_AGEMA_signal_9017), .Q (new_AGEMA_signal_9018) ) ;
    buf_clk new_AGEMA_reg_buffer_5561 ( .C (clk), .D (new_AGEMA_signal_9025), .Q (new_AGEMA_signal_9026) ) ;
    buf_clk new_AGEMA_reg_buffer_5569 ( .C (clk), .D (new_AGEMA_signal_9033), .Q (new_AGEMA_signal_9034) ) ;
    buf_clk new_AGEMA_reg_buffer_5577 ( .C (clk), .D (new_AGEMA_signal_9041), .Q (new_AGEMA_signal_9042) ) ;
    buf_clk new_AGEMA_reg_buffer_5585 ( .C (clk), .D (new_AGEMA_signal_9049), .Q (new_AGEMA_signal_9050) ) ;
    buf_clk new_AGEMA_reg_buffer_5593 ( .C (clk), .D (new_AGEMA_signal_9057), .Q (new_AGEMA_signal_9058) ) ;
    buf_clk new_AGEMA_reg_buffer_5601 ( .C (clk), .D (new_AGEMA_signal_9065), .Q (new_AGEMA_signal_9066) ) ;
    buf_clk new_AGEMA_reg_buffer_5609 ( .C (clk), .D (new_AGEMA_signal_9073), .Q (new_AGEMA_signal_9074) ) ;
    buf_clk new_AGEMA_reg_buffer_5617 ( .C (clk), .D (new_AGEMA_signal_9081), .Q (new_AGEMA_signal_9082) ) ;
    buf_clk new_AGEMA_reg_buffer_5625 ( .C (clk), .D (new_AGEMA_signal_9089), .Q (new_AGEMA_signal_9090) ) ;
    buf_clk new_AGEMA_reg_buffer_5633 ( .C (clk), .D (new_AGEMA_signal_9097), .Q (new_AGEMA_signal_9098) ) ;
    buf_clk new_AGEMA_reg_buffer_5641 ( .C (clk), .D (new_AGEMA_signal_9105), .Q (new_AGEMA_signal_9106) ) ;
    buf_clk new_AGEMA_reg_buffer_5649 ( .C (clk), .D (new_AGEMA_signal_9113), .Q (new_AGEMA_signal_9114) ) ;
    buf_clk new_AGEMA_reg_buffer_5657 ( .C (clk), .D (new_AGEMA_signal_9121), .Q (new_AGEMA_signal_9122) ) ;
    buf_clk new_AGEMA_reg_buffer_5665 ( .C (clk), .D (new_AGEMA_signal_9129), .Q (new_AGEMA_signal_9130) ) ;
    buf_clk new_AGEMA_reg_buffer_5673 ( .C (clk), .D (new_AGEMA_signal_9137), .Q (new_AGEMA_signal_9138) ) ;
    buf_clk new_AGEMA_reg_buffer_5681 ( .C (clk), .D (new_AGEMA_signal_9145), .Q (new_AGEMA_signal_9146) ) ;
    buf_clk new_AGEMA_reg_buffer_5689 ( .C (clk), .D (new_AGEMA_signal_9153), .Q (new_AGEMA_signal_9154) ) ;
    buf_clk new_AGEMA_reg_buffer_5697 ( .C (clk), .D (new_AGEMA_signal_9161), .Q (new_AGEMA_signal_9162) ) ;
    buf_clk new_AGEMA_reg_buffer_5705 ( .C (clk), .D (new_AGEMA_signal_9169), .Q (new_AGEMA_signal_9170) ) ;
    buf_clk new_AGEMA_reg_buffer_5713 ( .C (clk), .D (new_AGEMA_signal_9177), .Q (new_AGEMA_signal_9178) ) ;
    buf_clk new_AGEMA_reg_buffer_5721 ( .C (clk), .D (new_AGEMA_signal_9185), .Q (new_AGEMA_signal_9186) ) ;
    buf_clk new_AGEMA_reg_buffer_5729 ( .C (clk), .D (new_AGEMA_signal_9193), .Q (new_AGEMA_signal_9194) ) ;
    buf_clk new_AGEMA_reg_buffer_5737 ( .C (clk), .D (new_AGEMA_signal_9201), .Q (new_AGEMA_signal_9202) ) ;
    buf_clk new_AGEMA_reg_buffer_5745 ( .C (clk), .D (new_AGEMA_signal_9209), .Q (new_AGEMA_signal_9210) ) ;
    buf_clk new_AGEMA_reg_buffer_5753 ( .C (clk), .D (new_AGEMA_signal_9217), .Q (new_AGEMA_signal_9218) ) ;
    buf_clk new_AGEMA_reg_buffer_5761 ( .C (clk), .D (new_AGEMA_signal_9225), .Q (new_AGEMA_signal_9226) ) ;
    buf_clk new_AGEMA_reg_buffer_5769 ( .C (clk), .D (new_AGEMA_signal_9233), .Q (new_AGEMA_signal_9234) ) ;
    buf_clk new_AGEMA_reg_buffer_5777 ( .C (clk), .D (new_AGEMA_signal_9241), .Q (new_AGEMA_signal_9242) ) ;
    buf_clk new_AGEMA_reg_buffer_5785 ( .C (clk), .D (new_AGEMA_signal_9249), .Q (new_AGEMA_signal_9250) ) ;
    buf_clk new_AGEMA_reg_buffer_5793 ( .C (clk), .D (new_AGEMA_signal_9257), .Q (new_AGEMA_signal_9258) ) ;
    buf_clk new_AGEMA_reg_buffer_5801 ( .C (clk), .D (new_AGEMA_signal_9265), .Q (new_AGEMA_signal_9266) ) ;
    buf_clk new_AGEMA_reg_buffer_5809 ( .C (clk), .D (new_AGEMA_signal_9273), .Q (new_AGEMA_signal_9274) ) ;
    buf_clk new_AGEMA_reg_buffer_5817 ( .C (clk), .D (new_AGEMA_signal_9281), .Q (new_AGEMA_signal_9282) ) ;
    buf_clk new_AGEMA_reg_buffer_5825 ( .C (clk), .D (new_AGEMA_signal_9289), .Q (new_AGEMA_signal_9290) ) ;
    buf_clk new_AGEMA_reg_buffer_5833 ( .C (clk), .D (new_AGEMA_signal_9297), .Q (new_AGEMA_signal_9298) ) ;
    buf_clk new_AGEMA_reg_buffer_5841 ( .C (clk), .D (new_AGEMA_signal_9305), .Q (new_AGEMA_signal_9306) ) ;
    buf_clk new_AGEMA_reg_buffer_5849 ( .C (clk), .D (new_AGEMA_signal_9313), .Q (new_AGEMA_signal_9314) ) ;
    buf_clk new_AGEMA_reg_buffer_5857 ( .C (clk), .D (new_AGEMA_signal_9321), .Q (new_AGEMA_signal_9322) ) ;
    buf_clk new_AGEMA_reg_buffer_5865 ( .C (clk), .D (new_AGEMA_signal_9329), .Q (new_AGEMA_signal_9330) ) ;
    buf_clk new_AGEMA_reg_buffer_5873 ( .C (clk), .D (new_AGEMA_signal_9337), .Q (new_AGEMA_signal_9338) ) ;
    buf_clk new_AGEMA_reg_buffer_5881 ( .C (clk), .D (new_AGEMA_signal_9345), .Q (new_AGEMA_signal_9346) ) ;
    buf_clk new_AGEMA_reg_buffer_5889 ( .C (clk), .D (new_AGEMA_signal_9353), .Q (new_AGEMA_signal_9354) ) ;
    buf_clk new_AGEMA_reg_buffer_5897 ( .C (clk), .D (new_AGEMA_signal_9361), .Q (new_AGEMA_signal_9362) ) ;
    buf_clk new_AGEMA_reg_buffer_5905 ( .C (clk), .D (new_AGEMA_signal_9369), .Q (new_AGEMA_signal_9370) ) ;
    buf_clk new_AGEMA_reg_buffer_5913 ( .C (clk), .D (new_AGEMA_signal_9377), .Q (new_AGEMA_signal_9378) ) ;
    buf_clk new_AGEMA_reg_buffer_5921 ( .C (clk), .D (new_AGEMA_signal_9385), .Q (new_AGEMA_signal_9386) ) ;
    buf_clk new_AGEMA_reg_buffer_5929 ( .C (clk), .D (new_AGEMA_signal_9393), .Q (new_AGEMA_signal_9394) ) ;
    buf_clk new_AGEMA_reg_buffer_5937 ( .C (clk), .D (new_AGEMA_signal_9401), .Q (new_AGEMA_signal_9402) ) ;
    buf_clk new_AGEMA_reg_buffer_5945 ( .C (clk), .D (new_AGEMA_signal_9409), .Q (new_AGEMA_signal_9410) ) ;
    buf_clk new_AGEMA_reg_buffer_5953 ( .C (clk), .D (new_AGEMA_signal_9417), .Q (new_AGEMA_signal_9418) ) ;
    buf_clk new_AGEMA_reg_buffer_5961 ( .C (clk), .D (new_AGEMA_signal_9425), .Q (new_AGEMA_signal_9426) ) ;
    buf_clk new_AGEMA_reg_buffer_5969 ( .C (clk), .D (new_AGEMA_signal_9433), .Q (new_AGEMA_signal_9434) ) ;
    buf_clk new_AGEMA_reg_buffer_5977 ( .C (clk), .D (new_AGEMA_signal_9441), .Q (new_AGEMA_signal_9442) ) ;
    buf_clk new_AGEMA_reg_buffer_5985 ( .C (clk), .D (new_AGEMA_signal_9449), .Q (new_AGEMA_signal_9450) ) ;
    buf_clk new_AGEMA_reg_buffer_5993 ( .C (clk), .D (new_AGEMA_signal_9457), .Q (new_AGEMA_signal_9458) ) ;
    buf_clk new_AGEMA_reg_buffer_6001 ( .C (clk), .D (new_AGEMA_signal_9465), .Q (new_AGEMA_signal_9466) ) ;
    buf_clk new_AGEMA_reg_buffer_6009 ( .C (clk), .D (new_AGEMA_signal_9473), .Q (new_AGEMA_signal_9474) ) ;
    buf_clk new_AGEMA_reg_buffer_6017 ( .C (clk), .D (new_AGEMA_signal_9481), .Q (new_AGEMA_signal_9482) ) ;
    buf_clk new_AGEMA_reg_buffer_6025 ( .C (clk), .D (new_AGEMA_signal_9489), .Q (new_AGEMA_signal_9490) ) ;
    buf_clk new_AGEMA_reg_buffer_6033 ( .C (clk), .D (new_AGEMA_signal_9497), .Q (new_AGEMA_signal_9498) ) ;
    buf_clk new_AGEMA_reg_buffer_6041 ( .C (clk), .D (new_AGEMA_signal_9505), .Q (new_AGEMA_signal_9506) ) ;
    buf_clk new_AGEMA_reg_buffer_6049 ( .C (clk), .D (new_AGEMA_signal_9513), .Q (new_AGEMA_signal_9514) ) ;
    buf_clk new_AGEMA_reg_buffer_6057 ( .C (clk), .D (new_AGEMA_signal_9521), .Q (new_AGEMA_signal_9522) ) ;
    buf_clk new_AGEMA_reg_buffer_6065 ( .C (clk), .D (new_AGEMA_signal_9529), .Q (new_AGEMA_signal_9530) ) ;
    buf_clk new_AGEMA_reg_buffer_6073 ( .C (clk), .D (new_AGEMA_signal_9537), .Q (new_AGEMA_signal_9538) ) ;
    buf_clk new_AGEMA_reg_buffer_6081 ( .C (clk), .D (new_AGEMA_signal_9545), .Q (new_AGEMA_signal_9546) ) ;
    buf_clk new_AGEMA_reg_buffer_6089 ( .C (clk), .D (new_AGEMA_signal_9553), .Q (new_AGEMA_signal_9554) ) ;
    buf_clk new_AGEMA_reg_buffer_6097 ( .C (clk), .D (new_AGEMA_signal_9561), .Q (new_AGEMA_signal_9562) ) ;
    buf_clk new_AGEMA_reg_buffer_6105 ( .C (clk), .D (new_AGEMA_signal_9569), .Q (new_AGEMA_signal_9570) ) ;
    buf_clk new_AGEMA_reg_buffer_6113 ( .C (clk), .D (new_AGEMA_signal_9577), .Q (new_AGEMA_signal_9578) ) ;
    buf_clk new_AGEMA_reg_buffer_6121 ( .C (clk), .D (new_AGEMA_signal_9585), .Q (new_AGEMA_signal_9586) ) ;
    buf_clk new_AGEMA_reg_buffer_6129 ( .C (clk), .D (new_AGEMA_signal_9593), .Q (new_AGEMA_signal_9594) ) ;
    buf_clk new_AGEMA_reg_buffer_6137 ( .C (clk), .D (new_AGEMA_signal_9601), .Q (new_AGEMA_signal_9602) ) ;
    buf_clk new_AGEMA_reg_buffer_6145 ( .C (clk), .D (new_AGEMA_signal_9609), .Q (new_AGEMA_signal_9610) ) ;
    buf_clk new_AGEMA_reg_buffer_6153 ( .C (clk), .D (new_AGEMA_signal_9617), .Q (new_AGEMA_signal_9618) ) ;
    buf_clk new_AGEMA_reg_buffer_6161 ( .C (clk), .D (new_AGEMA_signal_9625), .Q (new_AGEMA_signal_9626) ) ;
    buf_clk new_AGEMA_reg_buffer_6169 ( .C (clk), .D (new_AGEMA_signal_9633), .Q (new_AGEMA_signal_9634) ) ;
    buf_clk new_AGEMA_reg_buffer_6173 ( .C (clk), .D (new_AGEMA_signal_7039), .Q (new_AGEMA_signal_9638) ) ;
    buf_clk new_AGEMA_reg_buffer_6175 ( .C (clk), .D (new_AGEMA_signal_7041), .Q (new_AGEMA_signal_9640) ) ;
    buf_clk new_AGEMA_reg_buffer_6177 ( .C (clk), .D (new_AGEMA_signal_7043), .Q (new_AGEMA_signal_9642) ) ;
    buf_clk new_AGEMA_reg_buffer_6181 ( .C (clk), .D (new_AGEMA_signal_9645), .Q (new_AGEMA_signal_9646) ) ;
    buf_clk new_AGEMA_reg_buffer_6185 ( .C (clk), .D (new_AGEMA_signal_9649), .Q (new_AGEMA_signal_9650) ) ;
    buf_clk new_AGEMA_reg_buffer_6189 ( .C (clk), .D (new_AGEMA_signal_9653), .Q (new_AGEMA_signal_9654) ) ;
    buf_clk new_AGEMA_reg_buffer_6191 ( .C (clk), .D (new_AGEMA_signal_7057), .Q (new_AGEMA_signal_9656) ) ;
    buf_clk new_AGEMA_reg_buffer_6193 ( .C (clk), .D (new_AGEMA_signal_7059), .Q (new_AGEMA_signal_9658) ) ;
    buf_clk new_AGEMA_reg_buffer_6195 ( .C (clk), .D (new_AGEMA_signal_7061), .Q (new_AGEMA_signal_9660) ) ;
    buf_clk new_AGEMA_reg_buffer_6199 ( .C (clk), .D (new_AGEMA_signal_9663), .Q (new_AGEMA_signal_9664) ) ;
    buf_clk new_AGEMA_reg_buffer_6203 ( .C (clk), .D (new_AGEMA_signal_9667), .Q (new_AGEMA_signal_9668) ) ;
    buf_clk new_AGEMA_reg_buffer_6207 ( .C (clk), .D (new_AGEMA_signal_9671), .Q (new_AGEMA_signal_9672) ) ;
    buf_clk new_AGEMA_reg_buffer_6209 ( .C (clk), .D (new_AGEMA_signal_7075), .Q (new_AGEMA_signal_9674) ) ;
    buf_clk new_AGEMA_reg_buffer_6211 ( .C (clk), .D (new_AGEMA_signal_7077), .Q (new_AGEMA_signal_9676) ) ;
    buf_clk new_AGEMA_reg_buffer_6213 ( .C (clk), .D (new_AGEMA_signal_7079), .Q (new_AGEMA_signal_9678) ) ;
    buf_clk new_AGEMA_reg_buffer_6217 ( .C (clk), .D (new_AGEMA_signal_9681), .Q (new_AGEMA_signal_9682) ) ;
    buf_clk new_AGEMA_reg_buffer_6221 ( .C (clk), .D (new_AGEMA_signal_9685), .Q (new_AGEMA_signal_9686) ) ;
    buf_clk new_AGEMA_reg_buffer_6225 ( .C (clk), .D (new_AGEMA_signal_9689), .Q (new_AGEMA_signal_9690) ) ;
    buf_clk new_AGEMA_reg_buffer_6227 ( .C (clk), .D (new_AGEMA_signal_7093), .Q (new_AGEMA_signal_9692) ) ;
    buf_clk new_AGEMA_reg_buffer_6229 ( .C (clk), .D (new_AGEMA_signal_7095), .Q (new_AGEMA_signal_9694) ) ;
    buf_clk new_AGEMA_reg_buffer_6231 ( .C (clk), .D (new_AGEMA_signal_7097), .Q (new_AGEMA_signal_9696) ) ;
    buf_clk new_AGEMA_reg_buffer_6235 ( .C (clk), .D (new_AGEMA_signal_9699), .Q (new_AGEMA_signal_9700) ) ;
    buf_clk new_AGEMA_reg_buffer_6239 ( .C (clk), .D (new_AGEMA_signal_9703), .Q (new_AGEMA_signal_9704) ) ;
    buf_clk new_AGEMA_reg_buffer_6243 ( .C (clk), .D (new_AGEMA_signal_9707), .Q (new_AGEMA_signal_9708) ) ;
    buf_clk new_AGEMA_reg_buffer_6245 ( .C (clk), .D (new_AGEMA_signal_7111), .Q (new_AGEMA_signal_9710) ) ;
    buf_clk new_AGEMA_reg_buffer_6247 ( .C (clk), .D (new_AGEMA_signal_7113), .Q (new_AGEMA_signal_9712) ) ;
    buf_clk new_AGEMA_reg_buffer_6249 ( .C (clk), .D (new_AGEMA_signal_7115), .Q (new_AGEMA_signal_9714) ) ;
    buf_clk new_AGEMA_reg_buffer_6253 ( .C (clk), .D (new_AGEMA_signal_9717), .Q (new_AGEMA_signal_9718) ) ;
    buf_clk new_AGEMA_reg_buffer_6257 ( .C (clk), .D (new_AGEMA_signal_9721), .Q (new_AGEMA_signal_9722) ) ;
    buf_clk new_AGEMA_reg_buffer_6261 ( .C (clk), .D (new_AGEMA_signal_9725), .Q (new_AGEMA_signal_9726) ) ;
    buf_clk new_AGEMA_reg_buffer_6263 ( .C (clk), .D (new_AGEMA_signal_7129), .Q (new_AGEMA_signal_9728) ) ;
    buf_clk new_AGEMA_reg_buffer_6265 ( .C (clk), .D (new_AGEMA_signal_7131), .Q (new_AGEMA_signal_9730) ) ;
    buf_clk new_AGEMA_reg_buffer_6267 ( .C (clk), .D (new_AGEMA_signal_7133), .Q (new_AGEMA_signal_9732) ) ;
    buf_clk new_AGEMA_reg_buffer_6271 ( .C (clk), .D (new_AGEMA_signal_9735), .Q (new_AGEMA_signal_9736) ) ;
    buf_clk new_AGEMA_reg_buffer_6275 ( .C (clk), .D (new_AGEMA_signal_9739), .Q (new_AGEMA_signal_9740) ) ;
    buf_clk new_AGEMA_reg_buffer_6279 ( .C (clk), .D (new_AGEMA_signal_9743), .Q (new_AGEMA_signal_9744) ) ;
    buf_clk new_AGEMA_reg_buffer_6281 ( .C (clk), .D (new_AGEMA_signal_7147), .Q (new_AGEMA_signal_9746) ) ;
    buf_clk new_AGEMA_reg_buffer_6283 ( .C (clk), .D (new_AGEMA_signal_7149), .Q (new_AGEMA_signal_9748) ) ;
    buf_clk new_AGEMA_reg_buffer_6285 ( .C (clk), .D (new_AGEMA_signal_7151), .Q (new_AGEMA_signal_9750) ) ;
    buf_clk new_AGEMA_reg_buffer_6289 ( .C (clk), .D (new_AGEMA_signal_9753), .Q (new_AGEMA_signal_9754) ) ;
    buf_clk new_AGEMA_reg_buffer_6293 ( .C (clk), .D (new_AGEMA_signal_9757), .Q (new_AGEMA_signal_9758) ) ;
    buf_clk new_AGEMA_reg_buffer_6297 ( .C (clk), .D (new_AGEMA_signal_9761), .Q (new_AGEMA_signal_9762) ) ;
    buf_clk new_AGEMA_reg_buffer_6299 ( .C (clk), .D (new_AGEMA_signal_7165), .Q (new_AGEMA_signal_9764) ) ;
    buf_clk new_AGEMA_reg_buffer_6301 ( .C (clk), .D (new_AGEMA_signal_7167), .Q (new_AGEMA_signal_9766) ) ;
    buf_clk new_AGEMA_reg_buffer_6303 ( .C (clk), .D (new_AGEMA_signal_7169), .Q (new_AGEMA_signal_9768) ) ;
    buf_clk new_AGEMA_reg_buffer_6307 ( .C (clk), .D (new_AGEMA_signal_9771), .Q (new_AGEMA_signal_9772) ) ;
    buf_clk new_AGEMA_reg_buffer_6311 ( .C (clk), .D (new_AGEMA_signal_9775), .Q (new_AGEMA_signal_9776) ) ;
    buf_clk new_AGEMA_reg_buffer_6315 ( .C (clk), .D (new_AGEMA_signal_9779), .Q (new_AGEMA_signal_9780) ) ;
    buf_clk new_AGEMA_reg_buffer_6317 ( .C (clk), .D (new_AGEMA_signal_7183), .Q (new_AGEMA_signal_9782) ) ;
    buf_clk new_AGEMA_reg_buffer_6319 ( .C (clk), .D (new_AGEMA_signal_7185), .Q (new_AGEMA_signal_9784) ) ;
    buf_clk new_AGEMA_reg_buffer_6321 ( .C (clk), .D (new_AGEMA_signal_7187), .Q (new_AGEMA_signal_9786) ) ;
    buf_clk new_AGEMA_reg_buffer_6325 ( .C (clk), .D (new_AGEMA_signal_9789), .Q (new_AGEMA_signal_9790) ) ;
    buf_clk new_AGEMA_reg_buffer_6329 ( .C (clk), .D (new_AGEMA_signal_9793), .Q (new_AGEMA_signal_9794) ) ;
    buf_clk new_AGEMA_reg_buffer_6333 ( .C (clk), .D (new_AGEMA_signal_9797), .Q (new_AGEMA_signal_9798) ) ;
    buf_clk new_AGEMA_reg_buffer_6335 ( .C (clk), .D (new_AGEMA_signal_7201), .Q (new_AGEMA_signal_9800) ) ;
    buf_clk new_AGEMA_reg_buffer_6337 ( .C (clk), .D (new_AGEMA_signal_7203), .Q (new_AGEMA_signal_9802) ) ;
    buf_clk new_AGEMA_reg_buffer_6339 ( .C (clk), .D (new_AGEMA_signal_7205), .Q (new_AGEMA_signal_9804) ) ;
    buf_clk new_AGEMA_reg_buffer_6343 ( .C (clk), .D (new_AGEMA_signal_9807), .Q (new_AGEMA_signal_9808) ) ;
    buf_clk new_AGEMA_reg_buffer_6347 ( .C (clk), .D (new_AGEMA_signal_9811), .Q (new_AGEMA_signal_9812) ) ;
    buf_clk new_AGEMA_reg_buffer_6351 ( .C (clk), .D (new_AGEMA_signal_9815), .Q (new_AGEMA_signal_9816) ) ;
    buf_clk new_AGEMA_reg_buffer_6353 ( .C (clk), .D (new_AGEMA_signal_7219), .Q (new_AGEMA_signal_9818) ) ;
    buf_clk new_AGEMA_reg_buffer_6355 ( .C (clk), .D (new_AGEMA_signal_7221), .Q (new_AGEMA_signal_9820) ) ;
    buf_clk new_AGEMA_reg_buffer_6357 ( .C (clk), .D (new_AGEMA_signal_7223), .Q (new_AGEMA_signal_9822) ) ;
    buf_clk new_AGEMA_reg_buffer_6361 ( .C (clk), .D (new_AGEMA_signal_9825), .Q (new_AGEMA_signal_9826) ) ;
    buf_clk new_AGEMA_reg_buffer_6365 ( .C (clk), .D (new_AGEMA_signal_9829), .Q (new_AGEMA_signal_9830) ) ;
    buf_clk new_AGEMA_reg_buffer_6369 ( .C (clk), .D (new_AGEMA_signal_9833), .Q (new_AGEMA_signal_9834) ) ;
    buf_clk new_AGEMA_reg_buffer_6371 ( .C (clk), .D (new_AGEMA_signal_7237), .Q (new_AGEMA_signal_9836) ) ;
    buf_clk new_AGEMA_reg_buffer_6373 ( .C (clk), .D (new_AGEMA_signal_7239), .Q (new_AGEMA_signal_9838) ) ;
    buf_clk new_AGEMA_reg_buffer_6375 ( .C (clk), .D (new_AGEMA_signal_7241), .Q (new_AGEMA_signal_9840) ) ;
    buf_clk new_AGEMA_reg_buffer_6379 ( .C (clk), .D (new_AGEMA_signal_9843), .Q (new_AGEMA_signal_9844) ) ;
    buf_clk new_AGEMA_reg_buffer_6383 ( .C (clk), .D (new_AGEMA_signal_9847), .Q (new_AGEMA_signal_9848) ) ;
    buf_clk new_AGEMA_reg_buffer_6387 ( .C (clk), .D (new_AGEMA_signal_9851), .Q (new_AGEMA_signal_9852) ) ;
    buf_clk new_AGEMA_reg_buffer_6389 ( .C (clk), .D (new_AGEMA_signal_7255), .Q (new_AGEMA_signal_9854) ) ;
    buf_clk new_AGEMA_reg_buffer_6391 ( .C (clk), .D (new_AGEMA_signal_7257), .Q (new_AGEMA_signal_9856) ) ;
    buf_clk new_AGEMA_reg_buffer_6393 ( .C (clk), .D (new_AGEMA_signal_7259), .Q (new_AGEMA_signal_9858) ) ;
    buf_clk new_AGEMA_reg_buffer_6397 ( .C (clk), .D (new_AGEMA_signal_9861), .Q (new_AGEMA_signal_9862) ) ;
    buf_clk new_AGEMA_reg_buffer_6401 ( .C (clk), .D (new_AGEMA_signal_9865), .Q (new_AGEMA_signal_9866) ) ;
    buf_clk new_AGEMA_reg_buffer_6405 ( .C (clk), .D (new_AGEMA_signal_9869), .Q (new_AGEMA_signal_9870) ) ;
    buf_clk new_AGEMA_reg_buffer_6407 ( .C (clk), .D (new_AGEMA_signal_7273), .Q (new_AGEMA_signal_9872) ) ;
    buf_clk new_AGEMA_reg_buffer_6409 ( .C (clk), .D (new_AGEMA_signal_7275), .Q (new_AGEMA_signal_9874) ) ;
    buf_clk new_AGEMA_reg_buffer_6411 ( .C (clk), .D (new_AGEMA_signal_7277), .Q (new_AGEMA_signal_9876) ) ;
    buf_clk new_AGEMA_reg_buffer_6415 ( .C (clk), .D (new_AGEMA_signal_9879), .Q (new_AGEMA_signal_9880) ) ;
    buf_clk new_AGEMA_reg_buffer_6419 ( .C (clk), .D (new_AGEMA_signal_9883), .Q (new_AGEMA_signal_9884) ) ;
    buf_clk new_AGEMA_reg_buffer_6423 ( .C (clk), .D (new_AGEMA_signal_9887), .Q (new_AGEMA_signal_9888) ) ;
    buf_clk new_AGEMA_reg_buffer_6425 ( .C (clk), .D (new_AGEMA_signal_7291), .Q (new_AGEMA_signal_9890) ) ;
    buf_clk new_AGEMA_reg_buffer_6427 ( .C (clk), .D (new_AGEMA_signal_7293), .Q (new_AGEMA_signal_9892) ) ;
    buf_clk new_AGEMA_reg_buffer_6429 ( .C (clk), .D (new_AGEMA_signal_7295), .Q (new_AGEMA_signal_9894) ) ;
    buf_clk new_AGEMA_reg_buffer_6433 ( .C (clk), .D (new_AGEMA_signal_9897), .Q (new_AGEMA_signal_9898) ) ;
    buf_clk new_AGEMA_reg_buffer_6437 ( .C (clk), .D (new_AGEMA_signal_9901), .Q (new_AGEMA_signal_9902) ) ;
    buf_clk new_AGEMA_reg_buffer_6441 ( .C (clk), .D (new_AGEMA_signal_9905), .Q (new_AGEMA_signal_9906) ) ;
    buf_clk new_AGEMA_reg_buffer_6443 ( .C (clk), .D (new_AGEMA_signal_7309), .Q (new_AGEMA_signal_9908) ) ;
    buf_clk new_AGEMA_reg_buffer_6445 ( .C (clk), .D (new_AGEMA_signal_7311), .Q (new_AGEMA_signal_9910) ) ;
    buf_clk new_AGEMA_reg_buffer_6447 ( .C (clk), .D (new_AGEMA_signal_7313), .Q (new_AGEMA_signal_9912) ) ;
    buf_clk new_AGEMA_reg_buffer_6451 ( .C (clk), .D (new_AGEMA_signal_9915), .Q (new_AGEMA_signal_9916) ) ;
    buf_clk new_AGEMA_reg_buffer_6455 ( .C (clk), .D (new_AGEMA_signal_9919), .Q (new_AGEMA_signal_9920) ) ;
    buf_clk new_AGEMA_reg_buffer_6459 ( .C (clk), .D (new_AGEMA_signal_9923), .Q (new_AGEMA_signal_9924) ) ;
    buf_clk new_AGEMA_reg_buffer_6467 ( .C (clk), .D (new_AGEMA_signal_9931), .Q (new_AGEMA_signal_9932) ) ;
    buf_clk new_AGEMA_reg_buffer_6475 ( .C (clk), .D (new_AGEMA_signal_9939), .Q (new_AGEMA_signal_9940) ) ;
    buf_clk new_AGEMA_reg_buffer_6483 ( .C (clk), .D (new_AGEMA_signal_9947), .Q (new_AGEMA_signal_9948) ) ;
    buf_clk new_AGEMA_reg_buffer_6491 ( .C (clk), .D (new_AGEMA_signal_9955), .Q (new_AGEMA_signal_9956) ) ;

    /* cells in depth 6 */
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U128 ( .a ({new_AGEMA_signal_5321, new_AGEMA_signal_5315, new_AGEMA_signal_5309}), .b ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, Midori_rounds_SR_Result[9]}), .c ({new_AGEMA_signal_4794, new_AGEMA_signal_4792, new_AGEMA_signal_4774}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U126 ( .a ({new_AGEMA_signal_5339, new_AGEMA_signal_5333, new_AGEMA_signal_5327}), .b ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, Midori_rounds_SR_Result[47]}), .c ({new_AGEMA_signal_4798, new_AGEMA_signal_4796, new_AGEMA_signal_4776}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U124 ( .a ({new_AGEMA_signal_5357, new_AGEMA_signal_5351, new_AGEMA_signal_5345}), .b ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, Midori_rounds_SR_Result[63]}), .c ({new_AGEMA_signal_4802, new_AGEMA_signal_4800, new_AGEMA_signal_4720}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U122 ( .a ({new_AGEMA_signal_5375, new_AGEMA_signal_5369, new_AGEMA_signal_5363}), .b ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, Midori_rounds_SR_Result[61]}), .c ({new_AGEMA_signal_4806, new_AGEMA_signal_4804, new_AGEMA_signal_4722}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U120 ( .a ({new_AGEMA_signal_5393, new_AGEMA_signal_5387, new_AGEMA_signal_5381}), .b ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, Midori_rounds_SR_Result[45]}), .c ({new_AGEMA_signal_4810, new_AGEMA_signal_4808, new_AGEMA_signal_4778}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U119 ( .a ({new_AGEMA_signal_5411, new_AGEMA_signal_5405, new_AGEMA_signal_5399}), .b ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, Midori_rounds_SR_Result[35]}), .c ({new_AGEMA_signal_4814, new_AGEMA_signal_4812, new_AGEMA_signal_4724}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U117 ( .a ({new_AGEMA_signal_5429, new_AGEMA_signal_5423, new_AGEMA_signal_5417}), .b ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, Midori_rounds_SR_Result[33]}), .c ({new_AGEMA_signal_4818, new_AGEMA_signal_4816, new_AGEMA_signal_4726}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U115 ( .a ({new_AGEMA_signal_5447, new_AGEMA_signal_5441, new_AGEMA_signal_5435}), .b ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, Midori_rounds_SR_Result[7]}), .c ({new_AGEMA_signal_4822, new_AGEMA_signal_4820, new_AGEMA_signal_4728}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U113 ( .a ({new_AGEMA_signal_5465, new_AGEMA_signal_5459, new_AGEMA_signal_5453}), .b ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, Midori_rounds_SR_Result[5]}), .c ({new_AGEMA_signal_4826, new_AGEMA_signal_4824, new_AGEMA_signal_4730}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U111 ( .a ({new_AGEMA_signal_5483, new_AGEMA_signal_5477, new_AGEMA_signal_5471}), .b ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, Midori_rounds_SR_Result[27]}), .c ({new_AGEMA_signal_4830, new_AGEMA_signal_4828, new_AGEMA_signal_4732}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U108 ( .a ({new_AGEMA_signal_5501, new_AGEMA_signal_5495, new_AGEMA_signal_5489}), .b ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, Midori_rounds_SR_Result[25]}), .c ({new_AGEMA_signal_4834, new_AGEMA_signal_4832, new_AGEMA_signal_4734}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U106 ( .a ({new_AGEMA_signal_5519, new_AGEMA_signal_5513, new_AGEMA_signal_5507}), .b ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, Midori_rounds_SR_Result[43]}), .c ({new_AGEMA_signal_4838, new_AGEMA_signal_4836, new_AGEMA_signal_4736}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U104 ( .a ({new_AGEMA_signal_5537, new_AGEMA_signal_5531, new_AGEMA_signal_5525}), .b ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, Midori_rounds_SR_Result[41]}), .c ({new_AGEMA_signal_4842, new_AGEMA_signal_4840, new_AGEMA_signal_4738}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U102 ( .a ({new_AGEMA_signal_5555, new_AGEMA_signal_5549, new_AGEMA_signal_5543}), .b ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, Midori_rounds_SR_Result[55]}), .c ({new_AGEMA_signal_4846, new_AGEMA_signal_4844, new_AGEMA_signal_4740}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U100 ( .a ({new_AGEMA_signal_5573, new_AGEMA_signal_5567, new_AGEMA_signal_5561}), .b ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, Midori_rounds_SR_Result[53]}), .c ({new_AGEMA_signal_4850, new_AGEMA_signal_4848, new_AGEMA_signal_4742}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U98 ( .a ({new_AGEMA_signal_5591, new_AGEMA_signal_5585, new_AGEMA_signal_5579}), .b ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, Midori_rounds_SR_Result[51]}), .c ({new_AGEMA_signal_4854, new_AGEMA_signal_4852, new_AGEMA_signal_4780}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U97 ( .a ({new_AGEMA_signal_5609, new_AGEMA_signal_5603, new_AGEMA_signal_5597}), .b ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, Midori_rounds_SR_Result[19]}), .c ({new_AGEMA_signal_4858, new_AGEMA_signal_4856, new_AGEMA_signal_4744}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U95 ( .a ({new_AGEMA_signal_5627, new_AGEMA_signal_5621, new_AGEMA_signal_5615}), .b ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, Midori_rounds_SR_Result[17]}), .c ({new_AGEMA_signal_4862, new_AGEMA_signal_4860, new_AGEMA_signal_4746}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U93 ( .a ({new_AGEMA_signal_5645, new_AGEMA_signal_5639, new_AGEMA_signal_5633}), .b ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, Midori_rounds_SR_Result[15]}), .c ({new_AGEMA_signal_4866, new_AGEMA_signal_4864, new_AGEMA_signal_4748}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U91 ( .a ({new_AGEMA_signal_5663, new_AGEMA_signal_5657, new_AGEMA_signal_5651}), .b ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, Midori_rounds_SR_Result[13]}), .c ({new_AGEMA_signal_4870, new_AGEMA_signal_4868, new_AGEMA_signal_4750}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U89 ( .a ({new_AGEMA_signal_5681, new_AGEMA_signal_5675, new_AGEMA_signal_5669}), .b ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, Midori_rounds_SR_Result[3]}), .c ({new_AGEMA_signal_4874, new_AGEMA_signal_4872, new_AGEMA_signal_4752}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U86 ( .a ({new_AGEMA_signal_5699, new_AGEMA_signal_5693, new_AGEMA_signal_5687}), .b ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, Midori_rounds_SR_Result[1]}), .c ({new_AGEMA_signal_4878, new_AGEMA_signal_4876, new_AGEMA_signal_4754}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U84 ( .a ({new_AGEMA_signal_5717, new_AGEMA_signal_5711, new_AGEMA_signal_5705}), .b ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, Midori_rounds_SR_Result[31]}), .c ({new_AGEMA_signal_4882, new_AGEMA_signal_4880, new_AGEMA_signal_4756}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U82 ( .a ({new_AGEMA_signal_5735, new_AGEMA_signal_5729, new_AGEMA_signal_5723}), .b ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, Midori_rounds_SR_Result[29]}), .c ({new_AGEMA_signal_4886, new_AGEMA_signal_4884, new_AGEMA_signal_4758}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U80 ( .a ({new_AGEMA_signal_5753, new_AGEMA_signal_5747, new_AGEMA_signal_5741}), .b ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, Midori_rounds_SR_Result[59]}), .c ({new_AGEMA_signal_4890, new_AGEMA_signal_4888, new_AGEMA_signal_4760}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U78 ( .a ({new_AGEMA_signal_5771, new_AGEMA_signal_5765, new_AGEMA_signal_5759}), .b ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, Midori_rounds_SR_Result[57]}), .c ({new_AGEMA_signal_4894, new_AGEMA_signal_4892, new_AGEMA_signal_4762}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U76 ( .a ({new_AGEMA_signal_5789, new_AGEMA_signal_5783, new_AGEMA_signal_5777}), .b ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, Midori_rounds_SR_Result[49]}), .c ({new_AGEMA_signal_4898, new_AGEMA_signal_4896, new_AGEMA_signal_4782}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U75 ( .a ({new_AGEMA_signal_5807, new_AGEMA_signal_5801, new_AGEMA_signal_5795}), .b ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, Midori_rounds_SR_Result[39]}), .c ({new_AGEMA_signal_4902, new_AGEMA_signal_4900, new_AGEMA_signal_4764}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U73 ( .a ({new_AGEMA_signal_5825, new_AGEMA_signal_5819, new_AGEMA_signal_5813}), .b ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, Midori_rounds_SR_Result[37]}), .c ({new_AGEMA_signal_4906, new_AGEMA_signal_4904, new_AGEMA_signal_4766}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U71 ( .a ({new_AGEMA_signal_5843, new_AGEMA_signal_5837, new_AGEMA_signal_5831}), .b ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, Midori_rounds_SR_Result[23]}), .c ({new_AGEMA_signal_4910, new_AGEMA_signal_4908, new_AGEMA_signal_4768}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U69 ( .a ({new_AGEMA_signal_5861, new_AGEMA_signal_5855, new_AGEMA_signal_5849}), .b ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, Midori_rounds_SR_Result[21]}), .c ({new_AGEMA_signal_4914, new_AGEMA_signal_4912, new_AGEMA_signal_4770}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U67 ( .a ({new_AGEMA_signal_5879, new_AGEMA_signal_5873, new_AGEMA_signal_5867}), .b ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, Midori_rounds_SR_Result[11]}), .c ({new_AGEMA_signal_4918, new_AGEMA_signal_4916, new_AGEMA_signal_4772}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U144 ( .a ({new_AGEMA_signal_5897, new_AGEMA_signal_5891, new_AGEMA_signal_5885}), .b ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, Midori_rounds_SR_Result[9]}), .c ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, Midori_rounds_sub_ResultXORkey[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U142 ( .a ({new_AGEMA_signal_5915, new_AGEMA_signal_5909, new_AGEMA_signal_5903}), .b ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, Midori_rounds_SR_Result[47]}), .c ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, Midori_rounds_sub_ResultXORkey[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U140 ( .a ({new_AGEMA_signal_5933, new_AGEMA_signal_5927, new_AGEMA_signal_5921}), .b ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, Midori_rounds_SR_Result[63]}), .c ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, Midori_rounds_sub_ResultXORkey[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U138 ( .a ({new_AGEMA_signal_5951, new_AGEMA_signal_5945, new_AGEMA_signal_5939}), .b ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, Midori_rounds_SR_Result[61]}), .c ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, Midori_rounds_sub_ResultXORkey[61]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U136 ( .a ({new_AGEMA_signal_5969, new_AGEMA_signal_5963, new_AGEMA_signal_5957}), .b ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, Midori_rounds_SR_Result[45]}), .c ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, Midori_rounds_sub_ResultXORkey[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U135 ( .a ({new_AGEMA_signal_5987, new_AGEMA_signal_5981, new_AGEMA_signal_5975}), .b ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, Midori_rounds_SR_Result[35]}), .c ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, Midori_rounds_sub_ResultXORkey[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U133 ( .a ({new_AGEMA_signal_6005, new_AGEMA_signal_5999, new_AGEMA_signal_5993}), .b ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, Midori_rounds_SR_Result[33]}), .c ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, Midori_rounds_sub_ResultXORkey[57]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U131 ( .a ({new_AGEMA_signal_6023, new_AGEMA_signal_6017, new_AGEMA_signal_6011}), .b ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, Midori_rounds_SR_Result[7]}), .c ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, Midori_rounds_sub_ResultXORkey[55]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U129 ( .a ({new_AGEMA_signal_6041, new_AGEMA_signal_6035, new_AGEMA_signal_6029}), .b ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, Midori_rounds_SR_Result[5]}), .c ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, Midori_rounds_sub_ResultXORkey[53]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U127 ( .a ({new_AGEMA_signal_6059, new_AGEMA_signal_6053, new_AGEMA_signal_6047}), .b ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, Midori_rounds_SR_Result[27]}), .c ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, Midori_rounds_sub_ResultXORkey[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U124 ( .a ({new_AGEMA_signal_6077, new_AGEMA_signal_6071, new_AGEMA_signal_6065}), .b ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, Midori_rounds_SR_Result[25]}), .c ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, Midori_rounds_sub_ResultXORkey[49]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U122 ( .a ({new_AGEMA_signal_6095, new_AGEMA_signal_6089, new_AGEMA_signal_6083}), .b ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, Midori_rounds_SR_Result[43]}), .c ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, Midori_rounds_sub_ResultXORkey[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U120 ( .a ({new_AGEMA_signal_6113, new_AGEMA_signal_6107, new_AGEMA_signal_6101}), .b ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, Midori_rounds_SR_Result[41]}), .c ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, Midori_rounds_sub_ResultXORkey[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U118 ( .a ({new_AGEMA_signal_6131, new_AGEMA_signal_6125, new_AGEMA_signal_6119}), .b ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, Midori_rounds_SR_Result[55]}), .c ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, Midori_rounds_sub_ResultXORkey[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U116 ( .a ({new_AGEMA_signal_6149, new_AGEMA_signal_6143, new_AGEMA_signal_6137}), .b ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, Midori_rounds_SR_Result[53]}), .c ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, Midori_rounds_sub_ResultXORkey[41]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U114 ( .a ({new_AGEMA_signal_6167, new_AGEMA_signal_6161, new_AGEMA_signal_6155}), .b ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, Midori_rounds_SR_Result[51]}), .c ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, Midori_rounds_sub_ResultXORkey[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U113 ( .a ({new_AGEMA_signal_6185, new_AGEMA_signal_6179, new_AGEMA_signal_6173}), .b ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, Midori_rounds_SR_Result[19]}), .c ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, Midori_rounds_sub_ResultXORkey[39]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U111 ( .a ({new_AGEMA_signal_6203, new_AGEMA_signal_6197, new_AGEMA_signal_6191}), .b ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, Midori_rounds_SR_Result[17]}), .c ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, Midori_rounds_sub_ResultXORkey[37]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U109 ( .a ({new_AGEMA_signal_6221, new_AGEMA_signal_6215, new_AGEMA_signal_6209}), .b ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, Midori_rounds_SR_Result[15]}), .c ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, Midori_rounds_sub_ResultXORkey[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U107 ( .a ({new_AGEMA_signal_6239, new_AGEMA_signal_6233, new_AGEMA_signal_6227}), .b ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, Midori_rounds_SR_Result[13]}), .c ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, Midori_rounds_sub_ResultXORkey[33]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U105 ( .a ({new_AGEMA_signal_6257, new_AGEMA_signal_6251, new_AGEMA_signal_6245}), .b ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, Midori_rounds_SR_Result[3]}), .c ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, Midori_rounds_sub_ResultXORkey[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U102 ( .a ({new_AGEMA_signal_6275, new_AGEMA_signal_6269, new_AGEMA_signal_6263}), .b ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, Midori_rounds_SR_Result[1]}), .c ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, Midori_rounds_sub_ResultXORkey[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U100 ( .a ({new_AGEMA_signal_6293, new_AGEMA_signal_6287, new_AGEMA_signal_6281}), .b ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, Midori_rounds_SR_Result[31]}), .c ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, Midori_rounds_sub_ResultXORkey[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U98 ( .a ({new_AGEMA_signal_6311, new_AGEMA_signal_6305, new_AGEMA_signal_6299}), .b ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, Midori_rounds_SR_Result[29]}), .c ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, Midori_rounds_sub_ResultXORkey[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U96 ( .a ({new_AGEMA_signal_6329, new_AGEMA_signal_6323, new_AGEMA_signal_6317}), .b ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, Midori_rounds_SR_Result[59]}), .c ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, Midori_rounds_sub_ResultXORkey[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U94 ( .a ({new_AGEMA_signal_6347, new_AGEMA_signal_6341, new_AGEMA_signal_6335}), .b ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, Midori_rounds_SR_Result[57]}), .c ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, Midori_rounds_sub_ResultXORkey[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U92 ( .a ({new_AGEMA_signal_6365, new_AGEMA_signal_6359, new_AGEMA_signal_6353}), .b ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, Midori_rounds_SR_Result[49]}), .c ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, Midori_rounds_sub_ResultXORkey[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U91 ( .a ({new_AGEMA_signal_6383, new_AGEMA_signal_6377, new_AGEMA_signal_6371}), .b ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, Midori_rounds_SR_Result[39]}), .c ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, Midori_rounds_sub_ResultXORkey[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U89 ( .a ({new_AGEMA_signal_6401, new_AGEMA_signal_6395, new_AGEMA_signal_6389}), .b ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, Midori_rounds_SR_Result[37]}), .c ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, Midori_rounds_sub_ResultXORkey[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U87 ( .a ({new_AGEMA_signal_6419, new_AGEMA_signal_6413, new_AGEMA_signal_6407}), .b ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, Midori_rounds_SR_Result[23]}), .c ({new_AGEMA_signal_3175, new_AGEMA_signal_3174, Midori_rounds_sub_ResultXORkey[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U85 ( .a ({new_AGEMA_signal_6437, new_AGEMA_signal_6431, new_AGEMA_signal_6425}), .b ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, Midori_rounds_SR_Result[21]}), .c ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, Midori_rounds_sub_ResultXORkey[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U83 ( .a ({new_AGEMA_signal_6455, new_AGEMA_signal_6449, new_AGEMA_signal_6443}), .b ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, Midori_rounds_SR_Result[11]}), .c ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, Midori_rounds_sub_ResultXORkey[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U80 ( .a ({new_AGEMA_signal_5897, new_AGEMA_signal_5891, new_AGEMA_signal_5885}), .b ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, Midori_rounds_SR_Inv_Result[9]}), .c ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, Midori_rounds_mul_ResultXORkey[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U77 ( .a ({new_AGEMA_signal_5915, new_AGEMA_signal_5909, new_AGEMA_signal_5903}), .b ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, Midori_rounds_SR_Inv_Result[55]}), .c ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, Midori_rounds_mul_ResultXORkey[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U75 ( .a ({new_AGEMA_signal_5933, new_AGEMA_signal_5927, new_AGEMA_signal_5921}), .b ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, Midori_rounds_SR_Inv_Result[63]}), .c ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, Midori_rounds_mul_ResultXORkey[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U73 ( .a ({new_AGEMA_signal_5951, new_AGEMA_signal_5945, new_AGEMA_signal_5939}), .b ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, Midori_rounds_SR_Inv_Result[61]}), .c ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, Midori_rounds_mul_ResultXORkey[61]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U70 ( .a ({new_AGEMA_signal_5969, new_AGEMA_signal_5963, new_AGEMA_signal_5957}), .b ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, Midori_rounds_SR_Inv_Result[53]}), .c ({new_AGEMA_signal_3439, new_AGEMA_signal_3438, Midori_rounds_mul_ResultXORkey[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U69 ( .a ({new_AGEMA_signal_5987, new_AGEMA_signal_5981, new_AGEMA_signal_5975}), .b ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, Midori_rounds_SR_Inv_Result[23]}), .c ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, Midori_rounds_mul_ResultXORkey[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U67 ( .a ({new_AGEMA_signal_6005, new_AGEMA_signal_5999, new_AGEMA_signal_5993}), .b ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, Midori_rounds_SR_Inv_Result[21]}), .c ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, Midori_rounds_mul_ResultXORkey[57]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U64 ( .a ({new_AGEMA_signal_6023, new_AGEMA_signal_6017, new_AGEMA_signal_6011}), .b ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, Midori_rounds_SR_Inv_Result[43]}), .c ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, Midori_rounds_mul_ResultXORkey[55]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U62 ( .a ({new_AGEMA_signal_6041, new_AGEMA_signal_6035, new_AGEMA_signal_6029}), .b ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, Midori_rounds_SR_Inv_Result[41]}), .c ({new_AGEMA_signal_3451, new_AGEMA_signal_3450, Midori_rounds_mul_ResultXORkey[53]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U59 ( .a ({new_AGEMA_signal_6059, new_AGEMA_signal_6053, new_AGEMA_signal_6047}), .b ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, Midori_rounds_SR_Inv_Result[3]}), .c ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, Midori_rounds_mul_ResultXORkey[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U55 ( .a ({new_AGEMA_signal_6077, new_AGEMA_signal_6071, new_AGEMA_signal_6065}), .b ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, Midori_rounds_SR_Inv_Result[1]}), .c ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, Midori_rounds_mul_ResultXORkey[49]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U52 ( .a ({new_AGEMA_signal_6095, new_AGEMA_signal_6089, new_AGEMA_signal_6083}), .b ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, Midori_rounds_SR_Inv_Result[7]}), .c ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, Midori_rounds_mul_ResultXORkey[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U50 ( .a ({new_AGEMA_signal_6113, new_AGEMA_signal_6107, new_AGEMA_signal_6101}), .b ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, Midori_rounds_SR_Inv_Result[5]}), .c ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, Midori_rounds_mul_ResultXORkey[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U47 ( .a ({new_AGEMA_signal_6131, new_AGEMA_signal_6125, new_AGEMA_signal_6119}), .b ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, Midori_rounds_SR_Inv_Result[47]}), .c ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, Midori_rounds_mul_ResultXORkey[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U45 ( .a ({new_AGEMA_signal_6149, new_AGEMA_signal_6143, new_AGEMA_signal_6137}), .b ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, Midori_rounds_SR_Inv_Result[45]}), .c ({new_AGEMA_signal_3471, new_AGEMA_signal_3470, Midori_rounds_mul_ResultXORkey[41]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U42 ( .a ({new_AGEMA_signal_6167, new_AGEMA_signal_6161, new_AGEMA_signal_6155}), .b ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, Midori_rounds_SR_Inv_Result[31]}), .c ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, Midori_rounds_mul_ResultXORkey[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U41 ( .a ({new_AGEMA_signal_6185, new_AGEMA_signal_6179, new_AGEMA_signal_6173}), .b ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, Midori_rounds_SR_Inv_Result[19]}), .c ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, Midori_rounds_mul_ResultXORkey[39]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U39 ( .a ({new_AGEMA_signal_6203, new_AGEMA_signal_6197, new_AGEMA_signal_6191}), .b ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, Midori_rounds_SR_Inv_Result[17]}), .c ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, Midori_rounds_mul_ResultXORkey[37]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U36 ( .a ({new_AGEMA_signal_6221, new_AGEMA_signal_6215, new_AGEMA_signal_6209}), .b ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, Midori_rounds_SR_Inv_Result[59]}), .c ({new_AGEMA_signal_3483, new_AGEMA_signal_3482, Midori_rounds_mul_ResultXORkey[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U34 ( .a ({new_AGEMA_signal_6239, new_AGEMA_signal_6233, new_AGEMA_signal_6227}), .b ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, Midori_rounds_SR_Inv_Result[57]}), .c ({new_AGEMA_signal_3487, new_AGEMA_signal_3486, Midori_rounds_mul_ResultXORkey[33]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U31 ( .a ({new_AGEMA_signal_6257, new_AGEMA_signal_6251, new_AGEMA_signal_6245}), .b ({new_AGEMA_signal_3391, new_AGEMA_signal_3390, Midori_rounds_SR_Inv_Result[27]}), .c ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, Midori_rounds_mul_ResultXORkey[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U28 ( .a ({new_AGEMA_signal_6275, new_AGEMA_signal_6269, new_AGEMA_signal_6263}), .b ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, Midori_rounds_SR_Inv_Result[25]}), .c ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, Midori_rounds_mul_ResultXORkey[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U25 ( .a ({new_AGEMA_signal_6293, new_AGEMA_signal_6287, new_AGEMA_signal_6281}), .b ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, Midori_rounds_SR_Inv_Result[51]}), .c ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, Midori_rounds_mul_ResultXORkey[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U23 ( .a ({new_AGEMA_signal_6311, new_AGEMA_signal_6305, new_AGEMA_signal_6299}), .b ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, Midori_rounds_SR_Inv_Result[49]}), .c ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, Midori_rounds_mul_ResultXORkey[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U20 ( .a ({new_AGEMA_signal_6329, new_AGEMA_signal_6323, new_AGEMA_signal_6317}), .b ({new_AGEMA_signal_3379, new_AGEMA_signal_3378, Midori_rounds_SR_Inv_Result[15]}), .c ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, Midori_rounds_mul_ResultXORkey[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U18 ( .a ({new_AGEMA_signal_6347, new_AGEMA_signal_6341, new_AGEMA_signal_6335}), .b ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, Midori_rounds_SR_Inv_Result[13]}), .c ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, Midori_rounds_mul_ResultXORkey[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U15 ( .a ({new_AGEMA_signal_6365, new_AGEMA_signal_6359, new_AGEMA_signal_6353}), .b ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, Midori_rounds_SR_Inv_Result[29]}), .c ({new_AGEMA_signal_3511, new_AGEMA_signal_3510, Midori_rounds_mul_ResultXORkey[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U14 ( .a ({new_AGEMA_signal_6383, new_AGEMA_signal_6377, new_AGEMA_signal_6371}), .b ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, Midori_rounds_SR_Inv_Result[39]}), .c ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, Midori_rounds_mul_ResultXORkey[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U12 ( .a ({new_AGEMA_signal_6401, new_AGEMA_signal_6395, new_AGEMA_signal_6389}), .b ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, Midori_rounds_SR_Inv_Result[37]}), .c ({new_AGEMA_signal_3517, new_AGEMA_signal_3516, Midori_rounds_mul_ResultXORkey[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U9 ( .a ({new_AGEMA_signal_6419, new_AGEMA_signal_6413, new_AGEMA_signal_6407}), .b ({new_AGEMA_signal_3415, new_AGEMA_signal_3414, Midori_rounds_SR_Inv_Result[35]}), .c ({new_AGEMA_signal_3519, new_AGEMA_signal_3518, Midori_rounds_mul_ResultXORkey[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U7 ( .a ({new_AGEMA_signal_6437, new_AGEMA_signal_6431, new_AGEMA_signal_6425}), .b ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, Midori_rounds_SR_Inv_Result[33]}), .c ({new_AGEMA_signal_3523, new_AGEMA_signal_3522, Midori_rounds_mul_ResultXORkey[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U4 ( .a ({new_AGEMA_signal_6455, new_AGEMA_signal_6449, new_AGEMA_signal_6443}), .b ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, Midori_rounds_SR_Inv_Result[11]}), .c ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, Midori_rounds_mul_ResultXORkey[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, Midori_rounds_round_Result[1]}), .a ({new_AGEMA_signal_6479, new_AGEMA_signal_6473, new_AGEMA_signal_6467}), .c ({new_AGEMA_signal_3675, new_AGEMA_signal_3674, Midori_rounds_roundResult_Reg_SFF_1_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, Midori_rounds_round_Result[3]}), .a ({new_AGEMA_signal_6497, new_AGEMA_signal_6491, new_AGEMA_signal_6485}), .c ({new_AGEMA_signal_3679, new_AGEMA_signal_3678, Midori_rounds_roundResult_Reg_SFF_3_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, Midori_rounds_round_Result[5]}), .a ({new_AGEMA_signal_6515, new_AGEMA_signal_6509, new_AGEMA_signal_6503}), .c ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, Midori_rounds_roundResult_Reg_SFF_5_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, Midori_rounds_round_Result[7]}), .a ({new_AGEMA_signal_6533, new_AGEMA_signal_6527, new_AGEMA_signal_6521}), .c ({new_AGEMA_signal_3685, new_AGEMA_signal_3684, Midori_rounds_roundResult_Reg_SFF_7_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, Midori_rounds_round_Result[9]}), .a ({new_AGEMA_signal_6551, new_AGEMA_signal_6545, new_AGEMA_signal_6539}), .c ({new_AGEMA_signal_3687, new_AGEMA_signal_3686, Midori_rounds_roundResult_Reg_SFF_9_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, Midori_rounds_round_Result[11]}), .a ({new_AGEMA_signal_6569, new_AGEMA_signal_6563, new_AGEMA_signal_6557}), .c ({new_AGEMA_signal_3691, new_AGEMA_signal_3690, Midori_rounds_roundResult_Reg_SFF_11_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, Midori_rounds_round_Result[13]}), .a ({new_AGEMA_signal_6587, new_AGEMA_signal_6581, new_AGEMA_signal_6575}), .c ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, Midori_rounds_roundResult_Reg_SFF_13_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, Midori_rounds_round_Result[15]}), .a ({new_AGEMA_signal_6605, new_AGEMA_signal_6599, new_AGEMA_signal_6593}), .c ({new_AGEMA_signal_3697, new_AGEMA_signal_3696, Midori_rounds_roundResult_Reg_SFF_15_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, Midori_rounds_round_Result[17]}), .a ({new_AGEMA_signal_6623, new_AGEMA_signal_6617, new_AGEMA_signal_6611}), .c ({new_AGEMA_signal_3699, new_AGEMA_signal_3698, Midori_rounds_roundResult_Reg_SFF_17_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, Midori_rounds_round_Result[19]}), .a ({new_AGEMA_signal_6641, new_AGEMA_signal_6635, new_AGEMA_signal_6629}), .c ({new_AGEMA_signal_3703, new_AGEMA_signal_3702, Midori_rounds_roundResult_Reg_SFF_19_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, Midori_rounds_round_Result[21]}), .a ({new_AGEMA_signal_6659, new_AGEMA_signal_6653, new_AGEMA_signal_6647}), .c ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, Midori_rounds_roundResult_Reg_SFF_21_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, Midori_rounds_round_Result[23]}), .a ({new_AGEMA_signal_6677, new_AGEMA_signal_6671, new_AGEMA_signal_6665}), .c ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, Midori_rounds_roundResult_Reg_SFF_23_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, Midori_rounds_round_Result[25]}), .a ({new_AGEMA_signal_6695, new_AGEMA_signal_6689, new_AGEMA_signal_6683}), .c ({new_AGEMA_signal_3711, new_AGEMA_signal_3710, Midori_rounds_roundResult_Reg_SFF_25_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, Midori_rounds_round_Result[27]}), .a ({new_AGEMA_signal_6713, new_AGEMA_signal_6707, new_AGEMA_signal_6701}), .c ({new_AGEMA_signal_3715, new_AGEMA_signal_3714, Midori_rounds_roundResult_Reg_SFF_27_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, Midori_rounds_round_Result[29]}), .a ({new_AGEMA_signal_6731, new_AGEMA_signal_6725, new_AGEMA_signal_6719}), .c ({new_AGEMA_signal_3717, new_AGEMA_signal_3716, Midori_rounds_roundResult_Reg_SFF_29_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, Midori_rounds_round_Result[31]}), .a ({new_AGEMA_signal_6749, new_AGEMA_signal_6743, new_AGEMA_signal_6737}), .c ({new_AGEMA_signal_3721, new_AGEMA_signal_3720, Midori_rounds_roundResult_Reg_SFF_31_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, Midori_rounds_round_Result[33]}), .a ({new_AGEMA_signal_6767, new_AGEMA_signal_6761, new_AGEMA_signal_6755}), .c ({new_AGEMA_signal_3723, new_AGEMA_signal_3722, Midori_rounds_roundResult_Reg_SFF_33_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, Midori_rounds_round_Result[35]}), .a ({new_AGEMA_signal_6785, new_AGEMA_signal_6779, new_AGEMA_signal_6773}), .c ({new_AGEMA_signal_3727, new_AGEMA_signal_3726, Midori_rounds_roundResult_Reg_SFF_35_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, Midori_rounds_round_Result[37]}), .a ({new_AGEMA_signal_6803, new_AGEMA_signal_6797, new_AGEMA_signal_6791}), .c ({new_AGEMA_signal_3729, new_AGEMA_signal_3728, Midori_rounds_roundResult_Reg_SFF_37_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, Midori_rounds_round_Result[39]}), .a ({new_AGEMA_signal_6821, new_AGEMA_signal_6815, new_AGEMA_signal_6809}), .c ({new_AGEMA_signal_3733, new_AGEMA_signal_3732, Midori_rounds_roundResult_Reg_SFF_39_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, Midori_rounds_round_Result[41]}), .a ({new_AGEMA_signal_6839, new_AGEMA_signal_6833, new_AGEMA_signal_6827}), .c ({new_AGEMA_signal_3735, new_AGEMA_signal_3734, Midori_rounds_roundResult_Reg_SFF_41_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, Midori_rounds_round_Result[43]}), .a ({new_AGEMA_signal_6857, new_AGEMA_signal_6851, new_AGEMA_signal_6845}), .c ({new_AGEMA_signal_3739, new_AGEMA_signal_3738, Midori_rounds_roundResult_Reg_SFF_43_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3623, new_AGEMA_signal_3622, Midori_rounds_round_Result[45]}), .a ({new_AGEMA_signal_6875, new_AGEMA_signal_6869, new_AGEMA_signal_6863}), .c ({new_AGEMA_signal_3741, new_AGEMA_signal_3740, Midori_rounds_roundResult_Reg_SFF_45_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3627, new_AGEMA_signal_3626, Midori_rounds_round_Result[47]}), .a ({new_AGEMA_signal_6893, new_AGEMA_signal_6887, new_AGEMA_signal_6881}), .c ({new_AGEMA_signal_3745, new_AGEMA_signal_3744, Midori_rounds_roundResult_Reg_SFF_47_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, Midori_rounds_round_Result[49]}), .a ({new_AGEMA_signal_6911, new_AGEMA_signal_6905, new_AGEMA_signal_6899}), .c ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, Midori_rounds_roundResult_Reg_SFF_49_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, Midori_rounds_round_Result[51]}), .a ({new_AGEMA_signal_6929, new_AGEMA_signal_6923, new_AGEMA_signal_6917}), .c ({new_AGEMA_signal_3751, new_AGEMA_signal_3750, Midori_rounds_roundResult_Reg_SFF_51_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3635, new_AGEMA_signal_3634, Midori_rounds_round_Result[53]}), .a ({new_AGEMA_signal_6947, new_AGEMA_signal_6941, new_AGEMA_signal_6935}), .c ({new_AGEMA_signal_3753, new_AGEMA_signal_3752, Midori_rounds_roundResult_Reg_SFF_53_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3639, new_AGEMA_signal_3638, Midori_rounds_round_Result[55]}), .a ({new_AGEMA_signal_6965, new_AGEMA_signal_6959, new_AGEMA_signal_6953}), .c ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, Midori_rounds_roundResult_Reg_SFF_55_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, Midori_rounds_round_Result[57]}), .a ({new_AGEMA_signal_6983, new_AGEMA_signal_6977, new_AGEMA_signal_6971}), .c ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, Midori_rounds_roundResult_Reg_SFF_57_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, Midori_rounds_round_Result[59]}), .a ({new_AGEMA_signal_7001, new_AGEMA_signal_6995, new_AGEMA_signal_6989}), .c ({new_AGEMA_signal_3763, new_AGEMA_signal_3762, Midori_rounds_roundResult_Reg_SFF_59_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3647, new_AGEMA_signal_3646, Midori_rounds_round_Result[61]}), .a ({new_AGEMA_signal_7019, new_AGEMA_signal_7013, new_AGEMA_signal_7007}), .c ({new_AGEMA_signal_3765, new_AGEMA_signal_3764, Midori_rounds_roundResult_Reg_SFF_61_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1 ( .s (new_AGEMA_signal_6461), .b ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, Midori_rounds_round_Result[63]}), .a ({new_AGEMA_signal_7037, new_AGEMA_signal_7031, new_AGEMA_signal_7025}), .c ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, Midori_rounds_roundResult_Reg_SFF_63_DQ}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U19 ( .a ({new_AGEMA_signal_7043, new_AGEMA_signal_7041, new_AGEMA_signal_7039}), .b ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, Midori_rounds_sub_sBox_PRINCE_0_n14}), .clk (clk), .r ({Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, Midori_rounds_SR_Result[51]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U16 ( .a ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, Midori_rounds_sub_sBox_PRINCE_0_n11}), .b ({new_AGEMA_signal_7049, new_AGEMA_signal_7047, new_AGEMA_signal_7045}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483]}), .c ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, Midori_rounds_sub_sBox_PRINCE_0_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U12 ( .a ({new_AGEMA_signal_7055, new_AGEMA_signal_7053, new_AGEMA_signal_7051}), .b ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, Midori_rounds_sub_sBox_PRINCE_0_n5}), .clk (clk), .r ({Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, Midori_rounds_SR_Result[49]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U7 ( .a ({new_AGEMA_signal_7049, new_AGEMA_signal_7047, new_AGEMA_signal_7045}), .b ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, Midori_rounds_sub_sBox_PRINCE_0_n2}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489]}), .c ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, Midori_rounds_sub_sBox_PRINCE_0_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U19 ( .a ({new_AGEMA_signal_7061, new_AGEMA_signal_7059, new_AGEMA_signal_7057}), .b ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, Midori_rounds_sub_sBox_PRINCE_1_n14}), .clk (clk), .r ({Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, Midori_rounds_SR_Result[47]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U16 ( .a ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, Midori_rounds_sub_sBox_PRINCE_1_n11}), .b ({new_AGEMA_signal_7067, new_AGEMA_signal_7065, new_AGEMA_signal_7063}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495]}), .c ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, Midori_rounds_sub_sBox_PRINCE_1_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U12 ( .a ({new_AGEMA_signal_7073, new_AGEMA_signal_7071, new_AGEMA_signal_7069}), .b ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, Midori_rounds_sub_sBox_PRINCE_1_n5}), .clk (clk), .r ({Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, Midori_rounds_SR_Result[45]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U7 ( .a ({new_AGEMA_signal_7067, new_AGEMA_signal_7065, new_AGEMA_signal_7063}), .b ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, Midori_rounds_sub_sBox_PRINCE_1_n2}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501]}), .c ({new_AGEMA_signal_2691, new_AGEMA_signal_2690, Midori_rounds_sub_sBox_PRINCE_1_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U19 ( .a ({new_AGEMA_signal_7079, new_AGEMA_signal_7077, new_AGEMA_signal_7075}), .b ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, Midori_rounds_sub_sBox_PRINCE_2_n14}), .clk (clk), .r ({Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, Midori_rounds_SR_Result[11]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U16 ( .a ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, Midori_rounds_sub_sBox_PRINCE_2_n11}), .b ({new_AGEMA_signal_7085, new_AGEMA_signal_7083, new_AGEMA_signal_7081}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507]}), .c ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, Midori_rounds_sub_sBox_PRINCE_2_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U12 ( .a ({new_AGEMA_signal_7091, new_AGEMA_signal_7089, new_AGEMA_signal_7087}), .b ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, Midori_rounds_sub_sBox_PRINCE_2_n5}), .clk (clk), .r ({Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, Midori_rounds_SR_Result[9]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U7 ( .a ({new_AGEMA_signal_7085, new_AGEMA_signal_7083, new_AGEMA_signal_7081}), .b ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, Midori_rounds_sub_sBox_PRINCE_2_n2}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513]}), .c ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, Midori_rounds_sub_sBox_PRINCE_2_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U19 ( .a ({new_AGEMA_signal_7097, new_AGEMA_signal_7095, new_AGEMA_signal_7093}), .b ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, Midori_rounds_sub_sBox_PRINCE_3_n14}), .clk (clk), .r ({Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, Midori_rounds_SR_Result[23]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U16 ( .a ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, Midori_rounds_sub_sBox_PRINCE_3_n11}), .b ({new_AGEMA_signal_7103, new_AGEMA_signal_7101, new_AGEMA_signal_7099}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519]}), .c ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, Midori_rounds_sub_sBox_PRINCE_3_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U12 ( .a ({new_AGEMA_signal_7109, new_AGEMA_signal_7107, new_AGEMA_signal_7105}), .b ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, Midori_rounds_sub_sBox_PRINCE_3_n5}), .clk (clk), .r ({Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, Midori_rounds_SR_Result[21]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U7 ( .a ({new_AGEMA_signal_7103, new_AGEMA_signal_7101, new_AGEMA_signal_7099}), .b ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, Midori_rounds_sub_sBox_PRINCE_3_n2}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525]}), .c ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, Midori_rounds_sub_sBox_PRINCE_3_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U19 ( .a ({new_AGEMA_signal_7115, new_AGEMA_signal_7113, new_AGEMA_signal_7111}), .b ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, Midori_rounds_sub_sBox_PRINCE_4_n14}), .clk (clk), .r ({Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, Midori_rounds_SR_Result[39]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U16 ( .a ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, Midori_rounds_sub_sBox_PRINCE_4_n11}), .b ({new_AGEMA_signal_7121, new_AGEMA_signal_7119, new_AGEMA_signal_7117}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531]}), .c ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, Midori_rounds_sub_sBox_PRINCE_4_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U12 ( .a ({new_AGEMA_signal_7127, new_AGEMA_signal_7125, new_AGEMA_signal_7123}), .b ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, Midori_rounds_sub_sBox_PRINCE_4_n5}), .clk (clk), .r ({Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, Midori_rounds_SR_Result[37]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U7 ( .a ({new_AGEMA_signal_7121, new_AGEMA_signal_7119, new_AGEMA_signal_7117}), .b ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, Midori_rounds_sub_sBox_PRINCE_4_n2}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537]}), .c ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, Midori_rounds_sub_sBox_PRINCE_4_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U19 ( .a ({new_AGEMA_signal_7133, new_AGEMA_signal_7131, new_AGEMA_signal_7129}), .b ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, Midori_rounds_sub_sBox_PRINCE_5_n14}), .clk (clk), .r ({Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, Midori_rounds_SR_Result[59]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U16 ( .a ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, Midori_rounds_sub_sBox_PRINCE_5_n11}), .b ({new_AGEMA_signal_7139, new_AGEMA_signal_7137, new_AGEMA_signal_7135}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543]}), .c ({new_AGEMA_signal_2727, new_AGEMA_signal_2726, Midori_rounds_sub_sBox_PRINCE_5_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U12 ( .a ({new_AGEMA_signal_7145, new_AGEMA_signal_7143, new_AGEMA_signal_7141}), .b ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, Midori_rounds_sub_sBox_PRINCE_5_n5}), .clk (clk), .r ({Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, Midori_rounds_SR_Result[57]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U7 ( .a ({new_AGEMA_signal_7139, new_AGEMA_signal_7137, new_AGEMA_signal_7135}), .b ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, Midori_rounds_sub_sBox_PRINCE_5_n2}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549]}), .c ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, Midori_rounds_sub_sBox_PRINCE_5_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U19 ( .a ({new_AGEMA_signal_7151, new_AGEMA_signal_7149, new_AGEMA_signal_7147}), .b ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, Midori_rounds_sub_sBox_PRINCE_6_n14}), .clk (clk), .r ({Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, Midori_rounds_SR_Result[31]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U16 ( .a ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, Midori_rounds_sub_sBox_PRINCE_6_n11}), .b ({new_AGEMA_signal_7157, new_AGEMA_signal_7155, new_AGEMA_signal_7153}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555]}), .c ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, Midori_rounds_sub_sBox_PRINCE_6_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U12 ( .a ({new_AGEMA_signal_7163, new_AGEMA_signal_7161, new_AGEMA_signal_7159}), .b ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, Midori_rounds_sub_sBox_PRINCE_6_n5}), .clk (clk), .r ({Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, Midori_rounds_SR_Result[29]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U7 ( .a ({new_AGEMA_signal_7157, new_AGEMA_signal_7155, new_AGEMA_signal_7153}), .b ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, Midori_rounds_sub_sBox_PRINCE_6_n2}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561]}), .c ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, Midori_rounds_sub_sBox_PRINCE_6_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U19 ( .a ({new_AGEMA_signal_7169, new_AGEMA_signal_7167, new_AGEMA_signal_7165}), .b ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, Midori_rounds_sub_sBox_PRINCE_7_n14}), .clk (clk), .r ({Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, Midori_rounds_SR_Result[3]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U16 ( .a ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, Midori_rounds_sub_sBox_PRINCE_7_n11}), .b ({new_AGEMA_signal_7175, new_AGEMA_signal_7173, new_AGEMA_signal_7171}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567]}), .c ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, Midori_rounds_sub_sBox_PRINCE_7_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U12 ( .a ({new_AGEMA_signal_7181, new_AGEMA_signal_7179, new_AGEMA_signal_7177}), .b ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, Midori_rounds_sub_sBox_PRINCE_7_n5}), .clk (clk), .r ({Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, Midori_rounds_SR_Result[1]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U7 ( .a ({new_AGEMA_signal_7175, new_AGEMA_signal_7173, new_AGEMA_signal_7171}), .b ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, Midori_rounds_sub_sBox_PRINCE_7_n2}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573]}), .c ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, Midori_rounds_sub_sBox_PRINCE_7_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U19 ( .a ({new_AGEMA_signal_7187, new_AGEMA_signal_7185, new_AGEMA_signal_7183}), .b ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, Midori_rounds_sub_sBox_PRINCE_8_n14}), .clk (clk), .r ({Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, Midori_rounds_SR_Result[15]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U16 ( .a ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, Midori_rounds_sub_sBox_PRINCE_8_n11}), .b ({new_AGEMA_signal_7193, new_AGEMA_signal_7191, new_AGEMA_signal_7189}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579]}), .c ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, Midori_rounds_sub_sBox_PRINCE_8_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U12 ( .a ({new_AGEMA_signal_7199, new_AGEMA_signal_7197, new_AGEMA_signal_7195}), .b ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, Midori_rounds_sub_sBox_PRINCE_8_n5}), .clk (clk), .r ({Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, Midori_rounds_SR_Result[13]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U7 ( .a ({new_AGEMA_signal_7193, new_AGEMA_signal_7191, new_AGEMA_signal_7189}), .b ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, Midori_rounds_sub_sBox_PRINCE_8_n2}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585]}), .c ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, Midori_rounds_sub_sBox_PRINCE_8_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U19 ( .a ({new_AGEMA_signal_7205, new_AGEMA_signal_7203, new_AGEMA_signal_7201}), .b ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, Midori_rounds_sub_sBox_PRINCE_9_n14}), .clk (clk), .r ({Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, Midori_rounds_SR_Result[19]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U16 ( .a ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, Midori_rounds_sub_sBox_PRINCE_9_n11}), .b ({new_AGEMA_signal_7211, new_AGEMA_signal_7209, new_AGEMA_signal_7207}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591]}), .c ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, Midori_rounds_sub_sBox_PRINCE_9_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U12 ( .a ({new_AGEMA_signal_7217, new_AGEMA_signal_7215, new_AGEMA_signal_7213}), .b ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, Midori_rounds_sub_sBox_PRINCE_9_n5}), .clk (clk), .r ({Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, Midori_rounds_SR_Result[17]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U7 ( .a ({new_AGEMA_signal_7211, new_AGEMA_signal_7209, new_AGEMA_signal_7207}), .b ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, Midori_rounds_sub_sBox_PRINCE_9_n2}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597]}), .c ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, Midori_rounds_sub_sBox_PRINCE_9_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U19 ( .a ({new_AGEMA_signal_7223, new_AGEMA_signal_7221, new_AGEMA_signal_7219}), .b ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, Midori_rounds_sub_sBox_PRINCE_10_n14}), .clk (clk), .r ({Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, Midori_rounds_SR_Result[55]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U16 ( .a ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, Midori_rounds_sub_sBox_PRINCE_10_n11}), .b ({new_AGEMA_signal_7229, new_AGEMA_signal_7227, new_AGEMA_signal_7225}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603]}), .c ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, Midori_rounds_sub_sBox_PRINCE_10_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U12 ( .a ({new_AGEMA_signal_7235, new_AGEMA_signal_7233, new_AGEMA_signal_7231}), .b ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, Midori_rounds_sub_sBox_PRINCE_10_n5}), .clk (clk), .r ({Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, Midori_rounds_SR_Result[53]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U7 ( .a ({new_AGEMA_signal_7229, new_AGEMA_signal_7227, new_AGEMA_signal_7225}), .b ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, Midori_rounds_sub_sBox_PRINCE_10_n2}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609]}), .c ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, Midori_rounds_sub_sBox_PRINCE_10_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U19 ( .a ({new_AGEMA_signal_7241, new_AGEMA_signal_7239, new_AGEMA_signal_7237}), .b ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, Midori_rounds_sub_sBox_PRINCE_11_n14}), .clk (clk), .r ({Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, Midori_rounds_SR_Result[43]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U16 ( .a ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, Midori_rounds_sub_sBox_PRINCE_11_n11}), .b ({new_AGEMA_signal_7247, new_AGEMA_signal_7245, new_AGEMA_signal_7243}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615]}), .c ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, Midori_rounds_sub_sBox_PRINCE_11_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U12 ( .a ({new_AGEMA_signal_7253, new_AGEMA_signal_7251, new_AGEMA_signal_7249}), .b ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, Midori_rounds_sub_sBox_PRINCE_11_n5}), .clk (clk), .r ({Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, Midori_rounds_SR_Result[41]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U7 ( .a ({new_AGEMA_signal_7247, new_AGEMA_signal_7245, new_AGEMA_signal_7243}), .b ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, Midori_rounds_sub_sBox_PRINCE_11_n2}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621]}), .c ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, Midori_rounds_sub_sBox_PRINCE_11_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U19 ( .a ({new_AGEMA_signal_7259, new_AGEMA_signal_7257, new_AGEMA_signal_7255}), .b ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, Midori_rounds_sub_sBox_PRINCE_12_n14}), .clk (clk), .r ({Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, Midori_rounds_SR_Result[27]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U16 ( .a ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, Midori_rounds_sub_sBox_PRINCE_12_n11}), .b ({new_AGEMA_signal_7265, new_AGEMA_signal_7263, new_AGEMA_signal_7261}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627]}), .c ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, Midori_rounds_sub_sBox_PRINCE_12_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U12 ( .a ({new_AGEMA_signal_7271, new_AGEMA_signal_7269, new_AGEMA_signal_7267}), .b ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, Midori_rounds_sub_sBox_PRINCE_12_n5}), .clk (clk), .r ({Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, Midori_rounds_SR_Result[25]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U7 ( .a ({new_AGEMA_signal_7265, new_AGEMA_signal_7263, new_AGEMA_signal_7261}), .b ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, Midori_rounds_sub_sBox_PRINCE_12_n2}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633]}), .c ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, Midori_rounds_sub_sBox_PRINCE_12_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U19 ( .a ({new_AGEMA_signal_7277, new_AGEMA_signal_7275, new_AGEMA_signal_7273}), .b ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, Midori_rounds_sub_sBox_PRINCE_13_n14}), .clk (clk), .r ({Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, Midori_rounds_SR_Result[7]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U16 ( .a ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, Midori_rounds_sub_sBox_PRINCE_13_n11}), .b ({new_AGEMA_signal_7283, new_AGEMA_signal_7281, new_AGEMA_signal_7279}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639]}), .c ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, Midori_rounds_sub_sBox_PRINCE_13_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U12 ( .a ({new_AGEMA_signal_7289, new_AGEMA_signal_7287, new_AGEMA_signal_7285}), .b ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, Midori_rounds_sub_sBox_PRINCE_13_n5}), .clk (clk), .r ({Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, Midori_rounds_SR_Result[5]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U7 ( .a ({new_AGEMA_signal_7283, new_AGEMA_signal_7281, new_AGEMA_signal_7279}), .b ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, Midori_rounds_sub_sBox_PRINCE_13_n2}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645]}), .c ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, Midori_rounds_sub_sBox_PRINCE_13_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U19 ( .a ({new_AGEMA_signal_7295, new_AGEMA_signal_7293, new_AGEMA_signal_7291}), .b ({new_AGEMA_signal_2815, new_AGEMA_signal_2814, Midori_rounds_sub_sBox_PRINCE_14_n14}), .clk (clk), .r ({Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, Midori_rounds_SR_Result[35]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U16 ( .a ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, Midori_rounds_sub_sBox_PRINCE_14_n11}), .b ({new_AGEMA_signal_7301, new_AGEMA_signal_7299, new_AGEMA_signal_7297}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651]}), .c ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, Midori_rounds_sub_sBox_PRINCE_14_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U12 ( .a ({new_AGEMA_signal_7307, new_AGEMA_signal_7305, new_AGEMA_signal_7303}), .b ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, Midori_rounds_sub_sBox_PRINCE_14_n5}), .clk (clk), .r ({Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, Midori_rounds_SR_Result[33]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U7 ( .a ({new_AGEMA_signal_7301, new_AGEMA_signal_7299, new_AGEMA_signal_7297}), .b ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, Midori_rounds_sub_sBox_PRINCE_14_n2}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657]}), .c ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, Midori_rounds_sub_sBox_PRINCE_14_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U19 ( .a ({new_AGEMA_signal_7313, new_AGEMA_signal_7311, new_AGEMA_signal_7309}), .b ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, Midori_rounds_sub_sBox_PRINCE_15_n14}), .clk (clk), .r ({Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, Midori_rounds_SR_Result[63]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U16 ( .a ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, Midori_rounds_sub_sBox_PRINCE_15_n11}), .b ({new_AGEMA_signal_7319, new_AGEMA_signal_7317, new_AGEMA_signal_7315}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663]}), .c ({new_AGEMA_signal_2827, new_AGEMA_signal_2826, Midori_rounds_sub_sBox_PRINCE_15_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U12 ( .a ({new_AGEMA_signal_7325, new_AGEMA_signal_7323, new_AGEMA_signal_7321}), .b ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, Midori_rounds_sub_sBox_PRINCE_15_n5}), .clk (clk), .r ({Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, Midori_rounds_SR_Result[61]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U7 ( .a ({new_AGEMA_signal_7319, new_AGEMA_signal_7317, new_AGEMA_signal_7315}), .b ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, Midori_rounds_sub_sBox_PRINCE_15_n2}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669]}), .c ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, Midori_rounds_sub_sBox_PRINCE_15_n3}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_1_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, Midori_rounds_SR_Result[1]}), .a ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, Midori_rounds_sub_ResultXORkey[1]}), .c ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, Midori_rounds_mul_input[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_3_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, Midori_rounds_SR_Result[3]}), .a ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, Midori_rounds_sub_ResultXORkey[3]}), .c ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, Midori_rounds_mul_input[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_5_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, Midori_rounds_SR_Result[5]}), .a ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, Midori_rounds_sub_ResultXORkey[5]}), .c ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, Midori_rounds_mul_input[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_7_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, Midori_rounds_SR_Result[7]}), .a ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, Midori_rounds_sub_ResultXORkey[7]}), .c ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, Midori_rounds_mul_input[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_9_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, Midori_rounds_SR_Result[9]}), .a ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, Midori_rounds_sub_ResultXORkey[9]}), .c ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, Midori_rounds_mul_input[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_11_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, Midori_rounds_SR_Result[11]}), .a ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, Midori_rounds_sub_ResultXORkey[11]}), .c ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, Midori_rounds_mul_input[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_13_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, Midori_rounds_SR_Result[13]}), .a ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, Midori_rounds_sub_ResultXORkey[13]}), .c ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, Midori_rounds_mul_input[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_15_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, Midori_rounds_SR_Result[15]}), .a ({new_AGEMA_signal_3175, new_AGEMA_signal_3174, Midori_rounds_sub_ResultXORkey[15]}), .c ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, Midori_rounds_mul_input[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_17_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, Midori_rounds_SR_Result[17]}), .a ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, Midori_rounds_sub_ResultXORkey[17]}), .c ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, Midori_rounds_mul_input[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_19_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, Midori_rounds_SR_Result[19]}), .a ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, Midori_rounds_sub_ResultXORkey[19]}), .c ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, Midori_rounds_mul_input[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_21_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, Midori_rounds_SR_Result[21]}), .a ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, Midori_rounds_sub_ResultXORkey[21]}), .c ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, Midori_rounds_mul_input[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_23_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, Midori_rounds_SR_Result[23]}), .a ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, Midori_rounds_sub_ResultXORkey[23]}), .c ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, Midori_rounds_mul_input[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_25_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, Midori_rounds_SR_Result[25]}), .a ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, Midori_rounds_sub_ResultXORkey[25]}), .c ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, Midori_rounds_mul_input[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_27_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, Midori_rounds_SR_Result[27]}), .a ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, Midori_rounds_sub_ResultXORkey[27]}), .c ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, Midori_rounds_mul_input[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_29_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, Midori_rounds_SR_Result[29]}), .a ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, Midori_rounds_sub_ResultXORkey[29]}), .c ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, Midori_rounds_mul_input[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_31_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, Midori_rounds_SR_Result[31]}), .a ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, Midori_rounds_sub_ResultXORkey[31]}), .c ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, Midori_rounds_mul_input[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_33_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, Midori_rounds_SR_Result[33]}), .a ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, Midori_rounds_sub_ResultXORkey[33]}), .c ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, Midori_rounds_mul_input[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_35_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, Midori_rounds_SR_Result[35]}), .a ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, Midori_rounds_sub_ResultXORkey[35]}), .c ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, Midori_rounds_mul_input[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_37_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, Midori_rounds_SR_Result[37]}), .a ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, Midori_rounds_sub_ResultXORkey[37]}), .c ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, Midori_rounds_mul_input[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_39_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, Midori_rounds_SR_Result[39]}), .a ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, Midori_rounds_sub_ResultXORkey[39]}), .c ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, Midori_rounds_mul_input[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_41_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, Midori_rounds_SR_Result[41]}), .a ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, Midori_rounds_sub_ResultXORkey[41]}), .c ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, Midori_rounds_mul_input[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_43_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, Midori_rounds_SR_Result[43]}), .a ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, Midori_rounds_sub_ResultXORkey[43]}), .c ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, Midori_rounds_mul_input[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_45_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, Midori_rounds_SR_Result[45]}), .a ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, Midori_rounds_sub_ResultXORkey[45]}), .c ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, Midori_rounds_mul_input[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_47_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, Midori_rounds_SR_Result[47]}), .a ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, Midori_rounds_sub_ResultXORkey[47]}), .c ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, Midori_rounds_mul_input[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_49_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, Midori_rounds_SR_Result[49]}), .a ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, Midori_rounds_sub_ResultXORkey[49]}), .c ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, Midori_rounds_mul_input[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_51_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, Midori_rounds_SR_Result[51]}), .a ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, Midori_rounds_sub_ResultXORkey[51]}), .c ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, Midori_rounds_mul_input[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_53_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, Midori_rounds_SR_Result[53]}), .a ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, Midori_rounds_sub_ResultXORkey[53]}), .c ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, Midori_rounds_mul_input[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_55_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, Midori_rounds_SR_Result[55]}), .a ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, Midori_rounds_sub_ResultXORkey[55]}), .c ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, Midori_rounds_mul_input[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_57_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, Midori_rounds_SR_Result[57]}), .a ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, Midori_rounds_sub_ResultXORkey[57]}), .c ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, Midori_rounds_mul_input[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_59_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, Midori_rounds_SR_Result[59]}), .a ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, Midori_rounds_sub_ResultXORkey[59]}), .c ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, Midori_rounds_mul_input[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_61_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, Midori_rounds_SR_Result[61]}), .a ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, Midori_rounds_sub_ResultXORkey[61]}), .c ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, Midori_rounds_mul_input[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_63_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, Midori_rounds_SR_Result[63]}), .a ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, Midori_rounds_sub_ResultXORkey[63]}), .c ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, Midori_rounds_mul_input[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U24 ( .a ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, Midori_rounds_mul_input[61]}), .b ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, Midori_rounds_mul_MC1_n8}), .c ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, Midori_rounds_SR_Inv_Result[21]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U22 ( .a ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, Midori_rounds_mul_input[51]}), .b ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, Midori_rounds_mul_MC1_n6}), .c ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, Midori_rounds_SR_Inv_Result[43]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U20 ( .a ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, Midori_rounds_mul_input[49]}), .b ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, Midori_rounds_mul_MC1_n4}), .c ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, Midori_rounds_SR_Inv_Result[41]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U18 ( .a ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, Midori_rounds_mul_input[55]}), .b ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, Midori_rounds_mul_MC1_n6}), .c ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, Midori_rounds_SR_Inv_Result[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U17 ( .a ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, Midori_rounds_mul_input[63]}), .b ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, Midori_rounds_mul_input[59]}), .c ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, Midori_rounds_mul_MC1_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U14 ( .a ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, Midori_rounds_mul_input[53]}), .b ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, Midori_rounds_mul_MC1_n4}), .c ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, Midori_rounds_SR_Inv_Result[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U13 ( .a ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, Midori_rounds_mul_input[57]}), .b ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, Midori_rounds_mul_input[61]}), .c ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, Midori_rounds_mul_MC1_n4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U12 ( .a ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, Midori_rounds_mul_input[59]}), .b ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, Midori_rounds_mul_MC1_n2}), .c ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, Midori_rounds_SR_Inv_Result[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U10 ( .a ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, Midori_rounds_mul_input[57]}), .b ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, Midori_rounds_mul_MC1_n8}), .c ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, Midori_rounds_SR_Inv_Result[61]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U9 ( .a ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, Midori_rounds_mul_input[49]}), .b ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, Midori_rounds_mul_input[53]}), .c ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, Midori_rounds_mul_MC1_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U6 ( .a ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, Midori_rounds_mul_input[63]}), .b ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, Midori_rounds_mul_MC1_n2}), .c ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, Midori_rounds_SR_Inv_Result[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U5 ( .a ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, Midori_rounds_mul_input[51]}), .b ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, Midori_rounds_mul_input[55]}), .c ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, Midori_rounds_mul_MC1_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U24 ( .a ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, Midori_rounds_mul_input[45]}), .b ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, Midori_rounds_mul_MC2_n8}), .c ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, Midori_rounds_SR_Inv_Result[45]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U22 ( .a ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, Midori_rounds_mul_input[35]}), .b ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, Midori_rounds_mul_MC2_n6}), .c ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, Midori_rounds_SR_Inv_Result[19]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U20 ( .a ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, Midori_rounds_mul_input[33]}), .b ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, Midori_rounds_mul_MC2_n4}), .c ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, Midori_rounds_SR_Inv_Result[17]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U18 ( .a ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, Midori_rounds_mul_input[39]}), .b ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, Midori_rounds_mul_MC2_n6}), .c ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, Midori_rounds_SR_Inv_Result[59]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U17 ( .a ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, Midori_rounds_mul_input[47]}), .b ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, Midori_rounds_mul_input[43]}), .c ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, Midori_rounds_mul_MC2_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U14 ( .a ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, Midori_rounds_mul_input[37]}), .b ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, Midori_rounds_mul_MC2_n4}), .c ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, Midori_rounds_SR_Inv_Result[57]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U13 ( .a ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, Midori_rounds_mul_input[41]}), .b ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, Midori_rounds_mul_input[45]}), .c ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, Midori_rounds_mul_MC2_n4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U12 ( .a ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, Midori_rounds_mul_input[43]}), .b ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, Midori_rounds_mul_MC2_n2}), .c ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, Midori_rounds_SR_Inv_Result[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U10 ( .a ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, Midori_rounds_mul_input[41]}), .b ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, Midori_rounds_mul_MC2_n8}), .c ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, Midori_rounds_SR_Inv_Result[5]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U9 ( .a ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, Midori_rounds_mul_input[33]}), .b ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, Midori_rounds_mul_input[37]}), .c ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, Midori_rounds_mul_MC2_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U6 ( .a ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, Midori_rounds_mul_input[47]}), .b ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, Midori_rounds_mul_MC2_n2}), .c ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, Midori_rounds_SR_Inv_Result[47]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U5 ( .a ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, Midori_rounds_mul_input[35]}), .b ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, Midori_rounds_mul_input[39]}), .c ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, Midori_rounds_mul_MC2_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U24 ( .a ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, Midori_rounds_mul_input[29]}), .b ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, Midori_rounds_mul_MC3_n8}), .c ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, Midori_rounds_SR_Inv_Result[49]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U22 ( .a ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, Midori_rounds_mul_input[19]}), .b ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, Midori_rounds_mul_MC3_n6}), .c ({new_AGEMA_signal_3379, new_AGEMA_signal_3378, Midori_rounds_SR_Inv_Result[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U20 ( .a ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, Midori_rounds_mul_input[17]}), .b ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, Midori_rounds_mul_MC3_n4}), .c ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, Midori_rounds_SR_Inv_Result[13]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U18 ( .a ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, Midori_rounds_mul_input[23]}), .b ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, Midori_rounds_mul_MC3_n6}), .c ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, Midori_rounds_SR_Inv_Result[39]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U17 ( .a ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, Midori_rounds_mul_input[31]}), .b ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, Midori_rounds_mul_input[27]}), .c ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, Midori_rounds_mul_MC3_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U14 ( .a ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, Midori_rounds_mul_input[21]}), .b ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, Midori_rounds_mul_MC3_n4}), .c ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, Midori_rounds_SR_Inv_Result[37]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U13 ( .a ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, Midori_rounds_mul_input[25]}), .b ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, Midori_rounds_mul_input[29]}), .c ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, Midori_rounds_mul_MC3_n4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U12 ( .a ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, Midori_rounds_mul_input[27]}), .b ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, Midori_rounds_mul_MC3_n2}), .c ({new_AGEMA_signal_3391, new_AGEMA_signal_3390, Midori_rounds_SR_Inv_Result[27]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U10 ( .a ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, Midori_rounds_mul_input[25]}), .b ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, Midori_rounds_mul_MC3_n8}), .c ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, Midori_rounds_SR_Inv_Result[25]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U9 ( .a ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, Midori_rounds_mul_input[17]}), .b ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, Midori_rounds_mul_input[21]}), .c ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, Midori_rounds_mul_MC3_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U6 ( .a ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, Midori_rounds_mul_input[31]}), .b ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, Midori_rounds_mul_MC3_n2}), .c ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, Midori_rounds_SR_Inv_Result[51]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U5 ( .a ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, Midori_rounds_mul_input[19]}), .b ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, Midori_rounds_mul_input[23]}), .c ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, Midori_rounds_mul_MC3_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U24 ( .a ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, Midori_rounds_mul_input[13]}), .b ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, Midori_rounds_mul_MC4_n8}), .c ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, Midori_rounds_SR_Inv_Result[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U22 ( .a ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, Midori_rounds_mul_input[3]}), .b ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, Midori_rounds_mul_MC4_n6}), .c ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, Midori_rounds_SR_Inv_Result[55]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U20 ( .a ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, Midori_rounds_mul_input[1]}), .b ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, Midori_rounds_mul_MC4_n4}), .c ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, Midori_rounds_SR_Inv_Result[53]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U18 ( .a ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, Midori_rounds_mul_input[7]}), .b ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, Midori_rounds_mul_MC4_n6}), .c ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, Midori_rounds_SR_Inv_Result[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U17 ( .a ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, Midori_rounds_mul_input[15]}), .b ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, Midori_rounds_mul_input[11]}), .c ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, Midori_rounds_mul_MC4_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U14 ( .a ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, Midori_rounds_mul_input[5]}), .b ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, Midori_rounds_mul_MC4_n4}), .c ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, Midori_rounds_SR_Inv_Result[29]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U13 ( .a ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, Midori_rounds_mul_input[9]}), .b ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, Midori_rounds_mul_input[13]}), .c ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, Midori_rounds_mul_MC4_n4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U12 ( .a ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, Midori_rounds_mul_input[11]}), .b ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, Midori_rounds_mul_MC4_n2}), .c ({new_AGEMA_signal_3415, new_AGEMA_signal_3414, Midori_rounds_SR_Inv_Result[35]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U10 ( .a ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, Midori_rounds_mul_input[9]}), .b ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, Midori_rounds_mul_MC4_n8}), .c ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, Midori_rounds_SR_Inv_Result[33]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U9 ( .a ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, Midori_rounds_mul_input[1]}), .b ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, Midori_rounds_mul_input[5]}), .c ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, Midori_rounds_mul_MC4_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U6 ( .a ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, Midori_rounds_mul_input[15]}), .b ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, Midori_rounds_mul_MC4_n2}), .c ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, Midori_rounds_SR_Inv_Result[11]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U5 ( .a ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, Midori_rounds_mul_input[3]}), .b ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, Midori_rounds_mul_input[7]}), .c ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, Midori_rounds_mul_MC4_n2}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_1_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3511, new_AGEMA_signal_3510, Midori_rounds_mul_ResultXORkey[1]}), .a ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, Midori_rounds_SR_Inv_Result[1]}), .c ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, Midori_rounds_round_Result[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_3_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, Midori_rounds_mul_ResultXORkey[3]}), .a ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, Midori_rounds_SR_Inv_Result[3]}), .c ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, Midori_rounds_round_Result[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_5_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3439, new_AGEMA_signal_3438, Midori_rounds_mul_ResultXORkey[5]}), .a ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, Midori_rounds_SR_Inv_Result[5]}), .c ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, Midori_rounds_round_Result[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_7_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, Midori_rounds_mul_ResultXORkey[7]}), .a ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, Midori_rounds_SR_Inv_Result[7]}), .c ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, Midori_rounds_round_Result[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_9_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, Midori_rounds_mul_ResultXORkey[9]}), .a ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, Midori_rounds_SR_Inv_Result[9]}), .c ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, Midori_rounds_round_Result[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_11_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, Midori_rounds_mul_ResultXORkey[11]}), .a ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, Midori_rounds_SR_Inv_Result[11]}), .c ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, Midori_rounds_round_Result[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_13_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3523, new_AGEMA_signal_3522, Midori_rounds_mul_ResultXORkey[13]}), .a ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, Midori_rounds_SR_Inv_Result[13]}), .c ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, Midori_rounds_round_Result[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_15_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3519, new_AGEMA_signal_3518, Midori_rounds_mul_ResultXORkey[15]}), .a ({new_AGEMA_signal_3379, new_AGEMA_signal_3378, Midori_rounds_SR_Inv_Result[15]}), .c ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, Midori_rounds_round_Result[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_17_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3517, new_AGEMA_signal_3516, Midori_rounds_mul_ResultXORkey[17]}), .a ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, Midori_rounds_SR_Inv_Result[17]}), .c ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, Midori_rounds_round_Result[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_19_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, Midori_rounds_mul_ResultXORkey[19]}), .a ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, Midori_rounds_SR_Inv_Result[19]}), .c ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, Midori_rounds_round_Result[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_21_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, Midori_rounds_mul_ResultXORkey[21]}), .a ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, Midori_rounds_SR_Inv_Result[21]}), .c ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, Midori_rounds_round_Result[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_23_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, Midori_rounds_mul_ResultXORkey[23]}), .a ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, Midori_rounds_SR_Inv_Result[23]}), .c ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, Midori_rounds_round_Result[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_25_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, Midori_rounds_mul_ResultXORkey[25]}), .a ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, Midori_rounds_SR_Inv_Result[25]}), .c ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, Midori_rounds_round_Result[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_27_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, Midori_rounds_mul_ResultXORkey[27]}), .a ({new_AGEMA_signal_3391, new_AGEMA_signal_3390, Midori_rounds_SR_Inv_Result[27]}), .c ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, Midori_rounds_round_Result[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_29_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, Midori_rounds_mul_ResultXORkey[29]}), .a ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, Midori_rounds_SR_Inv_Result[29]}), .c ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, Midori_rounds_round_Result[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_31_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, Midori_rounds_mul_ResultXORkey[31]}), .a ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, Midori_rounds_SR_Inv_Result[31]}), .c ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, Midori_rounds_round_Result[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_33_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3487, new_AGEMA_signal_3486, Midori_rounds_mul_ResultXORkey[33]}), .a ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, Midori_rounds_SR_Inv_Result[33]}), .c ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, Midori_rounds_round_Result[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_35_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3483, new_AGEMA_signal_3482, Midori_rounds_mul_ResultXORkey[35]}), .a ({new_AGEMA_signal_3415, new_AGEMA_signal_3414, Midori_rounds_SR_Inv_Result[35]}), .c ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, Midori_rounds_round_Result[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_37_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, Midori_rounds_mul_ResultXORkey[37]}), .a ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, Midori_rounds_SR_Inv_Result[37]}), .c ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, Midori_rounds_round_Result[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_39_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, Midori_rounds_mul_ResultXORkey[39]}), .a ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, Midori_rounds_SR_Inv_Result[39]}), .c ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, Midori_rounds_round_Result[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_41_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3471, new_AGEMA_signal_3470, Midori_rounds_mul_ResultXORkey[41]}), .a ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, Midori_rounds_SR_Inv_Result[41]}), .c ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, Midori_rounds_round_Result[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_43_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, Midori_rounds_mul_ResultXORkey[43]}), .a ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, Midori_rounds_SR_Inv_Result[43]}), .c ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, Midori_rounds_round_Result[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_45_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, Midori_rounds_mul_ResultXORkey[45]}), .a ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, Midori_rounds_SR_Inv_Result[45]}), .c ({new_AGEMA_signal_3623, new_AGEMA_signal_3622, Midori_rounds_round_Result[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_47_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, Midori_rounds_mul_ResultXORkey[47]}), .a ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, Midori_rounds_SR_Inv_Result[47]}), .c ({new_AGEMA_signal_3627, new_AGEMA_signal_3626, Midori_rounds_round_Result[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_49_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, Midori_rounds_mul_ResultXORkey[49]}), .a ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, Midori_rounds_SR_Inv_Result[49]}), .c ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, Midori_rounds_round_Result[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_51_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, Midori_rounds_mul_ResultXORkey[51]}), .a ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, Midori_rounds_SR_Inv_Result[51]}), .c ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, Midori_rounds_round_Result[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_53_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3451, new_AGEMA_signal_3450, Midori_rounds_mul_ResultXORkey[53]}), .a ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, Midori_rounds_SR_Inv_Result[53]}), .c ({new_AGEMA_signal_3635, new_AGEMA_signal_3634, Midori_rounds_round_Result[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_55_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, Midori_rounds_mul_ResultXORkey[55]}), .a ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, Midori_rounds_SR_Inv_Result[55]}), .c ({new_AGEMA_signal_3639, new_AGEMA_signal_3638, Midori_rounds_round_Result[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_57_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, Midori_rounds_mul_ResultXORkey[57]}), .a ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, Midori_rounds_SR_Inv_Result[57]}), .c ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, Midori_rounds_round_Result[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_59_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, Midori_rounds_mul_ResultXORkey[59]}), .a ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, Midori_rounds_SR_Inv_Result[59]}), .c ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, Midori_rounds_round_Result[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_61_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, Midori_rounds_mul_ResultXORkey[61]}), .a ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, Midori_rounds_SR_Inv_Result[61]}), .c ({new_AGEMA_signal_3647, new_AGEMA_signal_3646, Midori_rounds_round_Result[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_63_U1 ( .s (new_AGEMA_signal_7331), .b ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, Midori_rounds_mul_ResultXORkey[63]}), .a ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, Midori_rounds_SR_Inv_Result[63]}), .c ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, Midori_rounds_round_Result[63]}) ) ;
    buf_clk new_AGEMA_reg_buffer_1324 ( .C (clk), .D (new_AGEMA_signal_4789), .Q (new_AGEMA_signal_4790) ) ;
    buf_clk new_AGEMA_reg_buffer_1844 ( .C (clk), .D (new_AGEMA_signal_5308), .Q (new_AGEMA_signal_5309) ) ;
    buf_clk new_AGEMA_reg_buffer_1850 ( .C (clk), .D (new_AGEMA_signal_5314), .Q (new_AGEMA_signal_5315) ) ;
    buf_clk new_AGEMA_reg_buffer_1856 ( .C (clk), .D (new_AGEMA_signal_5320), .Q (new_AGEMA_signal_5321) ) ;
    buf_clk new_AGEMA_reg_buffer_1862 ( .C (clk), .D (new_AGEMA_signal_5326), .Q (new_AGEMA_signal_5327) ) ;
    buf_clk new_AGEMA_reg_buffer_1868 ( .C (clk), .D (new_AGEMA_signal_5332), .Q (new_AGEMA_signal_5333) ) ;
    buf_clk new_AGEMA_reg_buffer_1874 ( .C (clk), .D (new_AGEMA_signal_5338), .Q (new_AGEMA_signal_5339) ) ;
    buf_clk new_AGEMA_reg_buffer_1880 ( .C (clk), .D (new_AGEMA_signal_5344), .Q (new_AGEMA_signal_5345) ) ;
    buf_clk new_AGEMA_reg_buffer_1886 ( .C (clk), .D (new_AGEMA_signal_5350), .Q (new_AGEMA_signal_5351) ) ;
    buf_clk new_AGEMA_reg_buffer_1892 ( .C (clk), .D (new_AGEMA_signal_5356), .Q (new_AGEMA_signal_5357) ) ;
    buf_clk new_AGEMA_reg_buffer_1898 ( .C (clk), .D (new_AGEMA_signal_5362), .Q (new_AGEMA_signal_5363) ) ;
    buf_clk new_AGEMA_reg_buffer_1904 ( .C (clk), .D (new_AGEMA_signal_5368), .Q (new_AGEMA_signal_5369) ) ;
    buf_clk new_AGEMA_reg_buffer_1910 ( .C (clk), .D (new_AGEMA_signal_5374), .Q (new_AGEMA_signal_5375) ) ;
    buf_clk new_AGEMA_reg_buffer_1916 ( .C (clk), .D (new_AGEMA_signal_5380), .Q (new_AGEMA_signal_5381) ) ;
    buf_clk new_AGEMA_reg_buffer_1922 ( .C (clk), .D (new_AGEMA_signal_5386), .Q (new_AGEMA_signal_5387) ) ;
    buf_clk new_AGEMA_reg_buffer_1928 ( .C (clk), .D (new_AGEMA_signal_5392), .Q (new_AGEMA_signal_5393) ) ;
    buf_clk new_AGEMA_reg_buffer_1934 ( .C (clk), .D (new_AGEMA_signal_5398), .Q (new_AGEMA_signal_5399) ) ;
    buf_clk new_AGEMA_reg_buffer_1940 ( .C (clk), .D (new_AGEMA_signal_5404), .Q (new_AGEMA_signal_5405) ) ;
    buf_clk new_AGEMA_reg_buffer_1946 ( .C (clk), .D (new_AGEMA_signal_5410), .Q (new_AGEMA_signal_5411) ) ;
    buf_clk new_AGEMA_reg_buffer_1952 ( .C (clk), .D (new_AGEMA_signal_5416), .Q (new_AGEMA_signal_5417) ) ;
    buf_clk new_AGEMA_reg_buffer_1958 ( .C (clk), .D (new_AGEMA_signal_5422), .Q (new_AGEMA_signal_5423) ) ;
    buf_clk new_AGEMA_reg_buffer_1964 ( .C (clk), .D (new_AGEMA_signal_5428), .Q (new_AGEMA_signal_5429) ) ;
    buf_clk new_AGEMA_reg_buffer_1970 ( .C (clk), .D (new_AGEMA_signal_5434), .Q (new_AGEMA_signal_5435) ) ;
    buf_clk new_AGEMA_reg_buffer_1976 ( .C (clk), .D (new_AGEMA_signal_5440), .Q (new_AGEMA_signal_5441) ) ;
    buf_clk new_AGEMA_reg_buffer_1982 ( .C (clk), .D (new_AGEMA_signal_5446), .Q (new_AGEMA_signal_5447) ) ;
    buf_clk new_AGEMA_reg_buffer_1988 ( .C (clk), .D (new_AGEMA_signal_5452), .Q (new_AGEMA_signal_5453) ) ;
    buf_clk new_AGEMA_reg_buffer_1994 ( .C (clk), .D (new_AGEMA_signal_5458), .Q (new_AGEMA_signal_5459) ) ;
    buf_clk new_AGEMA_reg_buffer_2000 ( .C (clk), .D (new_AGEMA_signal_5464), .Q (new_AGEMA_signal_5465) ) ;
    buf_clk new_AGEMA_reg_buffer_2006 ( .C (clk), .D (new_AGEMA_signal_5470), .Q (new_AGEMA_signal_5471) ) ;
    buf_clk new_AGEMA_reg_buffer_2012 ( .C (clk), .D (new_AGEMA_signal_5476), .Q (new_AGEMA_signal_5477) ) ;
    buf_clk new_AGEMA_reg_buffer_2018 ( .C (clk), .D (new_AGEMA_signal_5482), .Q (new_AGEMA_signal_5483) ) ;
    buf_clk new_AGEMA_reg_buffer_2024 ( .C (clk), .D (new_AGEMA_signal_5488), .Q (new_AGEMA_signal_5489) ) ;
    buf_clk new_AGEMA_reg_buffer_2030 ( .C (clk), .D (new_AGEMA_signal_5494), .Q (new_AGEMA_signal_5495) ) ;
    buf_clk new_AGEMA_reg_buffer_2036 ( .C (clk), .D (new_AGEMA_signal_5500), .Q (new_AGEMA_signal_5501) ) ;
    buf_clk new_AGEMA_reg_buffer_2042 ( .C (clk), .D (new_AGEMA_signal_5506), .Q (new_AGEMA_signal_5507) ) ;
    buf_clk new_AGEMA_reg_buffer_2048 ( .C (clk), .D (new_AGEMA_signal_5512), .Q (new_AGEMA_signal_5513) ) ;
    buf_clk new_AGEMA_reg_buffer_2054 ( .C (clk), .D (new_AGEMA_signal_5518), .Q (new_AGEMA_signal_5519) ) ;
    buf_clk new_AGEMA_reg_buffer_2060 ( .C (clk), .D (new_AGEMA_signal_5524), .Q (new_AGEMA_signal_5525) ) ;
    buf_clk new_AGEMA_reg_buffer_2066 ( .C (clk), .D (new_AGEMA_signal_5530), .Q (new_AGEMA_signal_5531) ) ;
    buf_clk new_AGEMA_reg_buffer_2072 ( .C (clk), .D (new_AGEMA_signal_5536), .Q (new_AGEMA_signal_5537) ) ;
    buf_clk new_AGEMA_reg_buffer_2078 ( .C (clk), .D (new_AGEMA_signal_5542), .Q (new_AGEMA_signal_5543) ) ;
    buf_clk new_AGEMA_reg_buffer_2084 ( .C (clk), .D (new_AGEMA_signal_5548), .Q (new_AGEMA_signal_5549) ) ;
    buf_clk new_AGEMA_reg_buffer_2090 ( .C (clk), .D (new_AGEMA_signal_5554), .Q (new_AGEMA_signal_5555) ) ;
    buf_clk new_AGEMA_reg_buffer_2096 ( .C (clk), .D (new_AGEMA_signal_5560), .Q (new_AGEMA_signal_5561) ) ;
    buf_clk new_AGEMA_reg_buffer_2102 ( .C (clk), .D (new_AGEMA_signal_5566), .Q (new_AGEMA_signal_5567) ) ;
    buf_clk new_AGEMA_reg_buffer_2108 ( .C (clk), .D (new_AGEMA_signal_5572), .Q (new_AGEMA_signal_5573) ) ;
    buf_clk new_AGEMA_reg_buffer_2114 ( .C (clk), .D (new_AGEMA_signal_5578), .Q (new_AGEMA_signal_5579) ) ;
    buf_clk new_AGEMA_reg_buffer_2120 ( .C (clk), .D (new_AGEMA_signal_5584), .Q (new_AGEMA_signal_5585) ) ;
    buf_clk new_AGEMA_reg_buffer_2126 ( .C (clk), .D (new_AGEMA_signal_5590), .Q (new_AGEMA_signal_5591) ) ;
    buf_clk new_AGEMA_reg_buffer_2132 ( .C (clk), .D (new_AGEMA_signal_5596), .Q (new_AGEMA_signal_5597) ) ;
    buf_clk new_AGEMA_reg_buffer_2138 ( .C (clk), .D (new_AGEMA_signal_5602), .Q (new_AGEMA_signal_5603) ) ;
    buf_clk new_AGEMA_reg_buffer_2144 ( .C (clk), .D (new_AGEMA_signal_5608), .Q (new_AGEMA_signal_5609) ) ;
    buf_clk new_AGEMA_reg_buffer_2150 ( .C (clk), .D (new_AGEMA_signal_5614), .Q (new_AGEMA_signal_5615) ) ;
    buf_clk new_AGEMA_reg_buffer_2156 ( .C (clk), .D (new_AGEMA_signal_5620), .Q (new_AGEMA_signal_5621) ) ;
    buf_clk new_AGEMA_reg_buffer_2162 ( .C (clk), .D (new_AGEMA_signal_5626), .Q (new_AGEMA_signal_5627) ) ;
    buf_clk new_AGEMA_reg_buffer_2168 ( .C (clk), .D (new_AGEMA_signal_5632), .Q (new_AGEMA_signal_5633) ) ;
    buf_clk new_AGEMA_reg_buffer_2174 ( .C (clk), .D (new_AGEMA_signal_5638), .Q (new_AGEMA_signal_5639) ) ;
    buf_clk new_AGEMA_reg_buffer_2180 ( .C (clk), .D (new_AGEMA_signal_5644), .Q (new_AGEMA_signal_5645) ) ;
    buf_clk new_AGEMA_reg_buffer_2186 ( .C (clk), .D (new_AGEMA_signal_5650), .Q (new_AGEMA_signal_5651) ) ;
    buf_clk new_AGEMA_reg_buffer_2192 ( .C (clk), .D (new_AGEMA_signal_5656), .Q (new_AGEMA_signal_5657) ) ;
    buf_clk new_AGEMA_reg_buffer_2198 ( .C (clk), .D (new_AGEMA_signal_5662), .Q (new_AGEMA_signal_5663) ) ;
    buf_clk new_AGEMA_reg_buffer_2204 ( .C (clk), .D (new_AGEMA_signal_5668), .Q (new_AGEMA_signal_5669) ) ;
    buf_clk new_AGEMA_reg_buffer_2210 ( .C (clk), .D (new_AGEMA_signal_5674), .Q (new_AGEMA_signal_5675) ) ;
    buf_clk new_AGEMA_reg_buffer_2216 ( .C (clk), .D (new_AGEMA_signal_5680), .Q (new_AGEMA_signal_5681) ) ;
    buf_clk new_AGEMA_reg_buffer_2222 ( .C (clk), .D (new_AGEMA_signal_5686), .Q (new_AGEMA_signal_5687) ) ;
    buf_clk new_AGEMA_reg_buffer_2228 ( .C (clk), .D (new_AGEMA_signal_5692), .Q (new_AGEMA_signal_5693) ) ;
    buf_clk new_AGEMA_reg_buffer_2234 ( .C (clk), .D (new_AGEMA_signal_5698), .Q (new_AGEMA_signal_5699) ) ;
    buf_clk new_AGEMA_reg_buffer_2240 ( .C (clk), .D (new_AGEMA_signal_5704), .Q (new_AGEMA_signal_5705) ) ;
    buf_clk new_AGEMA_reg_buffer_2246 ( .C (clk), .D (new_AGEMA_signal_5710), .Q (new_AGEMA_signal_5711) ) ;
    buf_clk new_AGEMA_reg_buffer_2252 ( .C (clk), .D (new_AGEMA_signal_5716), .Q (new_AGEMA_signal_5717) ) ;
    buf_clk new_AGEMA_reg_buffer_2258 ( .C (clk), .D (new_AGEMA_signal_5722), .Q (new_AGEMA_signal_5723) ) ;
    buf_clk new_AGEMA_reg_buffer_2264 ( .C (clk), .D (new_AGEMA_signal_5728), .Q (new_AGEMA_signal_5729) ) ;
    buf_clk new_AGEMA_reg_buffer_2270 ( .C (clk), .D (new_AGEMA_signal_5734), .Q (new_AGEMA_signal_5735) ) ;
    buf_clk new_AGEMA_reg_buffer_2276 ( .C (clk), .D (new_AGEMA_signal_5740), .Q (new_AGEMA_signal_5741) ) ;
    buf_clk new_AGEMA_reg_buffer_2282 ( .C (clk), .D (new_AGEMA_signal_5746), .Q (new_AGEMA_signal_5747) ) ;
    buf_clk new_AGEMA_reg_buffer_2288 ( .C (clk), .D (new_AGEMA_signal_5752), .Q (new_AGEMA_signal_5753) ) ;
    buf_clk new_AGEMA_reg_buffer_2294 ( .C (clk), .D (new_AGEMA_signal_5758), .Q (new_AGEMA_signal_5759) ) ;
    buf_clk new_AGEMA_reg_buffer_2300 ( .C (clk), .D (new_AGEMA_signal_5764), .Q (new_AGEMA_signal_5765) ) ;
    buf_clk new_AGEMA_reg_buffer_2306 ( .C (clk), .D (new_AGEMA_signal_5770), .Q (new_AGEMA_signal_5771) ) ;
    buf_clk new_AGEMA_reg_buffer_2312 ( .C (clk), .D (new_AGEMA_signal_5776), .Q (new_AGEMA_signal_5777) ) ;
    buf_clk new_AGEMA_reg_buffer_2318 ( .C (clk), .D (new_AGEMA_signal_5782), .Q (new_AGEMA_signal_5783) ) ;
    buf_clk new_AGEMA_reg_buffer_2324 ( .C (clk), .D (new_AGEMA_signal_5788), .Q (new_AGEMA_signal_5789) ) ;
    buf_clk new_AGEMA_reg_buffer_2330 ( .C (clk), .D (new_AGEMA_signal_5794), .Q (new_AGEMA_signal_5795) ) ;
    buf_clk new_AGEMA_reg_buffer_2336 ( .C (clk), .D (new_AGEMA_signal_5800), .Q (new_AGEMA_signal_5801) ) ;
    buf_clk new_AGEMA_reg_buffer_2342 ( .C (clk), .D (new_AGEMA_signal_5806), .Q (new_AGEMA_signal_5807) ) ;
    buf_clk new_AGEMA_reg_buffer_2348 ( .C (clk), .D (new_AGEMA_signal_5812), .Q (new_AGEMA_signal_5813) ) ;
    buf_clk new_AGEMA_reg_buffer_2354 ( .C (clk), .D (new_AGEMA_signal_5818), .Q (new_AGEMA_signal_5819) ) ;
    buf_clk new_AGEMA_reg_buffer_2360 ( .C (clk), .D (new_AGEMA_signal_5824), .Q (new_AGEMA_signal_5825) ) ;
    buf_clk new_AGEMA_reg_buffer_2366 ( .C (clk), .D (new_AGEMA_signal_5830), .Q (new_AGEMA_signal_5831) ) ;
    buf_clk new_AGEMA_reg_buffer_2372 ( .C (clk), .D (new_AGEMA_signal_5836), .Q (new_AGEMA_signal_5837) ) ;
    buf_clk new_AGEMA_reg_buffer_2378 ( .C (clk), .D (new_AGEMA_signal_5842), .Q (new_AGEMA_signal_5843) ) ;
    buf_clk new_AGEMA_reg_buffer_2384 ( .C (clk), .D (new_AGEMA_signal_5848), .Q (new_AGEMA_signal_5849) ) ;
    buf_clk new_AGEMA_reg_buffer_2390 ( .C (clk), .D (new_AGEMA_signal_5854), .Q (new_AGEMA_signal_5855) ) ;
    buf_clk new_AGEMA_reg_buffer_2396 ( .C (clk), .D (new_AGEMA_signal_5860), .Q (new_AGEMA_signal_5861) ) ;
    buf_clk new_AGEMA_reg_buffer_2402 ( .C (clk), .D (new_AGEMA_signal_5866), .Q (new_AGEMA_signal_5867) ) ;
    buf_clk new_AGEMA_reg_buffer_2408 ( .C (clk), .D (new_AGEMA_signal_5872), .Q (new_AGEMA_signal_5873) ) ;
    buf_clk new_AGEMA_reg_buffer_2414 ( .C (clk), .D (new_AGEMA_signal_5878), .Q (new_AGEMA_signal_5879) ) ;
    buf_clk new_AGEMA_reg_buffer_2420 ( .C (clk), .D (new_AGEMA_signal_5884), .Q (new_AGEMA_signal_5885) ) ;
    buf_clk new_AGEMA_reg_buffer_2426 ( .C (clk), .D (new_AGEMA_signal_5890), .Q (new_AGEMA_signal_5891) ) ;
    buf_clk new_AGEMA_reg_buffer_2432 ( .C (clk), .D (new_AGEMA_signal_5896), .Q (new_AGEMA_signal_5897) ) ;
    buf_clk new_AGEMA_reg_buffer_2438 ( .C (clk), .D (new_AGEMA_signal_5902), .Q (new_AGEMA_signal_5903) ) ;
    buf_clk new_AGEMA_reg_buffer_2444 ( .C (clk), .D (new_AGEMA_signal_5908), .Q (new_AGEMA_signal_5909) ) ;
    buf_clk new_AGEMA_reg_buffer_2450 ( .C (clk), .D (new_AGEMA_signal_5914), .Q (new_AGEMA_signal_5915) ) ;
    buf_clk new_AGEMA_reg_buffer_2456 ( .C (clk), .D (new_AGEMA_signal_5920), .Q (new_AGEMA_signal_5921) ) ;
    buf_clk new_AGEMA_reg_buffer_2462 ( .C (clk), .D (new_AGEMA_signal_5926), .Q (new_AGEMA_signal_5927) ) ;
    buf_clk new_AGEMA_reg_buffer_2468 ( .C (clk), .D (new_AGEMA_signal_5932), .Q (new_AGEMA_signal_5933) ) ;
    buf_clk new_AGEMA_reg_buffer_2474 ( .C (clk), .D (new_AGEMA_signal_5938), .Q (new_AGEMA_signal_5939) ) ;
    buf_clk new_AGEMA_reg_buffer_2480 ( .C (clk), .D (new_AGEMA_signal_5944), .Q (new_AGEMA_signal_5945) ) ;
    buf_clk new_AGEMA_reg_buffer_2486 ( .C (clk), .D (new_AGEMA_signal_5950), .Q (new_AGEMA_signal_5951) ) ;
    buf_clk new_AGEMA_reg_buffer_2492 ( .C (clk), .D (new_AGEMA_signal_5956), .Q (new_AGEMA_signal_5957) ) ;
    buf_clk new_AGEMA_reg_buffer_2498 ( .C (clk), .D (new_AGEMA_signal_5962), .Q (new_AGEMA_signal_5963) ) ;
    buf_clk new_AGEMA_reg_buffer_2504 ( .C (clk), .D (new_AGEMA_signal_5968), .Q (new_AGEMA_signal_5969) ) ;
    buf_clk new_AGEMA_reg_buffer_2510 ( .C (clk), .D (new_AGEMA_signal_5974), .Q (new_AGEMA_signal_5975) ) ;
    buf_clk new_AGEMA_reg_buffer_2516 ( .C (clk), .D (new_AGEMA_signal_5980), .Q (new_AGEMA_signal_5981) ) ;
    buf_clk new_AGEMA_reg_buffer_2522 ( .C (clk), .D (new_AGEMA_signal_5986), .Q (new_AGEMA_signal_5987) ) ;
    buf_clk new_AGEMA_reg_buffer_2528 ( .C (clk), .D (new_AGEMA_signal_5992), .Q (new_AGEMA_signal_5993) ) ;
    buf_clk new_AGEMA_reg_buffer_2534 ( .C (clk), .D (new_AGEMA_signal_5998), .Q (new_AGEMA_signal_5999) ) ;
    buf_clk new_AGEMA_reg_buffer_2540 ( .C (clk), .D (new_AGEMA_signal_6004), .Q (new_AGEMA_signal_6005) ) ;
    buf_clk new_AGEMA_reg_buffer_2546 ( .C (clk), .D (new_AGEMA_signal_6010), .Q (new_AGEMA_signal_6011) ) ;
    buf_clk new_AGEMA_reg_buffer_2552 ( .C (clk), .D (new_AGEMA_signal_6016), .Q (new_AGEMA_signal_6017) ) ;
    buf_clk new_AGEMA_reg_buffer_2558 ( .C (clk), .D (new_AGEMA_signal_6022), .Q (new_AGEMA_signal_6023) ) ;
    buf_clk new_AGEMA_reg_buffer_2564 ( .C (clk), .D (new_AGEMA_signal_6028), .Q (new_AGEMA_signal_6029) ) ;
    buf_clk new_AGEMA_reg_buffer_2570 ( .C (clk), .D (new_AGEMA_signal_6034), .Q (new_AGEMA_signal_6035) ) ;
    buf_clk new_AGEMA_reg_buffer_2576 ( .C (clk), .D (new_AGEMA_signal_6040), .Q (new_AGEMA_signal_6041) ) ;
    buf_clk new_AGEMA_reg_buffer_2582 ( .C (clk), .D (new_AGEMA_signal_6046), .Q (new_AGEMA_signal_6047) ) ;
    buf_clk new_AGEMA_reg_buffer_2588 ( .C (clk), .D (new_AGEMA_signal_6052), .Q (new_AGEMA_signal_6053) ) ;
    buf_clk new_AGEMA_reg_buffer_2594 ( .C (clk), .D (new_AGEMA_signal_6058), .Q (new_AGEMA_signal_6059) ) ;
    buf_clk new_AGEMA_reg_buffer_2600 ( .C (clk), .D (new_AGEMA_signal_6064), .Q (new_AGEMA_signal_6065) ) ;
    buf_clk new_AGEMA_reg_buffer_2606 ( .C (clk), .D (new_AGEMA_signal_6070), .Q (new_AGEMA_signal_6071) ) ;
    buf_clk new_AGEMA_reg_buffer_2612 ( .C (clk), .D (new_AGEMA_signal_6076), .Q (new_AGEMA_signal_6077) ) ;
    buf_clk new_AGEMA_reg_buffer_2618 ( .C (clk), .D (new_AGEMA_signal_6082), .Q (new_AGEMA_signal_6083) ) ;
    buf_clk new_AGEMA_reg_buffer_2624 ( .C (clk), .D (new_AGEMA_signal_6088), .Q (new_AGEMA_signal_6089) ) ;
    buf_clk new_AGEMA_reg_buffer_2630 ( .C (clk), .D (new_AGEMA_signal_6094), .Q (new_AGEMA_signal_6095) ) ;
    buf_clk new_AGEMA_reg_buffer_2636 ( .C (clk), .D (new_AGEMA_signal_6100), .Q (new_AGEMA_signal_6101) ) ;
    buf_clk new_AGEMA_reg_buffer_2642 ( .C (clk), .D (new_AGEMA_signal_6106), .Q (new_AGEMA_signal_6107) ) ;
    buf_clk new_AGEMA_reg_buffer_2648 ( .C (clk), .D (new_AGEMA_signal_6112), .Q (new_AGEMA_signal_6113) ) ;
    buf_clk new_AGEMA_reg_buffer_2654 ( .C (clk), .D (new_AGEMA_signal_6118), .Q (new_AGEMA_signal_6119) ) ;
    buf_clk new_AGEMA_reg_buffer_2660 ( .C (clk), .D (new_AGEMA_signal_6124), .Q (new_AGEMA_signal_6125) ) ;
    buf_clk new_AGEMA_reg_buffer_2666 ( .C (clk), .D (new_AGEMA_signal_6130), .Q (new_AGEMA_signal_6131) ) ;
    buf_clk new_AGEMA_reg_buffer_2672 ( .C (clk), .D (new_AGEMA_signal_6136), .Q (new_AGEMA_signal_6137) ) ;
    buf_clk new_AGEMA_reg_buffer_2678 ( .C (clk), .D (new_AGEMA_signal_6142), .Q (new_AGEMA_signal_6143) ) ;
    buf_clk new_AGEMA_reg_buffer_2684 ( .C (clk), .D (new_AGEMA_signal_6148), .Q (new_AGEMA_signal_6149) ) ;
    buf_clk new_AGEMA_reg_buffer_2690 ( .C (clk), .D (new_AGEMA_signal_6154), .Q (new_AGEMA_signal_6155) ) ;
    buf_clk new_AGEMA_reg_buffer_2696 ( .C (clk), .D (new_AGEMA_signal_6160), .Q (new_AGEMA_signal_6161) ) ;
    buf_clk new_AGEMA_reg_buffer_2702 ( .C (clk), .D (new_AGEMA_signal_6166), .Q (new_AGEMA_signal_6167) ) ;
    buf_clk new_AGEMA_reg_buffer_2708 ( .C (clk), .D (new_AGEMA_signal_6172), .Q (new_AGEMA_signal_6173) ) ;
    buf_clk new_AGEMA_reg_buffer_2714 ( .C (clk), .D (new_AGEMA_signal_6178), .Q (new_AGEMA_signal_6179) ) ;
    buf_clk new_AGEMA_reg_buffer_2720 ( .C (clk), .D (new_AGEMA_signal_6184), .Q (new_AGEMA_signal_6185) ) ;
    buf_clk new_AGEMA_reg_buffer_2726 ( .C (clk), .D (new_AGEMA_signal_6190), .Q (new_AGEMA_signal_6191) ) ;
    buf_clk new_AGEMA_reg_buffer_2732 ( .C (clk), .D (new_AGEMA_signal_6196), .Q (new_AGEMA_signal_6197) ) ;
    buf_clk new_AGEMA_reg_buffer_2738 ( .C (clk), .D (new_AGEMA_signal_6202), .Q (new_AGEMA_signal_6203) ) ;
    buf_clk new_AGEMA_reg_buffer_2744 ( .C (clk), .D (new_AGEMA_signal_6208), .Q (new_AGEMA_signal_6209) ) ;
    buf_clk new_AGEMA_reg_buffer_2750 ( .C (clk), .D (new_AGEMA_signal_6214), .Q (new_AGEMA_signal_6215) ) ;
    buf_clk new_AGEMA_reg_buffer_2756 ( .C (clk), .D (new_AGEMA_signal_6220), .Q (new_AGEMA_signal_6221) ) ;
    buf_clk new_AGEMA_reg_buffer_2762 ( .C (clk), .D (new_AGEMA_signal_6226), .Q (new_AGEMA_signal_6227) ) ;
    buf_clk new_AGEMA_reg_buffer_2768 ( .C (clk), .D (new_AGEMA_signal_6232), .Q (new_AGEMA_signal_6233) ) ;
    buf_clk new_AGEMA_reg_buffer_2774 ( .C (clk), .D (new_AGEMA_signal_6238), .Q (new_AGEMA_signal_6239) ) ;
    buf_clk new_AGEMA_reg_buffer_2780 ( .C (clk), .D (new_AGEMA_signal_6244), .Q (new_AGEMA_signal_6245) ) ;
    buf_clk new_AGEMA_reg_buffer_2786 ( .C (clk), .D (new_AGEMA_signal_6250), .Q (new_AGEMA_signal_6251) ) ;
    buf_clk new_AGEMA_reg_buffer_2792 ( .C (clk), .D (new_AGEMA_signal_6256), .Q (new_AGEMA_signal_6257) ) ;
    buf_clk new_AGEMA_reg_buffer_2798 ( .C (clk), .D (new_AGEMA_signal_6262), .Q (new_AGEMA_signal_6263) ) ;
    buf_clk new_AGEMA_reg_buffer_2804 ( .C (clk), .D (new_AGEMA_signal_6268), .Q (new_AGEMA_signal_6269) ) ;
    buf_clk new_AGEMA_reg_buffer_2810 ( .C (clk), .D (new_AGEMA_signal_6274), .Q (new_AGEMA_signal_6275) ) ;
    buf_clk new_AGEMA_reg_buffer_2816 ( .C (clk), .D (new_AGEMA_signal_6280), .Q (new_AGEMA_signal_6281) ) ;
    buf_clk new_AGEMA_reg_buffer_2822 ( .C (clk), .D (new_AGEMA_signal_6286), .Q (new_AGEMA_signal_6287) ) ;
    buf_clk new_AGEMA_reg_buffer_2828 ( .C (clk), .D (new_AGEMA_signal_6292), .Q (new_AGEMA_signal_6293) ) ;
    buf_clk new_AGEMA_reg_buffer_2834 ( .C (clk), .D (new_AGEMA_signal_6298), .Q (new_AGEMA_signal_6299) ) ;
    buf_clk new_AGEMA_reg_buffer_2840 ( .C (clk), .D (new_AGEMA_signal_6304), .Q (new_AGEMA_signal_6305) ) ;
    buf_clk new_AGEMA_reg_buffer_2846 ( .C (clk), .D (new_AGEMA_signal_6310), .Q (new_AGEMA_signal_6311) ) ;
    buf_clk new_AGEMA_reg_buffer_2852 ( .C (clk), .D (new_AGEMA_signal_6316), .Q (new_AGEMA_signal_6317) ) ;
    buf_clk new_AGEMA_reg_buffer_2858 ( .C (clk), .D (new_AGEMA_signal_6322), .Q (new_AGEMA_signal_6323) ) ;
    buf_clk new_AGEMA_reg_buffer_2864 ( .C (clk), .D (new_AGEMA_signal_6328), .Q (new_AGEMA_signal_6329) ) ;
    buf_clk new_AGEMA_reg_buffer_2870 ( .C (clk), .D (new_AGEMA_signal_6334), .Q (new_AGEMA_signal_6335) ) ;
    buf_clk new_AGEMA_reg_buffer_2876 ( .C (clk), .D (new_AGEMA_signal_6340), .Q (new_AGEMA_signal_6341) ) ;
    buf_clk new_AGEMA_reg_buffer_2882 ( .C (clk), .D (new_AGEMA_signal_6346), .Q (new_AGEMA_signal_6347) ) ;
    buf_clk new_AGEMA_reg_buffer_2888 ( .C (clk), .D (new_AGEMA_signal_6352), .Q (new_AGEMA_signal_6353) ) ;
    buf_clk new_AGEMA_reg_buffer_2894 ( .C (clk), .D (new_AGEMA_signal_6358), .Q (new_AGEMA_signal_6359) ) ;
    buf_clk new_AGEMA_reg_buffer_2900 ( .C (clk), .D (new_AGEMA_signal_6364), .Q (new_AGEMA_signal_6365) ) ;
    buf_clk new_AGEMA_reg_buffer_2906 ( .C (clk), .D (new_AGEMA_signal_6370), .Q (new_AGEMA_signal_6371) ) ;
    buf_clk new_AGEMA_reg_buffer_2912 ( .C (clk), .D (new_AGEMA_signal_6376), .Q (new_AGEMA_signal_6377) ) ;
    buf_clk new_AGEMA_reg_buffer_2918 ( .C (clk), .D (new_AGEMA_signal_6382), .Q (new_AGEMA_signal_6383) ) ;
    buf_clk new_AGEMA_reg_buffer_2924 ( .C (clk), .D (new_AGEMA_signal_6388), .Q (new_AGEMA_signal_6389) ) ;
    buf_clk new_AGEMA_reg_buffer_2930 ( .C (clk), .D (new_AGEMA_signal_6394), .Q (new_AGEMA_signal_6395) ) ;
    buf_clk new_AGEMA_reg_buffer_2936 ( .C (clk), .D (new_AGEMA_signal_6400), .Q (new_AGEMA_signal_6401) ) ;
    buf_clk new_AGEMA_reg_buffer_2942 ( .C (clk), .D (new_AGEMA_signal_6406), .Q (new_AGEMA_signal_6407) ) ;
    buf_clk new_AGEMA_reg_buffer_2948 ( .C (clk), .D (new_AGEMA_signal_6412), .Q (new_AGEMA_signal_6413) ) ;
    buf_clk new_AGEMA_reg_buffer_2954 ( .C (clk), .D (new_AGEMA_signal_6418), .Q (new_AGEMA_signal_6419) ) ;
    buf_clk new_AGEMA_reg_buffer_2960 ( .C (clk), .D (new_AGEMA_signal_6424), .Q (new_AGEMA_signal_6425) ) ;
    buf_clk new_AGEMA_reg_buffer_2966 ( .C (clk), .D (new_AGEMA_signal_6430), .Q (new_AGEMA_signal_6431) ) ;
    buf_clk new_AGEMA_reg_buffer_2972 ( .C (clk), .D (new_AGEMA_signal_6436), .Q (new_AGEMA_signal_6437) ) ;
    buf_clk new_AGEMA_reg_buffer_2978 ( .C (clk), .D (new_AGEMA_signal_6442), .Q (new_AGEMA_signal_6443) ) ;
    buf_clk new_AGEMA_reg_buffer_2984 ( .C (clk), .D (new_AGEMA_signal_6448), .Q (new_AGEMA_signal_6449) ) ;
    buf_clk new_AGEMA_reg_buffer_2990 ( .C (clk), .D (new_AGEMA_signal_6454), .Q (new_AGEMA_signal_6455) ) ;
    buf_clk new_AGEMA_reg_buffer_2996 ( .C (clk), .D (new_AGEMA_signal_6460), .Q (new_AGEMA_signal_6461) ) ;
    buf_clk new_AGEMA_reg_buffer_3002 ( .C (clk), .D (new_AGEMA_signal_6466), .Q (new_AGEMA_signal_6467) ) ;
    buf_clk new_AGEMA_reg_buffer_3008 ( .C (clk), .D (new_AGEMA_signal_6472), .Q (new_AGEMA_signal_6473) ) ;
    buf_clk new_AGEMA_reg_buffer_3014 ( .C (clk), .D (new_AGEMA_signal_6478), .Q (new_AGEMA_signal_6479) ) ;
    buf_clk new_AGEMA_reg_buffer_3020 ( .C (clk), .D (new_AGEMA_signal_6484), .Q (new_AGEMA_signal_6485) ) ;
    buf_clk new_AGEMA_reg_buffer_3026 ( .C (clk), .D (new_AGEMA_signal_6490), .Q (new_AGEMA_signal_6491) ) ;
    buf_clk new_AGEMA_reg_buffer_3032 ( .C (clk), .D (new_AGEMA_signal_6496), .Q (new_AGEMA_signal_6497) ) ;
    buf_clk new_AGEMA_reg_buffer_3038 ( .C (clk), .D (new_AGEMA_signal_6502), .Q (new_AGEMA_signal_6503) ) ;
    buf_clk new_AGEMA_reg_buffer_3044 ( .C (clk), .D (new_AGEMA_signal_6508), .Q (new_AGEMA_signal_6509) ) ;
    buf_clk new_AGEMA_reg_buffer_3050 ( .C (clk), .D (new_AGEMA_signal_6514), .Q (new_AGEMA_signal_6515) ) ;
    buf_clk new_AGEMA_reg_buffer_3056 ( .C (clk), .D (new_AGEMA_signal_6520), .Q (new_AGEMA_signal_6521) ) ;
    buf_clk new_AGEMA_reg_buffer_3062 ( .C (clk), .D (new_AGEMA_signal_6526), .Q (new_AGEMA_signal_6527) ) ;
    buf_clk new_AGEMA_reg_buffer_3068 ( .C (clk), .D (new_AGEMA_signal_6532), .Q (new_AGEMA_signal_6533) ) ;
    buf_clk new_AGEMA_reg_buffer_3074 ( .C (clk), .D (new_AGEMA_signal_6538), .Q (new_AGEMA_signal_6539) ) ;
    buf_clk new_AGEMA_reg_buffer_3080 ( .C (clk), .D (new_AGEMA_signal_6544), .Q (new_AGEMA_signal_6545) ) ;
    buf_clk new_AGEMA_reg_buffer_3086 ( .C (clk), .D (new_AGEMA_signal_6550), .Q (new_AGEMA_signal_6551) ) ;
    buf_clk new_AGEMA_reg_buffer_3092 ( .C (clk), .D (new_AGEMA_signal_6556), .Q (new_AGEMA_signal_6557) ) ;
    buf_clk new_AGEMA_reg_buffer_3098 ( .C (clk), .D (new_AGEMA_signal_6562), .Q (new_AGEMA_signal_6563) ) ;
    buf_clk new_AGEMA_reg_buffer_3104 ( .C (clk), .D (new_AGEMA_signal_6568), .Q (new_AGEMA_signal_6569) ) ;
    buf_clk new_AGEMA_reg_buffer_3110 ( .C (clk), .D (new_AGEMA_signal_6574), .Q (new_AGEMA_signal_6575) ) ;
    buf_clk new_AGEMA_reg_buffer_3116 ( .C (clk), .D (new_AGEMA_signal_6580), .Q (new_AGEMA_signal_6581) ) ;
    buf_clk new_AGEMA_reg_buffer_3122 ( .C (clk), .D (new_AGEMA_signal_6586), .Q (new_AGEMA_signal_6587) ) ;
    buf_clk new_AGEMA_reg_buffer_3128 ( .C (clk), .D (new_AGEMA_signal_6592), .Q (new_AGEMA_signal_6593) ) ;
    buf_clk new_AGEMA_reg_buffer_3134 ( .C (clk), .D (new_AGEMA_signal_6598), .Q (new_AGEMA_signal_6599) ) ;
    buf_clk new_AGEMA_reg_buffer_3140 ( .C (clk), .D (new_AGEMA_signal_6604), .Q (new_AGEMA_signal_6605) ) ;
    buf_clk new_AGEMA_reg_buffer_3146 ( .C (clk), .D (new_AGEMA_signal_6610), .Q (new_AGEMA_signal_6611) ) ;
    buf_clk new_AGEMA_reg_buffer_3152 ( .C (clk), .D (new_AGEMA_signal_6616), .Q (new_AGEMA_signal_6617) ) ;
    buf_clk new_AGEMA_reg_buffer_3158 ( .C (clk), .D (new_AGEMA_signal_6622), .Q (new_AGEMA_signal_6623) ) ;
    buf_clk new_AGEMA_reg_buffer_3164 ( .C (clk), .D (new_AGEMA_signal_6628), .Q (new_AGEMA_signal_6629) ) ;
    buf_clk new_AGEMA_reg_buffer_3170 ( .C (clk), .D (new_AGEMA_signal_6634), .Q (new_AGEMA_signal_6635) ) ;
    buf_clk new_AGEMA_reg_buffer_3176 ( .C (clk), .D (new_AGEMA_signal_6640), .Q (new_AGEMA_signal_6641) ) ;
    buf_clk new_AGEMA_reg_buffer_3182 ( .C (clk), .D (new_AGEMA_signal_6646), .Q (new_AGEMA_signal_6647) ) ;
    buf_clk new_AGEMA_reg_buffer_3188 ( .C (clk), .D (new_AGEMA_signal_6652), .Q (new_AGEMA_signal_6653) ) ;
    buf_clk new_AGEMA_reg_buffer_3194 ( .C (clk), .D (new_AGEMA_signal_6658), .Q (new_AGEMA_signal_6659) ) ;
    buf_clk new_AGEMA_reg_buffer_3200 ( .C (clk), .D (new_AGEMA_signal_6664), .Q (new_AGEMA_signal_6665) ) ;
    buf_clk new_AGEMA_reg_buffer_3206 ( .C (clk), .D (new_AGEMA_signal_6670), .Q (new_AGEMA_signal_6671) ) ;
    buf_clk new_AGEMA_reg_buffer_3212 ( .C (clk), .D (new_AGEMA_signal_6676), .Q (new_AGEMA_signal_6677) ) ;
    buf_clk new_AGEMA_reg_buffer_3218 ( .C (clk), .D (new_AGEMA_signal_6682), .Q (new_AGEMA_signal_6683) ) ;
    buf_clk new_AGEMA_reg_buffer_3224 ( .C (clk), .D (new_AGEMA_signal_6688), .Q (new_AGEMA_signal_6689) ) ;
    buf_clk new_AGEMA_reg_buffer_3230 ( .C (clk), .D (new_AGEMA_signal_6694), .Q (new_AGEMA_signal_6695) ) ;
    buf_clk new_AGEMA_reg_buffer_3236 ( .C (clk), .D (new_AGEMA_signal_6700), .Q (new_AGEMA_signal_6701) ) ;
    buf_clk new_AGEMA_reg_buffer_3242 ( .C (clk), .D (new_AGEMA_signal_6706), .Q (new_AGEMA_signal_6707) ) ;
    buf_clk new_AGEMA_reg_buffer_3248 ( .C (clk), .D (new_AGEMA_signal_6712), .Q (new_AGEMA_signal_6713) ) ;
    buf_clk new_AGEMA_reg_buffer_3254 ( .C (clk), .D (new_AGEMA_signal_6718), .Q (new_AGEMA_signal_6719) ) ;
    buf_clk new_AGEMA_reg_buffer_3260 ( .C (clk), .D (new_AGEMA_signal_6724), .Q (new_AGEMA_signal_6725) ) ;
    buf_clk new_AGEMA_reg_buffer_3266 ( .C (clk), .D (new_AGEMA_signal_6730), .Q (new_AGEMA_signal_6731) ) ;
    buf_clk new_AGEMA_reg_buffer_3272 ( .C (clk), .D (new_AGEMA_signal_6736), .Q (new_AGEMA_signal_6737) ) ;
    buf_clk new_AGEMA_reg_buffer_3278 ( .C (clk), .D (new_AGEMA_signal_6742), .Q (new_AGEMA_signal_6743) ) ;
    buf_clk new_AGEMA_reg_buffer_3284 ( .C (clk), .D (new_AGEMA_signal_6748), .Q (new_AGEMA_signal_6749) ) ;
    buf_clk new_AGEMA_reg_buffer_3290 ( .C (clk), .D (new_AGEMA_signal_6754), .Q (new_AGEMA_signal_6755) ) ;
    buf_clk new_AGEMA_reg_buffer_3296 ( .C (clk), .D (new_AGEMA_signal_6760), .Q (new_AGEMA_signal_6761) ) ;
    buf_clk new_AGEMA_reg_buffer_3302 ( .C (clk), .D (new_AGEMA_signal_6766), .Q (new_AGEMA_signal_6767) ) ;
    buf_clk new_AGEMA_reg_buffer_3308 ( .C (clk), .D (new_AGEMA_signal_6772), .Q (new_AGEMA_signal_6773) ) ;
    buf_clk new_AGEMA_reg_buffer_3314 ( .C (clk), .D (new_AGEMA_signal_6778), .Q (new_AGEMA_signal_6779) ) ;
    buf_clk new_AGEMA_reg_buffer_3320 ( .C (clk), .D (new_AGEMA_signal_6784), .Q (new_AGEMA_signal_6785) ) ;
    buf_clk new_AGEMA_reg_buffer_3326 ( .C (clk), .D (new_AGEMA_signal_6790), .Q (new_AGEMA_signal_6791) ) ;
    buf_clk new_AGEMA_reg_buffer_3332 ( .C (clk), .D (new_AGEMA_signal_6796), .Q (new_AGEMA_signal_6797) ) ;
    buf_clk new_AGEMA_reg_buffer_3338 ( .C (clk), .D (new_AGEMA_signal_6802), .Q (new_AGEMA_signal_6803) ) ;
    buf_clk new_AGEMA_reg_buffer_3344 ( .C (clk), .D (new_AGEMA_signal_6808), .Q (new_AGEMA_signal_6809) ) ;
    buf_clk new_AGEMA_reg_buffer_3350 ( .C (clk), .D (new_AGEMA_signal_6814), .Q (new_AGEMA_signal_6815) ) ;
    buf_clk new_AGEMA_reg_buffer_3356 ( .C (clk), .D (new_AGEMA_signal_6820), .Q (new_AGEMA_signal_6821) ) ;
    buf_clk new_AGEMA_reg_buffer_3362 ( .C (clk), .D (new_AGEMA_signal_6826), .Q (new_AGEMA_signal_6827) ) ;
    buf_clk new_AGEMA_reg_buffer_3368 ( .C (clk), .D (new_AGEMA_signal_6832), .Q (new_AGEMA_signal_6833) ) ;
    buf_clk new_AGEMA_reg_buffer_3374 ( .C (clk), .D (new_AGEMA_signal_6838), .Q (new_AGEMA_signal_6839) ) ;
    buf_clk new_AGEMA_reg_buffer_3380 ( .C (clk), .D (new_AGEMA_signal_6844), .Q (new_AGEMA_signal_6845) ) ;
    buf_clk new_AGEMA_reg_buffer_3386 ( .C (clk), .D (new_AGEMA_signal_6850), .Q (new_AGEMA_signal_6851) ) ;
    buf_clk new_AGEMA_reg_buffer_3392 ( .C (clk), .D (new_AGEMA_signal_6856), .Q (new_AGEMA_signal_6857) ) ;
    buf_clk new_AGEMA_reg_buffer_3398 ( .C (clk), .D (new_AGEMA_signal_6862), .Q (new_AGEMA_signal_6863) ) ;
    buf_clk new_AGEMA_reg_buffer_3404 ( .C (clk), .D (new_AGEMA_signal_6868), .Q (new_AGEMA_signal_6869) ) ;
    buf_clk new_AGEMA_reg_buffer_3410 ( .C (clk), .D (new_AGEMA_signal_6874), .Q (new_AGEMA_signal_6875) ) ;
    buf_clk new_AGEMA_reg_buffer_3416 ( .C (clk), .D (new_AGEMA_signal_6880), .Q (new_AGEMA_signal_6881) ) ;
    buf_clk new_AGEMA_reg_buffer_3422 ( .C (clk), .D (new_AGEMA_signal_6886), .Q (new_AGEMA_signal_6887) ) ;
    buf_clk new_AGEMA_reg_buffer_3428 ( .C (clk), .D (new_AGEMA_signal_6892), .Q (new_AGEMA_signal_6893) ) ;
    buf_clk new_AGEMA_reg_buffer_3434 ( .C (clk), .D (new_AGEMA_signal_6898), .Q (new_AGEMA_signal_6899) ) ;
    buf_clk new_AGEMA_reg_buffer_3440 ( .C (clk), .D (new_AGEMA_signal_6904), .Q (new_AGEMA_signal_6905) ) ;
    buf_clk new_AGEMA_reg_buffer_3446 ( .C (clk), .D (new_AGEMA_signal_6910), .Q (new_AGEMA_signal_6911) ) ;
    buf_clk new_AGEMA_reg_buffer_3452 ( .C (clk), .D (new_AGEMA_signal_6916), .Q (new_AGEMA_signal_6917) ) ;
    buf_clk new_AGEMA_reg_buffer_3458 ( .C (clk), .D (new_AGEMA_signal_6922), .Q (new_AGEMA_signal_6923) ) ;
    buf_clk new_AGEMA_reg_buffer_3464 ( .C (clk), .D (new_AGEMA_signal_6928), .Q (new_AGEMA_signal_6929) ) ;
    buf_clk new_AGEMA_reg_buffer_3470 ( .C (clk), .D (new_AGEMA_signal_6934), .Q (new_AGEMA_signal_6935) ) ;
    buf_clk new_AGEMA_reg_buffer_3476 ( .C (clk), .D (new_AGEMA_signal_6940), .Q (new_AGEMA_signal_6941) ) ;
    buf_clk new_AGEMA_reg_buffer_3482 ( .C (clk), .D (new_AGEMA_signal_6946), .Q (new_AGEMA_signal_6947) ) ;
    buf_clk new_AGEMA_reg_buffer_3488 ( .C (clk), .D (new_AGEMA_signal_6952), .Q (new_AGEMA_signal_6953) ) ;
    buf_clk new_AGEMA_reg_buffer_3494 ( .C (clk), .D (new_AGEMA_signal_6958), .Q (new_AGEMA_signal_6959) ) ;
    buf_clk new_AGEMA_reg_buffer_3500 ( .C (clk), .D (new_AGEMA_signal_6964), .Q (new_AGEMA_signal_6965) ) ;
    buf_clk new_AGEMA_reg_buffer_3506 ( .C (clk), .D (new_AGEMA_signal_6970), .Q (new_AGEMA_signal_6971) ) ;
    buf_clk new_AGEMA_reg_buffer_3512 ( .C (clk), .D (new_AGEMA_signal_6976), .Q (new_AGEMA_signal_6977) ) ;
    buf_clk new_AGEMA_reg_buffer_3518 ( .C (clk), .D (new_AGEMA_signal_6982), .Q (new_AGEMA_signal_6983) ) ;
    buf_clk new_AGEMA_reg_buffer_3524 ( .C (clk), .D (new_AGEMA_signal_6988), .Q (new_AGEMA_signal_6989) ) ;
    buf_clk new_AGEMA_reg_buffer_3530 ( .C (clk), .D (new_AGEMA_signal_6994), .Q (new_AGEMA_signal_6995) ) ;
    buf_clk new_AGEMA_reg_buffer_3536 ( .C (clk), .D (new_AGEMA_signal_7000), .Q (new_AGEMA_signal_7001) ) ;
    buf_clk new_AGEMA_reg_buffer_3542 ( .C (clk), .D (new_AGEMA_signal_7006), .Q (new_AGEMA_signal_7007) ) ;
    buf_clk new_AGEMA_reg_buffer_3548 ( .C (clk), .D (new_AGEMA_signal_7012), .Q (new_AGEMA_signal_7013) ) ;
    buf_clk new_AGEMA_reg_buffer_3554 ( .C (clk), .D (new_AGEMA_signal_7018), .Q (new_AGEMA_signal_7019) ) ;
    buf_clk new_AGEMA_reg_buffer_3560 ( .C (clk), .D (new_AGEMA_signal_7024), .Q (new_AGEMA_signal_7025) ) ;
    buf_clk new_AGEMA_reg_buffer_3566 ( .C (clk), .D (new_AGEMA_signal_7030), .Q (new_AGEMA_signal_7031) ) ;
    buf_clk new_AGEMA_reg_buffer_3572 ( .C (clk), .D (new_AGEMA_signal_7036), .Q (new_AGEMA_signal_7037) ) ;
    buf_clk new_AGEMA_reg_buffer_3866 ( .C (clk), .D (new_AGEMA_signal_7330), .Q (new_AGEMA_signal_7331) ) ;
    buf_clk new_AGEMA_reg_buffer_3872 ( .C (clk), .D (new_AGEMA_signal_7336), .Q (new_AGEMA_signal_7337) ) ;
    buf_clk new_AGEMA_reg_buffer_3880 ( .C (clk), .D (new_AGEMA_signal_7344), .Q (new_AGEMA_signal_7345) ) ;
    buf_clk new_AGEMA_reg_buffer_3888 ( .C (clk), .D (new_AGEMA_signal_7352), .Q (new_AGEMA_signal_7353) ) ;
    buf_clk new_AGEMA_reg_buffer_3896 ( .C (clk), .D (new_AGEMA_signal_7360), .Q (new_AGEMA_signal_7361) ) ;
    buf_clk new_AGEMA_reg_buffer_3904 ( .C (clk), .D (new_AGEMA_signal_7368), .Q (new_AGEMA_signal_7369) ) ;
    buf_clk new_AGEMA_reg_buffer_3912 ( .C (clk), .D (new_AGEMA_signal_7376), .Q (new_AGEMA_signal_7377) ) ;
    buf_clk new_AGEMA_reg_buffer_3920 ( .C (clk), .D (new_AGEMA_signal_7384), .Q (new_AGEMA_signal_7385) ) ;
    buf_clk new_AGEMA_reg_buffer_3928 ( .C (clk), .D (new_AGEMA_signal_7392), .Q (new_AGEMA_signal_7393) ) ;
    buf_clk new_AGEMA_reg_buffer_3936 ( .C (clk), .D (new_AGEMA_signal_7400), .Q (new_AGEMA_signal_7401) ) ;
    buf_clk new_AGEMA_reg_buffer_3944 ( .C (clk), .D (new_AGEMA_signal_7408), .Q (new_AGEMA_signal_7409) ) ;
    buf_clk new_AGEMA_reg_buffer_3952 ( .C (clk), .D (new_AGEMA_signal_7416), .Q (new_AGEMA_signal_7417) ) ;
    buf_clk new_AGEMA_reg_buffer_3960 ( .C (clk), .D (new_AGEMA_signal_7424), .Q (new_AGEMA_signal_7425) ) ;
    buf_clk new_AGEMA_reg_buffer_3968 ( .C (clk), .D (new_AGEMA_signal_7432), .Q (new_AGEMA_signal_7433) ) ;
    buf_clk new_AGEMA_reg_buffer_3976 ( .C (clk), .D (new_AGEMA_signal_7440), .Q (new_AGEMA_signal_7441) ) ;
    buf_clk new_AGEMA_reg_buffer_3984 ( .C (clk), .D (new_AGEMA_signal_7448), .Q (new_AGEMA_signal_7449) ) ;
    buf_clk new_AGEMA_reg_buffer_3992 ( .C (clk), .D (new_AGEMA_signal_7456), .Q (new_AGEMA_signal_7457) ) ;
    buf_clk new_AGEMA_reg_buffer_4000 ( .C (clk), .D (new_AGEMA_signal_7464), .Q (new_AGEMA_signal_7465) ) ;
    buf_clk new_AGEMA_reg_buffer_4008 ( .C (clk), .D (new_AGEMA_signal_7472), .Q (new_AGEMA_signal_7473) ) ;
    buf_clk new_AGEMA_reg_buffer_4016 ( .C (clk), .D (new_AGEMA_signal_7480), .Q (new_AGEMA_signal_7481) ) ;
    buf_clk new_AGEMA_reg_buffer_4024 ( .C (clk), .D (new_AGEMA_signal_7488), .Q (new_AGEMA_signal_7489) ) ;
    buf_clk new_AGEMA_reg_buffer_4032 ( .C (clk), .D (new_AGEMA_signal_7496), .Q (new_AGEMA_signal_7497) ) ;
    buf_clk new_AGEMA_reg_buffer_4040 ( .C (clk), .D (new_AGEMA_signal_7504), .Q (new_AGEMA_signal_7505) ) ;
    buf_clk new_AGEMA_reg_buffer_4048 ( .C (clk), .D (new_AGEMA_signal_7512), .Q (new_AGEMA_signal_7513) ) ;
    buf_clk new_AGEMA_reg_buffer_4056 ( .C (clk), .D (new_AGEMA_signal_7520), .Q (new_AGEMA_signal_7521) ) ;
    buf_clk new_AGEMA_reg_buffer_4064 ( .C (clk), .D (new_AGEMA_signal_7528), .Q (new_AGEMA_signal_7529) ) ;
    buf_clk new_AGEMA_reg_buffer_4072 ( .C (clk), .D (new_AGEMA_signal_7536), .Q (new_AGEMA_signal_7537) ) ;
    buf_clk new_AGEMA_reg_buffer_4080 ( .C (clk), .D (new_AGEMA_signal_7544), .Q (new_AGEMA_signal_7545) ) ;
    buf_clk new_AGEMA_reg_buffer_4088 ( .C (clk), .D (new_AGEMA_signal_7552), .Q (new_AGEMA_signal_7553) ) ;
    buf_clk new_AGEMA_reg_buffer_4096 ( .C (clk), .D (new_AGEMA_signal_7560), .Q (new_AGEMA_signal_7561) ) ;
    buf_clk new_AGEMA_reg_buffer_4104 ( .C (clk), .D (new_AGEMA_signal_7568), .Q (new_AGEMA_signal_7569) ) ;
    buf_clk new_AGEMA_reg_buffer_4112 ( .C (clk), .D (new_AGEMA_signal_7576), .Q (new_AGEMA_signal_7577) ) ;
    buf_clk new_AGEMA_reg_buffer_4120 ( .C (clk), .D (new_AGEMA_signal_7584), .Q (new_AGEMA_signal_7585) ) ;
    buf_clk new_AGEMA_reg_buffer_4128 ( .C (clk), .D (new_AGEMA_signal_7592), .Q (new_AGEMA_signal_7593) ) ;
    buf_clk new_AGEMA_reg_buffer_4136 ( .C (clk), .D (new_AGEMA_signal_7600), .Q (new_AGEMA_signal_7601) ) ;
    buf_clk new_AGEMA_reg_buffer_4144 ( .C (clk), .D (new_AGEMA_signal_7608), .Q (new_AGEMA_signal_7609) ) ;
    buf_clk new_AGEMA_reg_buffer_4152 ( .C (clk), .D (new_AGEMA_signal_7616), .Q (new_AGEMA_signal_7617) ) ;
    buf_clk new_AGEMA_reg_buffer_4160 ( .C (clk), .D (new_AGEMA_signal_7624), .Q (new_AGEMA_signal_7625) ) ;
    buf_clk new_AGEMA_reg_buffer_4168 ( .C (clk), .D (new_AGEMA_signal_7632), .Q (new_AGEMA_signal_7633) ) ;
    buf_clk new_AGEMA_reg_buffer_4176 ( .C (clk), .D (new_AGEMA_signal_7640), .Q (new_AGEMA_signal_7641) ) ;
    buf_clk new_AGEMA_reg_buffer_4184 ( .C (clk), .D (new_AGEMA_signal_7648), .Q (new_AGEMA_signal_7649) ) ;
    buf_clk new_AGEMA_reg_buffer_4192 ( .C (clk), .D (new_AGEMA_signal_7656), .Q (new_AGEMA_signal_7657) ) ;
    buf_clk new_AGEMA_reg_buffer_4200 ( .C (clk), .D (new_AGEMA_signal_7664), .Q (new_AGEMA_signal_7665) ) ;
    buf_clk new_AGEMA_reg_buffer_4208 ( .C (clk), .D (new_AGEMA_signal_7672), .Q (new_AGEMA_signal_7673) ) ;
    buf_clk new_AGEMA_reg_buffer_4216 ( .C (clk), .D (new_AGEMA_signal_7680), .Q (new_AGEMA_signal_7681) ) ;
    buf_clk new_AGEMA_reg_buffer_4224 ( .C (clk), .D (new_AGEMA_signal_7688), .Q (new_AGEMA_signal_7689) ) ;
    buf_clk new_AGEMA_reg_buffer_4232 ( .C (clk), .D (new_AGEMA_signal_7696), .Q (new_AGEMA_signal_7697) ) ;
    buf_clk new_AGEMA_reg_buffer_4240 ( .C (clk), .D (new_AGEMA_signal_7704), .Q (new_AGEMA_signal_7705) ) ;
    buf_clk new_AGEMA_reg_buffer_4248 ( .C (clk), .D (new_AGEMA_signal_7712), .Q (new_AGEMA_signal_7713) ) ;
    buf_clk new_AGEMA_reg_buffer_4256 ( .C (clk), .D (new_AGEMA_signal_7720), .Q (new_AGEMA_signal_7721) ) ;
    buf_clk new_AGEMA_reg_buffer_4264 ( .C (clk), .D (new_AGEMA_signal_7728), .Q (new_AGEMA_signal_7729) ) ;
    buf_clk new_AGEMA_reg_buffer_4272 ( .C (clk), .D (new_AGEMA_signal_7736), .Q (new_AGEMA_signal_7737) ) ;
    buf_clk new_AGEMA_reg_buffer_4280 ( .C (clk), .D (new_AGEMA_signal_7744), .Q (new_AGEMA_signal_7745) ) ;
    buf_clk new_AGEMA_reg_buffer_4288 ( .C (clk), .D (new_AGEMA_signal_7752), .Q (new_AGEMA_signal_7753) ) ;
    buf_clk new_AGEMA_reg_buffer_4296 ( .C (clk), .D (new_AGEMA_signal_7760), .Q (new_AGEMA_signal_7761) ) ;
    buf_clk new_AGEMA_reg_buffer_4304 ( .C (clk), .D (new_AGEMA_signal_7768), .Q (new_AGEMA_signal_7769) ) ;
    buf_clk new_AGEMA_reg_buffer_4312 ( .C (clk), .D (new_AGEMA_signal_7776), .Q (new_AGEMA_signal_7777) ) ;
    buf_clk new_AGEMA_reg_buffer_4320 ( .C (clk), .D (new_AGEMA_signal_7784), .Q (new_AGEMA_signal_7785) ) ;
    buf_clk new_AGEMA_reg_buffer_4328 ( .C (clk), .D (new_AGEMA_signal_7792), .Q (new_AGEMA_signal_7793) ) ;
    buf_clk new_AGEMA_reg_buffer_4336 ( .C (clk), .D (new_AGEMA_signal_7800), .Q (new_AGEMA_signal_7801) ) ;
    buf_clk new_AGEMA_reg_buffer_4344 ( .C (clk), .D (new_AGEMA_signal_7808), .Q (new_AGEMA_signal_7809) ) ;
    buf_clk new_AGEMA_reg_buffer_4352 ( .C (clk), .D (new_AGEMA_signal_7816), .Q (new_AGEMA_signal_7817) ) ;
    buf_clk new_AGEMA_reg_buffer_4360 ( .C (clk), .D (new_AGEMA_signal_7824), .Q (new_AGEMA_signal_7825) ) ;
    buf_clk new_AGEMA_reg_buffer_4368 ( .C (clk), .D (new_AGEMA_signal_7832), .Q (new_AGEMA_signal_7833) ) ;
    buf_clk new_AGEMA_reg_buffer_4376 ( .C (clk), .D (new_AGEMA_signal_7840), .Q (new_AGEMA_signal_7841) ) ;
    buf_clk new_AGEMA_reg_buffer_4384 ( .C (clk), .D (new_AGEMA_signal_7848), .Q (new_AGEMA_signal_7849) ) ;
    buf_clk new_AGEMA_reg_buffer_4392 ( .C (clk), .D (new_AGEMA_signal_7856), .Q (new_AGEMA_signal_7857) ) ;
    buf_clk new_AGEMA_reg_buffer_4400 ( .C (clk), .D (new_AGEMA_signal_7864), .Q (new_AGEMA_signal_7865) ) ;
    buf_clk new_AGEMA_reg_buffer_4408 ( .C (clk), .D (new_AGEMA_signal_7872), .Q (new_AGEMA_signal_7873) ) ;
    buf_clk new_AGEMA_reg_buffer_4416 ( .C (clk), .D (new_AGEMA_signal_7880), .Q (new_AGEMA_signal_7881) ) ;
    buf_clk new_AGEMA_reg_buffer_4424 ( .C (clk), .D (new_AGEMA_signal_7888), .Q (new_AGEMA_signal_7889) ) ;
    buf_clk new_AGEMA_reg_buffer_4432 ( .C (clk), .D (new_AGEMA_signal_7896), .Q (new_AGEMA_signal_7897) ) ;
    buf_clk new_AGEMA_reg_buffer_4440 ( .C (clk), .D (new_AGEMA_signal_7904), .Q (new_AGEMA_signal_7905) ) ;
    buf_clk new_AGEMA_reg_buffer_4448 ( .C (clk), .D (new_AGEMA_signal_7912), .Q (new_AGEMA_signal_7913) ) ;
    buf_clk new_AGEMA_reg_buffer_4456 ( .C (clk), .D (new_AGEMA_signal_7920), .Q (new_AGEMA_signal_7921) ) ;
    buf_clk new_AGEMA_reg_buffer_4464 ( .C (clk), .D (new_AGEMA_signal_7928), .Q (new_AGEMA_signal_7929) ) ;
    buf_clk new_AGEMA_reg_buffer_4472 ( .C (clk), .D (new_AGEMA_signal_7936), .Q (new_AGEMA_signal_7937) ) ;
    buf_clk new_AGEMA_reg_buffer_4480 ( .C (clk), .D (new_AGEMA_signal_7944), .Q (new_AGEMA_signal_7945) ) ;
    buf_clk new_AGEMA_reg_buffer_4488 ( .C (clk), .D (new_AGEMA_signal_7952), .Q (new_AGEMA_signal_7953) ) ;
    buf_clk new_AGEMA_reg_buffer_4496 ( .C (clk), .D (new_AGEMA_signal_7960), .Q (new_AGEMA_signal_7961) ) ;
    buf_clk new_AGEMA_reg_buffer_4504 ( .C (clk), .D (new_AGEMA_signal_7968), .Q (new_AGEMA_signal_7969) ) ;
    buf_clk new_AGEMA_reg_buffer_4512 ( .C (clk), .D (new_AGEMA_signal_7976), .Q (new_AGEMA_signal_7977) ) ;
    buf_clk new_AGEMA_reg_buffer_4520 ( .C (clk), .D (new_AGEMA_signal_7984), .Q (new_AGEMA_signal_7985) ) ;
    buf_clk new_AGEMA_reg_buffer_4528 ( .C (clk), .D (new_AGEMA_signal_7992), .Q (new_AGEMA_signal_7993) ) ;
    buf_clk new_AGEMA_reg_buffer_4536 ( .C (clk), .D (new_AGEMA_signal_8000), .Q (new_AGEMA_signal_8001) ) ;
    buf_clk new_AGEMA_reg_buffer_4544 ( .C (clk), .D (new_AGEMA_signal_8008), .Q (new_AGEMA_signal_8009) ) ;
    buf_clk new_AGEMA_reg_buffer_4552 ( .C (clk), .D (new_AGEMA_signal_8016), .Q (new_AGEMA_signal_8017) ) ;
    buf_clk new_AGEMA_reg_buffer_4560 ( .C (clk), .D (new_AGEMA_signal_8024), .Q (new_AGEMA_signal_8025) ) ;
    buf_clk new_AGEMA_reg_buffer_4568 ( .C (clk), .D (new_AGEMA_signal_8032), .Q (new_AGEMA_signal_8033) ) ;
    buf_clk new_AGEMA_reg_buffer_4576 ( .C (clk), .D (new_AGEMA_signal_8040), .Q (new_AGEMA_signal_8041) ) ;
    buf_clk new_AGEMA_reg_buffer_4584 ( .C (clk), .D (new_AGEMA_signal_8048), .Q (new_AGEMA_signal_8049) ) ;
    buf_clk new_AGEMA_reg_buffer_4592 ( .C (clk), .D (new_AGEMA_signal_8056), .Q (new_AGEMA_signal_8057) ) ;
    buf_clk new_AGEMA_reg_buffer_4600 ( .C (clk), .D (new_AGEMA_signal_8064), .Q (new_AGEMA_signal_8065) ) ;
    buf_clk new_AGEMA_reg_buffer_4608 ( .C (clk), .D (new_AGEMA_signal_8072), .Q (new_AGEMA_signal_8073) ) ;
    buf_clk new_AGEMA_reg_buffer_4616 ( .C (clk), .D (new_AGEMA_signal_8080), .Q (new_AGEMA_signal_8081) ) ;
    buf_clk new_AGEMA_reg_buffer_4624 ( .C (clk), .D (new_AGEMA_signal_8088), .Q (new_AGEMA_signal_8089) ) ;
    buf_clk new_AGEMA_reg_buffer_4632 ( .C (clk), .D (new_AGEMA_signal_8096), .Q (new_AGEMA_signal_8097) ) ;
    buf_clk new_AGEMA_reg_buffer_4640 ( .C (clk), .D (new_AGEMA_signal_8104), .Q (new_AGEMA_signal_8105) ) ;
    buf_clk new_AGEMA_reg_buffer_4648 ( .C (clk), .D (new_AGEMA_signal_8112), .Q (new_AGEMA_signal_8113) ) ;
    buf_clk new_AGEMA_reg_buffer_4656 ( .C (clk), .D (new_AGEMA_signal_8120), .Q (new_AGEMA_signal_8121) ) ;
    buf_clk new_AGEMA_reg_buffer_4664 ( .C (clk), .D (new_AGEMA_signal_8128), .Q (new_AGEMA_signal_8129) ) ;
    buf_clk new_AGEMA_reg_buffer_4672 ( .C (clk), .D (new_AGEMA_signal_8136), .Q (new_AGEMA_signal_8137) ) ;
    buf_clk new_AGEMA_reg_buffer_4680 ( .C (clk), .D (new_AGEMA_signal_8144), .Q (new_AGEMA_signal_8145) ) ;
    buf_clk new_AGEMA_reg_buffer_4688 ( .C (clk), .D (new_AGEMA_signal_8152), .Q (new_AGEMA_signal_8153) ) ;
    buf_clk new_AGEMA_reg_buffer_4696 ( .C (clk), .D (new_AGEMA_signal_8160), .Q (new_AGEMA_signal_8161) ) ;
    buf_clk new_AGEMA_reg_buffer_4704 ( .C (clk), .D (new_AGEMA_signal_8168), .Q (new_AGEMA_signal_8169) ) ;
    buf_clk new_AGEMA_reg_buffer_4712 ( .C (clk), .D (new_AGEMA_signal_8176), .Q (new_AGEMA_signal_8177) ) ;
    buf_clk new_AGEMA_reg_buffer_4720 ( .C (clk), .D (new_AGEMA_signal_8184), .Q (new_AGEMA_signal_8185) ) ;
    buf_clk new_AGEMA_reg_buffer_4728 ( .C (clk), .D (new_AGEMA_signal_8192), .Q (new_AGEMA_signal_8193) ) ;
    buf_clk new_AGEMA_reg_buffer_4736 ( .C (clk), .D (new_AGEMA_signal_8200), .Q (new_AGEMA_signal_8201) ) ;
    buf_clk new_AGEMA_reg_buffer_4744 ( .C (clk), .D (new_AGEMA_signal_8208), .Q (new_AGEMA_signal_8209) ) ;
    buf_clk new_AGEMA_reg_buffer_4752 ( .C (clk), .D (new_AGEMA_signal_8216), .Q (new_AGEMA_signal_8217) ) ;
    buf_clk new_AGEMA_reg_buffer_4760 ( .C (clk), .D (new_AGEMA_signal_8224), .Q (new_AGEMA_signal_8225) ) ;
    buf_clk new_AGEMA_reg_buffer_4768 ( .C (clk), .D (new_AGEMA_signal_8232), .Q (new_AGEMA_signal_8233) ) ;
    buf_clk new_AGEMA_reg_buffer_4776 ( .C (clk), .D (new_AGEMA_signal_8240), .Q (new_AGEMA_signal_8241) ) ;
    buf_clk new_AGEMA_reg_buffer_4784 ( .C (clk), .D (new_AGEMA_signal_8248), .Q (new_AGEMA_signal_8249) ) ;
    buf_clk new_AGEMA_reg_buffer_4792 ( .C (clk), .D (new_AGEMA_signal_8256), .Q (new_AGEMA_signal_8257) ) ;
    buf_clk new_AGEMA_reg_buffer_4800 ( .C (clk), .D (new_AGEMA_signal_8264), .Q (new_AGEMA_signal_8265) ) ;
    buf_clk new_AGEMA_reg_buffer_4808 ( .C (clk), .D (new_AGEMA_signal_8272), .Q (new_AGEMA_signal_8273) ) ;
    buf_clk new_AGEMA_reg_buffer_4816 ( .C (clk), .D (new_AGEMA_signal_8280), .Q (new_AGEMA_signal_8281) ) ;
    buf_clk new_AGEMA_reg_buffer_4824 ( .C (clk), .D (new_AGEMA_signal_8288), .Q (new_AGEMA_signal_8289) ) ;
    buf_clk new_AGEMA_reg_buffer_4832 ( .C (clk), .D (new_AGEMA_signal_8296), .Q (new_AGEMA_signal_8297) ) ;
    buf_clk new_AGEMA_reg_buffer_4840 ( .C (clk), .D (new_AGEMA_signal_8304), .Q (new_AGEMA_signal_8305) ) ;
    buf_clk new_AGEMA_reg_buffer_4848 ( .C (clk), .D (new_AGEMA_signal_8312), .Q (new_AGEMA_signal_8313) ) ;
    buf_clk new_AGEMA_reg_buffer_4856 ( .C (clk), .D (new_AGEMA_signal_8320), .Q (new_AGEMA_signal_8321) ) ;
    buf_clk new_AGEMA_reg_buffer_4864 ( .C (clk), .D (new_AGEMA_signal_8328), .Q (new_AGEMA_signal_8329) ) ;
    buf_clk new_AGEMA_reg_buffer_4872 ( .C (clk), .D (new_AGEMA_signal_8336), .Q (new_AGEMA_signal_8337) ) ;
    buf_clk new_AGEMA_reg_buffer_4880 ( .C (clk), .D (new_AGEMA_signal_8344), .Q (new_AGEMA_signal_8345) ) ;
    buf_clk new_AGEMA_reg_buffer_4888 ( .C (clk), .D (new_AGEMA_signal_8352), .Q (new_AGEMA_signal_8353) ) ;
    buf_clk new_AGEMA_reg_buffer_4896 ( .C (clk), .D (new_AGEMA_signal_8360), .Q (new_AGEMA_signal_8361) ) ;
    buf_clk new_AGEMA_reg_buffer_4904 ( .C (clk), .D (new_AGEMA_signal_8368), .Q (new_AGEMA_signal_8369) ) ;
    buf_clk new_AGEMA_reg_buffer_4912 ( .C (clk), .D (new_AGEMA_signal_8376), .Q (new_AGEMA_signal_8377) ) ;
    buf_clk new_AGEMA_reg_buffer_4920 ( .C (clk), .D (new_AGEMA_signal_8384), .Q (new_AGEMA_signal_8385) ) ;
    buf_clk new_AGEMA_reg_buffer_4928 ( .C (clk), .D (new_AGEMA_signal_8392), .Q (new_AGEMA_signal_8393) ) ;
    buf_clk new_AGEMA_reg_buffer_4936 ( .C (clk), .D (new_AGEMA_signal_8400), .Q (new_AGEMA_signal_8401) ) ;
    buf_clk new_AGEMA_reg_buffer_4944 ( .C (clk), .D (new_AGEMA_signal_8408), .Q (new_AGEMA_signal_8409) ) ;
    buf_clk new_AGEMA_reg_buffer_4952 ( .C (clk), .D (new_AGEMA_signal_8416), .Q (new_AGEMA_signal_8417) ) ;
    buf_clk new_AGEMA_reg_buffer_4960 ( .C (clk), .D (new_AGEMA_signal_8424), .Q (new_AGEMA_signal_8425) ) ;
    buf_clk new_AGEMA_reg_buffer_4968 ( .C (clk), .D (new_AGEMA_signal_8432), .Q (new_AGEMA_signal_8433) ) ;
    buf_clk new_AGEMA_reg_buffer_4976 ( .C (clk), .D (new_AGEMA_signal_8440), .Q (new_AGEMA_signal_8441) ) ;
    buf_clk new_AGEMA_reg_buffer_4984 ( .C (clk), .D (new_AGEMA_signal_8448), .Q (new_AGEMA_signal_8449) ) ;
    buf_clk new_AGEMA_reg_buffer_4992 ( .C (clk), .D (new_AGEMA_signal_8456), .Q (new_AGEMA_signal_8457) ) ;
    buf_clk new_AGEMA_reg_buffer_5000 ( .C (clk), .D (new_AGEMA_signal_8464), .Q (new_AGEMA_signal_8465) ) ;
    buf_clk new_AGEMA_reg_buffer_5008 ( .C (clk), .D (new_AGEMA_signal_8472), .Q (new_AGEMA_signal_8473) ) ;
    buf_clk new_AGEMA_reg_buffer_5016 ( .C (clk), .D (new_AGEMA_signal_8480), .Q (new_AGEMA_signal_8481) ) ;
    buf_clk new_AGEMA_reg_buffer_5024 ( .C (clk), .D (new_AGEMA_signal_8488), .Q (new_AGEMA_signal_8489) ) ;
    buf_clk new_AGEMA_reg_buffer_5032 ( .C (clk), .D (new_AGEMA_signal_8496), .Q (new_AGEMA_signal_8497) ) ;
    buf_clk new_AGEMA_reg_buffer_5040 ( .C (clk), .D (new_AGEMA_signal_8504), .Q (new_AGEMA_signal_8505) ) ;
    buf_clk new_AGEMA_reg_buffer_5048 ( .C (clk), .D (new_AGEMA_signal_8512), .Q (new_AGEMA_signal_8513) ) ;
    buf_clk new_AGEMA_reg_buffer_5056 ( .C (clk), .D (new_AGEMA_signal_8520), .Q (new_AGEMA_signal_8521) ) ;
    buf_clk new_AGEMA_reg_buffer_5064 ( .C (clk), .D (new_AGEMA_signal_8528), .Q (new_AGEMA_signal_8529) ) ;
    buf_clk new_AGEMA_reg_buffer_5072 ( .C (clk), .D (new_AGEMA_signal_8536), .Q (new_AGEMA_signal_8537) ) ;
    buf_clk new_AGEMA_reg_buffer_5080 ( .C (clk), .D (new_AGEMA_signal_8544), .Q (new_AGEMA_signal_8545) ) ;
    buf_clk new_AGEMA_reg_buffer_5088 ( .C (clk), .D (new_AGEMA_signal_8552), .Q (new_AGEMA_signal_8553) ) ;
    buf_clk new_AGEMA_reg_buffer_5096 ( .C (clk), .D (new_AGEMA_signal_8560), .Q (new_AGEMA_signal_8561) ) ;
    buf_clk new_AGEMA_reg_buffer_5104 ( .C (clk), .D (new_AGEMA_signal_8568), .Q (new_AGEMA_signal_8569) ) ;
    buf_clk new_AGEMA_reg_buffer_5112 ( .C (clk), .D (new_AGEMA_signal_8576), .Q (new_AGEMA_signal_8577) ) ;
    buf_clk new_AGEMA_reg_buffer_5120 ( .C (clk), .D (new_AGEMA_signal_8584), .Q (new_AGEMA_signal_8585) ) ;
    buf_clk new_AGEMA_reg_buffer_5128 ( .C (clk), .D (new_AGEMA_signal_8592), .Q (new_AGEMA_signal_8593) ) ;
    buf_clk new_AGEMA_reg_buffer_5136 ( .C (clk), .D (new_AGEMA_signal_8600), .Q (new_AGEMA_signal_8601) ) ;
    buf_clk new_AGEMA_reg_buffer_5144 ( .C (clk), .D (new_AGEMA_signal_8608), .Q (new_AGEMA_signal_8609) ) ;
    buf_clk new_AGEMA_reg_buffer_5152 ( .C (clk), .D (new_AGEMA_signal_8616), .Q (new_AGEMA_signal_8617) ) ;
    buf_clk new_AGEMA_reg_buffer_5160 ( .C (clk), .D (new_AGEMA_signal_8624), .Q (new_AGEMA_signal_8625) ) ;
    buf_clk new_AGEMA_reg_buffer_5168 ( .C (clk), .D (new_AGEMA_signal_8632), .Q (new_AGEMA_signal_8633) ) ;
    buf_clk new_AGEMA_reg_buffer_5176 ( .C (clk), .D (new_AGEMA_signal_8640), .Q (new_AGEMA_signal_8641) ) ;
    buf_clk new_AGEMA_reg_buffer_5184 ( .C (clk), .D (new_AGEMA_signal_8648), .Q (new_AGEMA_signal_8649) ) ;
    buf_clk new_AGEMA_reg_buffer_5192 ( .C (clk), .D (new_AGEMA_signal_8656), .Q (new_AGEMA_signal_8657) ) ;
    buf_clk new_AGEMA_reg_buffer_5200 ( .C (clk), .D (new_AGEMA_signal_8664), .Q (new_AGEMA_signal_8665) ) ;
    buf_clk new_AGEMA_reg_buffer_5208 ( .C (clk), .D (new_AGEMA_signal_8672), .Q (new_AGEMA_signal_8673) ) ;
    buf_clk new_AGEMA_reg_buffer_5216 ( .C (clk), .D (new_AGEMA_signal_8680), .Q (new_AGEMA_signal_8681) ) ;
    buf_clk new_AGEMA_reg_buffer_5224 ( .C (clk), .D (new_AGEMA_signal_8688), .Q (new_AGEMA_signal_8689) ) ;
    buf_clk new_AGEMA_reg_buffer_5232 ( .C (clk), .D (new_AGEMA_signal_8696), .Q (new_AGEMA_signal_8697) ) ;
    buf_clk new_AGEMA_reg_buffer_5240 ( .C (clk), .D (new_AGEMA_signal_8704), .Q (new_AGEMA_signal_8705) ) ;
    buf_clk new_AGEMA_reg_buffer_5248 ( .C (clk), .D (new_AGEMA_signal_8712), .Q (new_AGEMA_signal_8713) ) ;
    buf_clk new_AGEMA_reg_buffer_5256 ( .C (clk), .D (new_AGEMA_signal_8720), .Q (new_AGEMA_signal_8721) ) ;
    buf_clk new_AGEMA_reg_buffer_5264 ( .C (clk), .D (new_AGEMA_signal_8728), .Q (new_AGEMA_signal_8729) ) ;
    buf_clk new_AGEMA_reg_buffer_5272 ( .C (clk), .D (new_AGEMA_signal_8736), .Q (new_AGEMA_signal_8737) ) ;
    buf_clk new_AGEMA_reg_buffer_5280 ( .C (clk), .D (new_AGEMA_signal_8744), .Q (new_AGEMA_signal_8745) ) ;
    buf_clk new_AGEMA_reg_buffer_5288 ( .C (clk), .D (new_AGEMA_signal_8752), .Q (new_AGEMA_signal_8753) ) ;
    buf_clk new_AGEMA_reg_buffer_5296 ( .C (clk), .D (new_AGEMA_signal_8760), .Q (new_AGEMA_signal_8761) ) ;
    buf_clk new_AGEMA_reg_buffer_5304 ( .C (clk), .D (new_AGEMA_signal_8768), .Q (new_AGEMA_signal_8769) ) ;
    buf_clk new_AGEMA_reg_buffer_5312 ( .C (clk), .D (new_AGEMA_signal_8776), .Q (new_AGEMA_signal_8777) ) ;
    buf_clk new_AGEMA_reg_buffer_5320 ( .C (clk), .D (new_AGEMA_signal_8784), .Q (new_AGEMA_signal_8785) ) ;
    buf_clk new_AGEMA_reg_buffer_5328 ( .C (clk), .D (new_AGEMA_signal_8792), .Q (new_AGEMA_signal_8793) ) ;
    buf_clk new_AGEMA_reg_buffer_5336 ( .C (clk), .D (new_AGEMA_signal_8800), .Q (new_AGEMA_signal_8801) ) ;
    buf_clk new_AGEMA_reg_buffer_5344 ( .C (clk), .D (new_AGEMA_signal_8808), .Q (new_AGEMA_signal_8809) ) ;
    buf_clk new_AGEMA_reg_buffer_5352 ( .C (clk), .D (new_AGEMA_signal_8816), .Q (new_AGEMA_signal_8817) ) ;
    buf_clk new_AGEMA_reg_buffer_5360 ( .C (clk), .D (new_AGEMA_signal_8824), .Q (new_AGEMA_signal_8825) ) ;
    buf_clk new_AGEMA_reg_buffer_5368 ( .C (clk), .D (new_AGEMA_signal_8832), .Q (new_AGEMA_signal_8833) ) ;
    buf_clk new_AGEMA_reg_buffer_5376 ( .C (clk), .D (new_AGEMA_signal_8840), .Q (new_AGEMA_signal_8841) ) ;
    buf_clk new_AGEMA_reg_buffer_5384 ( .C (clk), .D (new_AGEMA_signal_8848), .Q (new_AGEMA_signal_8849) ) ;
    buf_clk new_AGEMA_reg_buffer_5392 ( .C (clk), .D (new_AGEMA_signal_8856), .Q (new_AGEMA_signal_8857) ) ;
    buf_clk new_AGEMA_reg_buffer_5400 ( .C (clk), .D (new_AGEMA_signal_8864), .Q (new_AGEMA_signal_8865) ) ;
    buf_clk new_AGEMA_reg_buffer_5410 ( .C (clk), .D (new_AGEMA_signal_8874), .Q (new_AGEMA_signal_8875) ) ;
    buf_clk new_AGEMA_reg_buffer_5418 ( .C (clk), .D (new_AGEMA_signal_8882), .Q (new_AGEMA_signal_8883) ) ;
    buf_clk new_AGEMA_reg_buffer_5426 ( .C (clk), .D (new_AGEMA_signal_8890), .Q (new_AGEMA_signal_8891) ) ;
    buf_clk new_AGEMA_reg_buffer_5434 ( .C (clk), .D (new_AGEMA_signal_8898), .Q (new_AGEMA_signal_8899) ) ;
    buf_clk new_AGEMA_reg_buffer_5442 ( .C (clk), .D (new_AGEMA_signal_8906), .Q (new_AGEMA_signal_8907) ) ;
    buf_clk new_AGEMA_reg_buffer_5450 ( .C (clk), .D (new_AGEMA_signal_8914), .Q (new_AGEMA_signal_8915) ) ;
    buf_clk new_AGEMA_reg_buffer_5458 ( .C (clk), .D (new_AGEMA_signal_8922), .Q (new_AGEMA_signal_8923) ) ;
    buf_clk new_AGEMA_reg_buffer_5466 ( .C (clk), .D (new_AGEMA_signal_8930), .Q (new_AGEMA_signal_8931) ) ;
    buf_clk new_AGEMA_reg_buffer_5474 ( .C (clk), .D (new_AGEMA_signal_8938), .Q (new_AGEMA_signal_8939) ) ;
    buf_clk new_AGEMA_reg_buffer_5482 ( .C (clk), .D (new_AGEMA_signal_8946), .Q (new_AGEMA_signal_8947) ) ;
    buf_clk new_AGEMA_reg_buffer_5490 ( .C (clk), .D (new_AGEMA_signal_8954), .Q (new_AGEMA_signal_8955) ) ;
    buf_clk new_AGEMA_reg_buffer_5498 ( .C (clk), .D (new_AGEMA_signal_8962), .Q (new_AGEMA_signal_8963) ) ;
    buf_clk new_AGEMA_reg_buffer_5506 ( .C (clk), .D (new_AGEMA_signal_8970), .Q (new_AGEMA_signal_8971) ) ;
    buf_clk new_AGEMA_reg_buffer_5514 ( .C (clk), .D (new_AGEMA_signal_8978), .Q (new_AGEMA_signal_8979) ) ;
    buf_clk new_AGEMA_reg_buffer_5522 ( .C (clk), .D (new_AGEMA_signal_8986), .Q (new_AGEMA_signal_8987) ) ;
    buf_clk new_AGEMA_reg_buffer_5530 ( .C (clk), .D (new_AGEMA_signal_8994), .Q (new_AGEMA_signal_8995) ) ;
    buf_clk new_AGEMA_reg_buffer_5538 ( .C (clk), .D (new_AGEMA_signal_9002), .Q (new_AGEMA_signal_9003) ) ;
    buf_clk new_AGEMA_reg_buffer_5546 ( .C (clk), .D (new_AGEMA_signal_9010), .Q (new_AGEMA_signal_9011) ) ;
    buf_clk new_AGEMA_reg_buffer_5554 ( .C (clk), .D (new_AGEMA_signal_9018), .Q (new_AGEMA_signal_9019) ) ;
    buf_clk new_AGEMA_reg_buffer_5562 ( .C (clk), .D (new_AGEMA_signal_9026), .Q (new_AGEMA_signal_9027) ) ;
    buf_clk new_AGEMA_reg_buffer_5570 ( .C (clk), .D (new_AGEMA_signal_9034), .Q (new_AGEMA_signal_9035) ) ;
    buf_clk new_AGEMA_reg_buffer_5578 ( .C (clk), .D (new_AGEMA_signal_9042), .Q (new_AGEMA_signal_9043) ) ;
    buf_clk new_AGEMA_reg_buffer_5586 ( .C (clk), .D (new_AGEMA_signal_9050), .Q (new_AGEMA_signal_9051) ) ;
    buf_clk new_AGEMA_reg_buffer_5594 ( .C (clk), .D (new_AGEMA_signal_9058), .Q (new_AGEMA_signal_9059) ) ;
    buf_clk new_AGEMA_reg_buffer_5602 ( .C (clk), .D (new_AGEMA_signal_9066), .Q (new_AGEMA_signal_9067) ) ;
    buf_clk new_AGEMA_reg_buffer_5610 ( .C (clk), .D (new_AGEMA_signal_9074), .Q (new_AGEMA_signal_9075) ) ;
    buf_clk new_AGEMA_reg_buffer_5618 ( .C (clk), .D (new_AGEMA_signal_9082), .Q (new_AGEMA_signal_9083) ) ;
    buf_clk new_AGEMA_reg_buffer_5626 ( .C (clk), .D (new_AGEMA_signal_9090), .Q (new_AGEMA_signal_9091) ) ;
    buf_clk new_AGEMA_reg_buffer_5634 ( .C (clk), .D (new_AGEMA_signal_9098), .Q (new_AGEMA_signal_9099) ) ;
    buf_clk new_AGEMA_reg_buffer_5642 ( .C (clk), .D (new_AGEMA_signal_9106), .Q (new_AGEMA_signal_9107) ) ;
    buf_clk new_AGEMA_reg_buffer_5650 ( .C (clk), .D (new_AGEMA_signal_9114), .Q (new_AGEMA_signal_9115) ) ;
    buf_clk new_AGEMA_reg_buffer_5658 ( .C (clk), .D (new_AGEMA_signal_9122), .Q (new_AGEMA_signal_9123) ) ;
    buf_clk new_AGEMA_reg_buffer_5666 ( .C (clk), .D (new_AGEMA_signal_9130), .Q (new_AGEMA_signal_9131) ) ;
    buf_clk new_AGEMA_reg_buffer_5674 ( .C (clk), .D (new_AGEMA_signal_9138), .Q (new_AGEMA_signal_9139) ) ;
    buf_clk new_AGEMA_reg_buffer_5682 ( .C (clk), .D (new_AGEMA_signal_9146), .Q (new_AGEMA_signal_9147) ) ;
    buf_clk new_AGEMA_reg_buffer_5690 ( .C (clk), .D (new_AGEMA_signal_9154), .Q (new_AGEMA_signal_9155) ) ;
    buf_clk new_AGEMA_reg_buffer_5698 ( .C (clk), .D (new_AGEMA_signal_9162), .Q (new_AGEMA_signal_9163) ) ;
    buf_clk new_AGEMA_reg_buffer_5706 ( .C (clk), .D (new_AGEMA_signal_9170), .Q (new_AGEMA_signal_9171) ) ;
    buf_clk new_AGEMA_reg_buffer_5714 ( .C (clk), .D (new_AGEMA_signal_9178), .Q (new_AGEMA_signal_9179) ) ;
    buf_clk new_AGEMA_reg_buffer_5722 ( .C (clk), .D (new_AGEMA_signal_9186), .Q (new_AGEMA_signal_9187) ) ;
    buf_clk new_AGEMA_reg_buffer_5730 ( .C (clk), .D (new_AGEMA_signal_9194), .Q (new_AGEMA_signal_9195) ) ;
    buf_clk new_AGEMA_reg_buffer_5738 ( .C (clk), .D (new_AGEMA_signal_9202), .Q (new_AGEMA_signal_9203) ) ;
    buf_clk new_AGEMA_reg_buffer_5746 ( .C (clk), .D (new_AGEMA_signal_9210), .Q (new_AGEMA_signal_9211) ) ;
    buf_clk new_AGEMA_reg_buffer_5754 ( .C (clk), .D (new_AGEMA_signal_9218), .Q (new_AGEMA_signal_9219) ) ;
    buf_clk new_AGEMA_reg_buffer_5762 ( .C (clk), .D (new_AGEMA_signal_9226), .Q (new_AGEMA_signal_9227) ) ;
    buf_clk new_AGEMA_reg_buffer_5770 ( .C (clk), .D (new_AGEMA_signal_9234), .Q (new_AGEMA_signal_9235) ) ;
    buf_clk new_AGEMA_reg_buffer_5778 ( .C (clk), .D (new_AGEMA_signal_9242), .Q (new_AGEMA_signal_9243) ) ;
    buf_clk new_AGEMA_reg_buffer_5786 ( .C (clk), .D (new_AGEMA_signal_9250), .Q (new_AGEMA_signal_9251) ) ;
    buf_clk new_AGEMA_reg_buffer_5794 ( .C (clk), .D (new_AGEMA_signal_9258), .Q (new_AGEMA_signal_9259) ) ;
    buf_clk new_AGEMA_reg_buffer_5802 ( .C (clk), .D (new_AGEMA_signal_9266), .Q (new_AGEMA_signal_9267) ) ;
    buf_clk new_AGEMA_reg_buffer_5810 ( .C (clk), .D (new_AGEMA_signal_9274), .Q (new_AGEMA_signal_9275) ) ;
    buf_clk new_AGEMA_reg_buffer_5818 ( .C (clk), .D (new_AGEMA_signal_9282), .Q (new_AGEMA_signal_9283) ) ;
    buf_clk new_AGEMA_reg_buffer_5826 ( .C (clk), .D (new_AGEMA_signal_9290), .Q (new_AGEMA_signal_9291) ) ;
    buf_clk new_AGEMA_reg_buffer_5834 ( .C (clk), .D (new_AGEMA_signal_9298), .Q (new_AGEMA_signal_9299) ) ;
    buf_clk new_AGEMA_reg_buffer_5842 ( .C (clk), .D (new_AGEMA_signal_9306), .Q (new_AGEMA_signal_9307) ) ;
    buf_clk new_AGEMA_reg_buffer_5850 ( .C (clk), .D (new_AGEMA_signal_9314), .Q (new_AGEMA_signal_9315) ) ;
    buf_clk new_AGEMA_reg_buffer_5858 ( .C (clk), .D (new_AGEMA_signal_9322), .Q (new_AGEMA_signal_9323) ) ;
    buf_clk new_AGEMA_reg_buffer_5866 ( .C (clk), .D (new_AGEMA_signal_9330), .Q (new_AGEMA_signal_9331) ) ;
    buf_clk new_AGEMA_reg_buffer_5874 ( .C (clk), .D (new_AGEMA_signal_9338), .Q (new_AGEMA_signal_9339) ) ;
    buf_clk new_AGEMA_reg_buffer_5882 ( .C (clk), .D (new_AGEMA_signal_9346), .Q (new_AGEMA_signal_9347) ) ;
    buf_clk new_AGEMA_reg_buffer_5890 ( .C (clk), .D (new_AGEMA_signal_9354), .Q (new_AGEMA_signal_9355) ) ;
    buf_clk new_AGEMA_reg_buffer_5898 ( .C (clk), .D (new_AGEMA_signal_9362), .Q (new_AGEMA_signal_9363) ) ;
    buf_clk new_AGEMA_reg_buffer_5906 ( .C (clk), .D (new_AGEMA_signal_9370), .Q (new_AGEMA_signal_9371) ) ;
    buf_clk new_AGEMA_reg_buffer_5914 ( .C (clk), .D (new_AGEMA_signal_9378), .Q (new_AGEMA_signal_9379) ) ;
    buf_clk new_AGEMA_reg_buffer_5922 ( .C (clk), .D (new_AGEMA_signal_9386), .Q (new_AGEMA_signal_9387) ) ;
    buf_clk new_AGEMA_reg_buffer_5930 ( .C (clk), .D (new_AGEMA_signal_9394), .Q (new_AGEMA_signal_9395) ) ;
    buf_clk new_AGEMA_reg_buffer_5938 ( .C (clk), .D (new_AGEMA_signal_9402), .Q (new_AGEMA_signal_9403) ) ;
    buf_clk new_AGEMA_reg_buffer_5946 ( .C (clk), .D (new_AGEMA_signal_9410), .Q (new_AGEMA_signal_9411) ) ;
    buf_clk new_AGEMA_reg_buffer_5954 ( .C (clk), .D (new_AGEMA_signal_9418), .Q (new_AGEMA_signal_9419) ) ;
    buf_clk new_AGEMA_reg_buffer_5962 ( .C (clk), .D (new_AGEMA_signal_9426), .Q (new_AGEMA_signal_9427) ) ;
    buf_clk new_AGEMA_reg_buffer_5970 ( .C (clk), .D (new_AGEMA_signal_9434), .Q (new_AGEMA_signal_9435) ) ;
    buf_clk new_AGEMA_reg_buffer_5978 ( .C (clk), .D (new_AGEMA_signal_9442), .Q (new_AGEMA_signal_9443) ) ;
    buf_clk new_AGEMA_reg_buffer_5986 ( .C (clk), .D (new_AGEMA_signal_9450), .Q (new_AGEMA_signal_9451) ) ;
    buf_clk new_AGEMA_reg_buffer_5994 ( .C (clk), .D (new_AGEMA_signal_9458), .Q (new_AGEMA_signal_9459) ) ;
    buf_clk new_AGEMA_reg_buffer_6002 ( .C (clk), .D (new_AGEMA_signal_9466), .Q (new_AGEMA_signal_9467) ) ;
    buf_clk new_AGEMA_reg_buffer_6010 ( .C (clk), .D (new_AGEMA_signal_9474), .Q (new_AGEMA_signal_9475) ) ;
    buf_clk new_AGEMA_reg_buffer_6018 ( .C (clk), .D (new_AGEMA_signal_9482), .Q (new_AGEMA_signal_9483) ) ;
    buf_clk new_AGEMA_reg_buffer_6026 ( .C (clk), .D (new_AGEMA_signal_9490), .Q (new_AGEMA_signal_9491) ) ;
    buf_clk new_AGEMA_reg_buffer_6034 ( .C (clk), .D (new_AGEMA_signal_9498), .Q (new_AGEMA_signal_9499) ) ;
    buf_clk new_AGEMA_reg_buffer_6042 ( .C (clk), .D (new_AGEMA_signal_9506), .Q (new_AGEMA_signal_9507) ) ;
    buf_clk new_AGEMA_reg_buffer_6050 ( .C (clk), .D (new_AGEMA_signal_9514), .Q (new_AGEMA_signal_9515) ) ;
    buf_clk new_AGEMA_reg_buffer_6058 ( .C (clk), .D (new_AGEMA_signal_9522), .Q (new_AGEMA_signal_9523) ) ;
    buf_clk new_AGEMA_reg_buffer_6066 ( .C (clk), .D (new_AGEMA_signal_9530), .Q (new_AGEMA_signal_9531) ) ;
    buf_clk new_AGEMA_reg_buffer_6074 ( .C (clk), .D (new_AGEMA_signal_9538), .Q (new_AGEMA_signal_9539) ) ;
    buf_clk new_AGEMA_reg_buffer_6082 ( .C (clk), .D (new_AGEMA_signal_9546), .Q (new_AGEMA_signal_9547) ) ;
    buf_clk new_AGEMA_reg_buffer_6090 ( .C (clk), .D (new_AGEMA_signal_9554), .Q (new_AGEMA_signal_9555) ) ;
    buf_clk new_AGEMA_reg_buffer_6098 ( .C (clk), .D (new_AGEMA_signal_9562), .Q (new_AGEMA_signal_9563) ) ;
    buf_clk new_AGEMA_reg_buffer_6106 ( .C (clk), .D (new_AGEMA_signal_9570), .Q (new_AGEMA_signal_9571) ) ;
    buf_clk new_AGEMA_reg_buffer_6114 ( .C (clk), .D (new_AGEMA_signal_9578), .Q (new_AGEMA_signal_9579) ) ;
    buf_clk new_AGEMA_reg_buffer_6122 ( .C (clk), .D (new_AGEMA_signal_9586), .Q (new_AGEMA_signal_9587) ) ;
    buf_clk new_AGEMA_reg_buffer_6130 ( .C (clk), .D (new_AGEMA_signal_9594), .Q (new_AGEMA_signal_9595) ) ;
    buf_clk new_AGEMA_reg_buffer_6138 ( .C (clk), .D (new_AGEMA_signal_9602), .Q (new_AGEMA_signal_9603) ) ;
    buf_clk new_AGEMA_reg_buffer_6146 ( .C (clk), .D (new_AGEMA_signal_9610), .Q (new_AGEMA_signal_9611) ) ;
    buf_clk new_AGEMA_reg_buffer_6154 ( .C (clk), .D (new_AGEMA_signal_9618), .Q (new_AGEMA_signal_9619) ) ;
    buf_clk new_AGEMA_reg_buffer_6162 ( .C (clk), .D (new_AGEMA_signal_9626), .Q (new_AGEMA_signal_9627) ) ;
    buf_clk new_AGEMA_reg_buffer_6170 ( .C (clk), .D (new_AGEMA_signal_9634), .Q (new_AGEMA_signal_9635) ) ;
    buf_clk new_AGEMA_reg_buffer_6174 ( .C (clk), .D (new_AGEMA_signal_9638), .Q (new_AGEMA_signal_9639) ) ;
    buf_clk new_AGEMA_reg_buffer_6176 ( .C (clk), .D (new_AGEMA_signal_9640), .Q (new_AGEMA_signal_9641) ) ;
    buf_clk new_AGEMA_reg_buffer_6178 ( .C (clk), .D (new_AGEMA_signal_9642), .Q (new_AGEMA_signal_9643) ) ;
    buf_clk new_AGEMA_reg_buffer_6182 ( .C (clk), .D (new_AGEMA_signal_9646), .Q (new_AGEMA_signal_9647) ) ;
    buf_clk new_AGEMA_reg_buffer_6186 ( .C (clk), .D (new_AGEMA_signal_9650), .Q (new_AGEMA_signal_9651) ) ;
    buf_clk new_AGEMA_reg_buffer_6190 ( .C (clk), .D (new_AGEMA_signal_9654), .Q (new_AGEMA_signal_9655) ) ;
    buf_clk new_AGEMA_reg_buffer_6192 ( .C (clk), .D (new_AGEMA_signal_9656), .Q (new_AGEMA_signal_9657) ) ;
    buf_clk new_AGEMA_reg_buffer_6194 ( .C (clk), .D (new_AGEMA_signal_9658), .Q (new_AGEMA_signal_9659) ) ;
    buf_clk new_AGEMA_reg_buffer_6196 ( .C (clk), .D (new_AGEMA_signal_9660), .Q (new_AGEMA_signal_9661) ) ;
    buf_clk new_AGEMA_reg_buffer_6200 ( .C (clk), .D (new_AGEMA_signal_9664), .Q (new_AGEMA_signal_9665) ) ;
    buf_clk new_AGEMA_reg_buffer_6204 ( .C (clk), .D (new_AGEMA_signal_9668), .Q (new_AGEMA_signal_9669) ) ;
    buf_clk new_AGEMA_reg_buffer_6208 ( .C (clk), .D (new_AGEMA_signal_9672), .Q (new_AGEMA_signal_9673) ) ;
    buf_clk new_AGEMA_reg_buffer_6210 ( .C (clk), .D (new_AGEMA_signal_9674), .Q (new_AGEMA_signal_9675) ) ;
    buf_clk new_AGEMA_reg_buffer_6212 ( .C (clk), .D (new_AGEMA_signal_9676), .Q (new_AGEMA_signal_9677) ) ;
    buf_clk new_AGEMA_reg_buffer_6214 ( .C (clk), .D (new_AGEMA_signal_9678), .Q (new_AGEMA_signal_9679) ) ;
    buf_clk new_AGEMA_reg_buffer_6218 ( .C (clk), .D (new_AGEMA_signal_9682), .Q (new_AGEMA_signal_9683) ) ;
    buf_clk new_AGEMA_reg_buffer_6222 ( .C (clk), .D (new_AGEMA_signal_9686), .Q (new_AGEMA_signal_9687) ) ;
    buf_clk new_AGEMA_reg_buffer_6226 ( .C (clk), .D (new_AGEMA_signal_9690), .Q (new_AGEMA_signal_9691) ) ;
    buf_clk new_AGEMA_reg_buffer_6228 ( .C (clk), .D (new_AGEMA_signal_9692), .Q (new_AGEMA_signal_9693) ) ;
    buf_clk new_AGEMA_reg_buffer_6230 ( .C (clk), .D (new_AGEMA_signal_9694), .Q (new_AGEMA_signal_9695) ) ;
    buf_clk new_AGEMA_reg_buffer_6232 ( .C (clk), .D (new_AGEMA_signal_9696), .Q (new_AGEMA_signal_9697) ) ;
    buf_clk new_AGEMA_reg_buffer_6236 ( .C (clk), .D (new_AGEMA_signal_9700), .Q (new_AGEMA_signal_9701) ) ;
    buf_clk new_AGEMA_reg_buffer_6240 ( .C (clk), .D (new_AGEMA_signal_9704), .Q (new_AGEMA_signal_9705) ) ;
    buf_clk new_AGEMA_reg_buffer_6244 ( .C (clk), .D (new_AGEMA_signal_9708), .Q (new_AGEMA_signal_9709) ) ;
    buf_clk new_AGEMA_reg_buffer_6246 ( .C (clk), .D (new_AGEMA_signal_9710), .Q (new_AGEMA_signal_9711) ) ;
    buf_clk new_AGEMA_reg_buffer_6248 ( .C (clk), .D (new_AGEMA_signal_9712), .Q (new_AGEMA_signal_9713) ) ;
    buf_clk new_AGEMA_reg_buffer_6250 ( .C (clk), .D (new_AGEMA_signal_9714), .Q (new_AGEMA_signal_9715) ) ;
    buf_clk new_AGEMA_reg_buffer_6254 ( .C (clk), .D (new_AGEMA_signal_9718), .Q (new_AGEMA_signal_9719) ) ;
    buf_clk new_AGEMA_reg_buffer_6258 ( .C (clk), .D (new_AGEMA_signal_9722), .Q (new_AGEMA_signal_9723) ) ;
    buf_clk new_AGEMA_reg_buffer_6262 ( .C (clk), .D (new_AGEMA_signal_9726), .Q (new_AGEMA_signal_9727) ) ;
    buf_clk new_AGEMA_reg_buffer_6264 ( .C (clk), .D (new_AGEMA_signal_9728), .Q (new_AGEMA_signal_9729) ) ;
    buf_clk new_AGEMA_reg_buffer_6266 ( .C (clk), .D (new_AGEMA_signal_9730), .Q (new_AGEMA_signal_9731) ) ;
    buf_clk new_AGEMA_reg_buffer_6268 ( .C (clk), .D (new_AGEMA_signal_9732), .Q (new_AGEMA_signal_9733) ) ;
    buf_clk new_AGEMA_reg_buffer_6272 ( .C (clk), .D (new_AGEMA_signal_9736), .Q (new_AGEMA_signal_9737) ) ;
    buf_clk new_AGEMA_reg_buffer_6276 ( .C (clk), .D (new_AGEMA_signal_9740), .Q (new_AGEMA_signal_9741) ) ;
    buf_clk new_AGEMA_reg_buffer_6280 ( .C (clk), .D (new_AGEMA_signal_9744), .Q (new_AGEMA_signal_9745) ) ;
    buf_clk new_AGEMA_reg_buffer_6282 ( .C (clk), .D (new_AGEMA_signal_9746), .Q (new_AGEMA_signal_9747) ) ;
    buf_clk new_AGEMA_reg_buffer_6284 ( .C (clk), .D (new_AGEMA_signal_9748), .Q (new_AGEMA_signal_9749) ) ;
    buf_clk new_AGEMA_reg_buffer_6286 ( .C (clk), .D (new_AGEMA_signal_9750), .Q (new_AGEMA_signal_9751) ) ;
    buf_clk new_AGEMA_reg_buffer_6290 ( .C (clk), .D (new_AGEMA_signal_9754), .Q (new_AGEMA_signal_9755) ) ;
    buf_clk new_AGEMA_reg_buffer_6294 ( .C (clk), .D (new_AGEMA_signal_9758), .Q (new_AGEMA_signal_9759) ) ;
    buf_clk new_AGEMA_reg_buffer_6298 ( .C (clk), .D (new_AGEMA_signal_9762), .Q (new_AGEMA_signal_9763) ) ;
    buf_clk new_AGEMA_reg_buffer_6300 ( .C (clk), .D (new_AGEMA_signal_9764), .Q (new_AGEMA_signal_9765) ) ;
    buf_clk new_AGEMA_reg_buffer_6302 ( .C (clk), .D (new_AGEMA_signal_9766), .Q (new_AGEMA_signal_9767) ) ;
    buf_clk new_AGEMA_reg_buffer_6304 ( .C (clk), .D (new_AGEMA_signal_9768), .Q (new_AGEMA_signal_9769) ) ;
    buf_clk new_AGEMA_reg_buffer_6308 ( .C (clk), .D (new_AGEMA_signal_9772), .Q (new_AGEMA_signal_9773) ) ;
    buf_clk new_AGEMA_reg_buffer_6312 ( .C (clk), .D (new_AGEMA_signal_9776), .Q (new_AGEMA_signal_9777) ) ;
    buf_clk new_AGEMA_reg_buffer_6316 ( .C (clk), .D (new_AGEMA_signal_9780), .Q (new_AGEMA_signal_9781) ) ;
    buf_clk new_AGEMA_reg_buffer_6318 ( .C (clk), .D (new_AGEMA_signal_9782), .Q (new_AGEMA_signal_9783) ) ;
    buf_clk new_AGEMA_reg_buffer_6320 ( .C (clk), .D (new_AGEMA_signal_9784), .Q (new_AGEMA_signal_9785) ) ;
    buf_clk new_AGEMA_reg_buffer_6322 ( .C (clk), .D (new_AGEMA_signal_9786), .Q (new_AGEMA_signal_9787) ) ;
    buf_clk new_AGEMA_reg_buffer_6326 ( .C (clk), .D (new_AGEMA_signal_9790), .Q (new_AGEMA_signal_9791) ) ;
    buf_clk new_AGEMA_reg_buffer_6330 ( .C (clk), .D (new_AGEMA_signal_9794), .Q (new_AGEMA_signal_9795) ) ;
    buf_clk new_AGEMA_reg_buffer_6334 ( .C (clk), .D (new_AGEMA_signal_9798), .Q (new_AGEMA_signal_9799) ) ;
    buf_clk new_AGEMA_reg_buffer_6336 ( .C (clk), .D (new_AGEMA_signal_9800), .Q (new_AGEMA_signal_9801) ) ;
    buf_clk new_AGEMA_reg_buffer_6338 ( .C (clk), .D (new_AGEMA_signal_9802), .Q (new_AGEMA_signal_9803) ) ;
    buf_clk new_AGEMA_reg_buffer_6340 ( .C (clk), .D (new_AGEMA_signal_9804), .Q (new_AGEMA_signal_9805) ) ;
    buf_clk new_AGEMA_reg_buffer_6344 ( .C (clk), .D (new_AGEMA_signal_9808), .Q (new_AGEMA_signal_9809) ) ;
    buf_clk new_AGEMA_reg_buffer_6348 ( .C (clk), .D (new_AGEMA_signal_9812), .Q (new_AGEMA_signal_9813) ) ;
    buf_clk new_AGEMA_reg_buffer_6352 ( .C (clk), .D (new_AGEMA_signal_9816), .Q (new_AGEMA_signal_9817) ) ;
    buf_clk new_AGEMA_reg_buffer_6354 ( .C (clk), .D (new_AGEMA_signal_9818), .Q (new_AGEMA_signal_9819) ) ;
    buf_clk new_AGEMA_reg_buffer_6356 ( .C (clk), .D (new_AGEMA_signal_9820), .Q (new_AGEMA_signal_9821) ) ;
    buf_clk new_AGEMA_reg_buffer_6358 ( .C (clk), .D (new_AGEMA_signal_9822), .Q (new_AGEMA_signal_9823) ) ;
    buf_clk new_AGEMA_reg_buffer_6362 ( .C (clk), .D (new_AGEMA_signal_9826), .Q (new_AGEMA_signal_9827) ) ;
    buf_clk new_AGEMA_reg_buffer_6366 ( .C (clk), .D (new_AGEMA_signal_9830), .Q (new_AGEMA_signal_9831) ) ;
    buf_clk new_AGEMA_reg_buffer_6370 ( .C (clk), .D (new_AGEMA_signal_9834), .Q (new_AGEMA_signal_9835) ) ;
    buf_clk new_AGEMA_reg_buffer_6372 ( .C (clk), .D (new_AGEMA_signal_9836), .Q (new_AGEMA_signal_9837) ) ;
    buf_clk new_AGEMA_reg_buffer_6374 ( .C (clk), .D (new_AGEMA_signal_9838), .Q (new_AGEMA_signal_9839) ) ;
    buf_clk new_AGEMA_reg_buffer_6376 ( .C (clk), .D (new_AGEMA_signal_9840), .Q (new_AGEMA_signal_9841) ) ;
    buf_clk new_AGEMA_reg_buffer_6380 ( .C (clk), .D (new_AGEMA_signal_9844), .Q (new_AGEMA_signal_9845) ) ;
    buf_clk new_AGEMA_reg_buffer_6384 ( .C (clk), .D (new_AGEMA_signal_9848), .Q (new_AGEMA_signal_9849) ) ;
    buf_clk new_AGEMA_reg_buffer_6388 ( .C (clk), .D (new_AGEMA_signal_9852), .Q (new_AGEMA_signal_9853) ) ;
    buf_clk new_AGEMA_reg_buffer_6390 ( .C (clk), .D (new_AGEMA_signal_9854), .Q (new_AGEMA_signal_9855) ) ;
    buf_clk new_AGEMA_reg_buffer_6392 ( .C (clk), .D (new_AGEMA_signal_9856), .Q (new_AGEMA_signal_9857) ) ;
    buf_clk new_AGEMA_reg_buffer_6394 ( .C (clk), .D (new_AGEMA_signal_9858), .Q (new_AGEMA_signal_9859) ) ;
    buf_clk new_AGEMA_reg_buffer_6398 ( .C (clk), .D (new_AGEMA_signal_9862), .Q (new_AGEMA_signal_9863) ) ;
    buf_clk new_AGEMA_reg_buffer_6402 ( .C (clk), .D (new_AGEMA_signal_9866), .Q (new_AGEMA_signal_9867) ) ;
    buf_clk new_AGEMA_reg_buffer_6406 ( .C (clk), .D (new_AGEMA_signal_9870), .Q (new_AGEMA_signal_9871) ) ;
    buf_clk new_AGEMA_reg_buffer_6408 ( .C (clk), .D (new_AGEMA_signal_9872), .Q (new_AGEMA_signal_9873) ) ;
    buf_clk new_AGEMA_reg_buffer_6410 ( .C (clk), .D (new_AGEMA_signal_9874), .Q (new_AGEMA_signal_9875) ) ;
    buf_clk new_AGEMA_reg_buffer_6412 ( .C (clk), .D (new_AGEMA_signal_9876), .Q (new_AGEMA_signal_9877) ) ;
    buf_clk new_AGEMA_reg_buffer_6416 ( .C (clk), .D (new_AGEMA_signal_9880), .Q (new_AGEMA_signal_9881) ) ;
    buf_clk new_AGEMA_reg_buffer_6420 ( .C (clk), .D (new_AGEMA_signal_9884), .Q (new_AGEMA_signal_9885) ) ;
    buf_clk new_AGEMA_reg_buffer_6424 ( .C (clk), .D (new_AGEMA_signal_9888), .Q (new_AGEMA_signal_9889) ) ;
    buf_clk new_AGEMA_reg_buffer_6426 ( .C (clk), .D (new_AGEMA_signal_9890), .Q (new_AGEMA_signal_9891) ) ;
    buf_clk new_AGEMA_reg_buffer_6428 ( .C (clk), .D (new_AGEMA_signal_9892), .Q (new_AGEMA_signal_9893) ) ;
    buf_clk new_AGEMA_reg_buffer_6430 ( .C (clk), .D (new_AGEMA_signal_9894), .Q (new_AGEMA_signal_9895) ) ;
    buf_clk new_AGEMA_reg_buffer_6434 ( .C (clk), .D (new_AGEMA_signal_9898), .Q (new_AGEMA_signal_9899) ) ;
    buf_clk new_AGEMA_reg_buffer_6438 ( .C (clk), .D (new_AGEMA_signal_9902), .Q (new_AGEMA_signal_9903) ) ;
    buf_clk new_AGEMA_reg_buffer_6442 ( .C (clk), .D (new_AGEMA_signal_9906), .Q (new_AGEMA_signal_9907) ) ;
    buf_clk new_AGEMA_reg_buffer_6444 ( .C (clk), .D (new_AGEMA_signal_9908), .Q (new_AGEMA_signal_9909) ) ;
    buf_clk new_AGEMA_reg_buffer_6446 ( .C (clk), .D (new_AGEMA_signal_9910), .Q (new_AGEMA_signal_9911) ) ;
    buf_clk new_AGEMA_reg_buffer_6448 ( .C (clk), .D (new_AGEMA_signal_9912), .Q (new_AGEMA_signal_9913) ) ;
    buf_clk new_AGEMA_reg_buffer_6452 ( .C (clk), .D (new_AGEMA_signal_9916), .Q (new_AGEMA_signal_9917) ) ;
    buf_clk new_AGEMA_reg_buffer_6456 ( .C (clk), .D (new_AGEMA_signal_9920), .Q (new_AGEMA_signal_9921) ) ;
    buf_clk new_AGEMA_reg_buffer_6460 ( .C (clk), .D (new_AGEMA_signal_9924), .Q (new_AGEMA_signal_9925) ) ;
    buf_clk new_AGEMA_reg_buffer_6468 ( .C (clk), .D (new_AGEMA_signal_9932), .Q (new_AGEMA_signal_9933) ) ;
    buf_clk new_AGEMA_reg_buffer_6476 ( .C (clk), .D (new_AGEMA_signal_9940), .Q (new_AGEMA_signal_9941) ) ;
    buf_clk new_AGEMA_reg_buffer_6484 ( .C (clk), .D (new_AGEMA_signal_9948), .Q (new_AGEMA_signal_9949) ) ;
    buf_clk new_AGEMA_reg_buffer_6492 ( .C (clk), .D (new_AGEMA_signal_9956), .Q (new_AGEMA_signal_9957) ) ;

    /* cells in depth 7 */
    buf_clk new_AGEMA_reg_buffer_1255 ( .C (clk), .D (new_AGEMA_signal_4720), .Q (new_AGEMA_signal_4721) ) ;
    buf_clk new_AGEMA_reg_buffer_1257 ( .C (clk), .D (new_AGEMA_signal_4722), .Q (new_AGEMA_signal_4723) ) ;
    buf_clk new_AGEMA_reg_buffer_1259 ( .C (clk), .D (new_AGEMA_signal_4724), .Q (new_AGEMA_signal_4725) ) ;
    buf_clk new_AGEMA_reg_buffer_1261 ( .C (clk), .D (new_AGEMA_signal_4726), .Q (new_AGEMA_signal_4727) ) ;
    buf_clk new_AGEMA_reg_buffer_1263 ( .C (clk), .D (new_AGEMA_signal_4728), .Q (new_AGEMA_signal_4729) ) ;
    buf_clk new_AGEMA_reg_buffer_1265 ( .C (clk), .D (new_AGEMA_signal_4730), .Q (new_AGEMA_signal_4731) ) ;
    buf_clk new_AGEMA_reg_buffer_1267 ( .C (clk), .D (new_AGEMA_signal_4732), .Q (new_AGEMA_signal_4733) ) ;
    buf_clk new_AGEMA_reg_buffer_1269 ( .C (clk), .D (new_AGEMA_signal_4734), .Q (new_AGEMA_signal_4735) ) ;
    buf_clk new_AGEMA_reg_buffer_1271 ( .C (clk), .D (new_AGEMA_signal_4736), .Q (new_AGEMA_signal_4737) ) ;
    buf_clk new_AGEMA_reg_buffer_1273 ( .C (clk), .D (new_AGEMA_signal_4738), .Q (new_AGEMA_signal_4739) ) ;
    buf_clk new_AGEMA_reg_buffer_1275 ( .C (clk), .D (new_AGEMA_signal_4740), .Q (new_AGEMA_signal_4741) ) ;
    buf_clk new_AGEMA_reg_buffer_1277 ( .C (clk), .D (new_AGEMA_signal_4742), .Q (new_AGEMA_signal_4743) ) ;
    buf_clk new_AGEMA_reg_buffer_1279 ( .C (clk), .D (new_AGEMA_signal_4744), .Q (new_AGEMA_signal_4745) ) ;
    buf_clk new_AGEMA_reg_buffer_1281 ( .C (clk), .D (new_AGEMA_signal_4746), .Q (new_AGEMA_signal_4747) ) ;
    buf_clk new_AGEMA_reg_buffer_1283 ( .C (clk), .D (new_AGEMA_signal_4748), .Q (new_AGEMA_signal_4749) ) ;
    buf_clk new_AGEMA_reg_buffer_1285 ( .C (clk), .D (new_AGEMA_signal_4750), .Q (new_AGEMA_signal_4751) ) ;
    buf_clk new_AGEMA_reg_buffer_1287 ( .C (clk), .D (new_AGEMA_signal_4752), .Q (new_AGEMA_signal_4753) ) ;
    buf_clk new_AGEMA_reg_buffer_1289 ( .C (clk), .D (new_AGEMA_signal_4754), .Q (new_AGEMA_signal_4755) ) ;
    buf_clk new_AGEMA_reg_buffer_1291 ( .C (clk), .D (new_AGEMA_signal_4756), .Q (new_AGEMA_signal_4757) ) ;
    buf_clk new_AGEMA_reg_buffer_1293 ( .C (clk), .D (new_AGEMA_signal_4758), .Q (new_AGEMA_signal_4759) ) ;
    buf_clk new_AGEMA_reg_buffer_1295 ( .C (clk), .D (new_AGEMA_signal_4760), .Q (new_AGEMA_signal_4761) ) ;
    buf_clk new_AGEMA_reg_buffer_1297 ( .C (clk), .D (new_AGEMA_signal_4762), .Q (new_AGEMA_signal_4763) ) ;
    buf_clk new_AGEMA_reg_buffer_1299 ( .C (clk), .D (new_AGEMA_signal_4764), .Q (new_AGEMA_signal_4765) ) ;
    buf_clk new_AGEMA_reg_buffer_1301 ( .C (clk), .D (new_AGEMA_signal_4766), .Q (new_AGEMA_signal_4767) ) ;
    buf_clk new_AGEMA_reg_buffer_1303 ( .C (clk), .D (new_AGEMA_signal_4768), .Q (new_AGEMA_signal_4769) ) ;
    buf_clk new_AGEMA_reg_buffer_1305 ( .C (clk), .D (new_AGEMA_signal_4770), .Q (new_AGEMA_signal_4771) ) ;
    buf_clk new_AGEMA_reg_buffer_1307 ( .C (clk), .D (new_AGEMA_signal_4772), .Q (new_AGEMA_signal_4773) ) ;
    buf_clk new_AGEMA_reg_buffer_1309 ( .C (clk), .D (new_AGEMA_signal_4774), .Q (new_AGEMA_signal_4775) ) ;
    buf_clk new_AGEMA_reg_buffer_1311 ( .C (clk), .D (new_AGEMA_signal_4776), .Q (new_AGEMA_signal_4777) ) ;
    buf_clk new_AGEMA_reg_buffer_1313 ( .C (clk), .D (new_AGEMA_signal_4778), .Q (new_AGEMA_signal_4779) ) ;
    buf_clk new_AGEMA_reg_buffer_1315 ( .C (clk), .D (new_AGEMA_signal_4780), .Q (new_AGEMA_signal_4781) ) ;
    buf_clk new_AGEMA_reg_buffer_1317 ( .C (clk), .D (new_AGEMA_signal_4782), .Q (new_AGEMA_signal_4783) ) ;
    buf_clk new_AGEMA_reg_buffer_1325 ( .C (clk), .D (new_AGEMA_signal_4790), .Q (new_AGEMA_signal_4791) ) ;
    buf_clk new_AGEMA_reg_buffer_1327 ( .C (clk), .D (new_AGEMA_signal_4792), .Q (new_AGEMA_signal_4793) ) ;
    buf_clk new_AGEMA_reg_buffer_1329 ( .C (clk), .D (new_AGEMA_signal_4794), .Q (new_AGEMA_signal_4795) ) ;
    buf_clk new_AGEMA_reg_buffer_1331 ( .C (clk), .D (new_AGEMA_signal_4796), .Q (new_AGEMA_signal_4797) ) ;
    buf_clk new_AGEMA_reg_buffer_1333 ( .C (clk), .D (new_AGEMA_signal_4798), .Q (new_AGEMA_signal_4799) ) ;
    buf_clk new_AGEMA_reg_buffer_1335 ( .C (clk), .D (new_AGEMA_signal_4800), .Q (new_AGEMA_signal_4801) ) ;
    buf_clk new_AGEMA_reg_buffer_1337 ( .C (clk), .D (new_AGEMA_signal_4802), .Q (new_AGEMA_signal_4803) ) ;
    buf_clk new_AGEMA_reg_buffer_1339 ( .C (clk), .D (new_AGEMA_signal_4804), .Q (new_AGEMA_signal_4805) ) ;
    buf_clk new_AGEMA_reg_buffer_1341 ( .C (clk), .D (new_AGEMA_signal_4806), .Q (new_AGEMA_signal_4807) ) ;
    buf_clk new_AGEMA_reg_buffer_1343 ( .C (clk), .D (new_AGEMA_signal_4808), .Q (new_AGEMA_signal_4809) ) ;
    buf_clk new_AGEMA_reg_buffer_1345 ( .C (clk), .D (new_AGEMA_signal_4810), .Q (new_AGEMA_signal_4811) ) ;
    buf_clk new_AGEMA_reg_buffer_1347 ( .C (clk), .D (new_AGEMA_signal_4812), .Q (new_AGEMA_signal_4813) ) ;
    buf_clk new_AGEMA_reg_buffer_1349 ( .C (clk), .D (new_AGEMA_signal_4814), .Q (new_AGEMA_signal_4815) ) ;
    buf_clk new_AGEMA_reg_buffer_1351 ( .C (clk), .D (new_AGEMA_signal_4816), .Q (new_AGEMA_signal_4817) ) ;
    buf_clk new_AGEMA_reg_buffer_1353 ( .C (clk), .D (new_AGEMA_signal_4818), .Q (new_AGEMA_signal_4819) ) ;
    buf_clk new_AGEMA_reg_buffer_1355 ( .C (clk), .D (new_AGEMA_signal_4820), .Q (new_AGEMA_signal_4821) ) ;
    buf_clk new_AGEMA_reg_buffer_1357 ( .C (clk), .D (new_AGEMA_signal_4822), .Q (new_AGEMA_signal_4823) ) ;
    buf_clk new_AGEMA_reg_buffer_1359 ( .C (clk), .D (new_AGEMA_signal_4824), .Q (new_AGEMA_signal_4825) ) ;
    buf_clk new_AGEMA_reg_buffer_1361 ( .C (clk), .D (new_AGEMA_signal_4826), .Q (new_AGEMA_signal_4827) ) ;
    buf_clk new_AGEMA_reg_buffer_1363 ( .C (clk), .D (new_AGEMA_signal_4828), .Q (new_AGEMA_signal_4829) ) ;
    buf_clk new_AGEMA_reg_buffer_1365 ( .C (clk), .D (new_AGEMA_signal_4830), .Q (new_AGEMA_signal_4831) ) ;
    buf_clk new_AGEMA_reg_buffer_1367 ( .C (clk), .D (new_AGEMA_signal_4832), .Q (new_AGEMA_signal_4833) ) ;
    buf_clk new_AGEMA_reg_buffer_1369 ( .C (clk), .D (new_AGEMA_signal_4834), .Q (new_AGEMA_signal_4835) ) ;
    buf_clk new_AGEMA_reg_buffer_1371 ( .C (clk), .D (new_AGEMA_signal_4836), .Q (new_AGEMA_signal_4837) ) ;
    buf_clk new_AGEMA_reg_buffer_1373 ( .C (clk), .D (new_AGEMA_signal_4838), .Q (new_AGEMA_signal_4839) ) ;
    buf_clk new_AGEMA_reg_buffer_1375 ( .C (clk), .D (new_AGEMA_signal_4840), .Q (new_AGEMA_signal_4841) ) ;
    buf_clk new_AGEMA_reg_buffer_1377 ( .C (clk), .D (new_AGEMA_signal_4842), .Q (new_AGEMA_signal_4843) ) ;
    buf_clk new_AGEMA_reg_buffer_1379 ( .C (clk), .D (new_AGEMA_signal_4844), .Q (new_AGEMA_signal_4845) ) ;
    buf_clk new_AGEMA_reg_buffer_1381 ( .C (clk), .D (new_AGEMA_signal_4846), .Q (new_AGEMA_signal_4847) ) ;
    buf_clk new_AGEMA_reg_buffer_1383 ( .C (clk), .D (new_AGEMA_signal_4848), .Q (new_AGEMA_signal_4849) ) ;
    buf_clk new_AGEMA_reg_buffer_1385 ( .C (clk), .D (new_AGEMA_signal_4850), .Q (new_AGEMA_signal_4851) ) ;
    buf_clk new_AGEMA_reg_buffer_1387 ( .C (clk), .D (new_AGEMA_signal_4852), .Q (new_AGEMA_signal_4853) ) ;
    buf_clk new_AGEMA_reg_buffer_1389 ( .C (clk), .D (new_AGEMA_signal_4854), .Q (new_AGEMA_signal_4855) ) ;
    buf_clk new_AGEMA_reg_buffer_1391 ( .C (clk), .D (new_AGEMA_signal_4856), .Q (new_AGEMA_signal_4857) ) ;
    buf_clk new_AGEMA_reg_buffer_1393 ( .C (clk), .D (new_AGEMA_signal_4858), .Q (new_AGEMA_signal_4859) ) ;
    buf_clk new_AGEMA_reg_buffer_1395 ( .C (clk), .D (new_AGEMA_signal_4860), .Q (new_AGEMA_signal_4861) ) ;
    buf_clk new_AGEMA_reg_buffer_1397 ( .C (clk), .D (new_AGEMA_signal_4862), .Q (new_AGEMA_signal_4863) ) ;
    buf_clk new_AGEMA_reg_buffer_1399 ( .C (clk), .D (new_AGEMA_signal_4864), .Q (new_AGEMA_signal_4865) ) ;
    buf_clk new_AGEMA_reg_buffer_1401 ( .C (clk), .D (new_AGEMA_signal_4866), .Q (new_AGEMA_signal_4867) ) ;
    buf_clk new_AGEMA_reg_buffer_1403 ( .C (clk), .D (new_AGEMA_signal_4868), .Q (new_AGEMA_signal_4869) ) ;
    buf_clk new_AGEMA_reg_buffer_1405 ( .C (clk), .D (new_AGEMA_signal_4870), .Q (new_AGEMA_signal_4871) ) ;
    buf_clk new_AGEMA_reg_buffer_1407 ( .C (clk), .D (new_AGEMA_signal_4872), .Q (new_AGEMA_signal_4873) ) ;
    buf_clk new_AGEMA_reg_buffer_1409 ( .C (clk), .D (new_AGEMA_signal_4874), .Q (new_AGEMA_signal_4875) ) ;
    buf_clk new_AGEMA_reg_buffer_1411 ( .C (clk), .D (new_AGEMA_signal_4876), .Q (new_AGEMA_signal_4877) ) ;
    buf_clk new_AGEMA_reg_buffer_1413 ( .C (clk), .D (new_AGEMA_signal_4878), .Q (new_AGEMA_signal_4879) ) ;
    buf_clk new_AGEMA_reg_buffer_1415 ( .C (clk), .D (new_AGEMA_signal_4880), .Q (new_AGEMA_signal_4881) ) ;
    buf_clk new_AGEMA_reg_buffer_1417 ( .C (clk), .D (new_AGEMA_signal_4882), .Q (new_AGEMA_signal_4883) ) ;
    buf_clk new_AGEMA_reg_buffer_1419 ( .C (clk), .D (new_AGEMA_signal_4884), .Q (new_AGEMA_signal_4885) ) ;
    buf_clk new_AGEMA_reg_buffer_1421 ( .C (clk), .D (new_AGEMA_signal_4886), .Q (new_AGEMA_signal_4887) ) ;
    buf_clk new_AGEMA_reg_buffer_1423 ( .C (clk), .D (new_AGEMA_signal_4888), .Q (new_AGEMA_signal_4889) ) ;
    buf_clk new_AGEMA_reg_buffer_1425 ( .C (clk), .D (new_AGEMA_signal_4890), .Q (new_AGEMA_signal_4891) ) ;
    buf_clk new_AGEMA_reg_buffer_1427 ( .C (clk), .D (new_AGEMA_signal_4892), .Q (new_AGEMA_signal_4893) ) ;
    buf_clk new_AGEMA_reg_buffer_1429 ( .C (clk), .D (new_AGEMA_signal_4894), .Q (new_AGEMA_signal_4895) ) ;
    buf_clk new_AGEMA_reg_buffer_1431 ( .C (clk), .D (new_AGEMA_signal_4896), .Q (new_AGEMA_signal_4897) ) ;
    buf_clk new_AGEMA_reg_buffer_1433 ( .C (clk), .D (new_AGEMA_signal_4898), .Q (new_AGEMA_signal_4899) ) ;
    buf_clk new_AGEMA_reg_buffer_1435 ( .C (clk), .D (new_AGEMA_signal_4900), .Q (new_AGEMA_signal_4901) ) ;
    buf_clk new_AGEMA_reg_buffer_1437 ( .C (clk), .D (new_AGEMA_signal_4902), .Q (new_AGEMA_signal_4903) ) ;
    buf_clk new_AGEMA_reg_buffer_1439 ( .C (clk), .D (new_AGEMA_signal_4904), .Q (new_AGEMA_signal_4905) ) ;
    buf_clk new_AGEMA_reg_buffer_1441 ( .C (clk), .D (new_AGEMA_signal_4906), .Q (new_AGEMA_signal_4907) ) ;
    buf_clk new_AGEMA_reg_buffer_1443 ( .C (clk), .D (new_AGEMA_signal_4908), .Q (new_AGEMA_signal_4909) ) ;
    buf_clk new_AGEMA_reg_buffer_1445 ( .C (clk), .D (new_AGEMA_signal_4910), .Q (new_AGEMA_signal_4911) ) ;
    buf_clk new_AGEMA_reg_buffer_1447 ( .C (clk), .D (new_AGEMA_signal_4912), .Q (new_AGEMA_signal_4913) ) ;
    buf_clk new_AGEMA_reg_buffer_1449 ( .C (clk), .D (new_AGEMA_signal_4914), .Q (new_AGEMA_signal_4915) ) ;
    buf_clk new_AGEMA_reg_buffer_1451 ( .C (clk), .D (new_AGEMA_signal_4916), .Q (new_AGEMA_signal_4917) ) ;
    buf_clk new_AGEMA_reg_buffer_1453 ( .C (clk), .D (new_AGEMA_signal_4918), .Q (new_AGEMA_signal_4919) ) ;
    buf_clk new_AGEMA_reg_buffer_3873 ( .C (clk), .D (new_AGEMA_signal_7337), .Q (new_AGEMA_signal_7338) ) ;
    buf_clk new_AGEMA_reg_buffer_3881 ( .C (clk), .D (new_AGEMA_signal_7345), .Q (new_AGEMA_signal_7346) ) ;
    buf_clk new_AGEMA_reg_buffer_3889 ( .C (clk), .D (new_AGEMA_signal_7353), .Q (new_AGEMA_signal_7354) ) ;
    buf_clk new_AGEMA_reg_buffer_3897 ( .C (clk), .D (new_AGEMA_signal_7361), .Q (new_AGEMA_signal_7362) ) ;
    buf_clk new_AGEMA_reg_buffer_3905 ( .C (clk), .D (new_AGEMA_signal_7369), .Q (new_AGEMA_signal_7370) ) ;
    buf_clk new_AGEMA_reg_buffer_3913 ( .C (clk), .D (new_AGEMA_signal_7377), .Q (new_AGEMA_signal_7378) ) ;
    buf_clk new_AGEMA_reg_buffer_3921 ( .C (clk), .D (new_AGEMA_signal_7385), .Q (new_AGEMA_signal_7386) ) ;
    buf_clk new_AGEMA_reg_buffer_3929 ( .C (clk), .D (new_AGEMA_signal_7393), .Q (new_AGEMA_signal_7394) ) ;
    buf_clk new_AGEMA_reg_buffer_3937 ( .C (clk), .D (new_AGEMA_signal_7401), .Q (new_AGEMA_signal_7402) ) ;
    buf_clk new_AGEMA_reg_buffer_3945 ( .C (clk), .D (new_AGEMA_signal_7409), .Q (new_AGEMA_signal_7410) ) ;
    buf_clk new_AGEMA_reg_buffer_3953 ( .C (clk), .D (new_AGEMA_signal_7417), .Q (new_AGEMA_signal_7418) ) ;
    buf_clk new_AGEMA_reg_buffer_3961 ( .C (clk), .D (new_AGEMA_signal_7425), .Q (new_AGEMA_signal_7426) ) ;
    buf_clk new_AGEMA_reg_buffer_3969 ( .C (clk), .D (new_AGEMA_signal_7433), .Q (new_AGEMA_signal_7434) ) ;
    buf_clk new_AGEMA_reg_buffer_3977 ( .C (clk), .D (new_AGEMA_signal_7441), .Q (new_AGEMA_signal_7442) ) ;
    buf_clk new_AGEMA_reg_buffer_3985 ( .C (clk), .D (new_AGEMA_signal_7449), .Q (new_AGEMA_signal_7450) ) ;
    buf_clk new_AGEMA_reg_buffer_3993 ( .C (clk), .D (new_AGEMA_signal_7457), .Q (new_AGEMA_signal_7458) ) ;
    buf_clk new_AGEMA_reg_buffer_4001 ( .C (clk), .D (new_AGEMA_signal_7465), .Q (new_AGEMA_signal_7466) ) ;
    buf_clk new_AGEMA_reg_buffer_4009 ( .C (clk), .D (new_AGEMA_signal_7473), .Q (new_AGEMA_signal_7474) ) ;
    buf_clk new_AGEMA_reg_buffer_4017 ( .C (clk), .D (new_AGEMA_signal_7481), .Q (new_AGEMA_signal_7482) ) ;
    buf_clk new_AGEMA_reg_buffer_4025 ( .C (clk), .D (new_AGEMA_signal_7489), .Q (new_AGEMA_signal_7490) ) ;
    buf_clk new_AGEMA_reg_buffer_4033 ( .C (clk), .D (new_AGEMA_signal_7497), .Q (new_AGEMA_signal_7498) ) ;
    buf_clk new_AGEMA_reg_buffer_4041 ( .C (clk), .D (new_AGEMA_signal_7505), .Q (new_AGEMA_signal_7506) ) ;
    buf_clk new_AGEMA_reg_buffer_4049 ( .C (clk), .D (new_AGEMA_signal_7513), .Q (new_AGEMA_signal_7514) ) ;
    buf_clk new_AGEMA_reg_buffer_4057 ( .C (clk), .D (new_AGEMA_signal_7521), .Q (new_AGEMA_signal_7522) ) ;
    buf_clk new_AGEMA_reg_buffer_4065 ( .C (clk), .D (new_AGEMA_signal_7529), .Q (new_AGEMA_signal_7530) ) ;
    buf_clk new_AGEMA_reg_buffer_4073 ( .C (clk), .D (new_AGEMA_signal_7537), .Q (new_AGEMA_signal_7538) ) ;
    buf_clk new_AGEMA_reg_buffer_4081 ( .C (clk), .D (new_AGEMA_signal_7545), .Q (new_AGEMA_signal_7546) ) ;
    buf_clk new_AGEMA_reg_buffer_4089 ( .C (clk), .D (new_AGEMA_signal_7553), .Q (new_AGEMA_signal_7554) ) ;
    buf_clk new_AGEMA_reg_buffer_4097 ( .C (clk), .D (new_AGEMA_signal_7561), .Q (new_AGEMA_signal_7562) ) ;
    buf_clk new_AGEMA_reg_buffer_4105 ( .C (clk), .D (new_AGEMA_signal_7569), .Q (new_AGEMA_signal_7570) ) ;
    buf_clk new_AGEMA_reg_buffer_4113 ( .C (clk), .D (new_AGEMA_signal_7577), .Q (new_AGEMA_signal_7578) ) ;
    buf_clk new_AGEMA_reg_buffer_4121 ( .C (clk), .D (new_AGEMA_signal_7585), .Q (new_AGEMA_signal_7586) ) ;
    buf_clk new_AGEMA_reg_buffer_4129 ( .C (clk), .D (new_AGEMA_signal_7593), .Q (new_AGEMA_signal_7594) ) ;
    buf_clk new_AGEMA_reg_buffer_4137 ( .C (clk), .D (new_AGEMA_signal_7601), .Q (new_AGEMA_signal_7602) ) ;
    buf_clk new_AGEMA_reg_buffer_4145 ( .C (clk), .D (new_AGEMA_signal_7609), .Q (new_AGEMA_signal_7610) ) ;
    buf_clk new_AGEMA_reg_buffer_4153 ( .C (clk), .D (new_AGEMA_signal_7617), .Q (new_AGEMA_signal_7618) ) ;
    buf_clk new_AGEMA_reg_buffer_4161 ( .C (clk), .D (new_AGEMA_signal_7625), .Q (new_AGEMA_signal_7626) ) ;
    buf_clk new_AGEMA_reg_buffer_4169 ( .C (clk), .D (new_AGEMA_signal_7633), .Q (new_AGEMA_signal_7634) ) ;
    buf_clk new_AGEMA_reg_buffer_4177 ( .C (clk), .D (new_AGEMA_signal_7641), .Q (new_AGEMA_signal_7642) ) ;
    buf_clk new_AGEMA_reg_buffer_4185 ( .C (clk), .D (new_AGEMA_signal_7649), .Q (new_AGEMA_signal_7650) ) ;
    buf_clk new_AGEMA_reg_buffer_4193 ( .C (clk), .D (new_AGEMA_signal_7657), .Q (new_AGEMA_signal_7658) ) ;
    buf_clk new_AGEMA_reg_buffer_4201 ( .C (clk), .D (new_AGEMA_signal_7665), .Q (new_AGEMA_signal_7666) ) ;
    buf_clk new_AGEMA_reg_buffer_4209 ( .C (clk), .D (new_AGEMA_signal_7673), .Q (new_AGEMA_signal_7674) ) ;
    buf_clk new_AGEMA_reg_buffer_4217 ( .C (clk), .D (new_AGEMA_signal_7681), .Q (new_AGEMA_signal_7682) ) ;
    buf_clk new_AGEMA_reg_buffer_4225 ( .C (clk), .D (new_AGEMA_signal_7689), .Q (new_AGEMA_signal_7690) ) ;
    buf_clk new_AGEMA_reg_buffer_4233 ( .C (clk), .D (new_AGEMA_signal_7697), .Q (new_AGEMA_signal_7698) ) ;
    buf_clk new_AGEMA_reg_buffer_4241 ( .C (clk), .D (new_AGEMA_signal_7705), .Q (new_AGEMA_signal_7706) ) ;
    buf_clk new_AGEMA_reg_buffer_4249 ( .C (clk), .D (new_AGEMA_signal_7713), .Q (new_AGEMA_signal_7714) ) ;
    buf_clk new_AGEMA_reg_buffer_4257 ( .C (clk), .D (new_AGEMA_signal_7721), .Q (new_AGEMA_signal_7722) ) ;
    buf_clk new_AGEMA_reg_buffer_4265 ( .C (clk), .D (new_AGEMA_signal_7729), .Q (new_AGEMA_signal_7730) ) ;
    buf_clk new_AGEMA_reg_buffer_4273 ( .C (clk), .D (new_AGEMA_signal_7737), .Q (new_AGEMA_signal_7738) ) ;
    buf_clk new_AGEMA_reg_buffer_4281 ( .C (clk), .D (new_AGEMA_signal_7745), .Q (new_AGEMA_signal_7746) ) ;
    buf_clk new_AGEMA_reg_buffer_4289 ( .C (clk), .D (new_AGEMA_signal_7753), .Q (new_AGEMA_signal_7754) ) ;
    buf_clk new_AGEMA_reg_buffer_4297 ( .C (clk), .D (new_AGEMA_signal_7761), .Q (new_AGEMA_signal_7762) ) ;
    buf_clk new_AGEMA_reg_buffer_4305 ( .C (clk), .D (new_AGEMA_signal_7769), .Q (new_AGEMA_signal_7770) ) ;
    buf_clk new_AGEMA_reg_buffer_4313 ( .C (clk), .D (new_AGEMA_signal_7777), .Q (new_AGEMA_signal_7778) ) ;
    buf_clk new_AGEMA_reg_buffer_4321 ( .C (clk), .D (new_AGEMA_signal_7785), .Q (new_AGEMA_signal_7786) ) ;
    buf_clk new_AGEMA_reg_buffer_4329 ( .C (clk), .D (new_AGEMA_signal_7793), .Q (new_AGEMA_signal_7794) ) ;
    buf_clk new_AGEMA_reg_buffer_4337 ( .C (clk), .D (new_AGEMA_signal_7801), .Q (new_AGEMA_signal_7802) ) ;
    buf_clk new_AGEMA_reg_buffer_4345 ( .C (clk), .D (new_AGEMA_signal_7809), .Q (new_AGEMA_signal_7810) ) ;
    buf_clk new_AGEMA_reg_buffer_4353 ( .C (clk), .D (new_AGEMA_signal_7817), .Q (new_AGEMA_signal_7818) ) ;
    buf_clk new_AGEMA_reg_buffer_4361 ( .C (clk), .D (new_AGEMA_signal_7825), .Q (new_AGEMA_signal_7826) ) ;
    buf_clk new_AGEMA_reg_buffer_4369 ( .C (clk), .D (new_AGEMA_signal_7833), .Q (new_AGEMA_signal_7834) ) ;
    buf_clk new_AGEMA_reg_buffer_4377 ( .C (clk), .D (new_AGEMA_signal_7841), .Q (new_AGEMA_signal_7842) ) ;
    buf_clk new_AGEMA_reg_buffer_4385 ( .C (clk), .D (new_AGEMA_signal_7849), .Q (new_AGEMA_signal_7850) ) ;
    buf_clk new_AGEMA_reg_buffer_4393 ( .C (clk), .D (new_AGEMA_signal_7857), .Q (new_AGEMA_signal_7858) ) ;
    buf_clk new_AGEMA_reg_buffer_4401 ( .C (clk), .D (new_AGEMA_signal_7865), .Q (new_AGEMA_signal_7866) ) ;
    buf_clk new_AGEMA_reg_buffer_4409 ( .C (clk), .D (new_AGEMA_signal_7873), .Q (new_AGEMA_signal_7874) ) ;
    buf_clk new_AGEMA_reg_buffer_4417 ( .C (clk), .D (new_AGEMA_signal_7881), .Q (new_AGEMA_signal_7882) ) ;
    buf_clk new_AGEMA_reg_buffer_4425 ( .C (clk), .D (new_AGEMA_signal_7889), .Q (new_AGEMA_signal_7890) ) ;
    buf_clk new_AGEMA_reg_buffer_4433 ( .C (clk), .D (new_AGEMA_signal_7897), .Q (new_AGEMA_signal_7898) ) ;
    buf_clk new_AGEMA_reg_buffer_4441 ( .C (clk), .D (new_AGEMA_signal_7905), .Q (new_AGEMA_signal_7906) ) ;
    buf_clk new_AGEMA_reg_buffer_4449 ( .C (clk), .D (new_AGEMA_signal_7913), .Q (new_AGEMA_signal_7914) ) ;
    buf_clk new_AGEMA_reg_buffer_4457 ( .C (clk), .D (new_AGEMA_signal_7921), .Q (new_AGEMA_signal_7922) ) ;
    buf_clk new_AGEMA_reg_buffer_4465 ( .C (clk), .D (new_AGEMA_signal_7929), .Q (new_AGEMA_signal_7930) ) ;
    buf_clk new_AGEMA_reg_buffer_4473 ( .C (clk), .D (new_AGEMA_signal_7937), .Q (new_AGEMA_signal_7938) ) ;
    buf_clk new_AGEMA_reg_buffer_4481 ( .C (clk), .D (new_AGEMA_signal_7945), .Q (new_AGEMA_signal_7946) ) ;
    buf_clk new_AGEMA_reg_buffer_4489 ( .C (clk), .D (new_AGEMA_signal_7953), .Q (new_AGEMA_signal_7954) ) ;
    buf_clk new_AGEMA_reg_buffer_4497 ( .C (clk), .D (new_AGEMA_signal_7961), .Q (new_AGEMA_signal_7962) ) ;
    buf_clk new_AGEMA_reg_buffer_4505 ( .C (clk), .D (new_AGEMA_signal_7969), .Q (new_AGEMA_signal_7970) ) ;
    buf_clk new_AGEMA_reg_buffer_4513 ( .C (clk), .D (new_AGEMA_signal_7977), .Q (new_AGEMA_signal_7978) ) ;
    buf_clk new_AGEMA_reg_buffer_4521 ( .C (clk), .D (new_AGEMA_signal_7985), .Q (new_AGEMA_signal_7986) ) ;
    buf_clk new_AGEMA_reg_buffer_4529 ( .C (clk), .D (new_AGEMA_signal_7993), .Q (new_AGEMA_signal_7994) ) ;
    buf_clk new_AGEMA_reg_buffer_4537 ( .C (clk), .D (new_AGEMA_signal_8001), .Q (new_AGEMA_signal_8002) ) ;
    buf_clk new_AGEMA_reg_buffer_4545 ( .C (clk), .D (new_AGEMA_signal_8009), .Q (new_AGEMA_signal_8010) ) ;
    buf_clk new_AGEMA_reg_buffer_4553 ( .C (clk), .D (new_AGEMA_signal_8017), .Q (new_AGEMA_signal_8018) ) ;
    buf_clk new_AGEMA_reg_buffer_4561 ( .C (clk), .D (new_AGEMA_signal_8025), .Q (new_AGEMA_signal_8026) ) ;
    buf_clk new_AGEMA_reg_buffer_4569 ( .C (clk), .D (new_AGEMA_signal_8033), .Q (new_AGEMA_signal_8034) ) ;
    buf_clk new_AGEMA_reg_buffer_4577 ( .C (clk), .D (new_AGEMA_signal_8041), .Q (new_AGEMA_signal_8042) ) ;
    buf_clk new_AGEMA_reg_buffer_4585 ( .C (clk), .D (new_AGEMA_signal_8049), .Q (new_AGEMA_signal_8050) ) ;
    buf_clk new_AGEMA_reg_buffer_4593 ( .C (clk), .D (new_AGEMA_signal_8057), .Q (new_AGEMA_signal_8058) ) ;
    buf_clk new_AGEMA_reg_buffer_4601 ( .C (clk), .D (new_AGEMA_signal_8065), .Q (new_AGEMA_signal_8066) ) ;
    buf_clk new_AGEMA_reg_buffer_4609 ( .C (clk), .D (new_AGEMA_signal_8073), .Q (new_AGEMA_signal_8074) ) ;
    buf_clk new_AGEMA_reg_buffer_4617 ( .C (clk), .D (new_AGEMA_signal_8081), .Q (new_AGEMA_signal_8082) ) ;
    buf_clk new_AGEMA_reg_buffer_4625 ( .C (clk), .D (new_AGEMA_signal_8089), .Q (new_AGEMA_signal_8090) ) ;
    buf_clk new_AGEMA_reg_buffer_4633 ( .C (clk), .D (new_AGEMA_signal_8097), .Q (new_AGEMA_signal_8098) ) ;
    buf_clk new_AGEMA_reg_buffer_4641 ( .C (clk), .D (new_AGEMA_signal_8105), .Q (new_AGEMA_signal_8106) ) ;
    buf_clk new_AGEMA_reg_buffer_4649 ( .C (clk), .D (new_AGEMA_signal_8113), .Q (new_AGEMA_signal_8114) ) ;
    buf_clk new_AGEMA_reg_buffer_4657 ( .C (clk), .D (new_AGEMA_signal_8121), .Q (new_AGEMA_signal_8122) ) ;
    buf_clk new_AGEMA_reg_buffer_4665 ( .C (clk), .D (new_AGEMA_signal_8129), .Q (new_AGEMA_signal_8130) ) ;
    buf_clk new_AGEMA_reg_buffer_4673 ( .C (clk), .D (new_AGEMA_signal_8137), .Q (new_AGEMA_signal_8138) ) ;
    buf_clk new_AGEMA_reg_buffer_4681 ( .C (clk), .D (new_AGEMA_signal_8145), .Q (new_AGEMA_signal_8146) ) ;
    buf_clk new_AGEMA_reg_buffer_4689 ( .C (clk), .D (new_AGEMA_signal_8153), .Q (new_AGEMA_signal_8154) ) ;
    buf_clk new_AGEMA_reg_buffer_4697 ( .C (clk), .D (new_AGEMA_signal_8161), .Q (new_AGEMA_signal_8162) ) ;
    buf_clk new_AGEMA_reg_buffer_4705 ( .C (clk), .D (new_AGEMA_signal_8169), .Q (new_AGEMA_signal_8170) ) ;
    buf_clk new_AGEMA_reg_buffer_4713 ( .C (clk), .D (new_AGEMA_signal_8177), .Q (new_AGEMA_signal_8178) ) ;
    buf_clk new_AGEMA_reg_buffer_4721 ( .C (clk), .D (new_AGEMA_signal_8185), .Q (new_AGEMA_signal_8186) ) ;
    buf_clk new_AGEMA_reg_buffer_4729 ( .C (clk), .D (new_AGEMA_signal_8193), .Q (new_AGEMA_signal_8194) ) ;
    buf_clk new_AGEMA_reg_buffer_4737 ( .C (clk), .D (new_AGEMA_signal_8201), .Q (new_AGEMA_signal_8202) ) ;
    buf_clk new_AGEMA_reg_buffer_4745 ( .C (clk), .D (new_AGEMA_signal_8209), .Q (new_AGEMA_signal_8210) ) ;
    buf_clk new_AGEMA_reg_buffer_4753 ( .C (clk), .D (new_AGEMA_signal_8217), .Q (new_AGEMA_signal_8218) ) ;
    buf_clk new_AGEMA_reg_buffer_4761 ( .C (clk), .D (new_AGEMA_signal_8225), .Q (new_AGEMA_signal_8226) ) ;
    buf_clk new_AGEMA_reg_buffer_4769 ( .C (clk), .D (new_AGEMA_signal_8233), .Q (new_AGEMA_signal_8234) ) ;
    buf_clk new_AGEMA_reg_buffer_4777 ( .C (clk), .D (new_AGEMA_signal_8241), .Q (new_AGEMA_signal_8242) ) ;
    buf_clk new_AGEMA_reg_buffer_4785 ( .C (clk), .D (new_AGEMA_signal_8249), .Q (new_AGEMA_signal_8250) ) ;
    buf_clk new_AGEMA_reg_buffer_4793 ( .C (clk), .D (new_AGEMA_signal_8257), .Q (new_AGEMA_signal_8258) ) ;
    buf_clk new_AGEMA_reg_buffer_4801 ( .C (clk), .D (new_AGEMA_signal_8265), .Q (new_AGEMA_signal_8266) ) ;
    buf_clk new_AGEMA_reg_buffer_4809 ( .C (clk), .D (new_AGEMA_signal_8273), .Q (new_AGEMA_signal_8274) ) ;
    buf_clk new_AGEMA_reg_buffer_4817 ( .C (clk), .D (new_AGEMA_signal_8281), .Q (new_AGEMA_signal_8282) ) ;
    buf_clk new_AGEMA_reg_buffer_4825 ( .C (clk), .D (new_AGEMA_signal_8289), .Q (new_AGEMA_signal_8290) ) ;
    buf_clk new_AGEMA_reg_buffer_4833 ( .C (clk), .D (new_AGEMA_signal_8297), .Q (new_AGEMA_signal_8298) ) ;
    buf_clk new_AGEMA_reg_buffer_4841 ( .C (clk), .D (new_AGEMA_signal_8305), .Q (new_AGEMA_signal_8306) ) ;
    buf_clk new_AGEMA_reg_buffer_4849 ( .C (clk), .D (new_AGEMA_signal_8313), .Q (new_AGEMA_signal_8314) ) ;
    buf_clk new_AGEMA_reg_buffer_4857 ( .C (clk), .D (new_AGEMA_signal_8321), .Q (new_AGEMA_signal_8322) ) ;
    buf_clk new_AGEMA_reg_buffer_4865 ( .C (clk), .D (new_AGEMA_signal_8329), .Q (new_AGEMA_signal_8330) ) ;
    buf_clk new_AGEMA_reg_buffer_4873 ( .C (clk), .D (new_AGEMA_signal_8337), .Q (new_AGEMA_signal_8338) ) ;
    buf_clk new_AGEMA_reg_buffer_4881 ( .C (clk), .D (new_AGEMA_signal_8345), .Q (new_AGEMA_signal_8346) ) ;
    buf_clk new_AGEMA_reg_buffer_4889 ( .C (clk), .D (new_AGEMA_signal_8353), .Q (new_AGEMA_signal_8354) ) ;
    buf_clk new_AGEMA_reg_buffer_4897 ( .C (clk), .D (new_AGEMA_signal_8361), .Q (new_AGEMA_signal_8362) ) ;
    buf_clk new_AGEMA_reg_buffer_4905 ( .C (clk), .D (new_AGEMA_signal_8369), .Q (new_AGEMA_signal_8370) ) ;
    buf_clk new_AGEMA_reg_buffer_4913 ( .C (clk), .D (new_AGEMA_signal_8377), .Q (new_AGEMA_signal_8378) ) ;
    buf_clk new_AGEMA_reg_buffer_4921 ( .C (clk), .D (new_AGEMA_signal_8385), .Q (new_AGEMA_signal_8386) ) ;
    buf_clk new_AGEMA_reg_buffer_4929 ( .C (clk), .D (new_AGEMA_signal_8393), .Q (new_AGEMA_signal_8394) ) ;
    buf_clk new_AGEMA_reg_buffer_4937 ( .C (clk), .D (new_AGEMA_signal_8401), .Q (new_AGEMA_signal_8402) ) ;
    buf_clk new_AGEMA_reg_buffer_4945 ( .C (clk), .D (new_AGEMA_signal_8409), .Q (new_AGEMA_signal_8410) ) ;
    buf_clk new_AGEMA_reg_buffer_4953 ( .C (clk), .D (new_AGEMA_signal_8417), .Q (new_AGEMA_signal_8418) ) ;
    buf_clk new_AGEMA_reg_buffer_4961 ( .C (clk), .D (new_AGEMA_signal_8425), .Q (new_AGEMA_signal_8426) ) ;
    buf_clk new_AGEMA_reg_buffer_4969 ( .C (clk), .D (new_AGEMA_signal_8433), .Q (new_AGEMA_signal_8434) ) ;
    buf_clk new_AGEMA_reg_buffer_4977 ( .C (clk), .D (new_AGEMA_signal_8441), .Q (new_AGEMA_signal_8442) ) ;
    buf_clk new_AGEMA_reg_buffer_4985 ( .C (clk), .D (new_AGEMA_signal_8449), .Q (new_AGEMA_signal_8450) ) ;
    buf_clk new_AGEMA_reg_buffer_4993 ( .C (clk), .D (new_AGEMA_signal_8457), .Q (new_AGEMA_signal_8458) ) ;
    buf_clk new_AGEMA_reg_buffer_5001 ( .C (clk), .D (new_AGEMA_signal_8465), .Q (new_AGEMA_signal_8466) ) ;
    buf_clk new_AGEMA_reg_buffer_5009 ( .C (clk), .D (new_AGEMA_signal_8473), .Q (new_AGEMA_signal_8474) ) ;
    buf_clk new_AGEMA_reg_buffer_5017 ( .C (clk), .D (new_AGEMA_signal_8481), .Q (new_AGEMA_signal_8482) ) ;
    buf_clk new_AGEMA_reg_buffer_5025 ( .C (clk), .D (new_AGEMA_signal_8489), .Q (new_AGEMA_signal_8490) ) ;
    buf_clk new_AGEMA_reg_buffer_5033 ( .C (clk), .D (new_AGEMA_signal_8497), .Q (new_AGEMA_signal_8498) ) ;
    buf_clk new_AGEMA_reg_buffer_5041 ( .C (clk), .D (new_AGEMA_signal_8505), .Q (new_AGEMA_signal_8506) ) ;
    buf_clk new_AGEMA_reg_buffer_5049 ( .C (clk), .D (new_AGEMA_signal_8513), .Q (new_AGEMA_signal_8514) ) ;
    buf_clk new_AGEMA_reg_buffer_5057 ( .C (clk), .D (new_AGEMA_signal_8521), .Q (new_AGEMA_signal_8522) ) ;
    buf_clk new_AGEMA_reg_buffer_5065 ( .C (clk), .D (new_AGEMA_signal_8529), .Q (new_AGEMA_signal_8530) ) ;
    buf_clk new_AGEMA_reg_buffer_5073 ( .C (clk), .D (new_AGEMA_signal_8537), .Q (new_AGEMA_signal_8538) ) ;
    buf_clk new_AGEMA_reg_buffer_5081 ( .C (clk), .D (new_AGEMA_signal_8545), .Q (new_AGEMA_signal_8546) ) ;
    buf_clk new_AGEMA_reg_buffer_5089 ( .C (clk), .D (new_AGEMA_signal_8553), .Q (new_AGEMA_signal_8554) ) ;
    buf_clk new_AGEMA_reg_buffer_5097 ( .C (clk), .D (new_AGEMA_signal_8561), .Q (new_AGEMA_signal_8562) ) ;
    buf_clk new_AGEMA_reg_buffer_5105 ( .C (clk), .D (new_AGEMA_signal_8569), .Q (new_AGEMA_signal_8570) ) ;
    buf_clk new_AGEMA_reg_buffer_5113 ( .C (clk), .D (new_AGEMA_signal_8577), .Q (new_AGEMA_signal_8578) ) ;
    buf_clk new_AGEMA_reg_buffer_5121 ( .C (clk), .D (new_AGEMA_signal_8585), .Q (new_AGEMA_signal_8586) ) ;
    buf_clk new_AGEMA_reg_buffer_5129 ( .C (clk), .D (new_AGEMA_signal_8593), .Q (new_AGEMA_signal_8594) ) ;
    buf_clk new_AGEMA_reg_buffer_5137 ( .C (clk), .D (new_AGEMA_signal_8601), .Q (new_AGEMA_signal_8602) ) ;
    buf_clk new_AGEMA_reg_buffer_5145 ( .C (clk), .D (new_AGEMA_signal_8609), .Q (new_AGEMA_signal_8610) ) ;
    buf_clk new_AGEMA_reg_buffer_5153 ( .C (clk), .D (new_AGEMA_signal_8617), .Q (new_AGEMA_signal_8618) ) ;
    buf_clk new_AGEMA_reg_buffer_5161 ( .C (clk), .D (new_AGEMA_signal_8625), .Q (new_AGEMA_signal_8626) ) ;
    buf_clk new_AGEMA_reg_buffer_5169 ( .C (clk), .D (new_AGEMA_signal_8633), .Q (new_AGEMA_signal_8634) ) ;
    buf_clk new_AGEMA_reg_buffer_5177 ( .C (clk), .D (new_AGEMA_signal_8641), .Q (new_AGEMA_signal_8642) ) ;
    buf_clk new_AGEMA_reg_buffer_5185 ( .C (clk), .D (new_AGEMA_signal_8649), .Q (new_AGEMA_signal_8650) ) ;
    buf_clk new_AGEMA_reg_buffer_5193 ( .C (clk), .D (new_AGEMA_signal_8657), .Q (new_AGEMA_signal_8658) ) ;
    buf_clk new_AGEMA_reg_buffer_5201 ( .C (clk), .D (new_AGEMA_signal_8665), .Q (new_AGEMA_signal_8666) ) ;
    buf_clk new_AGEMA_reg_buffer_5209 ( .C (clk), .D (new_AGEMA_signal_8673), .Q (new_AGEMA_signal_8674) ) ;
    buf_clk new_AGEMA_reg_buffer_5217 ( .C (clk), .D (new_AGEMA_signal_8681), .Q (new_AGEMA_signal_8682) ) ;
    buf_clk new_AGEMA_reg_buffer_5225 ( .C (clk), .D (new_AGEMA_signal_8689), .Q (new_AGEMA_signal_8690) ) ;
    buf_clk new_AGEMA_reg_buffer_5233 ( .C (clk), .D (new_AGEMA_signal_8697), .Q (new_AGEMA_signal_8698) ) ;
    buf_clk new_AGEMA_reg_buffer_5241 ( .C (clk), .D (new_AGEMA_signal_8705), .Q (new_AGEMA_signal_8706) ) ;
    buf_clk new_AGEMA_reg_buffer_5249 ( .C (clk), .D (new_AGEMA_signal_8713), .Q (new_AGEMA_signal_8714) ) ;
    buf_clk new_AGEMA_reg_buffer_5257 ( .C (clk), .D (new_AGEMA_signal_8721), .Q (new_AGEMA_signal_8722) ) ;
    buf_clk new_AGEMA_reg_buffer_5265 ( .C (clk), .D (new_AGEMA_signal_8729), .Q (new_AGEMA_signal_8730) ) ;
    buf_clk new_AGEMA_reg_buffer_5273 ( .C (clk), .D (new_AGEMA_signal_8737), .Q (new_AGEMA_signal_8738) ) ;
    buf_clk new_AGEMA_reg_buffer_5281 ( .C (clk), .D (new_AGEMA_signal_8745), .Q (new_AGEMA_signal_8746) ) ;
    buf_clk new_AGEMA_reg_buffer_5289 ( .C (clk), .D (new_AGEMA_signal_8753), .Q (new_AGEMA_signal_8754) ) ;
    buf_clk new_AGEMA_reg_buffer_5297 ( .C (clk), .D (new_AGEMA_signal_8761), .Q (new_AGEMA_signal_8762) ) ;
    buf_clk new_AGEMA_reg_buffer_5305 ( .C (clk), .D (new_AGEMA_signal_8769), .Q (new_AGEMA_signal_8770) ) ;
    buf_clk new_AGEMA_reg_buffer_5313 ( .C (clk), .D (new_AGEMA_signal_8777), .Q (new_AGEMA_signal_8778) ) ;
    buf_clk new_AGEMA_reg_buffer_5321 ( .C (clk), .D (new_AGEMA_signal_8785), .Q (new_AGEMA_signal_8786) ) ;
    buf_clk new_AGEMA_reg_buffer_5329 ( .C (clk), .D (new_AGEMA_signal_8793), .Q (new_AGEMA_signal_8794) ) ;
    buf_clk new_AGEMA_reg_buffer_5337 ( .C (clk), .D (new_AGEMA_signal_8801), .Q (new_AGEMA_signal_8802) ) ;
    buf_clk new_AGEMA_reg_buffer_5345 ( .C (clk), .D (new_AGEMA_signal_8809), .Q (new_AGEMA_signal_8810) ) ;
    buf_clk new_AGEMA_reg_buffer_5353 ( .C (clk), .D (new_AGEMA_signal_8817), .Q (new_AGEMA_signal_8818) ) ;
    buf_clk new_AGEMA_reg_buffer_5361 ( .C (clk), .D (new_AGEMA_signal_8825), .Q (new_AGEMA_signal_8826) ) ;
    buf_clk new_AGEMA_reg_buffer_5369 ( .C (clk), .D (new_AGEMA_signal_8833), .Q (new_AGEMA_signal_8834) ) ;
    buf_clk new_AGEMA_reg_buffer_5377 ( .C (clk), .D (new_AGEMA_signal_8841), .Q (new_AGEMA_signal_8842) ) ;
    buf_clk new_AGEMA_reg_buffer_5385 ( .C (clk), .D (new_AGEMA_signal_8849), .Q (new_AGEMA_signal_8850) ) ;
    buf_clk new_AGEMA_reg_buffer_5393 ( .C (clk), .D (new_AGEMA_signal_8857), .Q (new_AGEMA_signal_8858) ) ;
    buf_clk new_AGEMA_reg_buffer_5401 ( .C (clk), .D (new_AGEMA_signal_8865), .Q (new_AGEMA_signal_8866) ) ;
    buf_clk new_AGEMA_reg_buffer_5403 ( .C (clk), .D (new_AGEMA_signal_6461), .Q (new_AGEMA_signal_8868) ) ;
    buf_clk new_AGEMA_reg_buffer_5411 ( .C (clk), .D (new_AGEMA_signal_8875), .Q (new_AGEMA_signal_8876) ) ;
    buf_clk new_AGEMA_reg_buffer_5419 ( .C (clk), .D (new_AGEMA_signal_8883), .Q (new_AGEMA_signal_8884) ) ;
    buf_clk new_AGEMA_reg_buffer_5427 ( .C (clk), .D (new_AGEMA_signal_8891), .Q (new_AGEMA_signal_8892) ) ;
    buf_clk new_AGEMA_reg_buffer_5435 ( .C (clk), .D (new_AGEMA_signal_8899), .Q (new_AGEMA_signal_8900) ) ;
    buf_clk new_AGEMA_reg_buffer_5443 ( .C (clk), .D (new_AGEMA_signal_8907), .Q (new_AGEMA_signal_8908) ) ;
    buf_clk new_AGEMA_reg_buffer_5451 ( .C (clk), .D (new_AGEMA_signal_8915), .Q (new_AGEMA_signal_8916) ) ;
    buf_clk new_AGEMA_reg_buffer_5459 ( .C (clk), .D (new_AGEMA_signal_8923), .Q (new_AGEMA_signal_8924) ) ;
    buf_clk new_AGEMA_reg_buffer_5467 ( .C (clk), .D (new_AGEMA_signal_8931), .Q (new_AGEMA_signal_8932) ) ;
    buf_clk new_AGEMA_reg_buffer_5475 ( .C (clk), .D (new_AGEMA_signal_8939), .Q (new_AGEMA_signal_8940) ) ;
    buf_clk new_AGEMA_reg_buffer_5483 ( .C (clk), .D (new_AGEMA_signal_8947), .Q (new_AGEMA_signal_8948) ) ;
    buf_clk new_AGEMA_reg_buffer_5491 ( .C (clk), .D (new_AGEMA_signal_8955), .Q (new_AGEMA_signal_8956) ) ;
    buf_clk new_AGEMA_reg_buffer_5499 ( .C (clk), .D (new_AGEMA_signal_8963), .Q (new_AGEMA_signal_8964) ) ;
    buf_clk new_AGEMA_reg_buffer_5507 ( .C (clk), .D (new_AGEMA_signal_8971), .Q (new_AGEMA_signal_8972) ) ;
    buf_clk new_AGEMA_reg_buffer_5515 ( .C (clk), .D (new_AGEMA_signal_8979), .Q (new_AGEMA_signal_8980) ) ;
    buf_clk new_AGEMA_reg_buffer_5523 ( .C (clk), .D (new_AGEMA_signal_8987), .Q (new_AGEMA_signal_8988) ) ;
    buf_clk new_AGEMA_reg_buffer_5531 ( .C (clk), .D (new_AGEMA_signal_8995), .Q (new_AGEMA_signal_8996) ) ;
    buf_clk new_AGEMA_reg_buffer_5539 ( .C (clk), .D (new_AGEMA_signal_9003), .Q (new_AGEMA_signal_9004) ) ;
    buf_clk new_AGEMA_reg_buffer_5547 ( .C (clk), .D (new_AGEMA_signal_9011), .Q (new_AGEMA_signal_9012) ) ;
    buf_clk new_AGEMA_reg_buffer_5555 ( .C (clk), .D (new_AGEMA_signal_9019), .Q (new_AGEMA_signal_9020) ) ;
    buf_clk new_AGEMA_reg_buffer_5563 ( .C (clk), .D (new_AGEMA_signal_9027), .Q (new_AGEMA_signal_9028) ) ;
    buf_clk new_AGEMA_reg_buffer_5571 ( .C (clk), .D (new_AGEMA_signal_9035), .Q (new_AGEMA_signal_9036) ) ;
    buf_clk new_AGEMA_reg_buffer_5579 ( .C (clk), .D (new_AGEMA_signal_9043), .Q (new_AGEMA_signal_9044) ) ;
    buf_clk new_AGEMA_reg_buffer_5587 ( .C (clk), .D (new_AGEMA_signal_9051), .Q (new_AGEMA_signal_9052) ) ;
    buf_clk new_AGEMA_reg_buffer_5595 ( .C (clk), .D (new_AGEMA_signal_9059), .Q (new_AGEMA_signal_9060) ) ;
    buf_clk new_AGEMA_reg_buffer_5603 ( .C (clk), .D (new_AGEMA_signal_9067), .Q (new_AGEMA_signal_9068) ) ;
    buf_clk new_AGEMA_reg_buffer_5611 ( .C (clk), .D (new_AGEMA_signal_9075), .Q (new_AGEMA_signal_9076) ) ;
    buf_clk new_AGEMA_reg_buffer_5619 ( .C (clk), .D (new_AGEMA_signal_9083), .Q (new_AGEMA_signal_9084) ) ;
    buf_clk new_AGEMA_reg_buffer_5627 ( .C (clk), .D (new_AGEMA_signal_9091), .Q (new_AGEMA_signal_9092) ) ;
    buf_clk new_AGEMA_reg_buffer_5635 ( .C (clk), .D (new_AGEMA_signal_9099), .Q (new_AGEMA_signal_9100) ) ;
    buf_clk new_AGEMA_reg_buffer_5643 ( .C (clk), .D (new_AGEMA_signal_9107), .Q (new_AGEMA_signal_9108) ) ;
    buf_clk new_AGEMA_reg_buffer_5651 ( .C (clk), .D (new_AGEMA_signal_9115), .Q (new_AGEMA_signal_9116) ) ;
    buf_clk new_AGEMA_reg_buffer_5659 ( .C (clk), .D (new_AGEMA_signal_9123), .Q (new_AGEMA_signal_9124) ) ;
    buf_clk new_AGEMA_reg_buffer_5667 ( .C (clk), .D (new_AGEMA_signal_9131), .Q (new_AGEMA_signal_9132) ) ;
    buf_clk new_AGEMA_reg_buffer_5675 ( .C (clk), .D (new_AGEMA_signal_9139), .Q (new_AGEMA_signal_9140) ) ;
    buf_clk new_AGEMA_reg_buffer_5683 ( .C (clk), .D (new_AGEMA_signal_9147), .Q (new_AGEMA_signal_9148) ) ;
    buf_clk new_AGEMA_reg_buffer_5691 ( .C (clk), .D (new_AGEMA_signal_9155), .Q (new_AGEMA_signal_9156) ) ;
    buf_clk new_AGEMA_reg_buffer_5699 ( .C (clk), .D (new_AGEMA_signal_9163), .Q (new_AGEMA_signal_9164) ) ;
    buf_clk new_AGEMA_reg_buffer_5707 ( .C (clk), .D (new_AGEMA_signal_9171), .Q (new_AGEMA_signal_9172) ) ;
    buf_clk new_AGEMA_reg_buffer_5715 ( .C (clk), .D (new_AGEMA_signal_9179), .Q (new_AGEMA_signal_9180) ) ;
    buf_clk new_AGEMA_reg_buffer_5723 ( .C (clk), .D (new_AGEMA_signal_9187), .Q (new_AGEMA_signal_9188) ) ;
    buf_clk new_AGEMA_reg_buffer_5731 ( .C (clk), .D (new_AGEMA_signal_9195), .Q (new_AGEMA_signal_9196) ) ;
    buf_clk new_AGEMA_reg_buffer_5739 ( .C (clk), .D (new_AGEMA_signal_9203), .Q (new_AGEMA_signal_9204) ) ;
    buf_clk new_AGEMA_reg_buffer_5747 ( .C (clk), .D (new_AGEMA_signal_9211), .Q (new_AGEMA_signal_9212) ) ;
    buf_clk new_AGEMA_reg_buffer_5755 ( .C (clk), .D (new_AGEMA_signal_9219), .Q (new_AGEMA_signal_9220) ) ;
    buf_clk new_AGEMA_reg_buffer_5763 ( .C (clk), .D (new_AGEMA_signal_9227), .Q (new_AGEMA_signal_9228) ) ;
    buf_clk new_AGEMA_reg_buffer_5771 ( .C (clk), .D (new_AGEMA_signal_9235), .Q (new_AGEMA_signal_9236) ) ;
    buf_clk new_AGEMA_reg_buffer_5779 ( .C (clk), .D (new_AGEMA_signal_9243), .Q (new_AGEMA_signal_9244) ) ;
    buf_clk new_AGEMA_reg_buffer_5787 ( .C (clk), .D (new_AGEMA_signal_9251), .Q (new_AGEMA_signal_9252) ) ;
    buf_clk new_AGEMA_reg_buffer_5795 ( .C (clk), .D (new_AGEMA_signal_9259), .Q (new_AGEMA_signal_9260) ) ;
    buf_clk new_AGEMA_reg_buffer_5803 ( .C (clk), .D (new_AGEMA_signal_9267), .Q (new_AGEMA_signal_9268) ) ;
    buf_clk new_AGEMA_reg_buffer_5811 ( .C (clk), .D (new_AGEMA_signal_9275), .Q (new_AGEMA_signal_9276) ) ;
    buf_clk new_AGEMA_reg_buffer_5819 ( .C (clk), .D (new_AGEMA_signal_9283), .Q (new_AGEMA_signal_9284) ) ;
    buf_clk new_AGEMA_reg_buffer_5827 ( .C (clk), .D (new_AGEMA_signal_9291), .Q (new_AGEMA_signal_9292) ) ;
    buf_clk new_AGEMA_reg_buffer_5835 ( .C (clk), .D (new_AGEMA_signal_9299), .Q (new_AGEMA_signal_9300) ) ;
    buf_clk new_AGEMA_reg_buffer_5843 ( .C (clk), .D (new_AGEMA_signal_9307), .Q (new_AGEMA_signal_9308) ) ;
    buf_clk new_AGEMA_reg_buffer_5851 ( .C (clk), .D (new_AGEMA_signal_9315), .Q (new_AGEMA_signal_9316) ) ;
    buf_clk new_AGEMA_reg_buffer_5859 ( .C (clk), .D (new_AGEMA_signal_9323), .Q (new_AGEMA_signal_9324) ) ;
    buf_clk new_AGEMA_reg_buffer_5867 ( .C (clk), .D (new_AGEMA_signal_9331), .Q (new_AGEMA_signal_9332) ) ;
    buf_clk new_AGEMA_reg_buffer_5875 ( .C (clk), .D (new_AGEMA_signal_9339), .Q (new_AGEMA_signal_9340) ) ;
    buf_clk new_AGEMA_reg_buffer_5883 ( .C (clk), .D (new_AGEMA_signal_9347), .Q (new_AGEMA_signal_9348) ) ;
    buf_clk new_AGEMA_reg_buffer_5891 ( .C (clk), .D (new_AGEMA_signal_9355), .Q (new_AGEMA_signal_9356) ) ;
    buf_clk new_AGEMA_reg_buffer_5899 ( .C (clk), .D (new_AGEMA_signal_9363), .Q (new_AGEMA_signal_9364) ) ;
    buf_clk new_AGEMA_reg_buffer_5907 ( .C (clk), .D (new_AGEMA_signal_9371), .Q (new_AGEMA_signal_9372) ) ;
    buf_clk new_AGEMA_reg_buffer_5915 ( .C (clk), .D (new_AGEMA_signal_9379), .Q (new_AGEMA_signal_9380) ) ;
    buf_clk new_AGEMA_reg_buffer_5923 ( .C (clk), .D (new_AGEMA_signal_9387), .Q (new_AGEMA_signal_9388) ) ;
    buf_clk new_AGEMA_reg_buffer_5931 ( .C (clk), .D (new_AGEMA_signal_9395), .Q (new_AGEMA_signal_9396) ) ;
    buf_clk new_AGEMA_reg_buffer_5939 ( .C (clk), .D (new_AGEMA_signal_9403), .Q (new_AGEMA_signal_9404) ) ;
    buf_clk new_AGEMA_reg_buffer_5947 ( .C (clk), .D (new_AGEMA_signal_9411), .Q (new_AGEMA_signal_9412) ) ;
    buf_clk new_AGEMA_reg_buffer_5955 ( .C (clk), .D (new_AGEMA_signal_9419), .Q (new_AGEMA_signal_9420) ) ;
    buf_clk new_AGEMA_reg_buffer_5963 ( .C (clk), .D (new_AGEMA_signal_9427), .Q (new_AGEMA_signal_9428) ) ;
    buf_clk new_AGEMA_reg_buffer_5971 ( .C (clk), .D (new_AGEMA_signal_9435), .Q (new_AGEMA_signal_9436) ) ;
    buf_clk new_AGEMA_reg_buffer_5979 ( .C (clk), .D (new_AGEMA_signal_9443), .Q (new_AGEMA_signal_9444) ) ;
    buf_clk new_AGEMA_reg_buffer_5987 ( .C (clk), .D (new_AGEMA_signal_9451), .Q (new_AGEMA_signal_9452) ) ;
    buf_clk new_AGEMA_reg_buffer_5995 ( .C (clk), .D (new_AGEMA_signal_9459), .Q (new_AGEMA_signal_9460) ) ;
    buf_clk new_AGEMA_reg_buffer_6003 ( .C (clk), .D (new_AGEMA_signal_9467), .Q (new_AGEMA_signal_9468) ) ;
    buf_clk new_AGEMA_reg_buffer_6011 ( .C (clk), .D (new_AGEMA_signal_9475), .Q (new_AGEMA_signal_9476) ) ;
    buf_clk new_AGEMA_reg_buffer_6019 ( .C (clk), .D (new_AGEMA_signal_9483), .Q (new_AGEMA_signal_9484) ) ;
    buf_clk new_AGEMA_reg_buffer_6027 ( .C (clk), .D (new_AGEMA_signal_9491), .Q (new_AGEMA_signal_9492) ) ;
    buf_clk new_AGEMA_reg_buffer_6035 ( .C (clk), .D (new_AGEMA_signal_9499), .Q (new_AGEMA_signal_9500) ) ;
    buf_clk new_AGEMA_reg_buffer_6043 ( .C (clk), .D (new_AGEMA_signal_9507), .Q (new_AGEMA_signal_9508) ) ;
    buf_clk new_AGEMA_reg_buffer_6051 ( .C (clk), .D (new_AGEMA_signal_9515), .Q (new_AGEMA_signal_9516) ) ;
    buf_clk new_AGEMA_reg_buffer_6059 ( .C (clk), .D (new_AGEMA_signal_9523), .Q (new_AGEMA_signal_9524) ) ;
    buf_clk new_AGEMA_reg_buffer_6067 ( .C (clk), .D (new_AGEMA_signal_9531), .Q (new_AGEMA_signal_9532) ) ;
    buf_clk new_AGEMA_reg_buffer_6075 ( .C (clk), .D (new_AGEMA_signal_9539), .Q (new_AGEMA_signal_9540) ) ;
    buf_clk new_AGEMA_reg_buffer_6083 ( .C (clk), .D (new_AGEMA_signal_9547), .Q (new_AGEMA_signal_9548) ) ;
    buf_clk new_AGEMA_reg_buffer_6091 ( .C (clk), .D (new_AGEMA_signal_9555), .Q (new_AGEMA_signal_9556) ) ;
    buf_clk new_AGEMA_reg_buffer_6099 ( .C (clk), .D (new_AGEMA_signal_9563), .Q (new_AGEMA_signal_9564) ) ;
    buf_clk new_AGEMA_reg_buffer_6107 ( .C (clk), .D (new_AGEMA_signal_9571), .Q (new_AGEMA_signal_9572) ) ;
    buf_clk new_AGEMA_reg_buffer_6115 ( .C (clk), .D (new_AGEMA_signal_9579), .Q (new_AGEMA_signal_9580) ) ;
    buf_clk new_AGEMA_reg_buffer_6123 ( .C (clk), .D (new_AGEMA_signal_9587), .Q (new_AGEMA_signal_9588) ) ;
    buf_clk new_AGEMA_reg_buffer_6131 ( .C (clk), .D (new_AGEMA_signal_9595), .Q (new_AGEMA_signal_9596) ) ;
    buf_clk new_AGEMA_reg_buffer_6139 ( .C (clk), .D (new_AGEMA_signal_9603), .Q (new_AGEMA_signal_9604) ) ;
    buf_clk new_AGEMA_reg_buffer_6147 ( .C (clk), .D (new_AGEMA_signal_9611), .Q (new_AGEMA_signal_9612) ) ;
    buf_clk new_AGEMA_reg_buffer_6155 ( .C (clk), .D (new_AGEMA_signal_9619), .Q (new_AGEMA_signal_9620) ) ;
    buf_clk new_AGEMA_reg_buffer_6163 ( .C (clk), .D (new_AGEMA_signal_9627), .Q (new_AGEMA_signal_9628) ) ;
    buf_clk new_AGEMA_reg_buffer_6171 ( .C (clk), .D (new_AGEMA_signal_9635), .Q (new_AGEMA_signal_9636) ) ;
    buf_clk new_AGEMA_reg_buffer_6461 ( .C (clk), .D (new_AGEMA_signal_7331), .Q (new_AGEMA_signal_9926) ) ;
    buf_clk new_AGEMA_reg_buffer_6469 ( .C (clk), .D (new_AGEMA_signal_9933), .Q (new_AGEMA_signal_9934) ) ;
    buf_clk new_AGEMA_reg_buffer_6477 ( .C (clk), .D (new_AGEMA_signal_9941), .Q (new_AGEMA_signal_9942) ) ;
    buf_clk new_AGEMA_reg_buffer_6485 ( .C (clk), .D (new_AGEMA_signal_9949), .Q (new_AGEMA_signal_9950) ) ;
    buf_clk new_AGEMA_reg_buffer_6493 ( .C (clk), .D (new_AGEMA_signal_9957), .Q (new_AGEMA_signal_9958) ) ;
    buf_clk new_AGEMA_reg_buffer_6495 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_1_DQ), .Q (new_AGEMA_signal_9960) ) ;
    buf_clk new_AGEMA_reg_buffer_6497 ( .C (clk), .D (new_AGEMA_signal_3674), .Q (new_AGEMA_signal_9962) ) ;
    buf_clk new_AGEMA_reg_buffer_6499 ( .C (clk), .D (new_AGEMA_signal_3675), .Q (new_AGEMA_signal_9964) ) ;
    buf_clk new_AGEMA_reg_buffer_6501 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_3_DQ), .Q (new_AGEMA_signal_9966) ) ;
    buf_clk new_AGEMA_reg_buffer_6503 ( .C (clk), .D (new_AGEMA_signal_3678), .Q (new_AGEMA_signal_9968) ) ;
    buf_clk new_AGEMA_reg_buffer_6505 ( .C (clk), .D (new_AGEMA_signal_3679), .Q (new_AGEMA_signal_9970) ) ;
    buf_clk new_AGEMA_reg_buffer_6507 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_5_DQ), .Q (new_AGEMA_signal_9972) ) ;
    buf_clk new_AGEMA_reg_buffer_6509 ( .C (clk), .D (new_AGEMA_signal_3680), .Q (new_AGEMA_signal_9974) ) ;
    buf_clk new_AGEMA_reg_buffer_6511 ( .C (clk), .D (new_AGEMA_signal_3681), .Q (new_AGEMA_signal_9976) ) ;
    buf_clk new_AGEMA_reg_buffer_6513 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_7_DQ), .Q (new_AGEMA_signal_9978) ) ;
    buf_clk new_AGEMA_reg_buffer_6515 ( .C (clk), .D (new_AGEMA_signal_3684), .Q (new_AGEMA_signal_9980) ) ;
    buf_clk new_AGEMA_reg_buffer_6517 ( .C (clk), .D (new_AGEMA_signal_3685), .Q (new_AGEMA_signal_9982) ) ;
    buf_clk new_AGEMA_reg_buffer_6519 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_9_DQ), .Q (new_AGEMA_signal_9984) ) ;
    buf_clk new_AGEMA_reg_buffer_6521 ( .C (clk), .D (new_AGEMA_signal_3686), .Q (new_AGEMA_signal_9986) ) ;
    buf_clk new_AGEMA_reg_buffer_6523 ( .C (clk), .D (new_AGEMA_signal_3687), .Q (new_AGEMA_signal_9988) ) ;
    buf_clk new_AGEMA_reg_buffer_6525 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_11_DQ), .Q (new_AGEMA_signal_9990) ) ;
    buf_clk new_AGEMA_reg_buffer_6527 ( .C (clk), .D (new_AGEMA_signal_3690), .Q (new_AGEMA_signal_9992) ) ;
    buf_clk new_AGEMA_reg_buffer_6529 ( .C (clk), .D (new_AGEMA_signal_3691), .Q (new_AGEMA_signal_9994) ) ;
    buf_clk new_AGEMA_reg_buffer_6531 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_13_DQ), .Q (new_AGEMA_signal_9996) ) ;
    buf_clk new_AGEMA_reg_buffer_6533 ( .C (clk), .D (new_AGEMA_signal_3692), .Q (new_AGEMA_signal_9998) ) ;
    buf_clk new_AGEMA_reg_buffer_6535 ( .C (clk), .D (new_AGEMA_signal_3693), .Q (new_AGEMA_signal_10000) ) ;
    buf_clk new_AGEMA_reg_buffer_6537 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_15_DQ), .Q (new_AGEMA_signal_10002) ) ;
    buf_clk new_AGEMA_reg_buffer_6539 ( .C (clk), .D (new_AGEMA_signal_3696), .Q (new_AGEMA_signal_10004) ) ;
    buf_clk new_AGEMA_reg_buffer_6541 ( .C (clk), .D (new_AGEMA_signal_3697), .Q (new_AGEMA_signal_10006) ) ;
    buf_clk new_AGEMA_reg_buffer_6543 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_17_DQ), .Q (new_AGEMA_signal_10008) ) ;
    buf_clk new_AGEMA_reg_buffer_6545 ( .C (clk), .D (new_AGEMA_signal_3698), .Q (new_AGEMA_signal_10010) ) ;
    buf_clk new_AGEMA_reg_buffer_6547 ( .C (clk), .D (new_AGEMA_signal_3699), .Q (new_AGEMA_signal_10012) ) ;
    buf_clk new_AGEMA_reg_buffer_6549 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_19_DQ), .Q (new_AGEMA_signal_10014) ) ;
    buf_clk new_AGEMA_reg_buffer_6551 ( .C (clk), .D (new_AGEMA_signal_3702), .Q (new_AGEMA_signal_10016) ) ;
    buf_clk new_AGEMA_reg_buffer_6553 ( .C (clk), .D (new_AGEMA_signal_3703), .Q (new_AGEMA_signal_10018) ) ;
    buf_clk new_AGEMA_reg_buffer_6555 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_21_DQ), .Q (new_AGEMA_signal_10020) ) ;
    buf_clk new_AGEMA_reg_buffer_6557 ( .C (clk), .D (new_AGEMA_signal_3704), .Q (new_AGEMA_signal_10022) ) ;
    buf_clk new_AGEMA_reg_buffer_6559 ( .C (clk), .D (new_AGEMA_signal_3705), .Q (new_AGEMA_signal_10024) ) ;
    buf_clk new_AGEMA_reg_buffer_6561 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_23_DQ), .Q (new_AGEMA_signal_10026) ) ;
    buf_clk new_AGEMA_reg_buffer_6563 ( .C (clk), .D (new_AGEMA_signal_3708), .Q (new_AGEMA_signal_10028) ) ;
    buf_clk new_AGEMA_reg_buffer_6565 ( .C (clk), .D (new_AGEMA_signal_3709), .Q (new_AGEMA_signal_10030) ) ;
    buf_clk new_AGEMA_reg_buffer_6567 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_25_DQ), .Q (new_AGEMA_signal_10032) ) ;
    buf_clk new_AGEMA_reg_buffer_6569 ( .C (clk), .D (new_AGEMA_signal_3710), .Q (new_AGEMA_signal_10034) ) ;
    buf_clk new_AGEMA_reg_buffer_6571 ( .C (clk), .D (new_AGEMA_signal_3711), .Q (new_AGEMA_signal_10036) ) ;
    buf_clk new_AGEMA_reg_buffer_6573 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_27_DQ), .Q (new_AGEMA_signal_10038) ) ;
    buf_clk new_AGEMA_reg_buffer_6575 ( .C (clk), .D (new_AGEMA_signal_3714), .Q (new_AGEMA_signal_10040) ) ;
    buf_clk new_AGEMA_reg_buffer_6577 ( .C (clk), .D (new_AGEMA_signal_3715), .Q (new_AGEMA_signal_10042) ) ;
    buf_clk new_AGEMA_reg_buffer_6579 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_29_DQ), .Q (new_AGEMA_signal_10044) ) ;
    buf_clk new_AGEMA_reg_buffer_6581 ( .C (clk), .D (new_AGEMA_signal_3716), .Q (new_AGEMA_signal_10046) ) ;
    buf_clk new_AGEMA_reg_buffer_6583 ( .C (clk), .D (new_AGEMA_signal_3717), .Q (new_AGEMA_signal_10048) ) ;
    buf_clk new_AGEMA_reg_buffer_6585 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_31_DQ), .Q (new_AGEMA_signal_10050) ) ;
    buf_clk new_AGEMA_reg_buffer_6587 ( .C (clk), .D (new_AGEMA_signal_3720), .Q (new_AGEMA_signal_10052) ) ;
    buf_clk new_AGEMA_reg_buffer_6589 ( .C (clk), .D (new_AGEMA_signal_3721), .Q (new_AGEMA_signal_10054) ) ;
    buf_clk new_AGEMA_reg_buffer_6591 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_33_DQ), .Q (new_AGEMA_signal_10056) ) ;
    buf_clk new_AGEMA_reg_buffer_6593 ( .C (clk), .D (new_AGEMA_signal_3722), .Q (new_AGEMA_signal_10058) ) ;
    buf_clk new_AGEMA_reg_buffer_6595 ( .C (clk), .D (new_AGEMA_signal_3723), .Q (new_AGEMA_signal_10060) ) ;
    buf_clk new_AGEMA_reg_buffer_6597 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_35_DQ), .Q (new_AGEMA_signal_10062) ) ;
    buf_clk new_AGEMA_reg_buffer_6599 ( .C (clk), .D (new_AGEMA_signal_3726), .Q (new_AGEMA_signal_10064) ) ;
    buf_clk new_AGEMA_reg_buffer_6601 ( .C (clk), .D (new_AGEMA_signal_3727), .Q (new_AGEMA_signal_10066) ) ;
    buf_clk new_AGEMA_reg_buffer_6603 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_37_DQ), .Q (new_AGEMA_signal_10068) ) ;
    buf_clk new_AGEMA_reg_buffer_6605 ( .C (clk), .D (new_AGEMA_signal_3728), .Q (new_AGEMA_signal_10070) ) ;
    buf_clk new_AGEMA_reg_buffer_6607 ( .C (clk), .D (new_AGEMA_signal_3729), .Q (new_AGEMA_signal_10072) ) ;
    buf_clk new_AGEMA_reg_buffer_6609 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_39_DQ), .Q (new_AGEMA_signal_10074) ) ;
    buf_clk new_AGEMA_reg_buffer_6611 ( .C (clk), .D (new_AGEMA_signal_3732), .Q (new_AGEMA_signal_10076) ) ;
    buf_clk new_AGEMA_reg_buffer_6613 ( .C (clk), .D (new_AGEMA_signal_3733), .Q (new_AGEMA_signal_10078) ) ;
    buf_clk new_AGEMA_reg_buffer_6615 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_41_DQ), .Q (new_AGEMA_signal_10080) ) ;
    buf_clk new_AGEMA_reg_buffer_6617 ( .C (clk), .D (new_AGEMA_signal_3734), .Q (new_AGEMA_signal_10082) ) ;
    buf_clk new_AGEMA_reg_buffer_6619 ( .C (clk), .D (new_AGEMA_signal_3735), .Q (new_AGEMA_signal_10084) ) ;
    buf_clk new_AGEMA_reg_buffer_6621 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_43_DQ), .Q (new_AGEMA_signal_10086) ) ;
    buf_clk new_AGEMA_reg_buffer_6623 ( .C (clk), .D (new_AGEMA_signal_3738), .Q (new_AGEMA_signal_10088) ) ;
    buf_clk new_AGEMA_reg_buffer_6625 ( .C (clk), .D (new_AGEMA_signal_3739), .Q (new_AGEMA_signal_10090) ) ;
    buf_clk new_AGEMA_reg_buffer_6627 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_45_DQ), .Q (new_AGEMA_signal_10092) ) ;
    buf_clk new_AGEMA_reg_buffer_6629 ( .C (clk), .D (new_AGEMA_signal_3740), .Q (new_AGEMA_signal_10094) ) ;
    buf_clk new_AGEMA_reg_buffer_6631 ( .C (clk), .D (new_AGEMA_signal_3741), .Q (new_AGEMA_signal_10096) ) ;
    buf_clk new_AGEMA_reg_buffer_6633 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_47_DQ), .Q (new_AGEMA_signal_10098) ) ;
    buf_clk new_AGEMA_reg_buffer_6635 ( .C (clk), .D (new_AGEMA_signal_3744), .Q (new_AGEMA_signal_10100) ) ;
    buf_clk new_AGEMA_reg_buffer_6637 ( .C (clk), .D (new_AGEMA_signal_3745), .Q (new_AGEMA_signal_10102) ) ;
    buf_clk new_AGEMA_reg_buffer_6639 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_49_DQ), .Q (new_AGEMA_signal_10104) ) ;
    buf_clk new_AGEMA_reg_buffer_6641 ( .C (clk), .D (new_AGEMA_signal_3746), .Q (new_AGEMA_signal_10106) ) ;
    buf_clk new_AGEMA_reg_buffer_6643 ( .C (clk), .D (new_AGEMA_signal_3747), .Q (new_AGEMA_signal_10108) ) ;
    buf_clk new_AGEMA_reg_buffer_6645 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_51_DQ), .Q (new_AGEMA_signal_10110) ) ;
    buf_clk new_AGEMA_reg_buffer_6647 ( .C (clk), .D (new_AGEMA_signal_3750), .Q (new_AGEMA_signal_10112) ) ;
    buf_clk new_AGEMA_reg_buffer_6649 ( .C (clk), .D (new_AGEMA_signal_3751), .Q (new_AGEMA_signal_10114) ) ;
    buf_clk new_AGEMA_reg_buffer_6651 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_53_DQ), .Q (new_AGEMA_signal_10116) ) ;
    buf_clk new_AGEMA_reg_buffer_6653 ( .C (clk), .D (new_AGEMA_signal_3752), .Q (new_AGEMA_signal_10118) ) ;
    buf_clk new_AGEMA_reg_buffer_6655 ( .C (clk), .D (new_AGEMA_signal_3753), .Q (new_AGEMA_signal_10120) ) ;
    buf_clk new_AGEMA_reg_buffer_6657 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_55_DQ), .Q (new_AGEMA_signal_10122) ) ;
    buf_clk new_AGEMA_reg_buffer_6659 ( .C (clk), .D (new_AGEMA_signal_3756), .Q (new_AGEMA_signal_10124) ) ;
    buf_clk new_AGEMA_reg_buffer_6661 ( .C (clk), .D (new_AGEMA_signal_3757), .Q (new_AGEMA_signal_10126) ) ;
    buf_clk new_AGEMA_reg_buffer_6663 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_57_DQ), .Q (new_AGEMA_signal_10128) ) ;
    buf_clk new_AGEMA_reg_buffer_6665 ( .C (clk), .D (new_AGEMA_signal_3758), .Q (new_AGEMA_signal_10130) ) ;
    buf_clk new_AGEMA_reg_buffer_6667 ( .C (clk), .D (new_AGEMA_signal_3759), .Q (new_AGEMA_signal_10132) ) ;
    buf_clk new_AGEMA_reg_buffer_6669 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_59_DQ), .Q (new_AGEMA_signal_10134) ) ;
    buf_clk new_AGEMA_reg_buffer_6671 ( .C (clk), .D (new_AGEMA_signal_3762), .Q (new_AGEMA_signal_10136) ) ;
    buf_clk new_AGEMA_reg_buffer_6673 ( .C (clk), .D (new_AGEMA_signal_3763), .Q (new_AGEMA_signal_10138) ) ;
    buf_clk new_AGEMA_reg_buffer_6675 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_61_DQ), .Q (new_AGEMA_signal_10140) ) ;
    buf_clk new_AGEMA_reg_buffer_6677 ( .C (clk), .D (new_AGEMA_signal_3764), .Q (new_AGEMA_signal_10142) ) ;
    buf_clk new_AGEMA_reg_buffer_6679 ( .C (clk), .D (new_AGEMA_signal_3765), .Q (new_AGEMA_signal_10144) ) ;
    buf_clk new_AGEMA_reg_buffer_6681 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_63_DQ), .Q (new_AGEMA_signal_10146) ) ;
    buf_clk new_AGEMA_reg_buffer_6683 ( .C (clk), .D (new_AGEMA_signal_3768), .Q (new_AGEMA_signal_10148) ) ;
    buf_clk new_AGEMA_reg_buffer_6685 ( .C (clk), .D (new_AGEMA_signal_3769), .Q (new_AGEMA_signal_10150) ) ;

    /* cells in depth 8 */
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U127 ( .a ({new_AGEMA_signal_7355, new_AGEMA_signal_7347, new_AGEMA_signal_7339}), .b ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, Midori_rounds_SR_Result[8]}), .c ({DataOut_s2[8], DataOut_s1[8], DataOut_s0[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U125 ( .a ({new_AGEMA_signal_7379, new_AGEMA_signal_7371, new_AGEMA_signal_7363}), .b ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, Midori_rounds_SR_Result[46]}), .c ({DataOut_s2[6], DataOut_s1[6], DataOut_s0[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U123 ( .a ({new_AGEMA_signal_7403, new_AGEMA_signal_7395, new_AGEMA_signal_7387}), .b ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, Midori_rounds_SR_Result[62]}), .c ({DataOut_s2[62], DataOut_s1[62], DataOut_s0[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U121 ( .a ({new_AGEMA_signal_7427, new_AGEMA_signal_7419, new_AGEMA_signal_7411}), .b ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, Midori_rounds_SR_Result[60]}), .c ({DataOut_s2[60], DataOut_s1[60], DataOut_s0[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U118 ( .a ({new_AGEMA_signal_7451, new_AGEMA_signal_7443, new_AGEMA_signal_7435}), .b ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, Midori_rounds_SR_Result[34]}), .c ({DataOut_s2[58], DataOut_s1[58], DataOut_s0[58]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U116 ( .a ({new_AGEMA_signal_7475, new_AGEMA_signal_7467, new_AGEMA_signal_7459}), .b ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, Midori_rounds_SR_Result[32]}), .c ({DataOut_s2[56], DataOut_s1[56], DataOut_s0[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U114 ( .a ({new_AGEMA_signal_7499, new_AGEMA_signal_7491, new_AGEMA_signal_7483}), .b ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, Midori_rounds_SR_Result[6]}), .c ({DataOut_s2[54], DataOut_s1[54], DataOut_s0[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U112 ( .a ({new_AGEMA_signal_7523, new_AGEMA_signal_7515, new_AGEMA_signal_7507}), .b ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, Midori_rounds_SR_Result[4]}), .c ({DataOut_s2[52], DataOut_s1[52], DataOut_s0[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U110 ( .a ({new_AGEMA_signal_7547, new_AGEMA_signal_7539, new_AGEMA_signal_7531}), .b ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, Midori_rounds_SR_Result[26]}), .c ({DataOut_s2[50], DataOut_s1[50], DataOut_s0[50]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U109 ( .a ({new_AGEMA_signal_7571, new_AGEMA_signal_7563, new_AGEMA_signal_7555}), .b ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, Midori_rounds_SR_Result[44]}), .c ({DataOut_s2[4], DataOut_s1[4], DataOut_s0[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U107 ( .a ({new_AGEMA_signal_7595, new_AGEMA_signal_7587, new_AGEMA_signal_7579}), .b ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, Midori_rounds_SR_Result[24]}), .c ({DataOut_s2[48], DataOut_s1[48], DataOut_s0[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U105 ( .a ({new_AGEMA_signal_7619, new_AGEMA_signal_7611, new_AGEMA_signal_7603}), .b ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, Midori_rounds_SR_Result[42]}), .c ({DataOut_s2[46], DataOut_s1[46], DataOut_s0[46]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U103 ( .a ({new_AGEMA_signal_7643, new_AGEMA_signal_7635, new_AGEMA_signal_7627}), .b ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, Midori_rounds_SR_Result[40]}), .c ({DataOut_s2[44], DataOut_s1[44], DataOut_s0[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U101 ( .a ({new_AGEMA_signal_7667, new_AGEMA_signal_7659, new_AGEMA_signal_7651}), .b ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, Midori_rounds_SR_Result[54]}), .c ({DataOut_s2[42], DataOut_s1[42], DataOut_s0[42]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U99 ( .a ({new_AGEMA_signal_7691, new_AGEMA_signal_7683, new_AGEMA_signal_7675}), .b ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, Midori_rounds_SR_Result[52]}), .c ({DataOut_s2[40], DataOut_s1[40], DataOut_s0[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U96 ( .a ({new_AGEMA_signal_7715, new_AGEMA_signal_7707, new_AGEMA_signal_7699}), .b ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, Midori_rounds_SR_Result[18]}), .c ({DataOut_s2[38], DataOut_s1[38], DataOut_s0[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U94 ( .a ({new_AGEMA_signal_7739, new_AGEMA_signal_7731, new_AGEMA_signal_7723}), .b ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, Midori_rounds_SR_Result[16]}), .c ({DataOut_s2[36], DataOut_s1[36], DataOut_s0[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U92 ( .a ({new_AGEMA_signal_7763, new_AGEMA_signal_7755, new_AGEMA_signal_7747}), .b ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, Midori_rounds_SR_Result[14]}), .c ({DataOut_s2[34], DataOut_s1[34], DataOut_s0[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U90 ( .a ({new_AGEMA_signal_7787, new_AGEMA_signal_7779, new_AGEMA_signal_7771}), .b ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, Midori_rounds_SR_Result[12]}), .c ({DataOut_s2[32], DataOut_s1[32], DataOut_s0[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U88 ( .a ({new_AGEMA_signal_7811, new_AGEMA_signal_7803, new_AGEMA_signal_7795}), .b ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, Midori_rounds_SR_Result[2]}), .c ({DataOut_s2[30], DataOut_s1[30], DataOut_s0[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U87 ( .a ({new_AGEMA_signal_7835, new_AGEMA_signal_7827, new_AGEMA_signal_7819}), .b ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, Midori_rounds_SR_Result[50]}), .c ({DataOut_s2[2], DataOut_s1[2], DataOut_s0[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U85 ( .a ({new_AGEMA_signal_7859, new_AGEMA_signal_7851, new_AGEMA_signal_7843}), .b ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, Midori_rounds_SR_Result[0]}), .c ({DataOut_s2[28], DataOut_s1[28], DataOut_s0[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U83 ( .a ({new_AGEMA_signal_7883, new_AGEMA_signal_7875, new_AGEMA_signal_7867}), .b ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, Midori_rounds_SR_Result[30]}), .c ({DataOut_s2[26], DataOut_s1[26], DataOut_s0[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U81 ( .a ({new_AGEMA_signal_7907, new_AGEMA_signal_7899, new_AGEMA_signal_7891}), .b ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, Midori_rounds_SR_Result[28]}), .c ({DataOut_s2[24], DataOut_s1[24], DataOut_s0[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U79 ( .a ({new_AGEMA_signal_7931, new_AGEMA_signal_7923, new_AGEMA_signal_7915}), .b ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, Midori_rounds_SR_Result[58]}), .c ({DataOut_s2[22], DataOut_s1[22], DataOut_s0[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U77 ( .a ({new_AGEMA_signal_7955, new_AGEMA_signal_7947, new_AGEMA_signal_7939}), .b ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, Midori_rounds_SR_Result[56]}), .c ({DataOut_s2[20], DataOut_s1[20], DataOut_s0[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U74 ( .a ({new_AGEMA_signal_7979, new_AGEMA_signal_7971, new_AGEMA_signal_7963}), .b ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, Midori_rounds_SR_Result[38]}), .c ({DataOut_s2[18], DataOut_s1[18], DataOut_s0[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U72 ( .a ({new_AGEMA_signal_8003, new_AGEMA_signal_7995, new_AGEMA_signal_7987}), .b ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, Midori_rounds_SR_Result[36]}), .c ({DataOut_s2[16], DataOut_s1[16], DataOut_s0[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U70 ( .a ({new_AGEMA_signal_8027, new_AGEMA_signal_8019, new_AGEMA_signal_8011}), .b ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, Midori_rounds_SR_Result[22]}), .c ({DataOut_s2[14], DataOut_s1[14], DataOut_s0[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U68 ( .a ({new_AGEMA_signal_8051, new_AGEMA_signal_8043, new_AGEMA_signal_8035}), .b ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, Midori_rounds_SR_Result[20]}), .c ({DataOut_s2[12], DataOut_s1[12], DataOut_s0[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U66 ( .a ({new_AGEMA_signal_8075, new_AGEMA_signal_8067, new_AGEMA_signal_8059}), .b ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, Midori_rounds_SR_Result[10]}), .c ({DataOut_s2[10], DataOut_s1[10], DataOut_s0[10]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_U65 ( .a ({new_AGEMA_signal_8099, new_AGEMA_signal_8091, new_AGEMA_signal_8083}), .b ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, Midori_rounds_SR_Result[48]}), .c ({DataOut_s2[0], DataOut_s1[0], DataOut_s0[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U143 ( .a ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, Midori_rounds_SR_Result[8]}), .b ({new_AGEMA_signal_8123, new_AGEMA_signal_8115, new_AGEMA_signal_8107}), .c ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, Midori_rounds_sub_ResultXORkey[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U141 ( .a ({new_AGEMA_signal_8147, new_AGEMA_signal_8139, new_AGEMA_signal_8131}), .b ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, Midori_rounds_SR_Result[46]}), .c ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, Midori_rounds_sub_ResultXORkey[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U139 ( .a ({new_AGEMA_signal_8171, new_AGEMA_signal_8163, new_AGEMA_signal_8155}), .b ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, Midori_rounds_SR_Result[62]}), .c ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, Midori_rounds_sub_ResultXORkey[62]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U137 ( .a ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, Midori_rounds_SR_Result[60]}), .b ({new_AGEMA_signal_8195, new_AGEMA_signal_8187, new_AGEMA_signal_8179}), .c ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, Midori_rounds_sub_ResultXORkey[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U134 ( .a ({new_AGEMA_signal_8219, new_AGEMA_signal_8211, new_AGEMA_signal_8203}), .b ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, Midori_rounds_SR_Result[34]}), .c ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, Midori_rounds_sub_ResultXORkey[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U132 ( .a ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, Midori_rounds_SR_Result[32]}), .b ({new_AGEMA_signal_8243, new_AGEMA_signal_8235, new_AGEMA_signal_8227}), .c ({new_AGEMA_signal_3655, new_AGEMA_signal_3654, Midori_rounds_sub_ResultXORkey[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U130 ( .a ({new_AGEMA_signal_8267, new_AGEMA_signal_8259, new_AGEMA_signal_8251}), .b ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, Midori_rounds_SR_Result[6]}), .c ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, Midori_rounds_sub_ResultXORkey[54]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U128 ( .a ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, Midori_rounds_SR_Result[4]}), .b ({new_AGEMA_signal_8291, new_AGEMA_signal_8283, new_AGEMA_signal_8275}), .c ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, Midori_rounds_sub_ResultXORkey[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U126 ( .a ({new_AGEMA_signal_8315, new_AGEMA_signal_8307, new_AGEMA_signal_8299}), .b ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, Midori_rounds_SR_Result[26]}), .c ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, Midori_rounds_sub_ResultXORkey[50]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U125 ( .a ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, Midori_rounds_SR_Result[44]}), .b ({new_AGEMA_signal_8339, new_AGEMA_signal_8331, new_AGEMA_signal_8323}), .c ({new_AGEMA_signal_3659, new_AGEMA_signal_3658, Midori_rounds_sub_ResultXORkey[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U123 ( .a ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, Midori_rounds_SR_Result[24]}), .b ({new_AGEMA_signal_8363, new_AGEMA_signal_8355, new_AGEMA_signal_8347}), .c ({new_AGEMA_signal_3803, new_AGEMA_signal_3802, Midori_rounds_sub_ResultXORkey[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U121 ( .a ({new_AGEMA_signal_8387, new_AGEMA_signal_8379, new_AGEMA_signal_8371}), .b ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, Midori_rounds_SR_Result[42]}), .c ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, Midori_rounds_sub_ResultXORkey[46]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U119 ( .a ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, Midori_rounds_SR_Result[40]}), .b ({new_AGEMA_signal_8411, new_AGEMA_signal_8403, new_AGEMA_signal_8395}), .c ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, Midori_rounds_sub_ResultXORkey[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U117 ( .a ({new_AGEMA_signal_8435, new_AGEMA_signal_8427, new_AGEMA_signal_8419}), .b ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, Midori_rounds_SR_Result[54]}), .c ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, Midori_rounds_sub_ResultXORkey[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U115 ( .a ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, Midori_rounds_SR_Result[52]}), .b ({new_AGEMA_signal_8459, new_AGEMA_signal_8451, new_AGEMA_signal_8443}), .c ({new_AGEMA_signal_3661, new_AGEMA_signal_3660, Midori_rounds_sub_ResultXORkey[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U112 ( .a ({new_AGEMA_signal_8483, new_AGEMA_signal_8475, new_AGEMA_signal_8467}), .b ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, Midori_rounds_SR_Result[18]}), .c ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, Midori_rounds_sub_ResultXORkey[38]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U110 ( .a ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, Midori_rounds_SR_Result[16]}), .b ({new_AGEMA_signal_8507, new_AGEMA_signal_8499, new_AGEMA_signal_8491}), .c ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, Midori_rounds_sub_ResultXORkey[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U108 ( .a ({new_AGEMA_signal_8531, new_AGEMA_signal_8523, new_AGEMA_signal_8515}), .b ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, Midori_rounds_SR_Result[14]}), .c ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, Midori_rounds_sub_ResultXORkey[34]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U106 ( .a ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, Midori_rounds_SR_Result[12]}), .b ({new_AGEMA_signal_8555, new_AGEMA_signal_8547, new_AGEMA_signal_8539}), .c ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, Midori_rounds_sub_ResultXORkey[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U104 ( .a ({new_AGEMA_signal_8579, new_AGEMA_signal_8571, new_AGEMA_signal_8563}), .b ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, Midori_rounds_SR_Result[2]}), .c ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, Midori_rounds_sub_ResultXORkey[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U103 ( .a ({new_AGEMA_signal_8603, new_AGEMA_signal_8595, new_AGEMA_signal_8587}), .b ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, Midori_rounds_SR_Result[50]}), .c ({new_AGEMA_signal_3151, new_AGEMA_signal_3150, Midori_rounds_sub_ResultXORkey[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U101 ( .a ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, Midori_rounds_SR_Result[0]}), .b ({new_AGEMA_signal_8627, new_AGEMA_signal_8619, new_AGEMA_signal_8611}), .c ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, Midori_rounds_sub_ResultXORkey[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U99 ( .a ({new_AGEMA_signal_8651, new_AGEMA_signal_8643, new_AGEMA_signal_8635}), .b ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, Midori_rounds_SR_Result[30]}), .c ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, Midori_rounds_sub_ResultXORkey[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U97 ( .a ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, Midori_rounds_SR_Result[28]}), .b ({new_AGEMA_signal_8675, new_AGEMA_signal_8667, new_AGEMA_signal_8659}), .c ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, Midori_rounds_sub_ResultXORkey[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U95 ( .a ({new_AGEMA_signal_8699, new_AGEMA_signal_8691, new_AGEMA_signal_8683}), .b ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, Midori_rounds_SR_Result[58]}), .c ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, Midori_rounds_sub_ResultXORkey[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U93 ( .a ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, Midori_rounds_SR_Result[56]}), .b ({new_AGEMA_signal_8723, new_AGEMA_signal_8715, new_AGEMA_signal_8707}), .c ({new_AGEMA_signal_3535, new_AGEMA_signal_3534, Midori_rounds_sub_ResultXORkey[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U90 ( .a ({new_AGEMA_signal_8747, new_AGEMA_signal_8739, new_AGEMA_signal_8731}), .b ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, Midori_rounds_SR_Result[38]}), .c ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, Midori_rounds_sub_ResultXORkey[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U88 ( .a ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, Midori_rounds_SR_Result[36]}), .b ({new_AGEMA_signal_8771, new_AGEMA_signal_8763, new_AGEMA_signal_8755}), .c ({new_AGEMA_signal_3667, new_AGEMA_signal_3666, Midori_rounds_sub_ResultXORkey[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U86 ( .a ({new_AGEMA_signal_8795, new_AGEMA_signal_8787, new_AGEMA_signal_8779}), .b ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, Midori_rounds_SR_Result[22]}), .c ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, Midori_rounds_sub_ResultXORkey[14]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U84 ( .a ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, Midori_rounds_SR_Result[20]}), .b ({new_AGEMA_signal_8819, new_AGEMA_signal_8811, new_AGEMA_signal_8803}), .c ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, Midori_rounds_sub_ResultXORkey[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U82 ( .a ({new_AGEMA_signal_8843, new_AGEMA_signal_8835, new_AGEMA_signal_8827}), .b ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, Midori_rounds_SR_Result[10]}), .c ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, Midori_rounds_sub_ResultXORkey[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U81 ( .a ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, Midori_rounds_SR_Result[48]}), .b ({new_AGEMA_signal_8867, new_AGEMA_signal_8859, new_AGEMA_signal_8851}), .c ({new_AGEMA_signal_3671, new_AGEMA_signal_3670, Midori_rounds_sub_ResultXORkey[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U79 ( .a ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, Midori_rounds_SR_Inv_Result[8]}), .b ({new_AGEMA_signal_8123, new_AGEMA_signal_8115, new_AGEMA_signal_8107}), .c ({new_AGEMA_signal_3845, new_AGEMA_signal_3844, Midori_rounds_mul_ResultXORkey[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U76 ( .a ({new_AGEMA_signal_8147, new_AGEMA_signal_8139, new_AGEMA_signal_8131}), .b ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, Midori_rounds_SR_Inv_Result[54]}), .c ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, Midori_rounds_mul_ResultXORkey[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U74 ( .a ({new_AGEMA_signal_8171, new_AGEMA_signal_8163, new_AGEMA_signal_8155}), .b ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, Midori_rounds_SR_Inv_Result[62]}), .c ({new_AGEMA_signal_3435, new_AGEMA_signal_3434, Midori_rounds_mul_ResultXORkey[62]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U72 ( .a ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, Midori_rounds_SR_Inv_Result[60]}), .b ({new_AGEMA_signal_8195, new_AGEMA_signal_8187, new_AGEMA_signal_8179}), .c ({new_AGEMA_signal_3907, new_AGEMA_signal_3906, Midori_rounds_mul_ResultXORkey[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U68 ( .a ({new_AGEMA_signal_8219, new_AGEMA_signal_8211, new_AGEMA_signal_8203}), .b ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, Midori_rounds_SR_Inv_Result[22]}), .c ({new_AGEMA_signal_3443, new_AGEMA_signal_3442, Midori_rounds_mul_ResultXORkey[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U66 ( .a ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, Midori_rounds_SR_Inv_Result[20]}), .b ({new_AGEMA_signal_8243, new_AGEMA_signal_8235, new_AGEMA_signal_8227}), .c ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, Midori_rounds_mul_ResultXORkey[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U63 ( .a ({new_AGEMA_signal_8267, new_AGEMA_signal_8259, new_AGEMA_signal_8251}), .b ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, Midori_rounds_SR_Inv_Result[42]}), .c ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, Midori_rounds_mul_ResultXORkey[54]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U61 ( .a ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, Midori_rounds_SR_Inv_Result[40]}), .b ({new_AGEMA_signal_8291, new_AGEMA_signal_8283, new_AGEMA_signal_8275}), .c ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, Midori_rounds_mul_ResultXORkey[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U58 ( .a ({new_AGEMA_signal_8315, new_AGEMA_signal_8307, new_AGEMA_signal_8299}), .b ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, Midori_rounds_SR_Inv_Result[2]}), .c ({new_AGEMA_signal_3455, new_AGEMA_signal_3454, Midori_rounds_mul_ResultXORkey[50]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U57 ( .a ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, Midori_rounds_SR_Inv_Result[52]}), .b ({new_AGEMA_signal_8339, new_AGEMA_signal_8331, new_AGEMA_signal_8323}), .c ({new_AGEMA_signal_3847, new_AGEMA_signal_3846, Midori_rounds_mul_ResultXORkey[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U54 ( .a ({new_AGEMA_signal_3821, new_AGEMA_signal_3820, Midori_rounds_SR_Inv_Result[0]}), .b ({new_AGEMA_signal_8363, new_AGEMA_signal_8355, new_AGEMA_signal_8347}), .c ({new_AGEMA_signal_3849, new_AGEMA_signal_3848, Midori_rounds_mul_ResultXORkey[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U51 ( .a ({new_AGEMA_signal_8387, new_AGEMA_signal_8379, new_AGEMA_signal_8371}), .b ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, Midori_rounds_SR_Inv_Result[6]}), .c ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, Midori_rounds_mul_ResultXORkey[46]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U49 ( .a ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, Midori_rounds_SR_Inv_Result[4]}), .b ({new_AGEMA_signal_8411, new_AGEMA_signal_8403, new_AGEMA_signal_8395}), .c ({new_AGEMA_signal_3851, new_AGEMA_signal_3850, Midori_rounds_mul_ResultXORkey[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U46 ( .a ({new_AGEMA_signal_8435, new_AGEMA_signal_8427, new_AGEMA_signal_8419}), .b ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, Midori_rounds_SR_Inv_Result[46]}), .c ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, Midori_rounds_mul_ResultXORkey[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U44 ( .a ({new_AGEMA_signal_3823, new_AGEMA_signal_3822, Midori_rounds_SR_Inv_Result[44]}), .b ({new_AGEMA_signal_8459, new_AGEMA_signal_8451, new_AGEMA_signal_8443}), .c ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, Midori_rounds_mul_ResultXORkey[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U40 ( .a ({new_AGEMA_signal_8483, new_AGEMA_signal_8475, new_AGEMA_signal_8467}), .b ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, Midori_rounds_SR_Inv_Result[18]}), .c ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, Midori_rounds_mul_ResultXORkey[38]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U38 ( .a ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, Midori_rounds_SR_Inv_Result[16]}), .b ({new_AGEMA_signal_8507, new_AGEMA_signal_8499, new_AGEMA_signal_8491}), .c ({new_AGEMA_signal_3855, new_AGEMA_signal_3854, Midori_rounds_mul_ResultXORkey[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U35 ( .a ({new_AGEMA_signal_8531, new_AGEMA_signal_8523, new_AGEMA_signal_8515}), .b ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, Midori_rounds_SR_Inv_Result[58]}), .c ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, Midori_rounds_mul_ResultXORkey[34]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U33 ( .a ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, Midori_rounds_SR_Inv_Result[56]}), .b ({new_AGEMA_signal_8555, new_AGEMA_signal_8547, new_AGEMA_signal_8539}), .c ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, Midori_rounds_mul_ResultXORkey[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U30 ( .a ({new_AGEMA_signal_8579, new_AGEMA_signal_8571, new_AGEMA_signal_8563}), .b ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, Midori_rounds_SR_Inv_Result[26]}), .c ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, Midori_rounds_mul_ResultXORkey[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U29 ( .a ({new_AGEMA_signal_8603, new_AGEMA_signal_8595, new_AGEMA_signal_8587}), .b ({new_AGEMA_signal_3411, new_AGEMA_signal_3410, Midori_rounds_SR_Inv_Result[30]}), .c ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, Midori_rounds_mul_ResultXORkey[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U27 ( .a ({new_AGEMA_signal_3833, new_AGEMA_signal_3832, Midori_rounds_SR_Inv_Result[24]}), .b ({new_AGEMA_signal_8627, new_AGEMA_signal_8619, new_AGEMA_signal_8611}), .c ({new_AGEMA_signal_3859, new_AGEMA_signal_3858, Midori_rounds_mul_ResultXORkey[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U24 ( .a ({new_AGEMA_signal_8651, new_AGEMA_signal_8643, new_AGEMA_signal_8635}), .b ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, Midori_rounds_SR_Inv_Result[50]}), .c ({new_AGEMA_signal_3499, new_AGEMA_signal_3498, Midori_rounds_mul_ResultXORkey[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U22 ( .a ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, Midori_rounds_SR_Inv_Result[48]}), .b ({new_AGEMA_signal_8675, new_AGEMA_signal_8667, new_AGEMA_signal_8659}), .c ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, Midori_rounds_mul_ResultXORkey[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U19 ( .a ({new_AGEMA_signal_8699, new_AGEMA_signal_8691, new_AGEMA_signal_8683}), .b ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, Midori_rounds_SR_Inv_Result[14]}), .c ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, Midori_rounds_mul_ResultXORkey[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U17 ( .a ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, Midori_rounds_SR_Inv_Result[12]}), .b ({new_AGEMA_signal_8723, new_AGEMA_signal_8715, new_AGEMA_signal_8707}), .c ({new_AGEMA_signal_3877, new_AGEMA_signal_3876, Midori_rounds_mul_ResultXORkey[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U13 ( .a ({new_AGEMA_signal_8747, new_AGEMA_signal_8739, new_AGEMA_signal_8731}), .b ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, Midori_rounds_SR_Inv_Result[38]}), .c ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, Midori_rounds_mul_ResultXORkey[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U11 ( .a ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, Midori_rounds_SR_Inv_Result[36]}), .b ({new_AGEMA_signal_8771, new_AGEMA_signal_8763, new_AGEMA_signal_8755}), .c ({new_AGEMA_signal_3879, new_AGEMA_signal_3878, Midori_rounds_mul_ResultXORkey[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U8 ( .a ({new_AGEMA_signal_8795, new_AGEMA_signal_8787, new_AGEMA_signal_8779}), .b ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, Midori_rounds_SR_Inv_Result[34]}), .c ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, Midori_rounds_mul_ResultXORkey[14]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U6 ( .a ({new_AGEMA_signal_3841, new_AGEMA_signal_3840, Midori_rounds_SR_Inv_Result[32]}), .b ({new_AGEMA_signal_8819, new_AGEMA_signal_8811, new_AGEMA_signal_8803}), .c ({new_AGEMA_signal_3863, new_AGEMA_signal_3862, Midori_rounds_mul_ResultXORkey[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U3 ( .a ({new_AGEMA_signal_8843, new_AGEMA_signal_8835, new_AGEMA_signal_8827}), .b ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, Midori_rounds_SR_Inv_Result[10]}), .c ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, Midori_rounds_mul_ResultXORkey[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_U2 ( .a ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, Midori_rounds_SR_Inv_Result[28]}), .b ({new_AGEMA_signal_8867, new_AGEMA_signal_8859, new_AGEMA_signal_8851}), .c ({new_AGEMA_signal_3865, new_AGEMA_signal_3864, Midori_rounds_mul_ResultXORkey[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, Midori_rounds_round_Result[0]}), .a ({new_AGEMA_signal_8893, new_AGEMA_signal_8885, new_AGEMA_signal_8877}), .c ({new_AGEMA_signal_3911, new_AGEMA_signal_3910, Midori_rounds_roundResult_Reg_SFF_0_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3559, new_AGEMA_signal_3558, Midori_rounds_round_Result[2]}), .a ({new_AGEMA_signal_8917, new_AGEMA_signal_8909, new_AGEMA_signal_8901}), .c ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, Midori_rounds_roundResult_Reg_SFF_2_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3887, new_AGEMA_signal_3886, Midori_rounds_round_Result[4]}), .a ({new_AGEMA_signal_8941, new_AGEMA_signal_8933, new_AGEMA_signal_8925}), .c ({new_AGEMA_signal_3913, new_AGEMA_signal_3912, Midori_rounds_roundResult_Reg_SFF_4_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, Midori_rounds_round_Result[6]}), .a ({new_AGEMA_signal_8965, new_AGEMA_signal_8957, new_AGEMA_signal_8949}), .c ({new_AGEMA_signal_3683, new_AGEMA_signal_3682, Midori_rounds_roundResult_Reg_SFF_6_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3889, new_AGEMA_signal_3888, Midori_rounds_round_Result[8]}), .a ({new_AGEMA_signal_8989, new_AGEMA_signal_8981, new_AGEMA_signal_8973}), .c ({new_AGEMA_signal_3915, new_AGEMA_signal_3914, Midori_rounds_roundResult_Reg_SFF_8_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3571, new_AGEMA_signal_3570, Midori_rounds_round_Result[10]}), .a ({new_AGEMA_signal_9013, new_AGEMA_signal_9005, new_AGEMA_signal_8997}), .c ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, Midori_rounds_roundResult_Reg_SFF_10_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, Midori_rounds_round_Result[12]}), .a ({new_AGEMA_signal_9037, new_AGEMA_signal_9029, new_AGEMA_signal_9021}), .c ({new_AGEMA_signal_3917, new_AGEMA_signal_3916, Midori_rounds_roundResult_Reg_SFF_12_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, Midori_rounds_round_Result[14]}), .a ({new_AGEMA_signal_9061, new_AGEMA_signal_9053, new_AGEMA_signal_9045}), .c ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, Midori_rounds_roundResult_Reg_SFF_14_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3933, new_AGEMA_signal_3932, Midori_rounds_round_Result[16]}), .a ({new_AGEMA_signal_9085, new_AGEMA_signal_9077, new_AGEMA_signal_9069}), .c ({new_AGEMA_signal_3939, new_AGEMA_signal_3938, Midori_rounds_roundResult_Reg_SFF_16_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, Midori_rounds_round_Result[18]}), .a ({new_AGEMA_signal_9109, new_AGEMA_signal_9101, new_AGEMA_signal_9093}), .c ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, Midori_rounds_roundResult_Reg_SFF_18_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3935, new_AGEMA_signal_3934, Midori_rounds_round_Result[20]}), .a ({new_AGEMA_signal_9133, new_AGEMA_signal_9125, new_AGEMA_signal_9117}), .c ({new_AGEMA_signal_3941, new_AGEMA_signal_3940, Midori_rounds_roundResult_Reg_SFF_20_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, Midori_rounds_round_Result[22]}), .a ({new_AGEMA_signal_9157, new_AGEMA_signal_9149, new_AGEMA_signal_9141}), .c ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, Midori_rounds_roundResult_Reg_SFF_22_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, Midori_rounds_round_Result[24]}), .a ({new_AGEMA_signal_9181, new_AGEMA_signal_9173, new_AGEMA_signal_9165}), .c ({new_AGEMA_signal_3919, new_AGEMA_signal_3918, Midori_rounds_roundResult_Reg_SFF_24_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3595, new_AGEMA_signal_3594, Midori_rounds_round_Result[26]}), .a ({new_AGEMA_signal_9205, new_AGEMA_signal_9197, new_AGEMA_signal_9189}), .c ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, Midori_rounds_roundResult_Reg_SFF_26_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3895, new_AGEMA_signal_3894, Midori_rounds_round_Result[28]}), .a ({new_AGEMA_signal_9229, new_AGEMA_signal_9221, new_AGEMA_signal_9213}), .c ({new_AGEMA_signal_3921, new_AGEMA_signal_3920, Midori_rounds_roundResult_Reg_SFF_28_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, Midori_rounds_round_Result[30]}), .a ({new_AGEMA_signal_9253, new_AGEMA_signal_9245, new_AGEMA_signal_9237}), .c ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, Midori_rounds_roundResult_Reg_SFF_30_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, Midori_rounds_round_Result[32]}), .a ({new_AGEMA_signal_9277, new_AGEMA_signal_9269, new_AGEMA_signal_9261}), .c ({new_AGEMA_signal_3923, new_AGEMA_signal_3922, Midori_rounds_roundResult_Reg_SFF_32_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3607, new_AGEMA_signal_3606, Midori_rounds_round_Result[34]}), .a ({new_AGEMA_signal_9301, new_AGEMA_signal_9293, new_AGEMA_signal_9285}), .c ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, Midori_rounds_roundResult_Reg_SFF_34_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3899, new_AGEMA_signal_3898, Midori_rounds_round_Result[36]}), .a ({new_AGEMA_signal_9325, new_AGEMA_signal_9317, new_AGEMA_signal_9309}), .c ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, Midori_rounds_roundResult_Reg_SFF_36_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, Midori_rounds_round_Result[38]}), .a ({new_AGEMA_signal_9349, new_AGEMA_signal_9341, new_AGEMA_signal_9333}), .c ({new_AGEMA_signal_3731, new_AGEMA_signal_3730, Midori_rounds_roundResult_Reg_SFF_38_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3901, new_AGEMA_signal_3900, Midori_rounds_round_Result[40]}), .a ({new_AGEMA_signal_9373, new_AGEMA_signal_9365, new_AGEMA_signal_9357}), .c ({new_AGEMA_signal_3927, new_AGEMA_signal_3926, Midori_rounds_roundResult_Reg_SFF_40_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3619, new_AGEMA_signal_3618, Midori_rounds_round_Result[42]}), .a ({new_AGEMA_signal_9397, new_AGEMA_signal_9389, new_AGEMA_signal_9381}), .c ({new_AGEMA_signal_3737, new_AGEMA_signal_3736, Midori_rounds_roundResult_Reg_SFF_42_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3903, new_AGEMA_signal_3902, Midori_rounds_round_Result[44]}), .a ({new_AGEMA_signal_9421, new_AGEMA_signal_9413, new_AGEMA_signal_9405}), .c ({new_AGEMA_signal_3929, new_AGEMA_signal_3928, Midori_rounds_roundResult_Reg_SFF_44_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3625, new_AGEMA_signal_3624, Midori_rounds_round_Result[46]}), .a ({new_AGEMA_signal_9445, new_AGEMA_signal_9437, new_AGEMA_signal_9429}), .c ({new_AGEMA_signal_3743, new_AGEMA_signal_3742, Midori_rounds_roundResult_Reg_SFF_46_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, Midori_rounds_round_Result[48]}), .a ({new_AGEMA_signal_9469, new_AGEMA_signal_9461, new_AGEMA_signal_9453}), .c ({new_AGEMA_signal_3931, new_AGEMA_signal_3930, Midori_rounds_roundResult_Reg_SFF_48_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3631, new_AGEMA_signal_3630, Midori_rounds_round_Result[50]}), .a ({new_AGEMA_signal_9493, new_AGEMA_signal_9485, new_AGEMA_signal_9477}), .c ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, Midori_rounds_roundResult_Reg_SFF_50_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3937, new_AGEMA_signal_3936, Midori_rounds_round_Result[52]}), .a ({new_AGEMA_signal_9517, new_AGEMA_signal_9509, new_AGEMA_signal_9501}), .c ({new_AGEMA_signal_3943, new_AGEMA_signal_3942, Midori_rounds_roundResult_Reg_SFF_52_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, Midori_rounds_round_Result[54]}), .a ({new_AGEMA_signal_9541, new_AGEMA_signal_9533, new_AGEMA_signal_9525}), .c ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, Midori_rounds_roundResult_Reg_SFF_54_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, Midori_rounds_round_Result[56]}), .a ({new_AGEMA_signal_9565, new_AGEMA_signal_9557, new_AGEMA_signal_9549}), .c ({new_AGEMA_signal_3949, new_AGEMA_signal_3948, Midori_rounds_roundResult_Reg_SFF_56_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3643, new_AGEMA_signal_3642, Midori_rounds_round_Result[58]}), .a ({new_AGEMA_signal_9589, new_AGEMA_signal_9581, new_AGEMA_signal_9573}), .c ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, Midori_rounds_roundResult_Reg_SFF_58_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3947, new_AGEMA_signal_3946, Midori_rounds_round_Result[60]}), .a ({new_AGEMA_signal_9613, new_AGEMA_signal_9605, new_AGEMA_signal_9597}), .c ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, Midori_rounds_roundResult_Reg_SFF_60_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1 ( .s (new_AGEMA_signal_8869), .b ({new_AGEMA_signal_3649, new_AGEMA_signal_3648, Midori_rounds_round_Result[62]}), .a ({new_AGEMA_signal_9637, new_AGEMA_signal_9629, new_AGEMA_signal_9621}), .c ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, Midori_rounds_roundResult_Reg_SFF_62_DQ}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U17 ( .a ({new_AGEMA_signal_9643, new_AGEMA_signal_9641, new_AGEMA_signal_9639}), .b ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, Midori_rounds_sub_sBox_PRINCE_0_n12}), .clk (clk), .r ({Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, Midori_rounds_SR_Result[50]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U8 ( .a ({new_AGEMA_signal_9655, new_AGEMA_signal_9651, new_AGEMA_signal_9647}), .b ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, Midori_rounds_sub_sBox_PRINCE_0_n3}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675]}), .c ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, Midori_rounds_SR_Result[48]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U17 ( .a ({new_AGEMA_signal_9661, new_AGEMA_signal_9659, new_AGEMA_signal_9657}), .b ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, Midori_rounds_sub_sBox_PRINCE_1_n12}), .clk (clk), .r ({Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, Midori_rounds_SR_Result[46]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U8 ( .a ({new_AGEMA_signal_9673, new_AGEMA_signal_9669, new_AGEMA_signal_9665}), .b ({new_AGEMA_signal_2691, new_AGEMA_signal_2690, Midori_rounds_sub_sBox_PRINCE_1_n3}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681]}), .c ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, Midori_rounds_SR_Result[44]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U17 ( .a ({new_AGEMA_signal_9679, new_AGEMA_signal_9677, new_AGEMA_signal_9675}), .b ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, Midori_rounds_sub_sBox_PRINCE_2_n12}), .clk (clk), .r ({Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, Midori_rounds_SR_Result[10]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U8 ( .a ({new_AGEMA_signal_9691, new_AGEMA_signal_9687, new_AGEMA_signal_9683}), .b ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, Midori_rounds_sub_sBox_PRINCE_2_n3}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687]}), .c ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, Midori_rounds_SR_Result[8]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U17 ( .a ({new_AGEMA_signal_9697, new_AGEMA_signal_9695, new_AGEMA_signal_9693}), .b ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, Midori_rounds_sub_sBox_PRINCE_3_n12}), .clk (clk), .r ({Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, Midori_rounds_SR_Result[22]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U8 ( .a ({new_AGEMA_signal_9709, new_AGEMA_signal_9705, new_AGEMA_signal_9701}), .b ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, Midori_rounds_sub_sBox_PRINCE_3_n3}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693]}), .c ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, Midori_rounds_SR_Result[20]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U17 ( .a ({new_AGEMA_signal_9715, new_AGEMA_signal_9713, new_AGEMA_signal_9711}), .b ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, Midori_rounds_sub_sBox_PRINCE_4_n12}), .clk (clk), .r ({Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, Midori_rounds_SR_Result[38]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U8 ( .a ({new_AGEMA_signal_9727, new_AGEMA_signal_9723, new_AGEMA_signal_9719}), .b ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, Midori_rounds_sub_sBox_PRINCE_4_n3}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699]}), .c ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, Midori_rounds_SR_Result[36]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U17 ( .a ({new_AGEMA_signal_9733, new_AGEMA_signal_9731, new_AGEMA_signal_9729}), .b ({new_AGEMA_signal_2727, new_AGEMA_signal_2726, Midori_rounds_sub_sBox_PRINCE_5_n12}), .clk (clk), .r ({Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, Midori_rounds_SR_Result[58]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U8 ( .a ({new_AGEMA_signal_9745, new_AGEMA_signal_9741, new_AGEMA_signal_9737}), .b ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, Midori_rounds_sub_sBox_PRINCE_5_n3}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705]}), .c ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, Midori_rounds_SR_Result[56]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U17 ( .a ({new_AGEMA_signal_9751, new_AGEMA_signal_9749, new_AGEMA_signal_9747}), .b ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, Midori_rounds_sub_sBox_PRINCE_6_n12}), .clk (clk), .r ({Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, Midori_rounds_SR_Result[30]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U8 ( .a ({new_AGEMA_signal_9763, new_AGEMA_signal_9759, new_AGEMA_signal_9755}), .b ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, Midori_rounds_sub_sBox_PRINCE_6_n3}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711]}), .c ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, Midori_rounds_SR_Result[28]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U17 ( .a ({new_AGEMA_signal_9769, new_AGEMA_signal_9767, new_AGEMA_signal_9765}), .b ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, Midori_rounds_sub_sBox_PRINCE_7_n12}), .clk (clk), .r ({Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, Midori_rounds_SR_Result[2]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U8 ( .a ({new_AGEMA_signal_9781, new_AGEMA_signal_9777, new_AGEMA_signal_9773}), .b ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, Midori_rounds_sub_sBox_PRINCE_7_n3}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717]}), .c ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, Midori_rounds_SR_Result[0]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U17 ( .a ({new_AGEMA_signal_9787, new_AGEMA_signal_9785, new_AGEMA_signal_9783}), .b ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, Midori_rounds_sub_sBox_PRINCE_8_n12}), .clk (clk), .r ({Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, Midori_rounds_SR_Result[14]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U8 ( .a ({new_AGEMA_signal_9799, new_AGEMA_signal_9795, new_AGEMA_signal_9791}), .b ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, Midori_rounds_sub_sBox_PRINCE_8_n3}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723]}), .c ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, Midori_rounds_SR_Result[12]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U17 ( .a ({new_AGEMA_signal_9805, new_AGEMA_signal_9803, new_AGEMA_signal_9801}), .b ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, Midori_rounds_sub_sBox_PRINCE_9_n12}), .clk (clk), .r ({Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, Midori_rounds_SR_Result[18]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U8 ( .a ({new_AGEMA_signal_9817, new_AGEMA_signal_9813, new_AGEMA_signal_9809}), .b ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, Midori_rounds_sub_sBox_PRINCE_9_n3}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729]}), .c ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, Midori_rounds_SR_Result[16]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U17 ( .a ({new_AGEMA_signal_9823, new_AGEMA_signal_9821, new_AGEMA_signal_9819}), .b ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, Midori_rounds_sub_sBox_PRINCE_10_n12}), .clk (clk), .r ({Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, Midori_rounds_SR_Result[54]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U8 ( .a ({new_AGEMA_signal_9835, new_AGEMA_signal_9831, new_AGEMA_signal_9827}), .b ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, Midori_rounds_sub_sBox_PRINCE_10_n3}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735]}), .c ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, Midori_rounds_SR_Result[52]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U17 ( .a ({new_AGEMA_signal_9841, new_AGEMA_signal_9839, new_AGEMA_signal_9837}), .b ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, Midori_rounds_sub_sBox_PRINCE_11_n12}), .clk (clk), .r ({Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, Midori_rounds_SR_Result[42]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U8 ( .a ({new_AGEMA_signal_9853, new_AGEMA_signal_9849, new_AGEMA_signal_9845}), .b ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, Midori_rounds_sub_sBox_PRINCE_11_n3}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741]}), .c ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, Midori_rounds_SR_Result[40]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U17 ( .a ({new_AGEMA_signal_9859, new_AGEMA_signal_9857, new_AGEMA_signal_9855}), .b ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, Midori_rounds_sub_sBox_PRINCE_12_n12}), .clk (clk), .r ({Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, Midori_rounds_SR_Result[26]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U8 ( .a ({new_AGEMA_signal_9871, new_AGEMA_signal_9867, new_AGEMA_signal_9863}), .b ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, Midori_rounds_sub_sBox_PRINCE_12_n3}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747]}), .c ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, Midori_rounds_SR_Result[24]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U17 ( .a ({new_AGEMA_signal_9877, new_AGEMA_signal_9875, new_AGEMA_signal_9873}), .b ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, Midori_rounds_sub_sBox_PRINCE_13_n12}), .clk (clk), .r ({Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, Midori_rounds_SR_Result[6]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U8 ( .a ({new_AGEMA_signal_9889, new_AGEMA_signal_9885, new_AGEMA_signal_9881}), .b ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, Midori_rounds_sub_sBox_PRINCE_13_n3}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753]}), .c ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, Midori_rounds_SR_Result[4]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U17 ( .a ({new_AGEMA_signal_9895, new_AGEMA_signal_9893, new_AGEMA_signal_9891}), .b ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, Midori_rounds_sub_sBox_PRINCE_14_n12}), .clk (clk), .r ({Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, Midori_rounds_SR_Result[34]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U8 ( .a ({new_AGEMA_signal_9907, new_AGEMA_signal_9903, new_AGEMA_signal_9899}), .b ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, Midori_rounds_sub_sBox_PRINCE_14_n3}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759]}), .c ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, Midori_rounds_SR_Result[32]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U17 ( .a ({new_AGEMA_signal_9913, new_AGEMA_signal_9911, new_AGEMA_signal_9909}), .b ({new_AGEMA_signal_2827, new_AGEMA_signal_2826, Midori_rounds_sub_sBox_PRINCE_15_n12}), .clk (clk), .r ({Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, Midori_rounds_SR_Result[62]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U8 ( .a ({new_AGEMA_signal_9925, new_AGEMA_signal_9921, new_AGEMA_signal_9917}), .b ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, Midori_rounds_sub_sBox_PRINCE_15_n3}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765]}), .c ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, Midori_rounds_SR_Result[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_0_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, Midori_rounds_SR_Result[0]}), .a ({new_AGEMA_signal_3671, new_AGEMA_signal_3670, Midori_rounds_sub_ResultXORkey[0]}), .c ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, Midori_rounds_mul_input[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_2_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, Midori_rounds_SR_Result[2]}), .a ({new_AGEMA_signal_3151, new_AGEMA_signal_3150, Midori_rounds_sub_ResultXORkey[2]}), .c ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, Midori_rounds_mul_input[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_4_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, Midori_rounds_SR_Result[4]}), .a ({new_AGEMA_signal_3659, new_AGEMA_signal_3658, Midori_rounds_sub_ResultXORkey[4]}), .c ({new_AGEMA_signal_3785, new_AGEMA_signal_3784, Midori_rounds_mul_input[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_6_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, Midori_rounds_SR_Result[6]}), .a ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, Midori_rounds_sub_ResultXORkey[6]}), .c ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, Midori_rounds_mul_input[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_8_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, Midori_rounds_SR_Result[8]}), .a ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, Midori_rounds_sub_ResultXORkey[8]}), .c ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, Midori_rounds_mul_input[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_10_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, Midori_rounds_SR_Result[10]}), .a ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, Midori_rounds_sub_ResultXORkey[10]}), .c ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, Midori_rounds_mul_input[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_12_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, Midori_rounds_SR_Result[12]}), .a ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, Midori_rounds_sub_ResultXORkey[12]}), .c ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, Midori_rounds_mul_input[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_14_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, Midori_rounds_SR_Result[14]}), .a ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, Midori_rounds_sub_ResultXORkey[14]}), .c ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, Midori_rounds_mul_input[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_16_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, Midori_rounds_SR_Result[16]}), .a ({new_AGEMA_signal_3667, new_AGEMA_signal_3666, Midori_rounds_sub_ResultXORkey[16]}), .c ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, Midori_rounds_mul_input[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_18_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, Midori_rounds_SR_Result[18]}), .a ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, Midori_rounds_sub_ResultXORkey[18]}), .c ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, Midori_rounds_mul_input[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_20_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, Midori_rounds_SR_Result[20]}), .a ({new_AGEMA_signal_3535, new_AGEMA_signal_3534, Midori_rounds_sub_ResultXORkey[20]}), .c ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, Midori_rounds_mul_input[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_22_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, Midori_rounds_SR_Result[22]}), .a ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, Midori_rounds_sub_ResultXORkey[22]}), .c ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, Midori_rounds_mul_input[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_24_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, Midori_rounds_SR_Result[24]}), .a ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, Midori_rounds_sub_ResultXORkey[24]}), .c ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, Midori_rounds_mul_input[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_26_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, Midori_rounds_SR_Result[26]}), .a ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, Midori_rounds_sub_ResultXORkey[26]}), .c ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, Midori_rounds_mul_input[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_28_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, Midori_rounds_SR_Result[28]}), .a ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, Midori_rounds_sub_ResultXORkey[28]}), .c ({new_AGEMA_signal_3805, new_AGEMA_signal_3804, Midori_rounds_mul_input[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_30_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, Midori_rounds_SR_Result[30]}), .a ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, Midori_rounds_sub_ResultXORkey[30]}), .c ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, Midori_rounds_mul_input[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_32_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, Midori_rounds_SR_Result[32]}), .a ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, Midori_rounds_sub_ResultXORkey[32]}), .c ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, Midori_rounds_mul_input[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_34_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, Midori_rounds_SR_Result[34]}), .a ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, Midori_rounds_sub_ResultXORkey[34]}), .c ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, Midori_rounds_mul_input[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_36_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, Midori_rounds_SR_Result[36]}), .a ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, Midori_rounds_sub_ResultXORkey[36]}), .c ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, Midori_rounds_mul_input[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_38_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, Midori_rounds_SR_Result[38]}), .a ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, Midori_rounds_sub_ResultXORkey[38]}), .c ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, Midori_rounds_mul_input[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_40_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, Midori_rounds_SR_Result[40]}), .a ({new_AGEMA_signal_3661, new_AGEMA_signal_3660, Midori_rounds_sub_ResultXORkey[40]}), .c ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, Midori_rounds_mul_input[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_42_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, Midori_rounds_SR_Result[42]}), .a ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, Midori_rounds_sub_ResultXORkey[42]}), .c ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, Midori_rounds_mul_input[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_44_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, Midori_rounds_SR_Result[44]}), .a ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, Midori_rounds_sub_ResultXORkey[44]}), .c ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, Midori_rounds_mul_input[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_46_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, Midori_rounds_SR_Result[46]}), .a ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, Midori_rounds_sub_ResultXORkey[46]}), .c ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, Midori_rounds_mul_input[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_48_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, Midori_rounds_SR_Result[48]}), .a ({new_AGEMA_signal_3803, new_AGEMA_signal_3802, Midori_rounds_sub_ResultXORkey[48]}), .c ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, Midori_rounds_mul_input[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_50_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, Midori_rounds_SR_Result[50]}), .a ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, Midori_rounds_sub_ResultXORkey[50]}), .c ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, Midori_rounds_mul_input[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_52_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, Midori_rounds_SR_Result[52]}), .a ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, Midori_rounds_sub_ResultXORkey[52]}), .c ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, Midori_rounds_mul_input[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_54_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, Midori_rounds_SR_Result[54]}), .a ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, Midori_rounds_sub_ResultXORkey[54]}), .c ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, Midori_rounds_mul_input[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_56_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, Midori_rounds_SR_Result[56]}), .a ({new_AGEMA_signal_3655, new_AGEMA_signal_3654, Midori_rounds_sub_ResultXORkey[56]}), .c ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, Midori_rounds_mul_input[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_58_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, Midori_rounds_SR_Result[58]}), .a ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, Midori_rounds_sub_ResultXORkey[58]}), .c ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, Midori_rounds_mul_input[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_60_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, Midori_rounds_SR_Result[60]}), .a ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, Midori_rounds_sub_ResultXORkey[60]}), .c ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, Midori_rounds_mul_input[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_62_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, Midori_rounds_SR_Result[62]}), .a ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, Midori_rounds_sub_ResultXORkey[62]}), .c ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, Midori_rounds_mul_input[62]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U23 ( .a ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, Midori_rounds_mul_input[60]}), .b ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, Midori_rounds_mul_MC1_n7}), .c ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, Midori_rounds_SR_Inv_Result[20]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U21 ( .a ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, Midori_rounds_mul_input[50]}), .b ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, Midori_rounds_mul_MC1_n5}), .c ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, Midori_rounds_SR_Inv_Result[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U19 ( .a ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, Midori_rounds_mul_input[48]}), .b ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, Midori_rounds_mul_MC1_n3}), .c ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, Midori_rounds_SR_Inv_Result[40]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U16 ( .a ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, Midori_rounds_mul_input[54]}), .b ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, Midori_rounds_mul_MC1_n5}), .c ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, Midori_rounds_SR_Inv_Result[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U15 ( .a ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, Midori_rounds_mul_input[62]}), .b ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, Midori_rounds_mul_input[58]}), .c ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, Midori_rounds_mul_MC1_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U11 ( .a ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, Midori_rounds_mul_input[58]}), .b ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, Midori_rounds_mul_MC1_n1}), .c ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, Midori_rounds_SR_Inv_Result[62]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U8 ( .a ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, Midori_rounds_mul_input[56]}), .b ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, Midori_rounds_mul_MC1_n7}), .c ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, Midori_rounds_SR_Inv_Result[60]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U7 ( .a ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, Midori_rounds_mul_input[52]}), .b ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, Midori_rounds_mul_input[48]}), .c ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, Midori_rounds_mul_MC1_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U4 ( .a ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, Midori_rounds_mul_input[62]}), .b ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, Midori_rounds_mul_MC1_n1}), .c ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, Midori_rounds_SR_Inv_Result[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U3 ( .a ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, Midori_rounds_mul_input[50]}), .b ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, Midori_rounds_mul_input[54]}), .c ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, Midori_rounds_mul_MC1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U2 ( .a ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, Midori_rounds_mul_input[52]}), .b ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, Midori_rounds_mul_MC1_n3}), .c ({new_AGEMA_signal_3821, new_AGEMA_signal_3820, Midori_rounds_SR_Inv_Result[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U1 ( .a ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, Midori_rounds_mul_input[60]}), .b ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, Midori_rounds_mul_input[56]}), .c ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, Midori_rounds_mul_MC1_n3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U23 ( .a ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, Midori_rounds_mul_input[44]}), .b ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, Midori_rounds_mul_MC2_n7}), .c ({new_AGEMA_signal_3823, new_AGEMA_signal_3822, Midori_rounds_SR_Inv_Result[44]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U21 ( .a ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, Midori_rounds_mul_input[34]}), .b ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, Midori_rounds_mul_MC2_n5}), .c ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, Midori_rounds_SR_Inv_Result[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U19 ( .a ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, Midori_rounds_mul_input[32]}), .b ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, Midori_rounds_mul_MC2_n3}), .c ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, Midori_rounds_SR_Inv_Result[16]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U16 ( .a ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, Midori_rounds_mul_input[38]}), .b ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, Midori_rounds_mul_MC2_n5}), .c ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, Midori_rounds_SR_Inv_Result[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U15 ( .a ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, Midori_rounds_mul_input[46]}), .b ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, Midori_rounds_mul_input[42]}), .c ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, Midori_rounds_mul_MC2_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U11 ( .a ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, Midori_rounds_mul_input[42]}), .b ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, Midori_rounds_mul_MC2_n1}), .c ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, Midori_rounds_SR_Inv_Result[6]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U8 ( .a ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, Midori_rounds_mul_input[40]}), .b ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, Midori_rounds_mul_MC2_n7}), .c ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, Midori_rounds_SR_Inv_Result[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U7 ( .a ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, Midori_rounds_mul_input[36]}), .b ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, Midori_rounds_mul_input[32]}), .c ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, Midori_rounds_mul_MC2_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U4 ( .a ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, Midori_rounds_mul_input[46]}), .b ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, Midori_rounds_mul_MC2_n1}), .c ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, Midori_rounds_SR_Inv_Result[46]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U3 ( .a ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, Midori_rounds_mul_input[34]}), .b ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, Midori_rounds_mul_input[38]}), .c ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, Midori_rounds_mul_MC2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U2 ( .a ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, Midori_rounds_mul_input[36]}), .b ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, Midori_rounds_mul_MC2_n3}), .c ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, Midori_rounds_SR_Inv_Result[56]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U1 ( .a ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, Midori_rounds_mul_input[44]}), .b ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, Midori_rounds_mul_input[40]}), .c ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, Midori_rounds_mul_MC2_n3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U23 ( .a ({new_AGEMA_signal_3805, new_AGEMA_signal_3804, Midori_rounds_mul_input[28]}), .b ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, Midori_rounds_mul_MC3_n7}), .c ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, Midori_rounds_SR_Inv_Result[48]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U21 ( .a ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, Midori_rounds_mul_input[18]}), .b ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, Midori_rounds_mul_MC3_n5}), .c ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, Midori_rounds_SR_Inv_Result[14]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U19 ( .a ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, Midori_rounds_mul_input[16]}), .b ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, Midori_rounds_mul_MC3_n3}), .c ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, Midori_rounds_SR_Inv_Result[12]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U16 ( .a ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, Midori_rounds_mul_input[22]}), .b ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, Midori_rounds_mul_MC3_n5}), .c ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, Midori_rounds_SR_Inv_Result[38]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U15 ( .a ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, Midori_rounds_mul_input[30]}), .b ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, Midori_rounds_mul_input[26]}), .c ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, Midori_rounds_mul_MC3_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U11 ( .a ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, Midori_rounds_mul_input[26]}), .b ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, Midori_rounds_mul_MC3_n1}), .c ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, Midori_rounds_SR_Inv_Result[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U8 ( .a ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, Midori_rounds_mul_input[24]}), .b ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, Midori_rounds_mul_MC3_n7}), .c ({new_AGEMA_signal_3833, new_AGEMA_signal_3832, Midori_rounds_SR_Inv_Result[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U7 ( .a ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, Midori_rounds_mul_input[20]}), .b ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, Midori_rounds_mul_input[16]}), .c ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, Midori_rounds_mul_MC3_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U4 ( .a ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, Midori_rounds_mul_input[30]}), .b ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, Midori_rounds_mul_MC3_n1}), .c ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, Midori_rounds_SR_Inv_Result[50]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U3 ( .a ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, Midori_rounds_mul_input[18]}), .b ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, Midori_rounds_mul_input[22]}), .c ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, Midori_rounds_mul_MC3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U2 ( .a ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, Midori_rounds_mul_input[20]}), .b ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, Midori_rounds_mul_MC3_n3}), .c ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, Midori_rounds_SR_Inv_Result[36]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U1 ( .a ({new_AGEMA_signal_3805, new_AGEMA_signal_3804, Midori_rounds_mul_input[28]}), .b ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, Midori_rounds_mul_input[24]}), .c ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, Midori_rounds_mul_MC3_n3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U23 ( .a ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, Midori_rounds_mul_input[12]}), .b ({new_AGEMA_signal_3815, new_AGEMA_signal_3814, Midori_rounds_mul_MC4_n7}), .c ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, Midori_rounds_SR_Inv_Result[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U21 ( .a ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, Midori_rounds_mul_input[2]}), .b ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, Midori_rounds_mul_MC4_n5}), .c ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, Midori_rounds_SR_Inv_Result[54]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U19 ( .a ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, Midori_rounds_mul_input[0]}), .b ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, Midori_rounds_mul_MC4_n3}), .c ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, Midori_rounds_SR_Inv_Result[52]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U16 ( .a ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, Midori_rounds_mul_input[6]}), .b ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, Midori_rounds_mul_MC4_n5}), .c ({new_AGEMA_signal_3411, new_AGEMA_signal_3410, Midori_rounds_SR_Inv_Result[30]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U15 ( .a ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, Midori_rounds_mul_input[14]}), .b ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, Midori_rounds_mul_input[10]}), .c ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, Midori_rounds_mul_MC4_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U11 ( .a ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, Midori_rounds_mul_input[10]}), .b ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, Midori_rounds_mul_MC4_n1}), .c ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, Midori_rounds_SR_Inv_Result[34]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U8 ( .a ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, Midori_rounds_mul_input[8]}), .b ({new_AGEMA_signal_3815, new_AGEMA_signal_3814, Midori_rounds_mul_MC4_n7}), .c ({new_AGEMA_signal_3841, new_AGEMA_signal_3840, Midori_rounds_SR_Inv_Result[32]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U7 ( .a ({new_AGEMA_signal_3785, new_AGEMA_signal_3784, Midori_rounds_mul_input[4]}), .b ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, Midori_rounds_mul_input[0]}), .c ({new_AGEMA_signal_3815, new_AGEMA_signal_3814, Midori_rounds_mul_MC4_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U4 ( .a ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, Midori_rounds_mul_input[14]}), .b ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, Midori_rounds_mul_MC4_n1}), .c ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, Midori_rounds_SR_Inv_Result[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U3 ( .a ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, Midori_rounds_mul_input[2]}), .b ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, Midori_rounds_mul_input[6]}), .c ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, Midori_rounds_mul_MC4_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U2 ( .a ({new_AGEMA_signal_3785, new_AGEMA_signal_3784, Midori_rounds_mul_input[4]}), .b ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, Midori_rounds_mul_MC4_n3}), .c ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, Midori_rounds_SR_Inv_Result[28]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U1 ( .a ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, Midori_rounds_mul_input[12]}), .b ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, Midori_rounds_mul_input[8]}), .c ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, Midori_rounds_mul_MC4_n3}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_0_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3865, new_AGEMA_signal_3864, Midori_rounds_mul_ResultXORkey[0]}), .a ({new_AGEMA_signal_3821, new_AGEMA_signal_3820, Midori_rounds_SR_Inv_Result[0]}), .c ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, Midori_rounds_round_Result[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_2_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, Midori_rounds_mul_ResultXORkey[2]}), .a ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, Midori_rounds_SR_Inv_Result[2]}), .c ({new_AGEMA_signal_3559, new_AGEMA_signal_3558, Midori_rounds_round_Result[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_4_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3847, new_AGEMA_signal_3846, Midori_rounds_mul_ResultXORkey[4]}), .a ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, Midori_rounds_SR_Inv_Result[4]}), .c ({new_AGEMA_signal_3887, new_AGEMA_signal_3886, Midori_rounds_round_Result[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_6_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, Midori_rounds_mul_ResultXORkey[6]}), .a ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, Midori_rounds_SR_Inv_Result[6]}), .c ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, Midori_rounds_round_Result[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_8_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3845, new_AGEMA_signal_3844, Midori_rounds_mul_ResultXORkey[8]}), .a ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, Midori_rounds_SR_Inv_Result[8]}), .c ({new_AGEMA_signal_3889, new_AGEMA_signal_3888, Midori_rounds_round_Result[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_10_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, Midori_rounds_mul_ResultXORkey[10]}), .a ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, Midori_rounds_SR_Inv_Result[10]}), .c ({new_AGEMA_signal_3571, new_AGEMA_signal_3570, Midori_rounds_round_Result[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_12_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3863, new_AGEMA_signal_3862, Midori_rounds_mul_ResultXORkey[12]}), .a ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, Midori_rounds_SR_Inv_Result[12]}), .c ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, Midori_rounds_round_Result[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_14_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, Midori_rounds_mul_ResultXORkey[14]}), .a ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, Midori_rounds_SR_Inv_Result[14]}), .c ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, Midori_rounds_round_Result[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_16_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3879, new_AGEMA_signal_3878, Midori_rounds_mul_ResultXORkey[16]}), .a ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, Midori_rounds_SR_Inv_Result[16]}), .c ({new_AGEMA_signal_3933, new_AGEMA_signal_3932, Midori_rounds_round_Result[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_18_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, Midori_rounds_mul_ResultXORkey[18]}), .a ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, Midori_rounds_SR_Inv_Result[18]}), .c ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, Midori_rounds_round_Result[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_20_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3877, new_AGEMA_signal_3876, Midori_rounds_mul_ResultXORkey[20]}), .a ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, Midori_rounds_SR_Inv_Result[20]}), .c ({new_AGEMA_signal_3935, new_AGEMA_signal_3934, Midori_rounds_round_Result[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_22_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, Midori_rounds_mul_ResultXORkey[22]}), .a ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, Midori_rounds_SR_Inv_Result[22]}), .c ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, Midori_rounds_round_Result[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_24_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, Midori_rounds_mul_ResultXORkey[24]}), .a ({new_AGEMA_signal_3833, new_AGEMA_signal_3832, Midori_rounds_SR_Inv_Result[24]}), .c ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, Midori_rounds_round_Result[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_26_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3499, new_AGEMA_signal_3498, Midori_rounds_mul_ResultXORkey[26]}), .a ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, Midori_rounds_SR_Inv_Result[26]}), .c ({new_AGEMA_signal_3595, new_AGEMA_signal_3594, Midori_rounds_round_Result[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_28_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3859, new_AGEMA_signal_3858, Midori_rounds_mul_ResultXORkey[28]}), .a ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, Midori_rounds_SR_Inv_Result[28]}), .c ({new_AGEMA_signal_3895, new_AGEMA_signal_3894, Midori_rounds_round_Result[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_30_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, Midori_rounds_mul_ResultXORkey[30]}), .a ({new_AGEMA_signal_3411, new_AGEMA_signal_3410, Midori_rounds_SR_Inv_Result[30]}), .c ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, Midori_rounds_round_Result[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_32_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, Midori_rounds_mul_ResultXORkey[32]}), .a ({new_AGEMA_signal_3841, new_AGEMA_signal_3840, Midori_rounds_SR_Inv_Result[32]}), .c ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, Midori_rounds_round_Result[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_34_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, Midori_rounds_mul_ResultXORkey[34]}), .a ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, Midori_rounds_SR_Inv_Result[34]}), .c ({new_AGEMA_signal_3607, new_AGEMA_signal_3606, Midori_rounds_round_Result[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_36_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3855, new_AGEMA_signal_3854, Midori_rounds_mul_ResultXORkey[36]}), .a ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, Midori_rounds_SR_Inv_Result[36]}), .c ({new_AGEMA_signal_3899, new_AGEMA_signal_3898, Midori_rounds_round_Result[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_38_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, Midori_rounds_mul_ResultXORkey[38]}), .a ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, Midori_rounds_SR_Inv_Result[38]}), .c ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, Midori_rounds_round_Result[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_40_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, Midori_rounds_mul_ResultXORkey[40]}), .a ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, Midori_rounds_SR_Inv_Result[40]}), .c ({new_AGEMA_signal_3901, new_AGEMA_signal_3900, Midori_rounds_round_Result[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_42_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, Midori_rounds_mul_ResultXORkey[42]}), .a ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, Midori_rounds_SR_Inv_Result[42]}), .c ({new_AGEMA_signal_3619, new_AGEMA_signal_3618, Midori_rounds_round_Result[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_44_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3851, new_AGEMA_signal_3850, Midori_rounds_mul_ResultXORkey[44]}), .a ({new_AGEMA_signal_3823, new_AGEMA_signal_3822, Midori_rounds_SR_Inv_Result[44]}), .c ({new_AGEMA_signal_3903, new_AGEMA_signal_3902, Midori_rounds_round_Result[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_46_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, Midori_rounds_mul_ResultXORkey[46]}), .a ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, Midori_rounds_SR_Inv_Result[46]}), .c ({new_AGEMA_signal_3625, new_AGEMA_signal_3624, Midori_rounds_round_Result[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_48_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3849, new_AGEMA_signal_3848, Midori_rounds_mul_ResultXORkey[48]}), .a ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, Midori_rounds_SR_Inv_Result[48]}), .c ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, Midori_rounds_round_Result[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_50_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3455, new_AGEMA_signal_3454, Midori_rounds_mul_ResultXORkey[50]}), .a ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, Midori_rounds_SR_Inv_Result[50]}), .c ({new_AGEMA_signal_3631, new_AGEMA_signal_3630, Midori_rounds_round_Result[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_52_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, Midori_rounds_mul_ResultXORkey[52]}), .a ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, Midori_rounds_SR_Inv_Result[52]}), .c ({new_AGEMA_signal_3937, new_AGEMA_signal_3936, Midori_rounds_round_Result[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_54_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, Midori_rounds_mul_ResultXORkey[54]}), .a ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, Midori_rounds_SR_Inv_Result[54]}), .c ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, Midori_rounds_round_Result[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_56_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, Midori_rounds_mul_ResultXORkey[56]}), .a ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, Midori_rounds_SR_Inv_Result[56]}), .c ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, Midori_rounds_round_Result[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_58_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3443, new_AGEMA_signal_3442, Midori_rounds_mul_ResultXORkey[58]}), .a ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, Midori_rounds_SR_Inv_Result[58]}), .c ({new_AGEMA_signal_3643, new_AGEMA_signal_3642, Midori_rounds_round_Result[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_60_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3907, new_AGEMA_signal_3906, Midori_rounds_mul_ResultXORkey[60]}), .a ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, Midori_rounds_SR_Inv_Result[60]}), .c ({new_AGEMA_signal_3947, new_AGEMA_signal_3946, Midori_rounds_round_Result[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_62_U1 ( .s (new_AGEMA_signal_9927), .b ({new_AGEMA_signal_3435, new_AGEMA_signal_3434, Midori_rounds_mul_ResultXORkey[62]}), .a ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, Midori_rounds_SR_Inv_Result[62]}), .c ({new_AGEMA_signal_3649, new_AGEMA_signal_3648, Midori_rounds_round_Result[62]}) ) ;
    buf_clk new_AGEMA_reg_buffer_1256 ( .C (clk), .D (new_AGEMA_signal_4721), .Q (DataOut_s0[63]) ) ;
    buf_clk new_AGEMA_reg_buffer_1258 ( .C (clk), .D (new_AGEMA_signal_4723), .Q (DataOut_s0[61]) ) ;
    buf_clk new_AGEMA_reg_buffer_1260 ( .C (clk), .D (new_AGEMA_signal_4725), .Q (DataOut_s0[59]) ) ;
    buf_clk new_AGEMA_reg_buffer_1262 ( .C (clk), .D (new_AGEMA_signal_4727), .Q (DataOut_s0[57]) ) ;
    buf_clk new_AGEMA_reg_buffer_1264 ( .C (clk), .D (new_AGEMA_signal_4729), .Q (DataOut_s0[55]) ) ;
    buf_clk new_AGEMA_reg_buffer_1266 ( .C (clk), .D (new_AGEMA_signal_4731), .Q (DataOut_s0[53]) ) ;
    buf_clk new_AGEMA_reg_buffer_1268 ( .C (clk), .D (new_AGEMA_signal_4733), .Q (DataOut_s0[51]) ) ;
    buf_clk new_AGEMA_reg_buffer_1270 ( .C (clk), .D (new_AGEMA_signal_4735), .Q (DataOut_s0[49]) ) ;
    buf_clk new_AGEMA_reg_buffer_1272 ( .C (clk), .D (new_AGEMA_signal_4737), .Q (DataOut_s0[47]) ) ;
    buf_clk new_AGEMA_reg_buffer_1274 ( .C (clk), .D (new_AGEMA_signal_4739), .Q (DataOut_s0[45]) ) ;
    buf_clk new_AGEMA_reg_buffer_1276 ( .C (clk), .D (new_AGEMA_signal_4741), .Q (DataOut_s0[43]) ) ;
    buf_clk new_AGEMA_reg_buffer_1278 ( .C (clk), .D (new_AGEMA_signal_4743), .Q (DataOut_s0[41]) ) ;
    buf_clk new_AGEMA_reg_buffer_1280 ( .C (clk), .D (new_AGEMA_signal_4745), .Q (DataOut_s0[39]) ) ;
    buf_clk new_AGEMA_reg_buffer_1282 ( .C (clk), .D (new_AGEMA_signal_4747), .Q (DataOut_s0[37]) ) ;
    buf_clk new_AGEMA_reg_buffer_1284 ( .C (clk), .D (new_AGEMA_signal_4749), .Q (DataOut_s0[35]) ) ;
    buf_clk new_AGEMA_reg_buffer_1286 ( .C (clk), .D (new_AGEMA_signal_4751), .Q (DataOut_s0[33]) ) ;
    buf_clk new_AGEMA_reg_buffer_1288 ( .C (clk), .D (new_AGEMA_signal_4753), .Q (DataOut_s0[31]) ) ;
    buf_clk new_AGEMA_reg_buffer_1290 ( .C (clk), .D (new_AGEMA_signal_4755), .Q (DataOut_s0[29]) ) ;
    buf_clk new_AGEMA_reg_buffer_1292 ( .C (clk), .D (new_AGEMA_signal_4757), .Q (DataOut_s0[27]) ) ;
    buf_clk new_AGEMA_reg_buffer_1294 ( .C (clk), .D (new_AGEMA_signal_4759), .Q (DataOut_s0[25]) ) ;
    buf_clk new_AGEMA_reg_buffer_1296 ( .C (clk), .D (new_AGEMA_signal_4761), .Q (DataOut_s0[23]) ) ;
    buf_clk new_AGEMA_reg_buffer_1298 ( .C (clk), .D (new_AGEMA_signal_4763), .Q (DataOut_s0[21]) ) ;
    buf_clk new_AGEMA_reg_buffer_1300 ( .C (clk), .D (new_AGEMA_signal_4765), .Q (DataOut_s0[19]) ) ;
    buf_clk new_AGEMA_reg_buffer_1302 ( .C (clk), .D (new_AGEMA_signal_4767), .Q (DataOut_s0[17]) ) ;
    buf_clk new_AGEMA_reg_buffer_1304 ( .C (clk), .D (new_AGEMA_signal_4769), .Q (DataOut_s0[15]) ) ;
    buf_clk new_AGEMA_reg_buffer_1306 ( .C (clk), .D (new_AGEMA_signal_4771), .Q (DataOut_s0[13]) ) ;
    buf_clk new_AGEMA_reg_buffer_1308 ( .C (clk), .D (new_AGEMA_signal_4773), .Q (DataOut_s0[11]) ) ;
    buf_clk new_AGEMA_reg_buffer_1310 ( .C (clk), .D (new_AGEMA_signal_4775), .Q (DataOut_s0[9]) ) ;
    buf_clk new_AGEMA_reg_buffer_1312 ( .C (clk), .D (new_AGEMA_signal_4777), .Q (DataOut_s0[7]) ) ;
    buf_clk new_AGEMA_reg_buffer_1314 ( .C (clk), .D (new_AGEMA_signal_4779), .Q (DataOut_s0[5]) ) ;
    buf_clk new_AGEMA_reg_buffer_1316 ( .C (clk), .D (new_AGEMA_signal_4781), .Q (DataOut_s0[3]) ) ;
    buf_clk new_AGEMA_reg_buffer_1318 ( .C (clk), .D (new_AGEMA_signal_4783), .Q (DataOut_s0[1]) ) ;
    buf_clk new_AGEMA_reg_buffer_1326 ( .C (clk), .D (new_AGEMA_signal_4791), .Q (done) ) ;
    buf_clk new_AGEMA_reg_buffer_1328 ( .C (clk), .D (new_AGEMA_signal_4793), .Q (DataOut_s1[9]) ) ;
    buf_clk new_AGEMA_reg_buffer_1330 ( .C (clk), .D (new_AGEMA_signal_4795), .Q (DataOut_s2[9]) ) ;
    buf_clk new_AGEMA_reg_buffer_1332 ( .C (clk), .D (new_AGEMA_signal_4797), .Q (DataOut_s1[7]) ) ;
    buf_clk new_AGEMA_reg_buffer_1334 ( .C (clk), .D (new_AGEMA_signal_4799), .Q (DataOut_s2[7]) ) ;
    buf_clk new_AGEMA_reg_buffer_1336 ( .C (clk), .D (new_AGEMA_signal_4801), .Q (DataOut_s1[63]) ) ;
    buf_clk new_AGEMA_reg_buffer_1338 ( .C (clk), .D (new_AGEMA_signal_4803), .Q (DataOut_s2[63]) ) ;
    buf_clk new_AGEMA_reg_buffer_1340 ( .C (clk), .D (new_AGEMA_signal_4805), .Q (DataOut_s1[61]) ) ;
    buf_clk new_AGEMA_reg_buffer_1342 ( .C (clk), .D (new_AGEMA_signal_4807), .Q (DataOut_s2[61]) ) ;
    buf_clk new_AGEMA_reg_buffer_1344 ( .C (clk), .D (new_AGEMA_signal_4809), .Q (DataOut_s1[5]) ) ;
    buf_clk new_AGEMA_reg_buffer_1346 ( .C (clk), .D (new_AGEMA_signal_4811), .Q (DataOut_s2[5]) ) ;
    buf_clk new_AGEMA_reg_buffer_1348 ( .C (clk), .D (new_AGEMA_signal_4813), .Q (DataOut_s1[59]) ) ;
    buf_clk new_AGEMA_reg_buffer_1350 ( .C (clk), .D (new_AGEMA_signal_4815), .Q (DataOut_s2[59]) ) ;
    buf_clk new_AGEMA_reg_buffer_1352 ( .C (clk), .D (new_AGEMA_signal_4817), .Q (DataOut_s1[57]) ) ;
    buf_clk new_AGEMA_reg_buffer_1354 ( .C (clk), .D (new_AGEMA_signal_4819), .Q (DataOut_s2[57]) ) ;
    buf_clk new_AGEMA_reg_buffer_1356 ( .C (clk), .D (new_AGEMA_signal_4821), .Q (DataOut_s1[55]) ) ;
    buf_clk new_AGEMA_reg_buffer_1358 ( .C (clk), .D (new_AGEMA_signal_4823), .Q (DataOut_s2[55]) ) ;
    buf_clk new_AGEMA_reg_buffer_1360 ( .C (clk), .D (new_AGEMA_signal_4825), .Q (DataOut_s1[53]) ) ;
    buf_clk new_AGEMA_reg_buffer_1362 ( .C (clk), .D (new_AGEMA_signal_4827), .Q (DataOut_s2[53]) ) ;
    buf_clk new_AGEMA_reg_buffer_1364 ( .C (clk), .D (new_AGEMA_signal_4829), .Q (DataOut_s1[51]) ) ;
    buf_clk new_AGEMA_reg_buffer_1366 ( .C (clk), .D (new_AGEMA_signal_4831), .Q (DataOut_s2[51]) ) ;
    buf_clk new_AGEMA_reg_buffer_1368 ( .C (clk), .D (new_AGEMA_signal_4833), .Q (DataOut_s1[49]) ) ;
    buf_clk new_AGEMA_reg_buffer_1370 ( .C (clk), .D (new_AGEMA_signal_4835), .Q (DataOut_s2[49]) ) ;
    buf_clk new_AGEMA_reg_buffer_1372 ( .C (clk), .D (new_AGEMA_signal_4837), .Q (DataOut_s1[47]) ) ;
    buf_clk new_AGEMA_reg_buffer_1374 ( .C (clk), .D (new_AGEMA_signal_4839), .Q (DataOut_s2[47]) ) ;
    buf_clk new_AGEMA_reg_buffer_1376 ( .C (clk), .D (new_AGEMA_signal_4841), .Q (DataOut_s1[45]) ) ;
    buf_clk new_AGEMA_reg_buffer_1378 ( .C (clk), .D (new_AGEMA_signal_4843), .Q (DataOut_s2[45]) ) ;
    buf_clk new_AGEMA_reg_buffer_1380 ( .C (clk), .D (new_AGEMA_signal_4845), .Q (DataOut_s1[43]) ) ;
    buf_clk new_AGEMA_reg_buffer_1382 ( .C (clk), .D (new_AGEMA_signal_4847), .Q (DataOut_s2[43]) ) ;
    buf_clk new_AGEMA_reg_buffer_1384 ( .C (clk), .D (new_AGEMA_signal_4849), .Q (DataOut_s1[41]) ) ;
    buf_clk new_AGEMA_reg_buffer_1386 ( .C (clk), .D (new_AGEMA_signal_4851), .Q (DataOut_s2[41]) ) ;
    buf_clk new_AGEMA_reg_buffer_1388 ( .C (clk), .D (new_AGEMA_signal_4853), .Q (DataOut_s1[3]) ) ;
    buf_clk new_AGEMA_reg_buffer_1390 ( .C (clk), .D (new_AGEMA_signal_4855), .Q (DataOut_s2[3]) ) ;
    buf_clk new_AGEMA_reg_buffer_1392 ( .C (clk), .D (new_AGEMA_signal_4857), .Q (DataOut_s1[39]) ) ;
    buf_clk new_AGEMA_reg_buffer_1394 ( .C (clk), .D (new_AGEMA_signal_4859), .Q (DataOut_s2[39]) ) ;
    buf_clk new_AGEMA_reg_buffer_1396 ( .C (clk), .D (new_AGEMA_signal_4861), .Q (DataOut_s1[37]) ) ;
    buf_clk new_AGEMA_reg_buffer_1398 ( .C (clk), .D (new_AGEMA_signal_4863), .Q (DataOut_s2[37]) ) ;
    buf_clk new_AGEMA_reg_buffer_1400 ( .C (clk), .D (new_AGEMA_signal_4865), .Q (DataOut_s1[35]) ) ;
    buf_clk new_AGEMA_reg_buffer_1402 ( .C (clk), .D (new_AGEMA_signal_4867), .Q (DataOut_s2[35]) ) ;
    buf_clk new_AGEMA_reg_buffer_1404 ( .C (clk), .D (new_AGEMA_signal_4869), .Q (DataOut_s1[33]) ) ;
    buf_clk new_AGEMA_reg_buffer_1406 ( .C (clk), .D (new_AGEMA_signal_4871), .Q (DataOut_s2[33]) ) ;
    buf_clk new_AGEMA_reg_buffer_1408 ( .C (clk), .D (new_AGEMA_signal_4873), .Q (DataOut_s1[31]) ) ;
    buf_clk new_AGEMA_reg_buffer_1410 ( .C (clk), .D (new_AGEMA_signal_4875), .Q (DataOut_s2[31]) ) ;
    buf_clk new_AGEMA_reg_buffer_1412 ( .C (clk), .D (new_AGEMA_signal_4877), .Q (DataOut_s1[29]) ) ;
    buf_clk new_AGEMA_reg_buffer_1414 ( .C (clk), .D (new_AGEMA_signal_4879), .Q (DataOut_s2[29]) ) ;
    buf_clk new_AGEMA_reg_buffer_1416 ( .C (clk), .D (new_AGEMA_signal_4881), .Q (DataOut_s1[27]) ) ;
    buf_clk new_AGEMA_reg_buffer_1418 ( .C (clk), .D (new_AGEMA_signal_4883), .Q (DataOut_s2[27]) ) ;
    buf_clk new_AGEMA_reg_buffer_1420 ( .C (clk), .D (new_AGEMA_signal_4885), .Q (DataOut_s1[25]) ) ;
    buf_clk new_AGEMA_reg_buffer_1422 ( .C (clk), .D (new_AGEMA_signal_4887), .Q (DataOut_s2[25]) ) ;
    buf_clk new_AGEMA_reg_buffer_1424 ( .C (clk), .D (new_AGEMA_signal_4889), .Q (DataOut_s1[23]) ) ;
    buf_clk new_AGEMA_reg_buffer_1426 ( .C (clk), .D (new_AGEMA_signal_4891), .Q (DataOut_s2[23]) ) ;
    buf_clk new_AGEMA_reg_buffer_1428 ( .C (clk), .D (new_AGEMA_signal_4893), .Q (DataOut_s1[21]) ) ;
    buf_clk new_AGEMA_reg_buffer_1430 ( .C (clk), .D (new_AGEMA_signal_4895), .Q (DataOut_s2[21]) ) ;
    buf_clk new_AGEMA_reg_buffer_1432 ( .C (clk), .D (new_AGEMA_signal_4897), .Q (DataOut_s1[1]) ) ;
    buf_clk new_AGEMA_reg_buffer_1434 ( .C (clk), .D (new_AGEMA_signal_4899), .Q (DataOut_s2[1]) ) ;
    buf_clk new_AGEMA_reg_buffer_1436 ( .C (clk), .D (new_AGEMA_signal_4901), .Q (DataOut_s1[19]) ) ;
    buf_clk new_AGEMA_reg_buffer_1438 ( .C (clk), .D (new_AGEMA_signal_4903), .Q (DataOut_s2[19]) ) ;
    buf_clk new_AGEMA_reg_buffer_1440 ( .C (clk), .D (new_AGEMA_signal_4905), .Q (DataOut_s1[17]) ) ;
    buf_clk new_AGEMA_reg_buffer_1442 ( .C (clk), .D (new_AGEMA_signal_4907), .Q (DataOut_s2[17]) ) ;
    buf_clk new_AGEMA_reg_buffer_1444 ( .C (clk), .D (new_AGEMA_signal_4909), .Q (DataOut_s1[15]) ) ;
    buf_clk new_AGEMA_reg_buffer_1446 ( .C (clk), .D (new_AGEMA_signal_4911), .Q (DataOut_s2[15]) ) ;
    buf_clk new_AGEMA_reg_buffer_1448 ( .C (clk), .D (new_AGEMA_signal_4913), .Q (DataOut_s1[13]) ) ;
    buf_clk new_AGEMA_reg_buffer_1450 ( .C (clk), .D (new_AGEMA_signal_4915), .Q (DataOut_s2[13]) ) ;
    buf_clk new_AGEMA_reg_buffer_1452 ( .C (clk), .D (new_AGEMA_signal_4917), .Q (DataOut_s1[11]) ) ;
    buf_clk new_AGEMA_reg_buffer_1454 ( .C (clk), .D (new_AGEMA_signal_4919), .Q (DataOut_s2[11]) ) ;
    buf_clk new_AGEMA_reg_buffer_3874 ( .C (clk), .D (new_AGEMA_signal_7338), .Q (new_AGEMA_signal_7339) ) ;
    buf_clk new_AGEMA_reg_buffer_3882 ( .C (clk), .D (new_AGEMA_signal_7346), .Q (new_AGEMA_signal_7347) ) ;
    buf_clk new_AGEMA_reg_buffer_3890 ( .C (clk), .D (new_AGEMA_signal_7354), .Q (new_AGEMA_signal_7355) ) ;
    buf_clk new_AGEMA_reg_buffer_3898 ( .C (clk), .D (new_AGEMA_signal_7362), .Q (new_AGEMA_signal_7363) ) ;
    buf_clk new_AGEMA_reg_buffer_3906 ( .C (clk), .D (new_AGEMA_signal_7370), .Q (new_AGEMA_signal_7371) ) ;
    buf_clk new_AGEMA_reg_buffer_3914 ( .C (clk), .D (new_AGEMA_signal_7378), .Q (new_AGEMA_signal_7379) ) ;
    buf_clk new_AGEMA_reg_buffer_3922 ( .C (clk), .D (new_AGEMA_signal_7386), .Q (new_AGEMA_signal_7387) ) ;
    buf_clk new_AGEMA_reg_buffer_3930 ( .C (clk), .D (new_AGEMA_signal_7394), .Q (new_AGEMA_signal_7395) ) ;
    buf_clk new_AGEMA_reg_buffer_3938 ( .C (clk), .D (new_AGEMA_signal_7402), .Q (new_AGEMA_signal_7403) ) ;
    buf_clk new_AGEMA_reg_buffer_3946 ( .C (clk), .D (new_AGEMA_signal_7410), .Q (new_AGEMA_signal_7411) ) ;
    buf_clk new_AGEMA_reg_buffer_3954 ( .C (clk), .D (new_AGEMA_signal_7418), .Q (new_AGEMA_signal_7419) ) ;
    buf_clk new_AGEMA_reg_buffer_3962 ( .C (clk), .D (new_AGEMA_signal_7426), .Q (new_AGEMA_signal_7427) ) ;
    buf_clk new_AGEMA_reg_buffer_3970 ( .C (clk), .D (new_AGEMA_signal_7434), .Q (new_AGEMA_signal_7435) ) ;
    buf_clk new_AGEMA_reg_buffer_3978 ( .C (clk), .D (new_AGEMA_signal_7442), .Q (new_AGEMA_signal_7443) ) ;
    buf_clk new_AGEMA_reg_buffer_3986 ( .C (clk), .D (new_AGEMA_signal_7450), .Q (new_AGEMA_signal_7451) ) ;
    buf_clk new_AGEMA_reg_buffer_3994 ( .C (clk), .D (new_AGEMA_signal_7458), .Q (new_AGEMA_signal_7459) ) ;
    buf_clk new_AGEMA_reg_buffer_4002 ( .C (clk), .D (new_AGEMA_signal_7466), .Q (new_AGEMA_signal_7467) ) ;
    buf_clk new_AGEMA_reg_buffer_4010 ( .C (clk), .D (new_AGEMA_signal_7474), .Q (new_AGEMA_signal_7475) ) ;
    buf_clk new_AGEMA_reg_buffer_4018 ( .C (clk), .D (new_AGEMA_signal_7482), .Q (new_AGEMA_signal_7483) ) ;
    buf_clk new_AGEMA_reg_buffer_4026 ( .C (clk), .D (new_AGEMA_signal_7490), .Q (new_AGEMA_signal_7491) ) ;
    buf_clk new_AGEMA_reg_buffer_4034 ( .C (clk), .D (new_AGEMA_signal_7498), .Q (new_AGEMA_signal_7499) ) ;
    buf_clk new_AGEMA_reg_buffer_4042 ( .C (clk), .D (new_AGEMA_signal_7506), .Q (new_AGEMA_signal_7507) ) ;
    buf_clk new_AGEMA_reg_buffer_4050 ( .C (clk), .D (new_AGEMA_signal_7514), .Q (new_AGEMA_signal_7515) ) ;
    buf_clk new_AGEMA_reg_buffer_4058 ( .C (clk), .D (new_AGEMA_signal_7522), .Q (new_AGEMA_signal_7523) ) ;
    buf_clk new_AGEMA_reg_buffer_4066 ( .C (clk), .D (new_AGEMA_signal_7530), .Q (new_AGEMA_signal_7531) ) ;
    buf_clk new_AGEMA_reg_buffer_4074 ( .C (clk), .D (new_AGEMA_signal_7538), .Q (new_AGEMA_signal_7539) ) ;
    buf_clk new_AGEMA_reg_buffer_4082 ( .C (clk), .D (new_AGEMA_signal_7546), .Q (new_AGEMA_signal_7547) ) ;
    buf_clk new_AGEMA_reg_buffer_4090 ( .C (clk), .D (new_AGEMA_signal_7554), .Q (new_AGEMA_signal_7555) ) ;
    buf_clk new_AGEMA_reg_buffer_4098 ( .C (clk), .D (new_AGEMA_signal_7562), .Q (new_AGEMA_signal_7563) ) ;
    buf_clk new_AGEMA_reg_buffer_4106 ( .C (clk), .D (new_AGEMA_signal_7570), .Q (new_AGEMA_signal_7571) ) ;
    buf_clk new_AGEMA_reg_buffer_4114 ( .C (clk), .D (new_AGEMA_signal_7578), .Q (new_AGEMA_signal_7579) ) ;
    buf_clk new_AGEMA_reg_buffer_4122 ( .C (clk), .D (new_AGEMA_signal_7586), .Q (new_AGEMA_signal_7587) ) ;
    buf_clk new_AGEMA_reg_buffer_4130 ( .C (clk), .D (new_AGEMA_signal_7594), .Q (new_AGEMA_signal_7595) ) ;
    buf_clk new_AGEMA_reg_buffer_4138 ( .C (clk), .D (new_AGEMA_signal_7602), .Q (new_AGEMA_signal_7603) ) ;
    buf_clk new_AGEMA_reg_buffer_4146 ( .C (clk), .D (new_AGEMA_signal_7610), .Q (new_AGEMA_signal_7611) ) ;
    buf_clk new_AGEMA_reg_buffer_4154 ( .C (clk), .D (new_AGEMA_signal_7618), .Q (new_AGEMA_signal_7619) ) ;
    buf_clk new_AGEMA_reg_buffer_4162 ( .C (clk), .D (new_AGEMA_signal_7626), .Q (new_AGEMA_signal_7627) ) ;
    buf_clk new_AGEMA_reg_buffer_4170 ( .C (clk), .D (new_AGEMA_signal_7634), .Q (new_AGEMA_signal_7635) ) ;
    buf_clk new_AGEMA_reg_buffer_4178 ( .C (clk), .D (new_AGEMA_signal_7642), .Q (new_AGEMA_signal_7643) ) ;
    buf_clk new_AGEMA_reg_buffer_4186 ( .C (clk), .D (new_AGEMA_signal_7650), .Q (new_AGEMA_signal_7651) ) ;
    buf_clk new_AGEMA_reg_buffer_4194 ( .C (clk), .D (new_AGEMA_signal_7658), .Q (new_AGEMA_signal_7659) ) ;
    buf_clk new_AGEMA_reg_buffer_4202 ( .C (clk), .D (new_AGEMA_signal_7666), .Q (new_AGEMA_signal_7667) ) ;
    buf_clk new_AGEMA_reg_buffer_4210 ( .C (clk), .D (new_AGEMA_signal_7674), .Q (new_AGEMA_signal_7675) ) ;
    buf_clk new_AGEMA_reg_buffer_4218 ( .C (clk), .D (new_AGEMA_signal_7682), .Q (new_AGEMA_signal_7683) ) ;
    buf_clk new_AGEMA_reg_buffer_4226 ( .C (clk), .D (new_AGEMA_signal_7690), .Q (new_AGEMA_signal_7691) ) ;
    buf_clk new_AGEMA_reg_buffer_4234 ( .C (clk), .D (new_AGEMA_signal_7698), .Q (new_AGEMA_signal_7699) ) ;
    buf_clk new_AGEMA_reg_buffer_4242 ( .C (clk), .D (new_AGEMA_signal_7706), .Q (new_AGEMA_signal_7707) ) ;
    buf_clk new_AGEMA_reg_buffer_4250 ( .C (clk), .D (new_AGEMA_signal_7714), .Q (new_AGEMA_signal_7715) ) ;
    buf_clk new_AGEMA_reg_buffer_4258 ( .C (clk), .D (new_AGEMA_signal_7722), .Q (new_AGEMA_signal_7723) ) ;
    buf_clk new_AGEMA_reg_buffer_4266 ( .C (clk), .D (new_AGEMA_signal_7730), .Q (new_AGEMA_signal_7731) ) ;
    buf_clk new_AGEMA_reg_buffer_4274 ( .C (clk), .D (new_AGEMA_signal_7738), .Q (new_AGEMA_signal_7739) ) ;
    buf_clk new_AGEMA_reg_buffer_4282 ( .C (clk), .D (new_AGEMA_signal_7746), .Q (new_AGEMA_signal_7747) ) ;
    buf_clk new_AGEMA_reg_buffer_4290 ( .C (clk), .D (new_AGEMA_signal_7754), .Q (new_AGEMA_signal_7755) ) ;
    buf_clk new_AGEMA_reg_buffer_4298 ( .C (clk), .D (new_AGEMA_signal_7762), .Q (new_AGEMA_signal_7763) ) ;
    buf_clk new_AGEMA_reg_buffer_4306 ( .C (clk), .D (new_AGEMA_signal_7770), .Q (new_AGEMA_signal_7771) ) ;
    buf_clk new_AGEMA_reg_buffer_4314 ( .C (clk), .D (new_AGEMA_signal_7778), .Q (new_AGEMA_signal_7779) ) ;
    buf_clk new_AGEMA_reg_buffer_4322 ( .C (clk), .D (new_AGEMA_signal_7786), .Q (new_AGEMA_signal_7787) ) ;
    buf_clk new_AGEMA_reg_buffer_4330 ( .C (clk), .D (new_AGEMA_signal_7794), .Q (new_AGEMA_signal_7795) ) ;
    buf_clk new_AGEMA_reg_buffer_4338 ( .C (clk), .D (new_AGEMA_signal_7802), .Q (new_AGEMA_signal_7803) ) ;
    buf_clk new_AGEMA_reg_buffer_4346 ( .C (clk), .D (new_AGEMA_signal_7810), .Q (new_AGEMA_signal_7811) ) ;
    buf_clk new_AGEMA_reg_buffer_4354 ( .C (clk), .D (new_AGEMA_signal_7818), .Q (new_AGEMA_signal_7819) ) ;
    buf_clk new_AGEMA_reg_buffer_4362 ( .C (clk), .D (new_AGEMA_signal_7826), .Q (new_AGEMA_signal_7827) ) ;
    buf_clk new_AGEMA_reg_buffer_4370 ( .C (clk), .D (new_AGEMA_signal_7834), .Q (new_AGEMA_signal_7835) ) ;
    buf_clk new_AGEMA_reg_buffer_4378 ( .C (clk), .D (new_AGEMA_signal_7842), .Q (new_AGEMA_signal_7843) ) ;
    buf_clk new_AGEMA_reg_buffer_4386 ( .C (clk), .D (new_AGEMA_signal_7850), .Q (new_AGEMA_signal_7851) ) ;
    buf_clk new_AGEMA_reg_buffer_4394 ( .C (clk), .D (new_AGEMA_signal_7858), .Q (new_AGEMA_signal_7859) ) ;
    buf_clk new_AGEMA_reg_buffer_4402 ( .C (clk), .D (new_AGEMA_signal_7866), .Q (new_AGEMA_signal_7867) ) ;
    buf_clk new_AGEMA_reg_buffer_4410 ( .C (clk), .D (new_AGEMA_signal_7874), .Q (new_AGEMA_signal_7875) ) ;
    buf_clk new_AGEMA_reg_buffer_4418 ( .C (clk), .D (new_AGEMA_signal_7882), .Q (new_AGEMA_signal_7883) ) ;
    buf_clk new_AGEMA_reg_buffer_4426 ( .C (clk), .D (new_AGEMA_signal_7890), .Q (new_AGEMA_signal_7891) ) ;
    buf_clk new_AGEMA_reg_buffer_4434 ( .C (clk), .D (new_AGEMA_signal_7898), .Q (new_AGEMA_signal_7899) ) ;
    buf_clk new_AGEMA_reg_buffer_4442 ( .C (clk), .D (new_AGEMA_signal_7906), .Q (new_AGEMA_signal_7907) ) ;
    buf_clk new_AGEMA_reg_buffer_4450 ( .C (clk), .D (new_AGEMA_signal_7914), .Q (new_AGEMA_signal_7915) ) ;
    buf_clk new_AGEMA_reg_buffer_4458 ( .C (clk), .D (new_AGEMA_signal_7922), .Q (new_AGEMA_signal_7923) ) ;
    buf_clk new_AGEMA_reg_buffer_4466 ( .C (clk), .D (new_AGEMA_signal_7930), .Q (new_AGEMA_signal_7931) ) ;
    buf_clk new_AGEMA_reg_buffer_4474 ( .C (clk), .D (new_AGEMA_signal_7938), .Q (new_AGEMA_signal_7939) ) ;
    buf_clk new_AGEMA_reg_buffer_4482 ( .C (clk), .D (new_AGEMA_signal_7946), .Q (new_AGEMA_signal_7947) ) ;
    buf_clk new_AGEMA_reg_buffer_4490 ( .C (clk), .D (new_AGEMA_signal_7954), .Q (new_AGEMA_signal_7955) ) ;
    buf_clk new_AGEMA_reg_buffer_4498 ( .C (clk), .D (new_AGEMA_signal_7962), .Q (new_AGEMA_signal_7963) ) ;
    buf_clk new_AGEMA_reg_buffer_4506 ( .C (clk), .D (new_AGEMA_signal_7970), .Q (new_AGEMA_signal_7971) ) ;
    buf_clk new_AGEMA_reg_buffer_4514 ( .C (clk), .D (new_AGEMA_signal_7978), .Q (new_AGEMA_signal_7979) ) ;
    buf_clk new_AGEMA_reg_buffer_4522 ( .C (clk), .D (new_AGEMA_signal_7986), .Q (new_AGEMA_signal_7987) ) ;
    buf_clk new_AGEMA_reg_buffer_4530 ( .C (clk), .D (new_AGEMA_signal_7994), .Q (new_AGEMA_signal_7995) ) ;
    buf_clk new_AGEMA_reg_buffer_4538 ( .C (clk), .D (new_AGEMA_signal_8002), .Q (new_AGEMA_signal_8003) ) ;
    buf_clk new_AGEMA_reg_buffer_4546 ( .C (clk), .D (new_AGEMA_signal_8010), .Q (new_AGEMA_signal_8011) ) ;
    buf_clk new_AGEMA_reg_buffer_4554 ( .C (clk), .D (new_AGEMA_signal_8018), .Q (new_AGEMA_signal_8019) ) ;
    buf_clk new_AGEMA_reg_buffer_4562 ( .C (clk), .D (new_AGEMA_signal_8026), .Q (new_AGEMA_signal_8027) ) ;
    buf_clk new_AGEMA_reg_buffer_4570 ( .C (clk), .D (new_AGEMA_signal_8034), .Q (new_AGEMA_signal_8035) ) ;
    buf_clk new_AGEMA_reg_buffer_4578 ( .C (clk), .D (new_AGEMA_signal_8042), .Q (new_AGEMA_signal_8043) ) ;
    buf_clk new_AGEMA_reg_buffer_4586 ( .C (clk), .D (new_AGEMA_signal_8050), .Q (new_AGEMA_signal_8051) ) ;
    buf_clk new_AGEMA_reg_buffer_4594 ( .C (clk), .D (new_AGEMA_signal_8058), .Q (new_AGEMA_signal_8059) ) ;
    buf_clk new_AGEMA_reg_buffer_4602 ( .C (clk), .D (new_AGEMA_signal_8066), .Q (new_AGEMA_signal_8067) ) ;
    buf_clk new_AGEMA_reg_buffer_4610 ( .C (clk), .D (new_AGEMA_signal_8074), .Q (new_AGEMA_signal_8075) ) ;
    buf_clk new_AGEMA_reg_buffer_4618 ( .C (clk), .D (new_AGEMA_signal_8082), .Q (new_AGEMA_signal_8083) ) ;
    buf_clk new_AGEMA_reg_buffer_4626 ( .C (clk), .D (new_AGEMA_signal_8090), .Q (new_AGEMA_signal_8091) ) ;
    buf_clk new_AGEMA_reg_buffer_4634 ( .C (clk), .D (new_AGEMA_signal_8098), .Q (new_AGEMA_signal_8099) ) ;
    buf_clk new_AGEMA_reg_buffer_4642 ( .C (clk), .D (new_AGEMA_signal_8106), .Q (new_AGEMA_signal_8107) ) ;
    buf_clk new_AGEMA_reg_buffer_4650 ( .C (clk), .D (new_AGEMA_signal_8114), .Q (new_AGEMA_signal_8115) ) ;
    buf_clk new_AGEMA_reg_buffer_4658 ( .C (clk), .D (new_AGEMA_signal_8122), .Q (new_AGEMA_signal_8123) ) ;
    buf_clk new_AGEMA_reg_buffer_4666 ( .C (clk), .D (new_AGEMA_signal_8130), .Q (new_AGEMA_signal_8131) ) ;
    buf_clk new_AGEMA_reg_buffer_4674 ( .C (clk), .D (new_AGEMA_signal_8138), .Q (new_AGEMA_signal_8139) ) ;
    buf_clk new_AGEMA_reg_buffer_4682 ( .C (clk), .D (new_AGEMA_signal_8146), .Q (new_AGEMA_signal_8147) ) ;
    buf_clk new_AGEMA_reg_buffer_4690 ( .C (clk), .D (new_AGEMA_signal_8154), .Q (new_AGEMA_signal_8155) ) ;
    buf_clk new_AGEMA_reg_buffer_4698 ( .C (clk), .D (new_AGEMA_signal_8162), .Q (new_AGEMA_signal_8163) ) ;
    buf_clk new_AGEMA_reg_buffer_4706 ( .C (clk), .D (new_AGEMA_signal_8170), .Q (new_AGEMA_signal_8171) ) ;
    buf_clk new_AGEMA_reg_buffer_4714 ( .C (clk), .D (new_AGEMA_signal_8178), .Q (new_AGEMA_signal_8179) ) ;
    buf_clk new_AGEMA_reg_buffer_4722 ( .C (clk), .D (new_AGEMA_signal_8186), .Q (new_AGEMA_signal_8187) ) ;
    buf_clk new_AGEMA_reg_buffer_4730 ( .C (clk), .D (new_AGEMA_signal_8194), .Q (new_AGEMA_signal_8195) ) ;
    buf_clk new_AGEMA_reg_buffer_4738 ( .C (clk), .D (new_AGEMA_signal_8202), .Q (new_AGEMA_signal_8203) ) ;
    buf_clk new_AGEMA_reg_buffer_4746 ( .C (clk), .D (new_AGEMA_signal_8210), .Q (new_AGEMA_signal_8211) ) ;
    buf_clk new_AGEMA_reg_buffer_4754 ( .C (clk), .D (new_AGEMA_signal_8218), .Q (new_AGEMA_signal_8219) ) ;
    buf_clk new_AGEMA_reg_buffer_4762 ( .C (clk), .D (new_AGEMA_signal_8226), .Q (new_AGEMA_signal_8227) ) ;
    buf_clk new_AGEMA_reg_buffer_4770 ( .C (clk), .D (new_AGEMA_signal_8234), .Q (new_AGEMA_signal_8235) ) ;
    buf_clk new_AGEMA_reg_buffer_4778 ( .C (clk), .D (new_AGEMA_signal_8242), .Q (new_AGEMA_signal_8243) ) ;
    buf_clk new_AGEMA_reg_buffer_4786 ( .C (clk), .D (new_AGEMA_signal_8250), .Q (new_AGEMA_signal_8251) ) ;
    buf_clk new_AGEMA_reg_buffer_4794 ( .C (clk), .D (new_AGEMA_signal_8258), .Q (new_AGEMA_signal_8259) ) ;
    buf_clk new_AGEMA_reg_buffer_4802 ( .C (clk), .D (new_AGEMA_signal_8266), .Q (new_AGEMA_signal_8267) ) ;
    buf_clk new_AGEMA_reg_buffer_4810 ( .C (clk), .D (new_AGEMA_signal_8274), .Q (new_AGEMA_signal_8275) ) ;
    buf_clk new_AGEMA_reg_buffer_4818 ( .C (clk), .D (new_AGEMA_signal_8282), .Q (new_AGEMA_signal_8283) ) ;
    buf_clk new_AGEMA_reg_buffer_4826 ( .C (clk), .D (new_AGEMA_signal_8290), .Q (new_AGEMA_signal_8291) ) ;
    buf_clk new_AGEMA_reg_buffer_4834 ( .C (clk), .D (new_AGEMA_signal_8298), .Q (new_AGEMA_signal_8299) ) ;
    buf_clk new_AGEMA_reg_buffer_4842 ( .C (clk), .D (new_AGEMA_signal_8306), .Q (new_AGEMA_signal_8307) ) ;
    buf_clk new_AGEMA_reg_buffer_4850 ( .C (clk), .D (new_AGEMA_signal_8314), .Q (new_AGEMA_signal_8315) ) ;
    buf_clk new_AGEMA_reg_buffer_4858 ( .C (clk), .D (new_AGEMA_signal_8322), .Q (new_AGEMA_signal_8323) ) ;
    buf_clk new_AGEMA_reg_buffer_4866 ( .C (clk), .D (new_AGEMA_signal_8330), .Q (new_AGEMA_signal_8331) ) ;
    buf_clk new_AGEMA_reg_buffer_4874 ( .C (clk), .D (new_AGEMA_signal_8338), .Q (new_AGEMA_signal_8339) ) ;
    buf_clk new_AGEMA_reg_buffer_4882 ( .C (clk), .D (new_AGEMA_signal_8346), .Q (new_AGEMA_signal_8347) ) ;
    buf_clk new_AGEMA_reg_buffer_4890 ( .C (clk), .D (new_AGEMA_signal_8354), .Q (new_AGEMA_signal_8355) ) ;
    buf_clk new_AGEMA_reg_buffer_4898 ( .C (clk), .D (new_AGEMA_signal_8362), .Q (new_AGEMA_signal_8363) ) ;
    buf_clk new_AGEMA_reg_buffer_4906 ( .C (clk), .D (new_AGEMA_signal_8370), .Q (new_AGEMA_signal_8371) ) ;
    buf_clk new_AGEMA_reg_buffer_4914 ( .C (clk), .D (new_AGEMA_signal_8378), .Q (new_AGEMA_signal_8379) ) ;
    buf_clk new_AGEMA_reg_buffer_4922 ( .C (clk), .D (new_AGEMA_signal_8386), .Q (new_AGEMA_signal_8387) ) ;
    buf_clk new_AGEMA_reg_buffer_4930 ( .C (clk), .D (new_AGEMA_signal_8394), .Q (new_AGEMA_signal_8395) ) ;
    buf_clk new_AGEMA_reg_buffer_4938 ( .C (clk), .D (new_AGEMA_signal_8402), .Q (new_AGEMA_signal_8403) ) ;
    buf_clk new_AGEMA_reg_buffer_4946 ( .C (clk), .D (new_AGEMA_signal_8410), .Q (new_AGEMA_signal_8411) ) ;
    buf_clk new_AGEMA_reg_buffer_4954 ( .C (clk), .D (new_AGEMA_signal_8418), .Q (new_AGEMA_signal_8419) ) ;
    buf_clk new_AGEMA_reg_buffer_4962 ( .C (clk), .D (new_AGEMA_signal_8426), .Q (new_AGEMA_signal_8427) ) ;
    buf_clk new_AGEMA_reg_buffer_4970 ( .C (clk), .D (new_AGEMA_signal_8434), .Q (new_AGEMA_signal_8435) ) ;
    buf_clk new_AGEMA_reg_buffer_4978 ( .C (clk), .D (new_AGEMA_signal_8442), .Q (new_AGEMA_signal_8443) ) ;
    buf_clk new_AGEMA_reg_buffer_4986 ( .C (clk), .D (new_AGEMA_signal_8450), .Q (new_AGEMA_signal_8451) ) ;
    buf_clk new_AGEMA_reg_buffer_4994 ( .C (clk), .D (new_AGEMA_signal_8458), .Q (new_AGEMA_signal_8459) ) ;
    buf_clk new_AGEMA_reg_buffer_5002 ( .C (clk), .D (new_AGEMA_signal_8466), .Q (new_AGEMA_signal_8467) ) ;
    buf_clk new_AGEMA_reg_buffer_5010 ( .C (clk), .D (new_AGEMA_signal_8474), .Q (new_AGEMA_signal_8475) ) ;
    buf_clk new_AGEMA_reg_buffer_5018 ( .C (clk), .D (new_AGEMA_signal_8482), .Q (new_AGEMA_signal_8483) ) ;
    buf_clk new_AGEMA_reg_buffer_5026 ( .C (clk), .D (new_AGEMA_signal_8490), .Q (new_AGEMA_signal_8491) ) ;
    buf_clk new_AGEMA_reg_buffer_5034 ( .C (clk), .D (new_AGEMA_signal_8498), .Q (new_AGEMA_signal_8499) ) ;
    buf_clk new_AGEMA_reg_buffer_5042 ( .C (clk), .D (new_AGEMA_signal_8506), .Q (new_AGEMA_signal_8507) ) ;
    buf_clk new_AGEMA_reg_buffer_5050 ( .C (clk), .D (new_AGEMA_signal_8514), .Q (new_AGEMA_signal_8515) ) ;
    buf_clk new_AGEMA_reg_buffer_5058 ( .C (clk), .D (new_AGEMA_signal_8522), .Q (new_AGEMA_signal_8523) ) ;
    buf_clk new_AGEMA_reg_buffer_5066 ( .C (clk), .D (new_AGEMA_signal_8530), .Q (new_AGEMA_signal_8531) ) ;
    buf_clk new_AGEMA_reg_buffer_5074 ( .C (clk), .D (new_AGEMA_signal_8538), .Q (new_AGEMA_signal_8539) ) ;
    buf_clk new_AGEMA_reg_buffer_5082 ( .C (clk), .D (new_AGEMA_signal_8546), .Q (new_AGEMA_signal_8547) ) ;
    buf_clk new_AGEMA_reg_buffer_5090 ( .C (clk), .D (new_AGEMA_signal_8554), .Q (new_AGEMA_signal_8555) ) ;
    buf_clk new_AGEMA_reg_buffer_5098 ( .C (clk), .D (new_AGEMA_signal_8562), .Q (new_AGEMA_signal_8563) ) ;
    buf_clk new_AGEMA_reg_buffer_5106 ( .C (clk), .D (new_AGEMA_signal_8570), .Q (new_AGEMA_signal_8571) ) ;
    buf_clk new_AGEMA_reg_buffer_5114 ( .C (clk), .D (new_AGEMA_signal_8578), .Q (new_AGEMA_signal_8579) ) ;
    buf_clk new_AGEMA_reg_buffer_5122 ( .C (clk), .D (new_AGEMA_signal_8586), .Q (new_AGEMA_signal_8587) ) ;
    buf_clk new_AGEMA_reg_buffer_5130 ( .C (clk), .D (new_AGEMA_signal_8594), .Q (new_AGEMA_signal_8595) ) ;
    buf_clk new_AGEMA_reg_buffer_5138 ( .C (clk), .D (new_AGEMA_signal_8602), .Q (new_AGEMA_signal_8603) ) ;
    buf_clk new_AGEMA_reg_buffer_5146 ( .C (clk), .D (new_AGEMA_signal_8610), .Q (new_AGEMA_signal_8611) ) ;
    buf_clk new_AGEMA_reg_buffer_5154 ( .C (clk), .D (new_AGEMA_signal_8618), .Q (new_AGEMA_signal_8619) ) ;
    buf_clk new_AGEMA_reg_buffer_5162 ( .C (clk), .D (new_AGEMA_signal_8626), .Q (new_AGEMA_signal_8627) ) ;
    buf_clk new_AGEMA_reg_buffer_5170 ( .C (clk), .D (new_AGEMA_signal_8634), .Q (new_AGEMA_signal_8635) ) ;
    buf_clk new_AGEMA_reg_buffer_5178 ( .C (clk), .D (new_AGEMA_signal_8642), .Q (new_AGEMA_signal_8643) ) ;
    buf_clk new_AGEMA_reg_buffer_5186 ( .C (clk), .D (new_AGEMA_signal_8650), .Q (new_AGEMA_signal_8651) ) ;
    buf_clk new_AGEMA_reg_buffer_5194 ( .C (clk), .D (new_AGEMA_signal_8658), .Q (new_AGEMA_signal_8659) ) ;
    buf_clk new_AGEMA_reg_buffer_5202 ( .C (clk), .D (new_AGEMA_signal_8666), .Q (new_AGEMA_signal_8667) ) ;
    buf_clk new_AGEMA_reg_buffer_5210 ( .C (clk), .D (new_AGEMA_signal_8674), .Q (new_AGEMA_signal_8675) ) ;
    buf_clk new_AGEMA_reg_buffer_5218 ( .C (clk), .D (new_AGEMA_signal_8682), .Q (new_AGEMA_signal_8683) ) ;
    buf_clk new_AGEMA_reg_buffer_5226 ( .C (clk), .D (new_AGEMA_signal_8690), .Q (new_AGEMA_signal_8691) ) ;
    buf_clk new_AGEMA_reg_buffer_5234 ( .C (clk), .D (new_AGEMA_signal_8698), .Q (new_AGEMA_signal_8699) ) ;
    buf_clk new_AGEMA_reg_buffer_5242 ( .C (clk), .D (new_AGEMA_signal_8706), .Q (new_AGEMA_signal_8707) ) ;
    buf_clk new_AGEMA_reg_buffer_5250 ( .C (clk), .D (new_AGEMA_signal_8714), .Q (new_AGEMA_signal_8715) ) ;
    buf_clk new_AGEMA_reg_buffer_5258 ( .C (clk), .D (new_AGEMA_signal_8722), .Q (new_AGEMA_signal_8723) ) ;
    buf_clk new_AGEMA_reg_buffer_5266 ( .C (clk), .D (new_AGEMA_signal_8730), .Q (new_AGEMA_signal_8731) ) ;
    buf_clk new_AGEMA_reg_buffer_5274 ( .C (clk), .D (new_AGEMA_signal_8738), .Q (new_AGEMA_signal_8739) ) ;
    buf_clk new_AGEMA_reg_buffer_5282 ( .C (clk), .D (new_AGEMA_signal_8746), .Q (new_AGEMA_signal_8747) ) ;
    buf_clk new_AGEMA_reg_buffer_5290 ( .C (clk), .D (new_AGEMA_signal_8754), .Q (new_AGEMA_signal_8755) ) ;
    buf_clk new_AGEMA_reg_buffer_5298 ( .C (clk), .D (new_AGEMA_signal_8762), .Q (new_AGEMA_signal_8763) ) ;
    buf_clk new_AGEMA_reg_buffer_5306 ( .C (clk), .D (new_AGEMA_signal_8770), .Q (new_AGEMA_signal_8771) ) ;
    buf_clk new_AGEMA_reg_buffer_5314 ( .C (clk), .D (new_AGEMA_signal_8778), .Q (new_AGEMA_signal_8779) ) ;
    buf_clk new_AGEMA_reg_buffer_5322 ( .C (clk), .D (new_AGEMA_signal_8786), .Q (new_AGEMA_signal_8787) ) ;
    buf_clk new_AGEMA_reg_buffer_5330 ( .C (clk), .D (new_AGEMA_signal_8794), .Q (new_AGEMA_signal_8795) ) ;
    buf_clk new_AGEMA_reg_buffer_5338 ( .C (clk), .D (new_AGEMA_signal_8802), .Q (new_AGEMA_signal_8803) ) ;
    buf_clk new_AGEMA_reg_buffer_5346 ( .C (clk), .D (new_AGEMA_signal_8810), .Q (new_AGEMA_signal_8811) ) ;
    buf_clk new_AGEMA_reg_buffer_5354 ( .C (clk), .D (new_AGEMA_signal_8818), .Q (new_AGEMA_signal_8819) ) ;
    buf_clk new_AGEMA_reg_buffer_5362 ( .C (clk), .D (new_AGEMA_signal_8826), .Q (new_AGEMA_signal_8827) ) ;
    buf_clk new_AGEMA_reg_buffer_5370 ( .C (clk), .D (new_AGEMA_signal_8834), .Q (new_AGEMA_signal_8835) ) ;
    buf_clk new_AGEMA_reg_buffer_5378 ( .C (clk), .D (new_AGEMA_signal_8842), .Q (new_AGEMA_signal_8843) ) ;
    buf_clk new_AGEMA_reg_buffer_5386 ( .C (clk), .D (new_AGEMA_signal_8850), .Q (new_AGEMA_signal_8851) ) ;
    buf_clk new_AGEMA_reg_buffer_5394 ( .C (clk), .D (new_AGEMA_signal_8858), .Q (new_AGEMA_signal_8859) ) ;
    buf_clk new_AGEMA_reg_buffer_5402 ( .C (clk), .D (new_AGEMA_signal_8866), .Q (new_AGEMA_signal_8867) ) ;
    buf_clk new_AGEMA_reg_buffer_5404 ( .C (clk), .D (new_AGEMA_signal_8868), .Q (new_AGEMA_signal_8869) ) ;
    buf_clk new_AGEMA_reg_buffer_5412 ( .C (clk), .D (new_AGEMA_signal_8876), .Q (new_AGEMA_signal_8877) ) ;
    buf_clk new_AGEMA_reg_buffer_5420 ( .C (clk), .D (new_AGEMA_signal_8884), .Q (new_AGEMA_signal_8885) ) ;
    buf_clk new_AGEMA_reg_buffer_5428 ( .C (clk), .D (new_AGEMA_signal_8892), .Q (new_AGEMA_signal_8893) ) ;
    buf_clk new_AGEMA_reg_buffer_5436 ( .C (clk), .D (new_AGEMA_signal_8900), .Q (new_AGEMA_signal_8901) ) ;
    buf_clk new_AGEMA_reg_buffer_5444 ( .C (clk), .D (new_AGEMA_signal_8908), .Q (new_AGEMA_signal_8909) ) ;
    buf_clk new_AGEMA_reg_buffer_5452 ( .C (clk), .D (new_AGEMA_signal_8916), .Q (new_AGEMA_signal_8917) ) ;
    buf_clk new_AGEMA_reg_buffer_5460 ( .C (clk), .D (new_AGEMA_signal_8924), .Q (new_AGEMA_signal_8925) ) ;
    buf_clk new_AGEMA_reg_buffer_5468 ( .C (clk), .D (new_AGEMA_signal_8932), .Q (new_AGEMA_signal_8933) ) ;
    buf_clk new_AGEMA_reg_buffer_5476 ( .C (clk), .D (new_AGEMA_signal_8940), .Q (new_AGEMA_signal_8941) ) ;
    buf_clk new_AGEMA_reg_buffer_5484 ( .C (clk), .D (new_AGEMA_signal_8948), .Q (new_AGEMA_signal_8949) ) ;
    buf_clk new_AGEMA_reg_buffer_5492 ( .C (clk), .D (new_AGEMA_signal_8956), .Q (new_AGEMA_signal_8957) ) ;
    buf_clk new_AGEMA_reg_buffer_5500 ( .C (clk), .D (new_AGEMA_signal_8964), .Q (new_AGEMA_signal_8965) ) ;
    buf_clk new_AGEMA_reg_buffer_5508 ( .C (clk), .D (new_AGEMA_signal_8972), .Q (new_AGEMA_signal_8973) ) ;
    buf_clk new_AGEMA_reg_buffer_5516 ( .C (clk), .D (new_AGEMA_signal_8980), .Q (new_AGEMA_signal_8981) ) ;
    buf_clk new_AGEMA_reg_buffer_5524 ( .C (clk), .D (new_AGEMA_signal_8988), .Q (new_AGEMA_signal_8989) ) ;
    buf_clk new_AGEMA_reg_buffer_5532 ( .C (clk), .D (new_AGEMA_signal_8996), .Q (new_AGEMA_signal_8997) ) ;
    buf_clk new_AGEMA_reg_buffer_5540 ( .C (clk), .D (new_AGEMA_signal_9004), .Q (new_AGEMA_signal_9005) ) ;
    buf_clk new_AGEMA_reg_buffer_5548 ( .C (clk), .D (new_AGEMA_signal_9012), .Q (new_AGEMA_signal_9013) ) ;
    buf_clk new_AGEMA_reg_buffer_5556 ( .C (clk), .D (new_AGEMA_signal_9020), .Q (new_AGEMA_signal_9021) ) ;
    buf_clk new_AGEMA_reg_buffer_5564 ( .C (clk), .D (new_AGEMA_signal_9028), .Q (new_AGEMA_signal_9029) ) ;
    buf_clk new_AGEMA_reg_buffer_5572 ( .C (clk), .D (new_AGEMA_signal_9036), .Q (new_AGEMA_signal_9037) ) ;
    buf_clk new_AGEMA_reg_buffer_5580 ( .C (clk), .D (new_AGEMA_signal_9044), .Q (new_AGEMA_signal_9045) ) ;
    buf_clk new_AGEMA_reg_buffer_5588 ( .C (clk), .D (new_AGEMA_signal_9052), .Q (new_AGEMA_signal_9053) ) ;
    buf_clk new_AGEMA_reg_buffer_5596 ( .C (clk), .D (new_AGEMA_signal_9060), .Q (new_AGEMA_signal_9061) ) ;
    buf_clk new_AGEMA_reg_buffer_5604 ( .C (clk), .D (new_AGEMA_signal_9068), .Q (new_AGEMA_signal_9069) ) ;
    buf_clk new_AGEMA_reg_buffer_5612 ( .C (clk), .D (new_AGEMA_signal_9076), .Q (new_AGEMA_signal_9077) ) ;
    buf_clk new_AGEMA_reg_buffer_5620 ( .C (clk), .D (new_AGEMA_signal_9084), .Q (new_AGEMA_signal_9085) ) ;
    buf_clk new_AGEMA_reg_buffer_5628 ( .C (clk), .D (new_AGEMA_signal_9092), .Q (new_AGEMA_signal_9093) ) ;
    buf_clk new_AGEMA_reg_buffer_5636 ( .C (clk), .D (new_AGEMA_signal_9100), .Q (new_AGEMA_signal_9101) ) ;
    buf_clk new_AGEMA_reg_buffer_5644 ( .C (clk), .D (new_AGEMA_signal_9108), .Q (new_AGEMA_signal_9109) ) ;
    buf_clk new_AGEMA_reg_buffer_5652 ( .C (clk), .D (new_AGEMA_signal_9116), .Q (new_AGEMA_signal_9117) ) ;
    buf_clk new_AGEMA_reg_buffer_5660 ( .C (clk), .D (new_AGEMA_signal_9124), .Q (new_AGEMA_signal_9125) ) ;
    buf_clk new_AGEMA_reg_buffer_5668 ( .C (clk), .D (new_AGEMA_signal_9132), .Q (new_AGEMA_signal_9133) ) ;
    buf_clk new_AGEMA_reg_buffer_5676 ( .C (clk), .D (new_AGEMA_signal_9140), .Q (new_AGEMA_signal_9141) ) ;
    buf_clk new_AGEMA_reg_buffer_5684 ( .C (clk), .D (new_AGEMA_signal_9148), .Q (new_AGEMA_signal_9149) ) ;
    buf_clk new_AGEMA_reg_buffer_5692 ( .C (clk), .D (new_AGEMA_signal_9156), .Q (new_AGEMA_signal_9157) ) ;
    buf_clk new_AGEMA_reg_buffer_5700 ( .C (clk), .D (new_AGEMA_signal_9164), .Q (new_AGEMA_signal_9165) ) ;
    buf_clk new_AGEMA_reg_buffer_5708 ( .C (clk), .D (new_AGEMA_signal_9172), .Q (new_AGEMA_signal_9173) ) ;
    buf_clk new_AGEMA_reg_buffer_5716 ( .C (clk), .D (new_AGEMA_signal_9180), .Q (new_AGEMA_signal_9181) ) ;
    buf_clk new_AGEMA_reg_buffer_5724 ( .C (clk), .D (new_AGEMA_signal_9188), .Q (new_AGEMA_signal_9189) ) ;
    buf_clk new_AGEMA_reg_buffer_5732 ( .C (clk), .D (new_AGEMA_signal_9196), .Q (new_AGEMA_signal_9197) ) ;
    buf_clk new_AGEMA_reg_buffer_5740 ( .C (clk), .D (new_AGEMA_signal_9204), .Q (new_AGEMA_signal_9205) ) ;
    buf_clk new_AGEMA_reg_buffer_5748 ( .C (clk), .D (new_AGEMA_signal_9212), .Q (new_AGEMA_signal_9213) ) ;
    buf_clk new_AGEMA_reg_buffer_5756 ( .C (clk), .D (new_AGEMA_signal_9220), .Q (new_AGEMA_signal_9221) ) ;
    buf_clk new_AGEMA_reg_buffer_5764 ( .C (clk), .D (new_AGEMA_signal_9228), .Q (new_AGEMA_signal_9229) ) ;
    buf_clk new_AGEMA_reg_buffer_5772 ( .C (clk), .D (new_AGEMA_signal_9236), .Q (new_AGEMA_signal_9237) ) ;
    buf_clk new_AGEMA_reg_buffer_5780 ( .C (clk), .D (new_AGEMA_signal_9244), .Q (new_AGEMA_signal_9245) ) ;
    buf_clk new_AGEMA_reg_buffer_5788 ( .C (clk), .D (new_AGEMA_signal_9252), .Q (new_AGEMA_signal_9253) ) ;
    buf_clk new_AGEMA_reg_buffer_5796 ( .C (clk), .D (new_AGEMA_signal_9260), .Q (new_AGEMA_signal_9261) ) ;
    buf_clk new_AGEMA_reg_buffer_5804 ( .C (clk), .D (new_AGEMA_signal_9268), .Q (new_AGEMA_signal_9269) ) ;
    buf_clk new_AGEMA_reg_buffer_5812 ( .C (clk), .D (new_AGEMA_signal_9276), .Q (new_AGEMA_signal_9277) ) ;
    buf_clk new_AGEMA_reg_buffer_5820 ( .C (clk), .D (new_AGEMA_signal_9284), .Q (new_AGEMA_signal_9285) ) ;
    buf_clk new_AGEMA_reg_buffer_5828 ( .C (clk), .D (new_AGEMA_signal_9292), .Q (new_AGEMA_signal_9293) ) ;
    buf_clk new_AGEMA_reg_buffer_5836 ( .C (clk), .D (new_AGEMA_signal_9300), .Q (new_AGEMA_signal_9301) ) ;
    buf_clk new_AGEMA_reg_buffer_5844 ( .C (clk), .D (new_AGEMA_signal_9308), .Q (new_AGEMA_signal_9309) ) ;
    buf_clk new_AGEMA_reg_buffer_5852 ( .C (clk), .D (new_AGEMA_signal_9316), .Q (new_AGEMA_signal_9317) ) ;
    buf_clk new_AGEMA_reg_buffer_5860 ( .C (clk), .D (new_AGEMA_signal_9324), .Q (new_AGEMA_signal_9325) ) ;
    buf_clk new_AGEMA_reg_buffer_5868 ( .C (clk), .D (new_AGEMA_signal_9332), .Q (new_AGEMA_signal_9333) ) ;
    buf_clk new_AGEMA_reg_buffer_5876 ( .C (clk), .D (new_AGEMA_signal_9340), .Q (new_AGEMA_signal_9341) ) ;
    buf_clk new_AGEMA_reg_buffer_5884 ( .C (clk), .D (new_AGEMA_signal_9348), .Q (new_AGEMA_signal_9349) ) ;
    buf_clk new_AGEMA_reg_buffer_5892 ( .C (clk), .D (new_AGEMA_signal_9356), .Q (new_AGEMA_signal_9357) ) ;
    buf_clk new_AGEMA_reg_buffer_5900 ( .C (clk), .D (new_AGEMA_signal_9364), .Q (new_AGEMA_signal_9365) ) ;
    buf_clk new_AGEMA_reg_buffer_5908 ( .C (clk), .D (new_AGEMA_signal_9372), .Q (new_AGEMA_signal_9373) ) ;
    buf_clk new_AGEMA_reg_buffer_5916 ( .C (clk), .D (new_AGEMA_signal_9380), .Q (new_AGEMA_signal_9381) ) ;
    buf_clk new_AGEMA_reg_buffer_5924 ( .C (clk), .D (new_AGEMA_signal_9388), .Q (new_AGEMA_signal_9389) ) ;
    buf_clk new_AGEMA_reg_buffer_5932 ( .C (clk), .D (new_AGEMA_signal_9396), .Q (new_AGEMA_signal_9397) ) ;
    buf_clk new_AGEMA_reg_buffer_5940 ( .C (clk), .D (new_AGEMA_signal_9404), .Q (new_AGEMA_signal_9405) ) ;
    buf_clk new_AGEMA_reg_buffer_5948 ( .C (clk), .D (new_AGEMA_signal_9412), .Q (new_AGEMA_signal_9413) ) ;
    buf_clk new_AGEMA_reg_buffer_5956 ( .C (clk), .D (new_AGEMA_signal_9420), .Q (new_AGEMA_signal_9421) ) ;
    buf_clk new_AGEMA_reg_buffer_5964 ( .C (clk), .D (new_AGEMA_signal_9428), .Q (new_AGEMA_signal_9429) ) ;
    buf_clk new_AGEMA_reg_buffer_5972 ( .C (clk), .D (new_AGEMA_signal_9436), .Q (new_AGEMA_signal_9437) ) ;
    buf_clk new_AGEMA_reg_buffer_5980 ( .C (clk), .D (new_AGEMA_signal_9444), .Q (new_AGEMA_signal_9445) ) ;
    buf_clk new_AGEMA_reg_buffer_5988 ( .C (clk), .D (new_AGEMA_signal_9452), .Q (new_AGEMA_signal_9453) ) ;
    buf_clk new_AGEMA_reg_buffer_5996 ( .C (clk), .D (new_AGEMA_signal_9460), .Q (new_AGEMA_signal_9461) ) ;
    buf_clk new_AGEMA_reg_buffer_6004 ( .C (clk), .D (new_AGEMA_signal_9468), .Q (new_AGEMA_signal_9469) ) ;
    buf_clk new_AGEMA_reg_buffer_6012 ( .C (clk), .D (new_AGEMA_signal_9476), .Q (new_AGEMA_signal_9477) ) ;
    buf_clk new_AGEMA_reg_buffer_6020 ( .C (clk), .D (new_AGEMA_signal_9484), .Q (new_AGEMA_signal_9485) ) ;
    buf_clk new_AGEMA_reg_buffer_6028 ( .C (clk), .D (new_AGEMA_signal_9492), .Q (new_AGEMA_signal_9493) ) ;
    buf_clk new_AGEMA_reg_buffer_6036 ( .C (clk), .D (new_AGEMA_signal_9500), .Q (new_AGEMA_signal_9501) ) ;
    buf_clk new_AGEMA_reg_buffer_6044 ( .C (clk), .D (new_AGEMA_signal_9508), .Q (new_AGEMA_signal_9509) ) ;
    buf_clk new_AGEMA_reg_buffer_6052 ( .C (clk), .D (new_AGEMA_signal_9516), .Q (new_AGEMA_signal_9517) ) ;
    buf_clk new_AGEMA_reg_buffer_6060 ( .C (clk), .D (new_AGEMA_signal_9524), .Q (new_AGEMA_signal_9525) ) ;
    buf_clk new_AGEMA_reg_buffer_6068 ( .C (clk), .D (new_AGEMA_signal_9532), .Q (new_AGEMA_signal_9533) ) ;
    buf_clk new_AGEMA_reg_buffer_6076 ( .C (clk), .D (new_AGEMA_signal_9540), .Q (new_AGEMA_signal_9541) ) ;
    buf_clk new_AGEMA_reg_buffer_6084 ( .C (clk), .D (new_AGEMA_signal_9548), .Q (new_AGEMA_signal_9549) ) ;
    buf_clk new_AGEMA_reg_buffer_6092 ( .C (clk), .D (new_AGEMA_signal_9556), .Q (new_AGEMA_signal_9557) ) ;
    buf_clk new_AGEMA_reg_buffer_6100 ( .C (clk), .D (new_AGEMA_signal_9564), .Q (new_AGEMA_signal_9565) ) ;
    buf_clk new_AGEMA_reg_buffer_6108 ( .C (clk), .D (new_AGEMA_signal_9572), .Q (new_AGEMA_signal_9573) ) ;
    buf_clk new_AGEMA_reg_buffer_6116 ( .C (clk), .D (new_AGEMA_signal_9580), .Q (new_AGEMA_signal_9581) ) ;
    buf_clk new_AGEMA_reg_buffer_6124 ( .C (clk), .D (new_AGEMA_signal_9588), .Q (new_AGEMA_signal_9589) ) ;
    buf_clk new_AGEMA_reg_buffer_6132 ( .C (clk), .D (new_AGEMA_signal_9596), .Q (new_AGEMA_signal_9597) ) ;
    buf_clk new_AGEMA_reg_buffer_6140 ( .C (clk), .D (new_AGEMA_signal_9604), .Q (new_AGEMA_signal_9605) ) ;
    buf_clk new_AGEMA_reg_buffer_6148 ( .C (clk), .D (new_AGEMA_signal_9612), .Q (new_AGEMA_signal_9613) ) ;
    buf_clk new_AGEMA_reg_buffer_6156 ( .C (clk), .D (new_AGEMA_signal_9620), .Q (new_AGEMA_signal_9621) ) ;
    buf_clk new_AGEMA_reg_buffer_6164 ( .C (clk), .D (new_AGEMA_signal_9628), .Q (new_AGEMA_signal_9629) ) ;
    buf_clk new_AGEMA_reg_buffer_6172 ( .C (clk), .D (new_AGEMA_signal_9636), .Q (new_AGEMA_signal_9637) ) ;
    buf_clk new_AGEMA_reg_buffer_6462 ( .C (clk), .D (new_AGEMA_signal_9926), .Q (new_AGEMA_signal_9927) ) ;
    buf_clk new_AGEMA_reg_buffer_6470 ( .C (clk), .D (new_AGEMA_signal_9934), .Q (new_AGEMA_signal_9935) ) ;
    buf_clk new_AGEMA_reg_buffer_6478 ( .C (clk), .D (new_AGEMA_signal_9942), .Q (new_AGEMA_signal_9943) ) ;
    buf_clk new_AGEMA_reg_buffer_6486 ( .C (clk), .D (new_AGEMA_signal_9950), .Q (new_AGEMA_signal_9951) ) ;
    buf_clk new_AGEMA_reg_buffer_6494 ( .C (clk), .D (new_AGEMA_signal_9958), .Q (new_AGEMA_signal_9959) ) ;
    buf_clk new_AGEMA_reg_buffer_6496 ( .C (clk), .D (new_AGEMA_signal_9960), .Q (new_AGEMA_signal_9961) ) ;
    buf_clk new_AGEMA_reg_buffer_6498 ( .C (clk), .D (new_AGEMA_signal_9962), .Q (new_AGEMA_signal_9963) ) ;
    buf_clk new_AGEMA_reg_buffer_6500 ( .C (clk), .D (new_AGEMA_signal_9964), .Q (new_AGEMA_signal_9965) ) ;
    buf_clk new_AGEMA_reg_buffer_6502 ( .C (clk), .D (new_AGEMA_signal_9966), .Q (new_AGEMA_signal_9967) ) ;
    buf_clk new_AGEMA_reg_buffer_6504 ( .C (clk), .D (new_AGEMA_signal_9968), .Q (new_AGEMA_signal_9969) ) ;
    buf_clk new_AGEMA_reg_buffer_6506 ( .C (clk), .D (new_AGEMA_signal_9970), .Q (new_AGEMA_signal_9971) ) ;
    buf_clk new_AGEMA_reg_buffer_6508 ( .C (clk), .D (new_AGEMA_signal_9972), .Q (new_AGEMA_signal_9973) ) ;
    buf_clk new_AGEMA_reg_buffer_6510 ( .C (clk), .D (new_AGEMA_signal_9974), .Q (new_AGEMA_signal_9975) ) ;
    buf_clk new_AGEMA_reg_buffer_6512 ( .C (clk), .D (new_AGEMA_signal_9976), .Q (new_AGEMA_signal_9977) ) ;
    buf_clk new_AGEMA_reg_buffer_6514 ( .C (clk), .D (new_AGEMA_signal_9978), .Q (new_AGEMA_signal_9979) ) ;
    buf_clk new_AGEMA_reg_buffer_6516 ( .C (clk), .D (new_AGEMA_signal_9980), .Q (new_AGEMA_signal_9981) ) ;
    buf_clk new_AGEMA_reg_buffer_6518 ( .C (clk), .D (new_AGEMA_signal_9982), .Q (new_AGEMA_signal_9983) ) ;
    buf_clk new_AGEMA_reg_buffer_6520 ( .C (clk), .D (new_AGEMA_signal_9984), .Q (new_AGEMA_signal_9985) ) ;
    buf_clk new_AGEMA_reg_buffer_6522 ( .C (clk), .D (new_AGEMA_signal_9986), .Q (new_AGEMA_signal_9987) ) ;
    buf_clk new_AGEMA_reg_buffer_6524 ( .C (clk), .D (new_AGEMA_signal_9988), .Q (new_AGEMA_signal_9989) ) ;
    buf_clk new_AGEMA_reg_buffer_6526 ( .C (clk), .D (new_AGEMA_signal_9990), .Q (new_AGEMA_signal_9991) ) ;
    buf_clk new_AGEMA_reg_buffer_6528 ( .C (clk), .D (new_AGEMA_signal_9992), .Q (new_AGEMA_signal_9993) ) ;
    buf_clk new_AGEMA_reg_buffer_6530 ( .C (clk), .D (new_AGEMA_signal_9994), .Q (new_AGEMA_signal_9995) ) ;
    buf_clk new_AGEMA_reg_buffer_6532 ( .C (clk), .D (new_AGEMA_signal_9996), .Q (new_AGEMA_signal_9997) ) ;
    buf_clk new_AGEMA_reg_buffer_6534 ( .C (clk), .D (new_AGEMA_signal_9998), .Q (new_AGEMA_signal_9999) ) ;
    buf_clk new_AGEMA_reg_buffer_6536 ( .C (clk), .D (new_AGEMA_signal_10000), .Q (new_AGEMA_signal_10001) ) ;
    buf_clk new_AGEMA_reg_buffer_6538 ( .C (clk), .D (new_AGEMA_signal_10002), .Q (new_AGEMA_signal_10003) ) ;
    buf_clk new_AGEMA_reg_buffer_6540 ( .C (clk), .D (new_AGEMA_signal_10004), .Q (new_AGEMA_signal_10005) ) ;
    buf_clk new_AGEMA_reg_buffer_6542 ( .C (clk), .D (new_AGEMA_signal_10006), .Q (new_AGEMA_signal_10007) ) ;
    buf_clk new_AGEMA_reg_buffer_6544 ( .C (clk), .D (new_AGEMA_signal_10008), .Q (new_AGEMA_signal_10009) ) ;
    buf_clk new_AGEMA_reg_buffer_6546 ( .C (clk), .D (new_AGEMA_signal_10010), .Q (new_AGEMA_signal_10011) ) ;
    buf_clk new_AGEMA_reg_buffer_6548 ( .C (clk), .D (new_AGEMA_signal_10012), .Q (new_AGEMA_signal_10013) ) ;
    buf_clk new_AGEMA_reg_buffer_6550 ( .C (clk), .D (new_AGEMA_signal_10014), .Q (new_AGEMA_signal_10015) ) ;
    buf_clk new_AGEMA_reg_buffer_6552 ( .C (clk), .D (new_AGEMA_signal_10016), .Q (new_AGEMA_signal_10017) ) ;
    buf_clk new_AGEMA_reg_buffer_6554 ( .C (clk), .D (new_AGEMA_signal_10018), .Q (new_AGEMA_signal_10019) ) ;
    buf_clk new_AGEMA_reg_buffer_6556 ( .C (clk), .D (new_AGEMA_signal_10020), .Q (new_AGEMA_signal_10021) ) ;
    buf_clk new_AGEMA_reg_buffer_6558 ( .C (clk), .D (new_AGEMA_signal_10022), .Q (new_AGEMA_signal_10023) ) ;
    buf_clk new_AGEMA_reg_buffer_6560 ( .C (clk), .D (new_AGEMA_signal_10024), .Q (new_AGEMA_signal_10025) ) ;
    buf_clk new_AGEMA_reg_buffer_6562 ( .C (clk), .D (new_AGEMA_signal_10026), .Q (new_AGEMA_signal_10027) ) ;
    buf_clk new_AGEMA_reg_buffer_6564 ( .C (clk), .D (new_AGEMA_signal_10028), .Q (new_AGEMA_signal_10029) ) ;
    buf_clk new_AGEMA_reg_buffer_6566 ( .C (clk), .D (new_AGEMA_signal_10030), .Q (new_AGEMA_signal_10031) ) ;
    buf_clk new_AGEMA_reg_buffer_6568 ( .C (clk), .D (new_AGEMA_signal_10032), .Q (new_AGEMA_signal_10033) ) ;
    buf_clk new_AGEMA_reg_buffer_6570 ( .C (clk), .D (new_AGEMA_signal_10034), .Q (new_AGEMA_signal_10035) ) ;
    buf_clk new_AGEMA_reg_buffer_6572 ( .C (clk), .D (new_AGEMA_signal_10036), .Q (new_AGEMA_signal_10037) ) ;
    buf_clk new_AGEMA_reg_buffer_6574 ( .C (clk), .D (new_AGEMA_signal_10038), .Q (new_AGEMA_signal_10039) ) ;
    buf_clk new_AGEMA_reg_buffer_6576 ( .C (clk), .D (new_AGEMA_signal_10040), .Q (new_AGEMA_signal_10041) ) ;
    buf_clk new_AGEMA_reg_buffer_6578 ( .C (clk), .D (new_AGEMA_signal_10042), .Q (new_AGEMA_signal_10043) ) ;
    buf_clk new_AGEMA_reg_buffer_6580 ( .C (clk), .D (new_AGEMA_signal_10044), .Q (new_AGEMA_signal_10045) ) ;
    buf_clk new_AGEMA_reg_buffer_6582 ( .C (clk), .D (new_AGEMA_signal_10046), .Q (new_AGEMA_signal_10047) ) ;
    buf_clk new_AGEMA_reg_buffer_6584 ( .C (clk), .D (new_AGEMA_signal_10048), .Q (new_AGEMA_signal_10049) ) ;
    buf_clk new_AGEMA_reg_buffer_6586 ( .C (clk), .D (new_AGEMA_signal_10050), .Q (new_AGEMA_signal_10051) ) ;
    buf_clk new_AGEMA_reg_buffer_6588 ( .C (clk), .D (new_AGEMA_signal_10052), .Q (new_AGEMA_signal_10053) ) ;
    buf_clk new_AGEMA_reg_buffer_6590 ( .C (clk), .D (new_AGEMA_signal_10054), .Q (new_AGEMA_signal_10055) ) ;
    buf_clk new_AGEMA_reg_buffer_6592 ( .C (clk), .D (new_AGEMA_signal_10056), .Q (new_AGEMA_signal_10057) ) ;
    buf_clk new_AGEMA_reg_buffer_6594 ( .C (clk), .D (new_AGEMA_signal_10058), .Q (new_AGEMA_signal_10059) ) ;
    buf_clk new_AGEMA_reg_buffer_6596 ( .C (clk), .D (new_AGEMA_signal_10060), .Q (new_AGEMA_signal_10061) ) ;
    buf_clk new_AGEMA_reg_buffer_6598 ( .C (clk), .D (new_AGEMA_signal_10062), .Q (new_AGEMA_signal_10063) ) ;
    buf_clk new_AGEMA_reg_buffer_6600 ( .C (clk), .D (new_AGEMA_signal_10064), .Q (new_AGEMA_signal_10065) ) ;
    buf_clk new_AGEMA_reg_buffer_6602 ( .C (clk), .D (new_AGEMA_signal_10066), .Q (new_AGEMA_signal_10067) ) ;
    buf_clk new_AGEMA_reg_buffer_6604 ( .C (clk), .D (new_AGEMA_signal_10068), .Q (new_AGEMA_signal_10069) ) ;
    buf_clk new_AGEMA_reg_buffer_6606 ( .C (clk), .D (new_AGEMA_signal_10070), .Q (new_AGEMA_signal_10071) ) ;
    buf_clk new_AGEMA_reg_buffer_6608 ( .C (clk), .D (new_AGEMA_signal_10072), .Q (new_AGEMA_signal_10073) ) ;
    buf_clk new_AGEMA_reg_buffer_6610 ( .C (clk), .D (new_AGEMA_signal_10074), .Q (new_AGEMA_signal_10075) ) ;
    buf_clk new_AGEMA_reg_buffer_6612 ( .C (clk), .D (new_AGEMA_signal_10076), .Q (new_AGEMA_signal_10077) ) ;
    buf_clk new_AGEMA_reg_buffer_6614 ( .C (clk), .D (new_AGEMA_signal_10078), .Q (new_AGEMA_signal_10079) ) ;
    buf_clk new_AGEMA_reg_buffer_6616 ( .C (clk), .D (new_AGEMA_signal_10080), .Q (new_AGEMA_signal_10081) ) ;
    buf_clk new_AGEMA_reg_buffer_6618 ( .C (clk), .D (new_AGEMA_signal_10082), .Q (new_AGEMA_signal_10083) ) ;
    buf_clk new_AGEMA_reg_buffer_6620 ( .C (clk), .D (new_AGEMA_signal_10084), .Q (new_AGEMA_signal_10085) ) ;
    buf_clk new_AGEMA_reg_buffer_6622 ( .C (clk), .D (new_AGEMA_signal_10086), .Q (new_AGEMA_signal_10087) ) ;
    buf_clk new_AGEMA_reg_buffer_6624 ( .C (clk), .D (new_AGEMA_signal_10088), .Q (new_AGEMA_signal_10089) ) ;
    buf_clk new_AGEMA_reg_buffer_6626 ( .C (clk), .D (new_AGEMA_signal_10090), .Q (new_AGEMA_signal_10091) ) ;
    buf_clk new_AGEMA_reg_buffer_6628 ( .C (clk), .D (new_AGEMA_signal_10092), .Q (new_AGEMA_signal_10093) ) ;
    buf_clk new_AGEMA_reg_buffer_6630 ( .C (clk), .D (new_AGEMA_signal_10094), .Q (new_AGEMA_signal_10095) ) ;
    buf_clk new_AGEMA_reg_buffer_6632 ( .C (clk), .D (new_AGEMA_signal_10096), .Q (new_AGEMA_signal_10097) ) ;
    buf_clk new_AGEMA_reg_buffer_6634 ( .C (clk), .D (new_AGEMA_signal_10098), .Q (new_AGEMA_signal_10099) ) ;
    buf_clk new_AGEMA_reg_buffer_6636 ( .C (clk), .D (new_AGEMA_signal_10100), .Q (new_AGEMA_signal_10101) ) ;
    buf_clk new_AGEMA_reg_buffer_6638 ( .C (clk), .D (new_AGEMA_signal_10102), .Q (new_AGEMA_signal_10103) ) ;
    buf_clk new_AGEMA_reg_buffer_6640 ( .C (clk), .D (new_AGEMA_signal_10104), .Q (new_AGEMA_signal_10105) ) ;
    buf_clk new_AGEMA_reg_buffer_6642 ( .C (clk), .D (new_AGEMA_signal_10106), .Q (new_AGEMA_signal_10107) ) ;
    buf_clk new_AGEMA_reg_buffer_6644 ( .C (clk), .D (new_AGEMA_signal_10108), .Q (new_AGEMA_signal_10109) ) ;
    buf_clk new_AGEMA_reg_buffer_6646 ( .C (clk), .D (new_AGEMA_signal_10110), .Q (new_AGEMA_signal_10111) ) ;
    buf_clk new_AGEMA_reg_buffer_6648 ( .C (clk), .D (new_AGEMA_signal_10112), .Q (new_AGEMA_signal_10113) ) ;
    buf_clk new_AGEMA_reg_buffer_6650 ( .C (clk), .D (new_AGEMA_signal_10114), .Q (new_AGEMA_signal_10115) ) ;
    buf_clk new_AGEMA_reg_buffer_6652 ( .C (clk), .D (new_AGEMA_signal_10116), .Q (new_AGEMA_signal_10117) ) ;
    buf_clk new_AGEMA_reg_buffer_6654 ( .C (clk), .D (new_AGEMA_signal_10118), .Q (new_AGEMA_signal_10119) ) ;
    buf_clk new_AGEMA_reg_buffer_6656 ( .C (clk), .D (new_AGEMA_signal_10120), .Q (new_AGEMA_signal_10121) ) ;
    buf_clk new_AGEMA_reg_buffer_6658 ( .C (clk), .D (new_AGEMA_signal_10122), .Q (new_AGEMA_signal_10123) ) ;
    buf_clk new_AGEMA_reg_buffer_6660 ( .C (clk), .D (new_AGEMA_signal_10124), .Q (new_AGEMA_signal_10125) ) ;
    buf_clk new_AGEMA_reg_buffer_6662 ( .C (clk), .D (new_AGEMA_signal_10126), .Q (new_AGEMA_signal_10127) ) ;
    buf_clk new_AGEMA_reg_buffer_6664 ( .C (clk), .D (new_AGEMA_signal_10128), .Q (new_AGEMA_signal_10129) ) ;
    buf_clk new_AGEMA_reg_buffer_6666 ( .C (clk), .D (new_AGEMA_signal_10130), .Q (new_AGEMA_signal_10131) ) ;
    buf_clk new_AGEMA_reg_buffer_6668 ( .C (clk), .D (new_AGEMA_signal_10132), .Q (new_AGEMA_signal_10133) ) ;
    buf_clk new_AGEMA_reg_buffer_6670 ( .C (clk), .D (new_AGEMA_signal_10134), .Q (new_AGEMA_signal_10135) ) ;
    buf_clk new_AGEMA_reg_buffer_6672 ( .C (clk), .D (new_AGEMA_signal_10136), .Q (new_AGEMA_signal_10137) ) ;
    buf_clk new_AGEMA_reg_buffer_6674 ( .C (clk), .D (new_AGEMA_signal_10138), .Q (new_AGEMA_signal_10139) ) ;
    buf_clk new_AGEMA_reg_buffer_6676 ( .C (clk), .D (new_AGEMA_signal_10140), .Q (new_AGEMA_signal_10141) ) ;
    buf_clk new_AGEMA_reg_buffer_6678 ( .C (clk), .D (new_AGEMA_signal_10142), .Q (new_AGEMA_signal_10143) ) ;
    buf_clk new_AGEMA_reg_buffer_6680 ( .C (clk), .D (new_AGEMA_signal_10144), .Q (new_AGEMA_signal_10145) ) ;
    buf_clk new_AGEMA_reg_buffer_6682 ( .C (clk), .D (new_AGEMA_signal_10146), .Q (new_AGEMA_signal_10147) ) ;
    buf_clk new_AGEMA_reg_buffer_6684 ( .C (clk), .D (new_AGEMA_signal_10148), .Q (new_AGEMA_signal_10149) ) ;
    buf_clk new_AGEMA_reg_buffer_6686 ( .C (clk), .D (new_AGEMA_signal_10150), .Q (new_AGEMA_signal_10151) ) ;

    /* register cells */
    DFF_X1 controller_roundCounter_count_reg_0__FF_FF ( .CK (clk), .D (new_AGEMA_signal_9935), .Q (round_Signal[0]), .QN () ) ;
    DFF_X1 controller_roundCounter_count_reg_1__FF_FF ( .CK (clk), .D (new_AGEMA_signal_9943), .Q (round_Signal[1]), .QN () ) ;
    DFF_X1 controller_roundCounter_count_reg_2__FF_FF ( .CK (clk), .D (new_AGEMA_signal_9951), .Q (round_Signal[2]), .QN () ) ;
    DFF_X1 controller_roundCounter_count_reg_3__FF_FF ( .CK (clk), .D (new_AGEMA_signal_9959), .Q (round_Signal[3]), .QN () ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3911, new_AGEMA_signal_3910, Midori_rounds_roundResult_Reg_SFF_0_DQ}), .Q ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, Midori_rounds_roundReg_out[0]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_9965, new_AGEMA_signal_9963, new_AGEMA_signal_9961}), .Q ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, Midori_rounds_roundReg_out[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, Midori_rounds_roundResult_Reg_SFF_2_DQ}), .Q ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, Midori_rounds_roundReg_out[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_9971, new_AGEMA_signal_9969, new_AGEMA_signal_9967}), .Q ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, Midori_rounds_roundReg_out[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3913, new_AGEMA_signal_3912, Midori_rounds_roundResult_Reg_SFF_4_DQ}), .Q ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, Midori_rounds_roundReg_out[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_9977, new_AGEMA_signal_9975, new_AGEMA_signal_9973}), .Q ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, Midori_rounds_roundReg_out[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3683, new_AGEMA_signal_3682, Midori_rounds_roundResult_Reg_SFF_6_DQ}), .Q ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, Midori_rounds_roundReg_out[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_9983, new_AGEMA_signal_9981, new_AGEMA_signal_9979}), .Q ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, Midori_rounds_roundReg_out[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_8_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3915, new_AGEMA_signal_3914, Midori_rounds_roundResult_Reg_SFF_8_DQ}), .Q ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, Midori_rounds_roundReg_out[8]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_9_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_9989, new_AGEMA_signal_9987, new_AGEMA_signal_9985}), .Q ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, Midori_rounds_roundReg_out[9]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_10_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, Midori_rounds_roundResult_Reg_SFF_10_DQ}), .Q ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, Midori_rounds_roundReg_out[10]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_11_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_9995, new_AGEMA_signal_9993, new_AGEMA_signal_9991}), .Q ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, Midori_rounds_roundReg_out[11]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_12_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3917, new_AGEMA_signal_3916, Midori_rounds_roundResult_Reg_SFF_12_DQ}), .Q ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, Midori_rounds_roundReg_out[12]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_13_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10001, new_AGEMA_signal_9999, new_AGEMA_signal_9997}), .Q ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, Midori_rounds_roundReg_out[13]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_14_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, Midori_rounds_roundResult_Reg_SFF_14_DQ}), .Q ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, Midori_rounds_roundReg_out[14]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_15_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10007, new_AGEMA_signal_10005, new_AGEMA_signal_10003}), .Q ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, Midori_rounds_roundReg_out[15]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_16_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3939, new_AGEMA_signal_3938, Midori_rounds_roundResult_Reg_SFF_16_DQ}), .Q ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, Midori_rounds_roundReg_out[16]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_17_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10013, new_AGEMA_signal_10011, new_AGEMA_signal_10009}), .Q ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, Midori_rounds_roundReg_out[17]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_18_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, Midori_rounds_roundResult_Reg_SFF_18_DQ}), .Q ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, Midori_rounds_roundReg_out[18]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_19_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10019, new_AGEMA_signal_10017, new_AGEMA_signal_10015}), .Q ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, Midori_rounds_roundReg_out[19]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_20_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3941, new_AGEMA_signal_3940, Midori_rounds_roundResult_Reg_SFF_20_DQ}), .Q ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, Midori_rounds_roundReg_out[20]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_21_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10025, new_AGEMA_signal_10023, new_AGEMA_signal_10021}), .Q ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, Midori_rounds_roundReg_out[21]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_22_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, Midori_rounds_roundResult_Reg_SFF_22_DQ}), .Q ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, Midori_rounds_roundReg_out[22]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_23_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10031, new_AGEMA_signal_10029, new_AGEMA_signal_10027}), .Q ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, Midori_rounds_roundReg_out[23]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_24_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3919, new_AGEMA_signal_3918, Midori_rounds_roundResult_Reg_SFF_24_DQ}), .Q ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, Midori_rounds_roundReg_out[24]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_25_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10037, new_AGEMA_signal_10035, new_AGEMA_signal_10033}), .Q ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, Midori_rounds_roundReg_out[25]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_26_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, Midori_rounds_roundResult_Reg_SFF_26_DQ}), .Q ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, Midori_rounds_roundReg_out[26]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_27_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10043, new_AGEMA_signal_10041, new_AGEMA_signal_10039}), .Q ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, Midori_rounds_roundReg_out[27]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_28_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3921, new_AGEMA_signal_3920, Midori_rounds_roundResult_Reg_SFF_28_DQ}), .Q ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, Midori_rounds_roundReg_out[28]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_29_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10049, new_AGEMA_signal_10047, new_AGEMA_signal_10045}), .Q ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, Midori_rounds_roundReg_out[29]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_30_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, Midori_rounds_roundResult_Reg_SFF_30_DQ}), .Q ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, Midori_rounds_roundReg_out[30]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_31_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10055, new_AGEMA_signal_10053, new_AGEMA_signal_10051}), .Q ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, Midori_rounds_roundReg_out[31]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_32_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3923, new_AGEMA_signal_3922, Midori_rounds_roundResult_Reg_SFF_32_DQ}), .Q ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, Midori_rounds_roundReg_out[32]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_33_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10061, new_AGEMA_signal_10059, new_AGEMA_signal_10057}), .Q ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, Midori_rounds_roundReg_out[33]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_34_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, Midori_rounds_roundResult_Reg_SFF_34_DQ}), .Q ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, Midori_rounds_roundReg_out[34]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_35_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10067, new_AGEMA_signal_10065, new_AGEMA_signal_10063}), .Q ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, Midori_rounds_roundReg_out[35]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_36_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, Midori_rounds_roundResult_Reg_SFF_36_DQ}), .Q ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, Midori_rounds_roundReg_out[36]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_37_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10073, new_AGEMA_signal_10071, new_AGEMA_signal_10069}), .Q ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, Midori_rounds_roundReg_out[37]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_38_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3731, new_AGEMA_signal_3730, Midori_rounds_roundResult_Reg_SFF_38_DQ}), .Q ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, Midori_rounds_roundReg_out[38]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_39_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10079, new_AGEMA_signal_10077, new_AGEMA_signal_10075}), .Q ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, Midori_rounds_roundReg_out[39]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_40_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3927, new_AGEMA_signal_3926, Midori_rounds_roundResult_Reg_SFF_40_DQ}), .Q ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, Midori_rounds_roundReg_out[40]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_41_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10085, new_AGEMA_signal_10083, new_AGEMA_signal_10081}), .Q ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, Midori_rounds_roundReg_out[41]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_42_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3737, new_AGEMA_signal_3736, Midori_rounds_roundResult_Reg_SFF_42_DQ}), .Q ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, Midori_rounds_roundReg_out[42]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_43_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10091, new_AGEMA_signal_10089, new_AGEMA_signal_10087}), .Q ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, Midori_rounds_roundReg_out[43]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_44_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3929, new_AGEMA_signal_3928, Midori_rounds_roundResult_Reg_SFF_44_DQ}), .Q ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, Midori_rounds_roundReg_out[44]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_45_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10097, new_AGEMA_signal_10095, new_AGEMA_signal_10093}), .Q ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, Midori_rounds_roundReg_out[45]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_46_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3743, new_AGEMA_signal_3742, Midori_rounds_roundResult_Reg_SFF_46_DQ}), .Q ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, Midori_rounds_roundReg_out[46]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_47_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10103, new_AGEMA_signal_10101, new_AGEMA_signal_10099}), .Q ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, Midori_rounds_roundReg_out[47]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_48_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3931, new_AGEMA_signal_3930, Midori_rounds_roundResult_Reg_SFF_48_DQ}), .Q ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, Midori_rounds_roundReg_out[48]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_49_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10109, new_AGEMA_signal_10107, new_AGEMA_signal_10105}), .Q ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, Midori_rounds_roundReg_out[49]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_50_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, Midori_rounds_roundResult_Reg_SFF_50_DQ}), .Q ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, Midori_rounds_roundReg_out[50]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_51_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10115, new_AGEMA_signal_10113, new_AGEMA_signal_10111}), .Q ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, Midori_rounds_roundReg_out[51]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_52_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3943, new_AGEMA_signal_3942, Midori_rounds_roundResult_Reg_SFF_52_DQ}), .Q ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, Midori_rounds_roundReg_out[52]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_53_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10121, new_AGEMA_signal_10119, new_AGEMA_signal_10117}), .Q ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, Midori_rounds_roundReg_out[53]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_54_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, Midori_rounds_roundResult_Reg_SFF_54_DQ}), .Q ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, Midori_rounds_roundReg_out[54]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_55_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10127, new_AGEMA_signal_10125, new_AGEMA_signal_10123}), .Q ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, Midori_rounds_roundReg_out[55]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_56_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3949, new_AGEMA_signal_3948, Midori_rounds_roundResult_Reg_SFF_56_DQ}), .Q ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, Midori_rounds_roundReg_out[56]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_57_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10133, new_AGEMA_signal_10131, new_AGEMA_signal_10129}), .Q ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, Midori_rounds_roundReg_out[57]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_58_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, Midori_rounds_roundResult_Reg_SFF_58_DQ}), .Q ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, Midori_rounds_roundReg_out[58]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_59_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10139, new_AGEMA_signal_10137, new_AGEMA_signal_10135}), .Q ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, Midori_rounds_roundReg_out[59]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_60_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, Midori_rounds_roundResult_Reg_SFF_60_DQ}), .Q ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, Midori_rounds_roundReg_out[60]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_61_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10145, new_AGEMA_signal_10143, new_AGEMA_signal_10141}), .Q ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, Midori_rounds_roundReg_out[61]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_62_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, Midori_rounds_roundResult_Reg_SFF_62_DQ}), .Q ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, Midori_rounds_roundReg_out[62]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_63_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10151, new_AGEMA_signal_10149, new_AGEMA_signal_10147}), .Q ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, Midori_rounds_roundReg_out[63]}) ) ;
endmodule
