////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module SkinnyTop in file /AGEMA/Designs/Skinny64_64_round-based/AGEMA/SkinnyTop.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module SkinnyTop_HPC2_Pipeline_d3 (Plaintext_s0, Key_s0, clk, rst, Key_s1, Key_s2, Key_s3, Plaintext_s1, Plaintext_s2, Plaintext_s3, Fresh, Ciphertext_s0, done, Ciphertext_s1, Ciphertext_s2, Ciphertext_s3);
    input [63:0] Plaintext_s0 ;
    input [63:0] Key_s0 ;
    input clk ;
    input rst ;
    input [63:0] Key_s1 ;
    input [63:0] Key_s2 ;
    input [63:0] Key_s3 ;
    input [63:0] Plaintext_s1 ;
    input [63:0] Plaintext_s2 ;
    input [63:0] Plaintext_s3 ;
    input [383:0] Fresh ;
    output [63:0] Ciphertext_s0 ;
    output done ;
    output [63:0] Ciphertext_s1 ;
    output [63:0] Ciphertext_s2 ;
    output [63:0] Ciphertext_s3 ;
    wire SubCellInst_SboxInst_0_n3 ;
    wire SubCellInst_SboxInst_0_YY_0_ ;
    wire SubCellInst_SboxInst_0_YY_1_ ;
    wire SubCellInst_SboxInst_0_L3 ;
    wire SubCellInst_SboxInst_0_YY_3 ;
    wire SubCellInst_SboxInst_0_L2 ;
    wire SubCellInst_SboxInst_0_T3 ;
    wire SubCellInst_SboxInst_0_Q7 ;
    wire SubCellInst_SboxInst_0_L1 ;
    wire SubCellInst_SboxInst_0_Q6 ;
    wire SubCellInst_SboxInst_0_L0 ;
    wire SubCellInst_SboxInst_0_T2 ;
    wire SubCellInst_SboxInst_0_Q4 ;
    wire SubCellInst_SboxInst_0_T1 ;
    wire SubCellInst_SboxInst_0_Q2 ;
    wire SubCellInst_SboxInst_0_T0 ;
    wire SubCellInst_SboxInst_0_Q1 ;
    wire SubCellInst_SboxInst_0_Q0 ;
    wire SubCellInst_SboxInst_0_XX_1_ ;
    wire SubCellInst_SboxInst_0_XX_2_ ;
    wire SubCellInst_SboxInst_1_n3 ;
    wire SubCellInst_SboxInst_1_YY_0_ ;
    wire SubCellInst_SboxInst_1_YY_1_ ;
    wire SubCellInst_SboxInst_1_L3 ;
    wire SubCellInst_SboxInst_1_YY_3 ;
    wire SubCellInst_SboxInst_1_L2 ;
    wire SubCellInst_SboxInst_1_T3 ;
    wire SubCellInst_SboxInst_1_Q7 ;
    wire SubCellInst_SboxInst_1_L1 ;
    wire SubCellInst_SboxInst_1_Q6 ;
    wire SubCellInst_SboxInst_1_L0 ;
    wire SubCellInst_SboxInst_1_T2 ;
    wire SubCellInst_SboxInst_1_Q4 ;
    wire SubCellInst_SboxInst_1_T1 ;
    wire SubCellInst_SboxInst_1_Q2 ;
    wire SubCellInst_SboxInst_1_T0 ;
    wire SubCellInst_SboxInst_1_Q1 ;
    wire SubCellInst_SboxInst_1_Q0 ;
    wire SubCellInst_SboxInst_1_XX_1_ ;
    wire SubCellInst_SboxInst_1_XX_2_ ;
    wire SubCellInst_SboxInst_2_n3 ;
    wire SubCellInst_SboxInst_2_YY_0_ ;
    wire SubCellInst_SboxInst_2_YY_1_ ;
    wire SubCellInst_SboxInst_2_L3 ;
    wire SubCellInst_SboxInst_2_YY_3 ;
    wire SubCellInst_SboxInst_2_L2 ;
    wire SubCellInst_SboxInst_2_T3 ;
    wire SubCellInst_SboxInst_2_Q7 ;
    wire SubCellInst_SboxInst_2_L1 ;
    wire SubCellInst_SboxInst_2_Q6 ;
    wire SubCellInst_SboxInst_2_L0 ;
    wire SubCellInst_SboxInst_2_T2 ;
    wire SubCellInst_SboxInst_2_Q4 ;
    wire SubCellInst_SboxInst_2_T1 ;
    wire SubCellInst_SboxInst_2_Q2 ;
    wire SubCellInst_SboxInst_2_T0 ;
    wire SubCellInst_SboxInst_2_Q1 ;
    wire SubCellInst_SboxInst_2_Q0 ;
    wire SubCellInst_SboxInst_2_XX_1_ ;
    wire SubCellInst_SboxInst_2_XX_2_ ;
    wire SubCellInst_SboxInst_3_n3 ;
    wire SubCellInst_SboxInst_3_YY_0_ ;
    wire SubCellInst_SboxInst_3_YY_1_ ;
    wire SubCellInst_SboxInst_3_L3 ;
    wire SubCellInst_SboxInst_3_YY_3 ;
    wire SubCellInst_SboxInst_3_L2 ;
    wire SubCellInst_SboxInst_3_T3 ;
    wire SubCellInst_SboxInst_3_Q7 ;
    wire SubCellInst_SboxInst_3_L1 ;
    wire SubCellInst_SboxInst_3_Q6 ;
    wire SubCellInst_SboxInst_3_L0 ;
    wire SubCellInst_SboxInst_3_T2 ;
    wire SubCellInst_SboxInst_3_Q4 ;
    wire SubCellInst_SboxInst_3_T1 ;
    wire SubCellInst_SboxInst_3_Q2 ;
    wire SubCellInst_SboxInst_3_T0 ;
    wire SubCellInst_SboxInst_3_Q1 ;
    wire SubCellInst_SboxInst_3_Q0 ;
    wire SubCellInst_SboxInst_3_XX_1_ ;
    wire SubCellInst_SboxInst_3_XX_2_ ;
    wire SubCellInst_SboxInst_4_n3 ;
    wire SubCellInst_SboxInst_4_YY_0_ ;
    wire SubCellInst_SboxInst_4_YY_1_ ;
    wire SubCellInst_SboxInst_4_L3 ;
    wire SubCellInst_SboxInst_4_YY_3 ;
    wire SubCellInst_SboxInst_4_L2 ;
    wire SubCellInst_SboxInst_4_T3 ;
    wire SubCellInst_SboxInst_4_Q7 ;
    wire SubCellInst_SboxInst_4_L1 ;
    wire SubCellInst_SboxInst_4_Q6 ;
    wire SubCellInst_SboxInst_4_L0 ;
    wire SubCellInst_SboxInst_4_T2 ;
    wire SubCellInst_SboxInst_4_Q4 ;
    wire SubCellInst_SboxInst_4_T1 ;
    wire SubCellInst_SboxInst_4_Q2 ;
    wire SubCellInst_SboxInst_4_T0 ;
    wire SubCellInst_SboxInst_4_Q1 ;
    wire SubCellInst_SboxInst_4_Q0 ;
    wire SubCellInst_SboxInst_4_XX_1_ ;
    wire SubCellInst_SboxInst_4_XX_2_ ;
    wire SubCellInst_SboxInst_5_n3 ;
    wire SubCellInst_SboxInst_5_YY_0_ ;
    wire SubCellInst_SboxInst_5_YY_1_ ;
    wire SubCellInst_SboxInst_5_L3 ;
    wire SubCellInst_SboxInst_5_YY_3 ;
    wire SubCellInst_SboxInst_5_L2 ;
    wire SubCellInst_SboxInst_5_T3 ;
    wire SubCellInst_SboxInst_5_Q7 ;
    wire SubCellInst_SboxInst_5_L1 ;
    wire SubCellInst_SboxInst_5_Q6 ;
    wire SubCellInst_SboxInst_5_L0 ;
    wire SubCellInst_SboxInst_5_T2 ;
    wire SubCellInst_SboxInst_5_Q4 ;
    wire SubCellInst_SboxInst_5_T1 ;
    wire SubCellInst_SboxInst_5_Q2 ;
    wire SubCellInst_SboxInst_5_T0 ;
    wire SubCellInst_SboxInst_5_Q1 ;
    wire SubCellInst_SboxInst_5_Q0 ;
    wire SubCellInst_SboxInst_5_XX_1_ ;
    wire SubCellInst_SboxInst_5_XX_2_ ;
    wire SubCellInst_SboxInst_6_n3 ;
    wire SubCellInst_SboxInst_6_YY_0_ ;
    wire SubCellInst_SboxInst_6_YY_1_ ;
    wire SubCellInst_SboxInst_6_L3 ;
    wire SubCellInst_SboxInst_6_YY_3 ;
    wire SubCellInst_SboxInst_6_L2 ;
    wire SubCellInst_SboxInst_6_T3 ;
    wire SubCellInst_SboxInst_6_Q7 ;
    wire SubCellInst_SboxInst_6_L1 ;
    wire SubCellInst_SboxInst_6_Q6 ;
    wire SubCellInst_SboxInst_6_L0 ;
    wire SubCellInst_SboxInst_6_T2 ;
    wire SubCellInst_SboxInst_6_Q4 ;
    wire SubCellInst_SboxInst_6_T1 ;
    wire SubCellInst_SboxInst_6_Q2 ;
    wire SubCellInst_SboxInst_6_T0 ;
    wire SubCellInst_SboxInst_6_Q1 ;
    wire SubCellInst_SboxInst_6_Q0 ;
    wire SubCellInst_SboxInst_6_XX_1_ ;
    wire SubCellInst_SboxInst_6_XX_2_ ;
    wire SubCellInst_SboxInst_7_n3 ;
    wire SubCellInst_SboxInst_7_YY_0_ ;
    wire SubCellInst_SboxInst_7_YY_1_ ;
    wire SubCellInst_SboxInst_7_L3 ;
    wire SubCellInst_SboxInst_7_YY_3 ;
    wire SubCellInst_SboxInst_7_L2 ;
    wire SubCellInst_SboxInst_7_T3 ;
    wire SubCellInst_SboxInst_7_Q7 ;
    wire SubCellInst_SboxInst_7_L1 ;
    wire SubCellInst_SboxInst_7_Q6 ;
    wire SubCellInst_SboxInst_7_L0 ;
    wire SubCellInst_SboxInst_7_T2 ;
    wire SubCellInst_SboxInst_7_Q4 ;
    wire SubCellInst_SboxInst_7_T1 ;
    wire SubCellInst_SboxInst_7_Q2 ;
    wire SubCellInst_SboxInst_7_T0 ;
    wire SubCellInst_SboxInst_7_Q1 ;
    wire SubCellInst_SboxInst_7_Q0 ;
    wire SubCellInst_SboxInst_7_XX_1_ ;
    wire SubCellInst_SboxInst_7_XX_2_ ;
    wire SubCellInst_SboxInst_8_n3 ;
    wire SubCellInst_SboxInst_8_YY_0_ ;
    wire SubCellInst_SboxInst_8_YY_1_ ;
    wire SubCellInst_SboxInst_8_L3 ;
    wire SubCellInst_SboxInst_8_YY_3 ;
    wire SubCellInst_SboxInst_8_L2 ;
    wire SubCellInst_SboxInst_8_T3 ;
    wire SubCellInst_SboxInst_8_Q7 ;
    wire SubCellInst_SboxInst_8_L1 ;
    wire SubCellInst_SboxInst_8_Q6 ;
    wire SubCellInst_SboxInst_8_L0 ;
    wire SubCellInst_SboxInst_8_T2 ;
    wire SubCellInst_SboxInst_8_Q4 ;
    wire SubCellInst_SboxInst_8_T1 ;
    wire SubCellInst_SboxInst_8_Q2 ;
    wire SubCellInst_SboxInst_8_T0 ;
    wire SubCellInst_SboxInst_8_Q1 ;
    wire SubCellInst_SboxInst_8_Q0 ;
    wire SubCellInst_SboxInst_8_XX_1_ ;
    wire SubCellInst_SboxInst_8_XX_2_ ;
    wire SubCellInst_SboxInst_9_n3 ;
    wire SubCellInst_SboxInst_9_YY_0_ ;
    wire SubCellInst_SboxInst_9_YY_1_ ;
    wire SubCellInst_SboxInst_9_L3 ;
    wire SubCellInst_SboxInst_9_YY_3 ;
    wire SubCellInst_SboxInst_9_L2 ;
    wire SubCellInst_SboxInst_9_T3 ;
    wire SubCellInst_SboxInst_9_Q7 ;
    wire SubCellInst_SboxInst_9_L1 ;
    wire SubCellInst_SboxInst_9_Q6 ;
    wire SubCellInst_SboxInst_9_L0 ;
    wire SubCellInst_SboxInst_9_T2 ;
    wire SubCellInst_SboxInst_9_Q4 ;
    wire SubCellInst_SboxInst_9_T1 ;
    wire SubCellInst_SboxInst_9_Q2 ;
    wire SubCellInst_SboxInst_9_T0 ;
    wire SubCellInst_SboxInst_9_Q1 ;
    wire SubCellInst_SboxInst_9_Q0 ;
    wire SubCellInst_SboxInst_9_XX_1_ ;
    wire SubCellInst_SboxInst_9_XX_2_ ;
    wire SubCellInst_SboxInst_10_n3 ;
    wire SubCellInst_SboxInst_10_YY_0_ ;
    wire SubCellInst_SboxInst_10_YY_1_ ;
    wire SubCellInst_SboxInst_10_L3 ;
    wire SubCellInst_SboxInst_10_YY_3 ;
    wire SubCellInst_SboxInst_10_L2 ;
    wire SubCellInst_SboxInst_10_T3 ;
    wire SubCellInst_SboxInst_10_Q7 ;
    wire SubCellInst_SboxInst_10_L1 ;
    wire SubCellInst_SboxInst_10_Q6 ;
    wire SubCellInst_SboxInst_10_L0 ;
    wire SubCellInst_SboxInst_10_T2 ;
    wire SubCellInst_SboxInst_10_Q4 ;
    wire SubCellInst_SboxInst_10_T1 ;
    wire SubCellInst_SboxInst_10_Q2 ;
    wire SubCellInst_SboxInst_10_T0 ;
    wire SubCellInst_SboxInst_10_Q1 ;
    wire SubCellInst_SboxInst_10_Q0 ;
    wire SubCellInst_SboxInst_10_XX_1_ ;
    wire SubCellInst_SboxInst_10_XX_2_ ;
    wire SubCellInst_SboxInst_11_n3 ;
    wire SubCellInst_SboxInst_11_YY_0_ ;
    wire SubCellInst_SboxInst_11_YY_1_ ;
    wire SubCellInst_SboxInst_11_L3 ;
    wire SubCellInst_SboxInst_11_YY_3 ;
    wire SubCellInst_SboxInst_11_L2 ;
    wire SubCellInst_SboxInst_11_T3 ;
    wire SubCellInst_SboxInst_11_Q7 ;
    wire SubCellInst_SboxInst_11_L1 ;
    wire SubCellInst_SboxInst_11_Q6 ;
    wire SubCellInst_SboxInst_11_L0 ;
    wire SubCellInst_SboxInst_11_T2 ;
    wire SubCellInst_SboxInst_11_Q4 ;
    wire SubCellInst_SboxInst_11_T1 ;
    wire SubCellInst_SboxInst_11_Q2 ;
    wire SubCellInst_SboxInst_11_T0 ;
    wire SubCellInst_SboxInst_11_Q1 ;
    wire SubCellInst_SboxInst_11_Q0 ;
    wire SubCellInst_SboxInst_11_XX_1_ ;
    wire SubCellInst_SboxInst_11_XX_2_ ;
    wire SubCellInst_SboxInst_12_n3 ;
    wire SubCellInst_SboxInst_12_YY_0_ ;
    wire SubCellInst_SboxInst_12_YY_1_ ;
    wire SubCellInst_SboxInst_12_L3 ;
    wire SubCellInst_SboxInst_12_YY_3 ;
    wire SubCellInst_SboxInst_12_L2 ;
    wire SubCellInst_SboxInst_12_T3 ;
    wire SubCellInst_SboxInst_12_Q7 ;
    wire SubCellInst_SboxInst_12_L1 ;
    wire SubCellInst_SboxInst_12_Q6 ;
    wire SubCellInst_SboxInst_12_L0 ;
    wire SubCellInst_SboxInst_12_T2 ;
    wire SubCellInst_SboxInst_12_Q4 ;
    wire SubCellInst_SboxInst_12_T1 ;
    wire SubCellInst_SboxInst_12_Q2 ;
    wire SubCellInst_SboxInst_12_T0 ;
    wire SubCellInst_SboxInst_12_Q1 ;
    wire SubCellInst_SboxInst_12_Q0 ;
    wire SubCellInst_SboxInst_12_XX_1_ ;
    wire SubCellInst_SboxInst_12_XX_2_ ;
    wire SubCellInst_SboxInst_13_n3 ;
    wire SubCellInst_SboxInst_13_YY_0_ ;
    wire SubCellInst_SboxInst_13_YY_1_ ;
    wire SubCellInst_SboxInst_13_L3 ;
    wire SubCellInst_SboxInst_13_YY_3 ;
    wire SubCellInst_SboxInst_13_L2 ;
    wire SubCellInst_SboxInst_13_T3 ;
    wire SubCellInst_SboxInst_13_Q7 ;
    wire SubCellInst_SboxInst_13_L1 ;
    wire SubCellInst_SboxInst_13_Q6 ;
    wire SubCellInst_SboxInst_13_L0 ;
    wire SubCellInst_SboxInst_13_T2 ;
    wire SubCellInst_SboxInst_13_Q4 ;
    wire SubCellInst_SboxInst_13_T1 ;
    wire SubCellInst_SboxInst_13_Q2 ;
    wire SubCellInst_SboxInst_13_T0 ;
    wire SubCellInst_SboxInst_13_Q1 ;
    wire SubCellInst_SboxInst_13_Q0 ;
    wire SubCellInst_SboxInst_13_XX_1_ ;
    wire SubCellInst_SboxInst_13_XX_2_ ;
    wire SubCellInst_SboxInst_14_n3 ;
    wire SubCellInst_SboxInst_14_YY_0_ ;
    wire SubCellInst_SboxInst_14_YY_1_ ;
    wire SubCellInst_SboxInst_14_L3 ;
    wire SubCellInst_SboxInst_14_YY_3 ;
    wire SubCellInst_SboxInst_14_L2 ;
    wire SubCellInst_SboxInst_14_T3 ;
    wire SubCellInst_SboxInst_14_Q7 ;
    wire SubCellInst_SboxInst_14_L1 ;
    wire SubCellInst_SboxInst_14_Q6 ;
    wire SubCellInst_SboxInst_14_L0 ;
    wire SubCellInst_SboxInst_14_T2 ;
    wire SubCellInst_SboxInst_14_Q4 ;
    wire SubCellInst_SboxInst_14_T1 ;
    wire SubCellInst_SboxInst_14_Q2 ;
    wire SubCellInst_SboxInst_14_T0 ;
    wire SubCellInst_SboxInst_14_Q1 ;
    wire SubCellInst_SboxInst_14_Q0 ;
    wire SubCellInst_SboxInst_14_XX_1_ ;
    wire SubCellInst_SboxInst_14_XX_2_ ;
    wire SubCellInst_SboxInst_15_n3 ;
    wire SubCellInst_SboxInst_15_YY_0_ ;
    wire SubCellInst_SboxInst_15_YY_1_ ;
    wire SubCellInst_SboxInst_15_L3 ;
    wire SubCellInst_SboxInst_15_YY_3 ;
    wire SubCellInst_SboxInst_15_L2 ;
    wire SubCellInst_SboxInst_15_T3 ;
    wire SubCellInst_SboxInst_15_Q7 ;
    wire SubCellInst_SboxInst_15_L1 ;
    wire SubCellInst_SboxInst_15_Q6 ;
    wire SubCellInst_SboxInst_15_L0 ;
    wire SubCellInst_SboxInst_15_T2 ;
    wire SubCellInst_SboxInst_15_Q4 ;
    wire SubCellInst_SboxInst_15_T1 ;
    wire SubCellInst_SboxInst_15_Q2 ;
    wire SubCellInst_SboxInst_15_T0 ;
    wire SubCellInst_SboxInst_15_Q1 ;
    wire SubCellInst_SboxInst_15_Q0 ;
    wire SubCellInst_SboxInst_15_XX_1_ ;
    wire SubCellInst_SboxInst_15_XX_2_ ;
    wire AddConstXOR_AddConstXOR_XORInst_0_0_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_0_1_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_0_2_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_0_3_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_0_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_1_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_2_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_3_n1 ;
    wire MCInst_MCR0_XORInst_0_0_n2 ;
    wire MCInst_MCR0_XORInst_0_0_n1 ;
    wire MCInst_MCR0_XORInst_0_1_n2 ;
    wire MCInst_MCR0_XORInst_0_1_n1 ;
    wire MCInst_MCR0_XORInst_0_2_n2 ;
    wire MCInst_MCR0_XORInst_0_2_n1 ;
    wire MCInst_MCR0_XORInst_0_3_n2 ;
    wire MCInst_MCR0_XORInst_0_3_n1 ;
    wire MCInst_MCR0_XORInst_1_0_n2 ;
    wire MCInst_MCR0_XORInst_1_0_n1 ;
    wire MCInst_MCR0_XORInst_1_1_n2 ;
    wire MCInst_MCR0_XORInst_1_1_n1 ;
    wire MCInst_MCR0_XORInst_1_2_n2 ;
    wire MCInst_MCR0_XORInst_1_2_n1 ;
    wire MCInst_MCR0_XORInst_1_3_n2 ;
    wire MCInst_MCR0_XORInst_1_3_n1 ;
    wire MCInst_MCR0_XORInst_2_0_n2 ;
    wire MCInst_MCR0_XORInst_2_0_n1 ;
    wire MCInst_MCR0_XORInst_2_1_n2 ;
    wire MCInst_MCR0_XORInst_2_1_n1 ;
    wire MCInst_MCR0_XORInst_2_2_n2 ;
    wire MCInst_MCR0_XORInst_2_2_n1 ;
    wire MCInst_MCR0_XORInst_2_3_n2 ;
    wire MCInst_MCR0_XORInst_2_3_n1 ;
    wire MCInst_MCR0_XORInst_3_0_n2 ;
    wire MCInst_MCR0_XORInst_3_0_n1 ;
    wire MCInst_MCR0_XORInst_3_1_n2 ;
    wire MCInst_MCR0_XORInst_3_1_n1 ;
    wire MCInst_MCR0_XORInst_3_2_n2 ;
    wire MCInst_MCR0_XORInst_3_2_n1 ;
    wire MCInst_MCR0_XORInst_3_3_n2 ;
    wire MCInst_MCR0_XORInst_3_3_n1 ;
    wire MCInst_MCR2_XORInst_0_0_n1 ;
    wire MCInst_MCR2_XORInst_0_1_n1 ;
    wire MCInst_MCR2_XORInst_0_2_n1 ;
    wire MCInst_MCR2_XORInst_0_3_n1 ;
    wire MCInst_MCR2_XORInst_1_0_n1 ;
    wire MCInst_MCR2_XORInst_1_1_n1 ;
    wire MCInst_MCR2_XORInst_1_2_n1 ;
    wire MCInst_MCR2_XORInst_1_3_n1 ;
    wire MCInst_MCR2_XORInst_2_0_n1 ;
    wire MCInst_MCR2_XORInst_2_1_n1 ;
    wire MCInst_MCR2_XORInst_2_2_n1 ;
    wire MCInst_MCR2_XORInst_2_3_n1 ;
    wire MCInst_MCR2_XORInst_3_0_n1 ;
    wire MCInst_MCR2_XORInst_3_1_n1 ;
    wire MCInst_MCR2_XORInst_3_2_n1 ;
    wire MCInst_MCR2_XORInst_3_3_n1 ;
    wire MCInst_MCR3_XORInst_0_0_n1 ;
    wire MCInst_MCR3_XORInst_0_1_n1 ;
    wire MCInst_MCR3_XORInst_0_2_n1 ;
    wire MCInst_MCR3_XORInst_0_3_n1 ;
    wire MCInst_MCR3_XORInst_1_0_n1 ;
    wire MCInst_MCR3_XORInst_1_1_n1 ;
    wire MCInst_MCR3_XORInst_1_2_n1 ;
    wire MCInst_MCR3_XORInst_1_3_n1 ;
    wire MCInst_MCR3_XORInst_2_0_n1 ;
    wire MCInst_MCR3_XORInst_2_1_n1 ;
    wire MCInst_MCR3_XORInst_2_2_n1 ;
    wire MCInst_MCR3_XORInst_2_3_n1 ;
    wire MCInst_MCR3_XORInst_3_0_n1 ;
    wire MCInst_MCR3_XORInst_3_1_n1 ;
    wire MCInst_MCR3_XORInst_3_2_n1 ;
    wire MCInst_MCR3_XORInst_3_3_n1 ;
    wire FSMUpdateInst_StateUpdateInst_0_n4 ;
    wire FSMUpdateInst_StateUpdateInst_0_n3 ;
    wire FSMUpdateInst_StateUpdateInst_0_n2 ;
    wire FSMUpdateInst_StateUpdateInst_0_n1 ;
    wire FSMUpdateInst_StateUpdateInst_2_n4 ;
    wire FSMUpdateInst_StateUpdateInst_2_n3 ;
    wire FSMUpdateInst_StateUpdateInst_2_n2 ;
    wire FSMUpdateInst_StateUpdateInst_2_n1 ;
    wire FSMUpdateInst_StateUpdateInst_5_n4 ;
    wire FSMUpdateInst_StateUpdateInst_5_n3 ;
    wire FSMUpdateInst_StateUpdateInst_5_n2 ;
    wire FSMUpdateInst_StateUpdateInst_5_n1 ;
    wire FSMSignalsInst_doneInst_n5 ;
    wire FSMSignalsInst_doneInst_n4 ;
    wire FSMSignalsInst_doneInst_n3 ;
    wire FSMSignalsInst_doneInst_n2 ;
    wire FSMSignalsInst_doneInst_n1 ;
    wire [63:0] MCOutput ;
    wire [63:0] StateRegInput ;
    wire [63:29] SubCellOutput ;
    wire [5:1] FSM ;
    wire [63:32] AddRoundConstantOutput ;
    wire [47:0] ShiftRowsOutput ;
    wire [5:0] FSMUpdate ;
    wire [5:0] FSMSelected ;
    wire [63:0] TweakeyGeneration_StateRegInput ;
    wire [63:0] TweakeyGeneration_key_Feedback ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4497 ;
    wire new_AGEMA_signal_4498 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5195 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5202 ;
    wire new_AGEMA_signal_5203 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5207 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5213 ;
    wire new_AGEMA_signal_5214 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5219 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5226 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5231 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5238 ;
    wire new_AGEMA_signal_5239 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5249 ;
    wire new_AGEMA_signal_5250 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5255 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5262 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5273 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5291 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5303 ;
    wire new_AGEMA_signal_5304 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5309 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6654 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;
    wire new_AGEMA_signal_6672 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6677 ;
    wire new_AGEMA_signal_6678 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6682 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6688 ;
    wire new_AGEMA_signal_6689 ;
    wire new_AGEMA_signal_6690 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6695 ;
    wire new_AGEMA_signal_6696 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6700 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6706 ;
    wire new_AGEMA_signal_6707 ;
    wire new_AGEMA_signal_6708 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6713 ;
    wire new_AGEMA_signal_6714 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6718 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6724 ;
    wire new_AGEMA_signal_6725 ;
    wire new_AGEMA_signal_6726 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7036 ;
    wire new_AGEMA_signal_7037 ;
    wire new_AGEMA_signal_7038 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7042 ;
    wire new_AGEMA_signal_7043 ;
    wire new_AGEMA_signal_7044 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7048 ;
    wire new_AGEMA_signal_7049 ;
    wire new_AGEMA_signal_7050 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7054 ;
    wire new_AGEMA_signal_7055 ;
    wire new_AGEMA_signal_7056 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7060 ;
    wire new_AGEMA_signal_7061 ;
    wire new_AGEMA_signal_7062 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7066 ;
    wire new_AGEMA_signal_7067 ;
    wire new_AGEMA_signal_7068 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7072 ;
    wire new_AGEMA_signal_7073 ;
    wire new_AGEMA_signal_7074 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7078 ;
    wire new_AGEMA_signal_7079 ;
    wire new_AGEMA_signal_7080 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7084 ;
    wire new_AGEMA_signal_7085 ;
    wire new_AGEMA_signal_7086 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7090 ;
    wire new_AGEMA_signal_7091 ;
    wire new_AGEMA_signal_7092 ;
    wire new_AGEMA_signal_7093 ;
    wire new_AGEMA_signal_7094 ;
    wire new_AGEMA_signal_7095 ;
    wire new_AGEMA_signal_7096 ;
    wire new_AGEMA_signal_7097 ;
    wire new_AGEMA_signal_7098 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7102 ;
    wire new_AGEMA_signal_7103 ;
    wire new_AGEMA_signal_7104 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7108 ;
    wire new_AGEMA_signal_7109 ;
    wire new_AGEMA_signal_7110 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7114 ;
    wire new_AGEMA_signal_7115 ;
    wire new_AGEMA_signal_7116 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7120 ;
    wire new_AGEMA_signal_7121 ;
    wire new_AGEMA_signal_7122 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7126 ;
    wire new_AGEMA_signal_7127 ;
    wire new_AGEMA_signal_7128 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7132 ;
    wire new_AGEMA_signal_7133 ;
    wire new_AGEMA_signal_7134 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7138 ;
    wire new_AGEMA_signal_7139 ;
    wire new_AGEMA_signal_7140 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7144 ;
    wire new_AGEMA_signal_7145 ;
    wire new_AGEMA_signal_7146 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7150 ;
    wire new_AGEMA_signal_7151 ;
    wire new_AGEMA_signal_7152 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7156 ;
    wire new_AGEMA_signal_7157 ;
    wire new_AGEMA_signal_7158 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7162 ;
    wire new_AGEMA_signal_7163 ;
    wire new_AGEMA_signal_7164 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7168 ;
    wire new_AGEMA_signal_7169 ;
    wire new_AGEMA_signal_7170 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7174 ;
    wire new_AGEMA_signal_7175 ;
    wire new_AGEMA_signal_7176 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7180 ;
    wire new_AGEMA_signal_7181 ;
    wire new_AGEMA_signal_7182 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7186 ;
    wire new_AGEMA_signal_7187 ;
    wire new_AGEMA_signal_7188 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7192 ;
    wire new_AGEMA_signal_7193 ;
    wire new_AGEMA_signal_7194 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7198 ;
    wire new_AGEMA_signal_7199 ;
    wire new_AGEMA_signal_7200 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7204 ;
    wire new_AGEMA_signal_7205 ;
    wire new_AGEMA_signal_7206 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7489 ;
    wire new_AGEMA_signal_7490 ;
    wire new_AGEMA_signal_7491 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7495 ;
    wire new_AGEMA_signal_7496 ;
    wire new_AGEMA_signal_7497 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7499 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7501 ;
    wire new_AGEMA_signal_7502 ;
    wire new_AGEMA_signal_7503 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7507 ;
    wire new_AGEMA_signal_7508 ;
    wire new_AGEMA_signal_7509 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7513 ;
    wire new_AGEMA_signal_7514 ;
    wire new_AGEMA_signal_7515 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7519 ;
    wire new_AGEMA_signal_7520 ;
    wire new_AGEMA_signal_7521 ;
    wire new_AGEMA_signal_7522 ;
    wire new_AGEMA_signal_7523 ;
    wire new_AGEMA_signal_7524 ;
    wire new_AGEMA_signal_7525 ;
    wire new_AGEMA_signal_7526 ;
    wire new_AGEMA_signal_7527 ;
    wire new_AGEMA_signal_7528 ;
    wire new_AGEMA_signal_7529 ;
    wire new_AGEMA_signal_7530 ;
    wire new_AGEMA_signal_7531 ;
    wire new_AGEMA_signal_7532 ;
    wire new_AGEMA_signal_7533 ;
    wire new_AGEMA_signal_7534 ;
    wire new_AGEMA_signal_7535 ;
    wire new_AGEMA_signal_7536 ;
    wire new_AGEMA_signal_7537 ;
    wire new_AGEMA_signal_7538 ;
    wire new_AGEMA_signal_7539 ;
    wire new_AGEMA_signal_7540 ;
    wire new_AGEMA_signal_7541 ;
    wire new_AGEMA_signal_7542 ;
    wire new_AGEMA_signal_7543 ;
    wire new_AGEMA_signal_7544 ;
    wire new_AGEMA_signal_7545 ;
    wire new_AGEMA_signal_7546 ;
    wire new_AGEMA_signal_7547 ;
    wire new_AGEMA_signal_7548 ;
    wire new_AGEMA_signal_7549 ;
    wire new_AGEMA_signal_7550 ;
    wire new_AGEMA_signal_7551 ;
    wire new_AGEMA_signal_7552 ;
    wire new_AGEMA_signal_7553 ;
    wire new_AGEMA_signal_7554 ;
    wire new_AGEMA_signal_7555 ;
    wire new_AGEMA_signal_7556 ;
    wire new_AGEMA_signal_7557 ;
    wire new_AGEMA_signal_7558 ;
    wire new_AGEMA_signal_7559 ;
    wire new_AGEMA_signal_7560 ;
    wire new_AGEMA_signal_7561 ;
    wire new_AGEMA_signal_7562 ;
    wire new_AGEMA_signal_7563 ;
    wire new_AGEMA_signal_7564 ;
    wire new_AGEMA_signal_7565 ;
    wire new_AGEMA_signal_7566 ;
    wire new_AGEMA_signal_7567 ;
    wire new_AGEMA_signal_7568 ;
    wire new_AGEMA_signal_7569 ;
    wire new_AGEMA_signal_7570 ;
    wire new_AGEMA_signal_7571 ;
    wire new_AGEMA_signal_7572 ;
    wire new_AGEMA_signal_7573 ;
    wire new_AGEMA_signal_7574 ;
    wire new_AGEMA_signal_7575 ;
    wire new_AGEMA_signal_7576 ;
    wire new_AGEMA_signal_7577 ;
    wire new_AGEMA_signal_7578 ;
    wire new_AGEMA_signal_7579 ;
    wire new_AGEMA_signal_7580 ;
    wire new_AGEMA_signal_7581 ;
    wire new_AGEMA_signal_7582 ;
    wire new_AGEMA_signal_7583 ;
    wire new_AGEMA_signal_7584 ;
    wire new_AGEMA_signal_7585 ;
    wire new_AGEMA_signal_7586 ;
    wire new_AGEMA_signal_7587 ;
    wire new_AGEMA_signal_7588 ;
    wire new_AGEMA_signal_7589 ;
    wire new_AGEMA_signal_7590 ;
    wire new_AGEMA_signal_7591 ;
    wire new_AGEMA_signal_7592 ;
    wire new_AGEMA_signal_7593 ;
    wire new_AGEMA_signal_7594 ;
    wire new_AGEMA_signal_7595 ;
    wire new_AGEMA_signal_7596 ;
    wire new_AGEMA_signal_7597 ;
    wire new_AGEMA_signal_7598 ;
    wire new_AGEMA_signal_7599 ;
    wire new_AGEMA_signal_7600 ;
    wire new_AGEMA_signal_7601 ;
    wire new_AGEMA_signal_7602 ;
    wire new_AGEMA_signal_7603 ;
    wire new_AGEMA_signal_7604 ;
    wire new_AGEMA_signal_7605 ;
    wire new_AGEMA_signal_7606 ;
    wire new_AGEMA_signal_7607 ;
    wire new_AGEMA_signal_7608 ;
    wire new_AGEMA_signal_7609 ;
    wire new_AGEMA_signal_7610 ;
    wire new_AGEMA_signal_7611 ;
    wire new_AGEMA_signal_7612 ;
    wire new_AGEMA_signal_7613 ;
    wire new_AGEMA_signal_7614 ;
    wire new_AGEMA_signal_7615 ;
    wire new_AGEMA_signal_7616 ;
    wire new_AGEMA_signal_7617 ;
    wire new_AGEMA_signal_7618 ;
    wire new_AGEMA_signal_7619 ;
    wire new_AGEMA_signal_7620 ;
    wire new_AGEMA_signal_7621 ;
    wire new_AGEMA_signal_7622 ;
    wire new_AGEMA_signal_7623 ;
    wire new_AGEMA_signal_7624 ;
    wire new_AGEMA_signal_7625 ;
    wire new_AGEMA_signal_7626 ;
    wire new_AGEMA_signal_7627 ;
    wire new_AGEMA_signal_7628 ;
    wire new_AGEMA_signal_7629 ;
    wire new_AGEMA_signal_7630 ;
    wire new_AGEMA_signal_7631 ;
    wire new_AGEMA_signal_7632 ;
    wire new_AGEMA_signal_7633 ;
    wire new_AGEMA_signal_7634 ;
    wire new_AGEMA_signal_7635 ;
    wire new_AGEMA_signal_7636 ;
    wire new_AGEMA_signal_7637 ;
    wire new_AGEMA_signal_7638 ;
    wire new_AGEMA_signal_7639 ;
    wire new_AGEMA_signal_7640 ;
    wire new_AGEMA_signal_7641 ;
    wire new_AGEMA_signal_7642 ;
    wire new_AGEMA_signal_7643 ;
    wire new_AGEMA_signal_7644 ;
    wire new_AGEMA_signal_7645 ;
    wire new_AGEMA_signal_7646 ;
    wire new_AGEMA_signal_7647 ;
    wire new_AGEMA_signal_7648 ;
    wire new_AGEMA_signal_7649 ;
    wire new_AGEMA_signal_7650 ;
    wire new_AGEMA_signal_7651 ;
    wire new_AGEMA_signal_7652 ;
    wire new_AGEMA_signal_7653 ;
    wire new_AGEMA_signal_7654 ;
    wire new_AGEMA_signal_7655 ;
    wire new_AGEMA_signal_7656 ;
    wire new_AGEMA_signal_7657 ;
    wire new_AGEMA_signal_7658 ;
    wire new_AGEMA_signal_7659 ;
    wire new_AGEMA_signal_7660 ;
    wire new_AGEMA_signal_7661 ;
    wire new_AGEMA_signal_7662 ;
    wire new_AGEMA_signal_7663 ;
    wire new_AGEMA_signal_7664 ;
    wire new_AGEMA_signal_7665 ;
    wire new_AGEMA_signal_7666 ;
    wire new_AGEMA_signal_7667 ;
    wire new_AGEMA_signal_7668 ;
    wire new_AGEMA_signal_7669 ;
    wire new_AGEMA_signal_7670 ;
    wire new_AGEMA_signal_7671 ;
    wire new_AGEMA_signal_7672 ;
    wire new_AGEMA_signal_7673 ;
    wire new_AGEMA_signal_7674 ;
    wire new_AGEMA_signal_7675 ;
    wire new_AGEMA_signal_7676 ;
    wire new_AGEMA_signal_7677 ;
    wire new_AGEMA_signal_7678 ;
    wire new_AGEMA_signal_7679 ;
    wire new_AGEMA_signal_7680 ;
    wire new_AGEMA_signal_7681 ;
    wire new_AGEMA_signal_7682 ;
    wire new_AGEMA_signal_7683 ;
    wire new_AGEMA_signal_7684 ;
    wire new_AGEMA_signal_7685 ;
    wire new_AGEMA_signal_7686 ;
    wire new_AGEMA_signal_7687 ;
    wire new_AGEMA_signal_7688 ;
    wire new_AGEMA_signal_7689 ;
    wire new_AGEMA_signal_7690 ;
    wire new_AGEMA_signal_7691 ;
    wire new_AGEMA_signal_7692 ;
    wire new_AGEMA_signal_7693 ;
    wire new_AGEMA_signal_7694 ;
    wire new_AGEMA_signal_7695 ;
    wire new_AGEMA_signal_7696 ;
    wire new_AGEMA_signal_7697 ;
    wire new_AGEMA_signal_7698 ;
    wire new_AGEMA_signal_7699 ;
    wire new_AGEMA_signal_7700 ;
    wire new_AGEMA_signal_7701 ;
    wire new_AGEMA_signal_7702 ;
    wire new_AGEMA_signal_7703 ;
    wire new_AGEMA_signal_7704 ;
    wire new_AGEMA_signal_7705 ;
    wire new_AGEMA_signal_7706 ;
    wire new_AGEMA_signal_7707 ;
    wire new_AGEMA_signal_7708 ;
    wire new_AGEMA_signal_7709 ;
    wire new_AGEMA_signal_7710 ;
    wire new_AGEMA_signal_7711 ;
    wire new_AGEMA_signal_7712 ;
    wire new_AGEMA_signal_7713 ;
    wire new_AGEMA_signal_7714 ;
    wire new_AGEMA_signal_7715 ;
    wire new_AGEMA_signal_7716 ;
    wire new_AGEMA_signal_7717 ;
    wire new_AGEMA_signal_7718 ;
    wire new_AGEMA_signal_7719 ;
    wire new_AGEMA_signal_7720 ;
    wire new_AGEMA_signal_7721 ;
    wire new_AGEMA_signal_7722 ;
    wire new_AGEMA_signal_7723 ;
    wire new_AGEMA_signal_7724 ;
    wire new_AGEMA_signal_7725 ;
    wire new_AGEMA_signal_7726 ;
    wire new_AGEMA_signal_7727 ;
    wire new_AGEMA_signal_7728 ;
    wire new_AGEMA_signal_7729 ;
    wire new_AGEMA_signal_7730 ;
    wire new_AGEMA_signal_7731 ;
    wire new_AGEMA_signal_7732 ;
    wire new_AGEMA_signal_7733 ;
    wire new_AGEMA_signal_7734 ;
    wire new_AGEMA_signal_7735 ;
    wire new_AGEMA_signal_7736 ;
    wire new_AGEMA_signal_7737 ;
    wire new_AGEMA_signal_7738 ;
    wire new_AGEMA_signal_7739 ;
    wire new_AGEMA_signal_7740 ;
    wire new_AGEMA_signal_7741 ;
    wire new_AGEMA_signal_7742 ;
    wire new_AGEMA_signal_7743 ;
    wire new_AGEMA_signal_7744 ;
    wire new_AGEMA_signal_7745 ;
    wire new_AGEMA_signal_7746 ;
    wire new_AGEMA_signal_7747 ;
    wire new_AGEMA_signal_7748 ;
    wire new_AGEMA_signal_7749 ;
    wire new_AGEMA_signal_7750 ;
    wire new_AGEMA_signal_7751 ;
    wire new_AGEMA_signal_7752 ;
    wire new_AGEMA_signal_7753 ;
    wire new_AGEMA_signal_7754 ;
    wire new_AGEMA_signal_7755 ;
    wire new_AGEMA_signal_7756 ;
    wire new_AGEMA_signal_7757 ;
    wire new_AGEMA_signal_7758 ;
    wire new_AGEMA_signal_7759 ;
    wire new_AGEMA_signal_7760 ;
    wire new_AGEMA_signal_7761 ;
    wire new_AGEMA_signal_7762 ;
    wire new_AGEMA_signal_7763 ;
    wire new_AGEMA_signal_7764 ;
    wire new_AGEMA_signal_7765 ;
    wire new_AGEMA_signal_7766 ;
    wire new_AGEMA_signal_7767 ;
    wire new_AGEMA_signal_7768 ;
    wire new_AGEMA_signal_7769 ;
    wire new_AGEMA_signal_7770 ;
    wire new_AGEMA_signal_7771 ;
    wire new_AGEMA_signal_7772 ;
    wire new_AGEMA_signal_7773 ;
    wire new_AGEMA_signal_7774 ;
    wire new_AGEMA_signal_7775 ;
    wire new_AGEMA_signal_7776 ;
    wire new_AGEMA_signal_7777 ;
    wire new_AGEMA_signal_7778 ;
    wire new_AGEMA_signal_7779 ;
    wire new_AGEMA_signal_7780 ;
    wire new_AGEMA_signal_7781 ;
    wire new_AGEMA_signal_7782 ;
    wire new_AGEMA_signal_7783 ;
    wire new_AGEMA_signal_7784 ;
    wire new_AGEMA_signal_7785 ;
    wire new_AGEMA_signal_7786 ;
    wire new_AGEMA_signal_7787 ;
    wire new_AGEMA_signal_7788 ;
    wire new_AGEMA_signal_7789 ;
    wire new_AGEMA_signal_7790 ;
    wire new_AGEMA_signal_7791 ;
    wire new_AGEMA_signal_7792 ;
    wire new_AGEMA_signal_7793 ;
    wire new_AGEMA_signal_7794 ;
    wire new_AGEMA_signal_7795 ;
    wire new_AGEMA_signal_7796 ;
    wire new_AGEMA_signal_7797 ;
    wire new_AGEMA_signal_7798 ;
    wire new_AGEMA_signal_7799 ;
    wire new_AGEMA_signal_7800 ;
    wire new_AGEMA_signal_7801 ;
    wire new_AGEMA_signal_7802 ;
    wire new_AGEMA_signal_7803 ;
    wire new_AGEMA_signal_7804 ;
    wire new_AGEMA_signal_7805 ;
    wire new_AGEMA_signal_7806 ;
    wire new_AGEMA_signal_7807 ;
    wire new_AGEMA_signal_7808 ;
    wire new_AGEMA_signal_7809 ;
    wire new_AGEMA_signal_7810 ;
    wire new_AGEMA_signal_7811 ;
    wire new_AGEMA_signal_7812 ;
    wire new_AGEMA_signal_7813 ;
    wire new_AGEMA_signal_7814 ;
    wire new_AGEMA_signal_7815 ;
    wire new_AGEMA_signal_7816 ;
    wire new_AGEMA_signal_7817 ;
    wire new_AGEMA_signal_7818 ;
    wire new_AGEMA_signal_7819 ;
    wire new_AGEMA_signal_7820 ;
    wire new_AGEMA_signal_7821 ;
    wire new_AGEMA_signal_7822 ;
    wire new_AGEMA_signal_7823 ;
    wire new_AGEMA_signal_7824 ;
    wire new_AGEMA_signal_7825 ;
    wire new_AGEMA_signal_7826 ;
    wire new_AGEMA_signal_7827 ;
    wire new_AGEMA_signal_7828 ;
    wire new_AGEMA_signal_7829 ;
    wire new_AGEMA_signal_7830 ;
    wire new_AGEMA_signal_7831 ;
    wire new_AGEMA_signal_7832 ;
    wire new_AGEMA_signal_7833 ;
    wire new_AGEMA_signal_7834 ;
    wire new_AGEMA_signal_7835 ;
    wire new_AGEMA_signal_7836 ;
    wire new_AGEMA_signal_7837 ;
    wire new_AGEMA_signal_7838 ;
    wire new_AGEMA_signal_7839 ;
    wire new_AGEMA_signal_7840 ;
    wire new_AGEMA_signal_7841 ;
    wire new_AGEMA_signal_7842 ;
    wire new_AGEMA_signal_7843 ;
    wire new_AGEMA_signal_7844 ;
    wire new_AGEMA_signal_7845 ;
    wire new_AGEMA_signal_7846 ;
    wire new_AGEMA_signal_7847 ;
    wire new_AGEMA_signal_7848 ;
    wire new_AGEMA_signal_7849 ;
    wire new_AGEMA_signal_7850 ;
    wire new_AGEMA_signal_7851 ;
    wire new_AGEMA_signal_7852 ;
    wire new_AGEMA_signal_7853 ;
    wire new_AGEMA_signal_7854 ;
    wire new_AGEMA_signal_7855 ;
    wire new_AGEMA_signal_7856 ;
    wire new_AGEMA_signal_7857 ;
    wire new_AGEMA_signal_7858 ;
    wire new_AGEMA_signal_7859 ;
    wire new_AGEMA_signal_7860 ;
    wire new_AGEMA_signal_7861 ;
    wire new_AGEMA_signal_7862 ;
    wire new_AGEMA_signal_7863 ;
    wire new_AGEMA_signal_7864 ;
    wire new_AGEMA_signal_7865 ;
    wire new_AGEMA_signal_7866 ;
    wire new_AGEMA_signal_7867 ;
    wire new_AGEMA_signal_7868 ;
    wire new_AGEMA_signal_7869 ;
    wire new_AGEMA_signal_7870 ;
    wire new_AGEMA_signal_7871 ;
    wire new_AGEMA_signal_7872 ;
    wire new_AGEMA_signal_7873 ;
    wire new_AGEMA_signal_7874 ;
    wire new_AGEMA_signal_7875 ;
    wire new_AGEMA_signal_7876 ;
    wire new_AGEMA_signal_7877 ;
    wire new_AGEMA_signal_7878 ;
    wire new_AGEMA_signal_7879 ;
    wire new_AGEMA_signal_7880 ;
    wire new_AGEMA_signal_7881 ;
    wire new_AGEMA_signal_7882 ;
    wire new_AGEMA_signal_7883 ;
    wire new_AGEMA_signal_7884 ;
    wire new_AGEMA_signal_7885 ;
    wire new_AGEMA_signal_7886 ;
    wire new_AGEMA_signal_7887 ;
    wire new_AGEMA_signal_7888 ;
    wire new_AGEMA_signal_7889 ;
    wire new_AGEMA_signal_7890 ;
    wire new_AGEMA_signal_7891 ;
    wire new_AGEMA_signal_7892 ;
    wire new_AGEMA_signal_7893 ;
    wire new_AGEMA_signal_7894 ;
    wire new_AGEMA_signal_7895 ;
    wire new_AGEMA_signal_7896 ;
    wire new_AGEMA_signal_7897 ;
    wire new_AGEMA_signal_7898 ;
    wire new_AGEMA_signal_7899 ;
    wire new_AGEMA_signal_7900 ;
    wire new_AGEMA_signal_7901 ;
    wire new_AGEMA_signal_7902 ;
    wire new_AGEMA_signal_7903 ;
    wire new_AGEMA_signal_7904 ;
    wire new_AGEMA_signal_7905 ;
    wire new_AGEMA_signal_7906 ;
    wire new_AGEMA_signal_7907 ;
    wire new_AGEMA_signal_7908 ;
    wire new_AGEMA_signal_7909 ;
    wire new_AGEMA_signal_7910 ;
    wire new_AGEMA_signal_7911 ;
    wire new_AGEMA_signal_7912 ;
    wire new_AGEMA_signal_7913 ;
    wire new_AGEMA_signal_7914 ;
    wire new_AGEMA_signal_7915 ;
    wire new_AGEMA_signal_7916 ;
    wire new_AGEMA_signal_7917 ;
    wire new_AGEMA_signal_7918 ;
    wire new_AGEMA_signal_7919 ;
    wire new_AGEMA_signal_7920 ;
    wire new_AGEMA_signal_7921 ;
    wire new_AGEMA_signal_7922 ;
    wire new_AGEMA_signal_7923 ;
    wire new_AGEMA_signal_7924 ;
    wire new_AGEMA_signal_7925 ;
    wire new_AGEMA_signal_7926 ;
    wire new_AGEMA_signal_7927 ;
    wire new_AGEMA_signal_7928 ;
    wire new_AGEMA_signal_7929 ;
    wire new_AGEMA_signal_7930 ;
    wire new_AGEMA_signal_7931 ;
    wire new_AGEMA_signal_7932 ;
    wire new_AGEMA_signal_7933 ;
    wire new_AGEMA_signal_7934 ;
    wire new_AGEMA_signal_7935 ;
    wire new_AGEMA_signal_7936 ;
    wire new_AGEMA_signal_7937 ;
    wire new_AGEMA_signal_7938 ;
    wire new_AGEMA_signal_7939 ;
    wire new_AGEMA_signal_7940 ;
    wire new_AGEMA_signal_7941 ;
    wire new_AGEMA_signal_7942 ;
    wire new_AGEMA_signal_7943 ;
    wire new_AGEMA_signal_7944 ;
    wire new_AGEMA_signal_7945 ;
    wire new_AGEMA_signal_7946 ;
    wire new_AGEMA_signal_7947 ;
    wire new_AGEMA_signal_7948 ;
    wire new_AGEMA_signal_7949 ;
    wire new_AGEMA_signal_7950 ;
    wire new_AGEMA_signal_7951 ;
    wire new_AGEMA_signal_7952 ;
    wire new_AGEMA_signal_7953 ;
    wire new_AGEMA_signal_7954 ;
    wire new_AGEMA_signal_7955 ;
    wire new_AGEMA_signal_7956 ;
    wire new_AGEMA_signal_7957 ;
    wire new_AGEMA_signal_7958 ;
    wire new_AGEMA_signal_7959 ;
    wire new_AGEMA_signal_7960 ;
    wire new_AGEMA_signal_7961 ;
    wire new_AGEMA_signal_7962 ;
    wire new_AGEMA_signal_7963 ;
    wire new_AGEMA_signal_7964 ;
    wire new_AGEMA_signal_7965 ;
    wire new_AGEMA_signal_7966 ;
    wire new_AGEMA_signal_7967 ;
    wire new_AGEMA_signal_7968 ;
    wire new_AGEMA_signal_7969 ;
    wire new_AGEMA_signal_7970 ;
    wire new_AGEMA_signal_7971 ;
    wire new_AGEMA_signal_7972 ;
    wire new_AGEMA_signal_7973 ;
    wire new_AGEMA_signal_7974 ;
    wire new_AGEMA_signal_7975 ;
    wire new_AGEMA_signal_7976 ;
    wire new_AGEMA_signal_7977 ;
    wire new_AGEMA_signal_7978 ;
    wire new_AGEMA_signal_7979 ;
    wire new_AGEMA_signal_7980 ;
    wire new_AGEMA_signal_7981 ;
    wire new_AGEMA_signal_7982 ;
    wire new_AGEMA_signal_7983 ;
    wire new_AGEMA_signal_7984 ;
    wire new_AGEMA_signal_7985 ;
    wire new_AGEMA_signal_7986 ;
    wire new_AGEMA_signal_7987 ;
    wire new_AGEMA_signal_7988 ;
    wire new_AGEMA_signal_7989 ;
    wire new_AGEMA_signal_7990 ;
    wire new_AGEMA_signal_7991 ;
    wire new_AGEMA_signal_7992 ;
    wire new_AGEMA_signal_7993 ;
    wire new_AGEMA_signal_7994 ;
    wire new_AGEMA_signal_7995 ;
    wire new_AGEMA_signal_7996 ;
    wire new_AGEMA_signal_7997 ;
    wire new_AGEMA_signal_7998 ;
    wire new_AGEMA_signal_7999 ;
    wire new_AGEMA_signal_8000 ;
    wire new_AGEMA_signal_8001 ;
    wire new_AGEMA_signal_8002 ;
    wire new_AGEMA_signal_8003 ;
    wire new_AGEMA_signal_8004 ;
    wire new_AGEMA_signal_8005 ;
    wire new_AGEMA_signal_8006 ;
    wire new_AGEMA_signal_8007 ;
    wire new_AGEMA_signal_8008 ;
    wire new_AGEMA_signal_8009 ;
    wire new_AGEMA_signal_8010 ;
    wire new_AGEMA_signal_8011 ;
    wire new_AGEMA_signal_8012 ;
    wire new_AGEMA_signal_8013 ;
    wire new_AGEMA_signal_8014 ;
    wire new_AGEMA_signal_8015 ;
    wire new_AGEMA_signal_8016 ;
    wire new_AGEMA_signal_8017 ;
    wire new_AGEMA_signal_8018 ;
    wire new_AGEMA_signal_8019 ;
    wire new_AGEMA_signal_8020 ;
    wire new_AGEMA_signal_8021 ;
    wire new_AGEMA_signal_8022 ;
    wire new_AGEMA_signal_8023 ;
    wire new_AGEMA_signal_8024 ;
    wire new_AGEMA_signal_8025 ;
    wire new_AGEMA_signal_8026 ;
    wire new_AGEMA_signal_8027 ;
    wire new_AGEMA_signal_8028 ;
    wire new_AGEMA_signal_8029 ;
    wire new_AGEMA_signal_8030 ;
    wire new_AGEMA_signal_8031 ;
    wire new_AGEMA_signal_8032 ;
    wire new_AGEMA_signal_8033 ;
    wire new_AGEMA_signal_8034 ;
    wire new_AGEMA_signal_8035 ;
    wire new_AGEMA_signal_8036 ;
    wire new_AGEMA_signal_8037 ;
    wire new_AGEMA_signal_8038 ;
    wire new_AGEMA_signal_8039 ;
    wire new_AGEMA_signal_8040 ;
    wire new_AGEMA_signal_8041 ;
    wire new_AGEMA_signal_8042 ;
    wire new_AGEMA_signal_8043 ;
    wire new_AGEMA_signal_8044 ;
    wire new_AGEMA_signal_8045 ;
    wire new_AGEMA_signal_8046 ;
    wire new_AGEMA_signal_8047 ;
    wire new_AGEMA_signal_8048 ;
    wire new_AGEMA_signal_8049 ;
    wire new_AGEMA_signal_8050 ;
    wire new_AGEMA_signal_8051 ;
    wire new_AGEMA_signal_8052 ;
    wire new_AGEMA_signal_8053 ;
    wire new_AGEMA_signal_8054 ;
    wire new_AGEMA_signal_8055 ;
    wire new_AGEMA_signal_8056 ;
    wire new_AGEMA_signal_8057 ;
    wire new_AGEMA_signal_8058 ;
    wire new_AGEMA_signal_8059 ;
    wire new_AGEMA_signal_8060 ;
    wire new_AGEMA_signal_8061 ;
    wire new_AGEMA_signal_8062 ;
    wire new_AGEMA_signal_8063 ;
    wire new_AGEMA_signal_8064 ;
    wire new_AGEMA_signal_8065 ;
    wire new_AGEMA_signal_8066 ;
    wire new_AGEMA_signal_8067 ;
    wire new_AGEMA_signal_8068 ;
    wire new_AGEMA_signal_8069 ;
    wire new_AGEMA_signal_8070 ;
    wire new_AGEMA_signal_8071 ;
    wire new_AGEMA_signal_8072 ;
    wire new_AGEMA_signal_8073 ;
    wire new_AGEMA_signal_8074 ;
    wire new_AGEMA_signal_8075 ;
    wire new_AGEMA_signal_8076 ;
    wire new_AGEMA_signal_8077 ;
    wire new_AGEMA_signal_8078 ;
    wire new_AGEMA_signal_8079 ;
    wire new_AGEMA_signal_8080 ;
    wire new_AGEMA_signal_8081 ;
    wire new_AGEMA_signal_8082 ;
    wire new_AGEMA_signal_8083 ;
    wire new_AGEMA_signal_8084 ;
    wire new_AGEMA_signal_8085 ;
    wire new_AGEMA_signal_8086 ;
    wire new_AGEMA_signal_8087 ;
    wire new_AGEMA_signal_8088 ;
    wire new_AGEMA_signal_8089 ;
    wire new_AGEMA_signal_8090 ;
    wire new_AGEMA_signal_8091 ;
    wire new_AGEMA_signal_8092 ;
    wire new_AGEMA_signal_8093 ;
    wire new_AGEMA_signal_8094 ;
    wire new_AGEMA_signal_8095 ;
    wire new_AGEMA_signal_8096 ;
    wire new_AGEMA_signal_8097 ;
    wire new_AGEMA_signal_8098 ;
    wire new_AGEMA_signal_8099 ;
    wire new_AGEMA_signal_8100 ;
    wire new_AGEMA_signal_8101 ;
    wire new_AGEMA_signal_8102 ;
    wire new_AGEMA_signal_8103 ;
    wire new_AGEMA_signal_8104 ;
    wire new_AGEMA_signal_8105 ;
    wire new_AGEMA_signal_8106 ;
    wire new_AGEMA_signal_8107 ;
    wire new_AGEMA_signal_8108 ;
    wire new_AGEMA_signal_8109 ;
    wire new_AGEMA_signal_8110 ;
    wire new_AGEMA_signal_8111 ;
    wire new_AGEMA_signal_8112 ;
    wire new_AGEMA_signal_8113 ;
    wire new_AGEMA_signal_8114 ;
    wire new_AGEMA_signal_8115 ;
    wire new_AGEMA_signal_8116 ;
    wire new_AGEMA_signal_8117 ;
    wire new_AGEMA_signal_8118 ;
    wire new_AGEMA_signal_8119 ;
    wire new_AGEMA_signal_8120 ;
    wire new_AGEMA_signal_8121 ;
    wire new_AGEMA_signal_8122 ;
    wire new_AGEMA_signal_8123 ;
    wire new_AGEMA_signal_8124 ;
    wire new_AGEMA_signal_8125 ;
    wire new_AGEMA_signal_8126 ;
    wire new_AGEMA_signal_8127 ;
    wire new_AGEMA_signal_8128 ;
    wire new_AGEMA_signal_8129 ;
    wire new_AGEMA_signal_8130 ;
    wire new_AGEMA_signal_8131 ;
    wire new_AGEMA_signal_8132 ;
    wire new_AGEMA_signal_8133 ;
    wire new_AGEMA_signal_8134 ;
    wire new_AGEMA_signal_8135 ;
    wire new_AGEMA_signal_8136 ;
    wire new_AGEMA_signal_8137 ;
    wire new_AGEMA_signal_8138 ;
    wire new_AGEMA_signal_8139 ;
    wire new_AGEMA_signal_8140 ;
    wire new_AGEMA_signal_8141 ;
    wire new_AGEMA_signal_8142 ;
    wire new_AGEMA_signal_8143 ;
    wire new_AGEMA_signal_8144 ;
    wire new_AGEMA_signal_8145 ;
    wire new_AGEMA_signal_8146 ;
    wire new_AGEMA_signal_8147 ;
    wire new_AGEMA_signal_8148 ;
    wire new_AGEMA_signal_8149 ;
    wire new_AGEMA_signal_8150 ;
    wire new_AGEMA_signal_8151 ;
    wire new_AGEMA_signal_8152 ;
    wire new_AGEMA_signal_8153 ;
    wire new_AGEMA_signal_8154 ;
    wire new_AGEMA_signal_8155 ;
    wire new_AGEMA_signal_8156 ;
    wire new_AGEMA_signal_8157 ;
    wire new_AGEMA_signal_8158 ;
    wire new_AGEMA_signal_8159 ;
    wire new_AGEMA_signal_8160 ;
    wire new_AGEMA_signal_8161 ;
    wire new_AGEMA_signal_8162 ;
    wire new_AGEMA_signal_8163 ;
    wire new_AGEMA_signal_8164 ;
    wire new_AGEMA_signal_8165 ;
    wire new_AGEMA_signal_8166 ;
    wire new_AGEMA_signal_8167 ;
    wire new_AGEMA_signal_8168 ;
    wire new_AGEMA_signal_8169 ;
    wire new_AGEMA_signal_8170 ;
    wire new_AGEMA_signal_8171 ;
    wire new_AGEMA_signal_8172 ;
    wire new_AGEMA_signal_8173 ;
    wire new_AGEMA_signal_8174 ;
    wire new_AGEMA_signal_8175 ;
    wire new_AGEMA_signal_8176 ;
    wire new_AGEMA_signal_8177 ;
    wire new_AGEMA_signal_8178 ;
    wire new_AGEMA_signal_8179 ;
    wire new_AGEMA_signal_8180 ;
    wire new_AGEMA_signal_8181 ;
    wire new_AGEMA_signal_8182 ;
    wire new_AGEMA_signal_8183 ;
    wire new_AGEMA_signal_8184 ;
    wire new_AGEMA_signal_8185 ;
    wire new_AGEMA_signal_8186 ;
    wire new_AGEMA_signal_8187 ;
    wire new_AGEMA_signal_8188 ;
    wire new_AGEMA_signal_8189 ;
    wire new_AGEMA_signal_8190 ;

    /* cells in depth 0 */
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_U1 ( .a ({Ciphertext_s3[2], Ciphertext_s2[2], Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, SubCellInst_SboxInst_0_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_XOR_i1_U1 ( .a ({Ciphertext_s3[2], Ciphertext_s2[2], Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({Ciphertext_s3[3], Ciphertext_s2[3], Ciphertext_s1[3], Ciphertext_s0[3]}), .c ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, new_AGEMA_signal_1173, SubCellInst_SboxInst_0_XX_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_XOR_i2_U1 ( .a ({Ciphertext_s3[0], Ciphertext_s2[0], Ciphertext_s1[0], Ciphertext_s0[0]}), .b ({Ciphertext_s3[2], Ciphertext_s2[2], Ciphertext_s1[2], Ciphertext_s0[2]}), .c ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, new_AGEMA_signal_1179, SubCellInst_SboxInst_0_XX_2_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_XOR0_U1 ( .a ({Ciphertext_s3[1], Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, new_AGEMA_signal_1179, SubCellInst_SboxInst_0_XX_2_}), .c ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, new_AGEMA_signal_2031, SubCellInst_SboxInst_0_Q0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_XOR1_U1 ( .a ({Ciphertext_s3[1], Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, new_AGEMA_signal_1173, SubCellInst_SboxInst_0_XX_1_}), .c ({new_AGEMA_signal_2036, new_AGEMA_signal_2035, new_AGEMA_signal_2034, SubCellInst_SboxInst_0_Q1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_XOR3_U1 ( .a ({Ciphertext_s3[1], Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, SubCellInst_SboxInst_0_n3}), .c ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, new_AGEMA_signal_2037, SubCellInst_SboxInst_0_Q4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_XOR5_U1 ( .a ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, new_AGEMA_signal_1179, SubCellInst_SboxInst_0_XX_2_}), .b ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, SubCellInst_SboxInst_0_n3}), .c ({new_AGEMA_signal_2042, new_AGEMA_signal_2041, new_AGEMA_signal_2040, SubCellInst_SboxInst_0_Q6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_XOR6_U1 ( .a ({new_AGEMA_signal_2036, new_AGEMA_signal_2035, new_AGEMA_signal_2034, SubCellInst_SboxInst_0_Q1}), .b ({new_AGEMA_signal_2042, new_AGEMA_signal_2041, new_AGEMA_signal_2040, SubCellInst_SboxInst_0_Q6}), .c ({new_AGEMA_signal_2324, new_AGEMA_signal_2323, new_AGEMA_signal_2322, SubCellInst_SboxInst_0_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_XOR8_U1 ( .a ({Ciphertext_s3[1], Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, SubCellInst_SboxInst_0_n3}), .c ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, new_AGEMA_signal_2043, SubCellInst_SboxInst_0_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_U1 ( .a ({Ciphertext_s3[6], Ciphertext_s2[6], Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, SubCellInst_SboxInst_1_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_XOR_i1_U1 ( .a ({Ciphertext_s3[6], Ciphertext_s2[6], Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({Ciphertext_s3[7], Ciphertext_s2[7], Ciphertext_s1[7], Ciphertext_s0[7]}), .c ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, SubCellInst_SboxInst_1_XX_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_XOR_i2_U1 ( .a ({Ciphertext_s3[4], Ciphertext_s2[4], Ciphertext_s1[4], Ciphertext_s0[4]}), .b ({Ciphertext_s3[6], Ciphertext_s2[6], Ciphertext_s1[6], Ciphertext_s0[6]}), .c ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, SubCellInst_SboxInst_1_XX_2_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_XOR0_U1 ( .a ({Ciphertext_s3[5], Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, SubCellInst_SboxInst_1_XX_2_}), .c ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, new_AGEMA_signal_2049, SubCellInst_SboxInst_1_Q0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_XOR1_U1 ( .a ({Ciphertext_s3[5], Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, SubCellInst_SboxInst_1_XX_1_}), .c ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, new_AGEMA_signal_2052, SubCellInst_SboxInst_1_Q1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_XOR3_U1 ( .a ({Ciphertext_s3[5], Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, SubCellInst_SboxInst_1_n3}), .c ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, new_AGEMA_signal_2055, SubCellInst_SboxInst_1_Q4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_XOR5_U1 ( .a ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, SubCellInst_SboxInst_1_XX_2_}), .b ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, SubCellInst_SboxInst_1_n3}), .c ({new_AGEMA_signal_2060, new_AGEMA_signal_2059, new_AGEMA_signal_2058, SubCellInst_SboxInst_1_Q6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_XOR6_U1 ( .a ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, new_AGEMA_signal_2052, SubCellInst_SboxInst_1_Q1}), .b ({new_AGEMA_signal_2060, new_AGEMA_signal_2059, new_AGEMA_signal_2058, SubCellInst_SboxInst_1_Q6}), .c ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, new_AGEMA_signal_2331, SubCellInst_SboxInst_1_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_XOR8_U1 ( .a ({Ciphertext_s3[5], Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, SubCellInst_SboxInst_1_n3}), .c ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, new_AGEMA_signal_2061, SubCellInst_SboxInst_1_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_U1 ( .a ({Ciphertext_s3[10], Ciphertext_s2[10], Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, SubCellInst_SboxInst_2_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_XOR_i1_U1 ( .a ({Ciphertext_s3[10], Ciphertext_s2[10], Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({Ciphertext_s3[11], Ciphertext_s2[11], Ciphertext_s1[11], Ciphertext_s0[11]}), .c ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, SubCellInst_SboxInst_2_XX_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_XOR_i2_U1 ( .a ({Ciphertext_s3[8], Ciphertext_s2[8], Ciphertext_s1[8], Ciphertext_s0[8]}), .b ({Ciphertext_s3[10], Ciphertext_s2[10], Ciphertext_s1[10], Ciphertext_s0[10]}), .c ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, new_AGEMA_signal_1215, SubCellInst_SboxInst_2_XX_2_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_XOR0_U1 ( .a ({Ciphertext_s3[9], Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, new_AGEMA_signal_1215, SubCellInst_SboxInst_2_XX_2_}), .c ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, new_AGEMA_signal_2067, SubCellInst_SboxInst_2_Q0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_XOR1_U1 ( .a ({Ciphertext_s3[9], Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, SubCellInst_SboxInst_2_XX_1_}), .c ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, new_AGEMA_signal_2070, SubCellInst_SboxInst_2_Q1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_XOR3_U1 ( .a ({Ciphertext_s3[9], Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, SubCellInst_SboxInst_2_n3}), .c ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, new_AGEMA_signal_2073, SubCellInst_SboxInst_2_Q4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_XOR5_U1 ( .a ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, new_AGEMA_signal_1215, SubCellInst_SboxInst_2_XX_2_}), .b ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, SubCellInst_SboxInst_2_n3}), .c ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, new_AGEMA_signal_2076, SubCellInst_SboxInst_2_Q6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_XOR6_U1 ( .a ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, new_AGEMA_signal_2070, SubCellInst_SboxInst_2_Q1}), .b ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, new_AGEMA_signal_2076, SubCellInst_SboxInst_2_Q6}), .c ({new_AGEMA_signal_2342, new_AGEMA_signal_2341, new_AGEMA_signal_2340, SubCellInst_SboxInst_2_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_XOR8_U1 ( .a ({Ciphertext_s3[9], Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, SubCellInst_SboxInst_2_n3}), .c ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, new_AGEMA_signal_2079, SubCellInst_SboxInst_2_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_U1 ( .a ({Ciphertext_s3[14], Ciphertext_s2[14], Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, SubCellInst_SboxInst_3_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_XOR_i1_U1 ( .a ({Ciphertext_s3[14], Ciphertext_s2[14], Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({Ciphertext_s3[15], Ciphertext_s2[15], Ciphertext_s1[15], Ciphertext_s0[15]}), .c ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, SubCellInst_SboxInst_3_XX_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_XOR_i2_U1 ( .a ({Ciphertext_s3[12], Ciphertext_s2[12], Ciphertext_s1[12], Ciphertext_s0[12]}), .b ({Ciphertext_s3[14], Ciphertext_s2[14], Ciphertext_s1[14], Ciphertext_s0[14]}), .c ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, SubCellInst_SboxInst_3_XX_2_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_XOR0_U1 ( .a ({Ciphertext_s3[13], Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, SubCellInst_SboxInst_3_XX_2_}), .c ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, new_AGEMA_signal_2085, SubCellInst_SboxInst_3_Q0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_XOR1_U1 ( .a ({Ciphertext_s3[13], Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, SubCellInst_SboxInst_3_XX_1_}), .c ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, SubCellInst_SboxInst_3_Q1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_XOR3_U1 ( .a ({Ciphertext_s3[13], Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, SubCellInst_SboxInst_3_n3}), .c ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, new_AGEMA_signal_2091, SubCellInst_SboxInst_3_Q4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_XOR5_U1 ( .a ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, SubCellInst_SboxInst_3_XX_2_}), .b ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, SubCellInst_SboxInst_3_n3}), .c ({new_AGEMA_signal_2096, new_AGEMA_signal_2095, new_AGEMA_signal_2094, SubCellInst_SboxInst_3_Q6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_XOR6_U1 ( .a ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, SubCellInst_SboxInst_3_Q1}), .b ({new_AGEMA_signal_2096, new_AGEMA_signal_2095, new_AGEMA_signal_2094, SubCellInst_SboxInst_3_Q6}), .c ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, new_AGEMA_signal_2349, SubCellInst_SboxInst_3_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_XOR8_U1 ( .a ({Ciphertext_s3[13], Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, SubCellInst_SboxInst_3_n3}), .c ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, new_AGEMA_signal_2097, SubCellInst_SboxInst_3_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_U1 ( .a ({Ciphertext_s3[18], Ciphertext_s2[18], Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_4_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_XOR_i1_U1 ( .a ({Ciphertext_s3[18], Ciphertext_s2[18], Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({Ciphertext_s3[19], Ciphertext_s2[19], Ciphertext_s1[19], Ciphertext_s0[19]}), .c ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, new_AGEMA_signal_1245, SubCellInst_SboxInst_4_XX_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_XOR_i2_U1 ( .a ({Ciphertext_s3[16], Ciphertext_s2[16], Ciphertext_s1[16], Ciphertext_s0[16]}), .b ({Ciphertext_s3[18], Ciphertext_s2[18], Ciphertext_s1[18], Ciphertext_s0[18]}), .c ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, SubCellInst_SboxInst_4_XX_2_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_XOR0_U1 ( .a ({Ciphertext_s3[17], Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, SubCellInst_SboxInst_4_XX_2_}), .c ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, new_AGEMA_signal_2103, SubCellInst_SboxInst_4_Q0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_XOR1_U1 ( .a ({Ciphertext_s3[17], Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, new_AGEMA_signal_1245, SubCellInst_SboxInst_4_XX_1_}), .c ({new_AGEMA_signal_2108, new_AGEMA_signal_2107, new_AGEMA_signal_2106, SubCellInst_SboxInst_4_Q1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_XOR3_U1 ( .a ({Ciphertext_s3[17], Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_4_n3}), .c ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, new_AGEMA_signal_2109, SubCellInst_SboxInst_4_Q4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_XOR5_U1 ( .a ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, SubCellInst_SboxInst_4_XX_2_}), .b ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_4_n3}), .c ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, new_AGEMA_signal_2112, SubCellInst_SboxInst_4_Q6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_XOR6_U1 ( .a ({new_AGEMA_signal_2108, new_AGEMA_signal_2107, new_AGEMA_signal_2106, SubCellInst_SboxInst_4_Q1}), .b ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, new_AGEMA_signal_2112, SubCellInst_SboxInst_4_Q6}), .c ({new_AGEMA_signal_2360, new_AGEMA_signal_2359, new_AGEMA_signal_2358, SubCellInst_SboxInst_4_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_XOR8_U1 ( .a ({Ciphertext_s3[17], Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_4_n3}), .c ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, new_AGEMA_signal_2115, SubCellInst_SboxInst_4_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_U1 ( .a ({Ciphertext_s3[22], Ciphertext_s2[22], Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_5_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_XOR_i1_U1 ( .a ({Ciphertext_s3[22], Ciphertext_s2[22], Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({Ciphertext_s3[23], Ciphertext_s2[23], Ciphertext_s1[23], Ciphertext_s0[23]}), .c ({new_AGEMA_signal_1265, new_AGEMA_signal_1264, new_AGEMA_signal_1263, SubCellInst_SboxInst_5_XX_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_XOR_i2_U1 ( .a ({Ciphertext_s3[20], Ciphertext_s2[20], Ciphertext_s1[20], Ciphertext_s0[20]}), .b ({Ciphertext_s3[22], Ciphertext_s2[22], Ciphertext_s1[22], Ciphertext_s0[22]}), .c ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, SubCellInst_SboxInst_5_XX_2_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_XOR0_U1 ( .a ({Ciphertext_s3[21], Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, SubCellInst_SboxInst_5_XX_2_}), .c ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, new_AGEMA_signal_2121, SubCellInst_SboxInst_5_Q0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_XOR1_U1 ( .a ({Ciphertext_s3[21], Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1265, new_AGEMA_signal_1264, new_AGEMA_signal_1263, SubCellInst_SboxInst_5_XX_1_}), .c ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, new_AGEMA_signal_2124, SubCellInst_SboxInst_5_Q1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_XOR3_U1 ( .a ({Ciphertext_s3[21], Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_5_n3}), .c ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, new_AGEMA_signal_2127, SubCellInst_SboxInst_5_Q4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_XOR5_U1 ( .a ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, SubCellInst_SboxInst_5_XX_2_}), .b ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_5_n3}), .c ({new_AGEMA_signal_2132, new_AGEMA_signal_2131, new_AGEMA_signal_2130, SubCellInst_SboxInst_5_Q6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_XOR6_U1 ( .a ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, new_AGEMA_signal_2124, SubCellInst_SboxInst_5_Q1}), .b ({new_AGEMA_signal_2132, new_AGEMA_signal_2131, new_AGEMA_signal_2130, SubCellInst_SboxInst_5_Q6}), .c ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, new_AGEMA_signal_2367, SubCellInst_SboxInst_5_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_XOR8_U1 ( .a ({Ciphertext_s3[21], Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_5_n3}), .c ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, new_AGEMA_signal_2133, SubCellInst_SboxInst_5_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_U1 ( .a ({Ciphertext_s3[26], Ciphertext_s2[26], Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_6_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_XOR_i1_U1 ( .a ({Ciphertext_s3[26], Ciphertext_s2[26], Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({Ciphertext_s3[27], Ciphertext_s2[27], Ciphertext_s1[27], Ciphertext_s0[27]}), .c ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, new_AGEMA_signal_1281, SubCellInst_SboxInst_6_XX_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_XOR_i2_U1 ( .a ({Ciphertext_s3[24], Ciphertext_s2[24], Ciphertext_s1[24], Ciphertext_s0[24]}), .b ({Ciphertext_s3[26], Ciphertext_s2[26], Ciphertext_s1[26], Ciphertext_s0[26]}), .c ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, SubCellInst_SboxInst_6_XX_2_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_XOR0_U1 ( .a ({Ciphertext_s3[25], Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, SubCellInst_SboxInst_6_XX_2_}), .c ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, new_AGEMA_signal_2139, SubCellInst_SboxInst_6_Q0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_XOR1_U1 ( .a ({Ciphertext_s3[25], Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, new_AGEMA_signal_1281, SubCellInst_SboxInst_6_XX_1_}), .c ({new_AGEMA_signal_2144, new_AGEMA_signal_2143, new_AGEMA_signal_2142, SubCellInst_SboxInst_6_Q1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_XOR3_U1 ( .a ({Ciphertext_s3[25], Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_6_n3}), .c ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, new_AGEMA_signal_2145, SubCellInst_SboxInst_6_Q4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_XOR5_U1 ( .a ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, SubCellInst_SboxInst_6_XX_2_}), .b ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_6_n3}), .c ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, new_AGEMA_signal_2148, SubCellInst_SboxInst_6_Q6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_XOR6_U1 ( .a ({new_AGEMA_signal_2144, new_AGEMA_signal_2143, new_AGEMA_signal_2142, SubCellInst_SboxInst_6_Q1}), .b ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, new_AGEMA_signal_2148, SubCellInst_SboxInst_6_Q6}), .c ({new_AGEMA_signal_2378, new_AGEMA_signal_2377, new_AGEMA_signal_2376, SubCellInst_SboxInst_6_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_XOR8_U1 ( .a ({Ciphertext_s3[25], Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_6_n3}), .c ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, new_AGEMA_signal_2151, SubCellInst_SboxInst_6_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_U1 ( .a ({Ciphertext_s3[30], Ciphertext_s2[30], Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, SubCellInst_SboxInst_7_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_XOR_i1_U1 ( .a ({Ciphertext_s3[30], Ciphertext_s2[30], Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({Ciphertext_s3[31], Ciphertext_s2[31], Ciphertext_s1[31], Ciphertext_s0[31]}), .c ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, SubCellInst_SboxInst_7_XX_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_XOR_i2_U1 ( .a ({Ciphertext_s3[28], Ciphertext_s2[28], Ciphertext_s1[28], Ciphertext_s0[28]}), .b ({Ciphertext_s3[30], Ciphertext_s2[30], Ciphertext_s1[30], Ciphertext_s0[30]}), .c ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, SubCellInst_SboxInst_7_XX_2_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_XOR0_U1 ( .a ({Ciphertext_s3[29], Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, SubCellInst_SboxInst_7_XX_2_}), .c ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, new_AGEMA_signal_2157, SubCellInst_SboxInst_7_Q0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_XOR1_U1 ( .a ({Ciphertext_s3[29], Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, SubCellInst_SboxInst_7_XX_1_}), .c ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, new_AGEMA_signal_2160, SubCellInst_SboxInst_7_Q1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_XOR3_U1 ( .a ({Ciphertext_s3[29], Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, SubCellInst_SboxInst_7_n3}), .c ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, new_AGEMA_signal_2163, SubCellInst_SboxInst_7_Q4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_XOR5_U1 ( .a ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, SubCellInst_SboxInst_7_XX_2_}), .b ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, SubCellInst_SboxInst_7_n3}), .c ({new_AGEMA_signal_2168, new_AGEMA_signal_2167, new_AGEMA_signal_2166, SubCellInst_SboxInst_7_Q6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_XOR6_U1 ( .a ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, new_AGEMA_signal_2160, SubCellInst_SboxInst_7_Q1}), .b ({new_AGEMA_signal_2168, new_AGEMA_signal_2167, new_AGEMA_signal_2166, SubCellInst_SboxInst_7_Q6}), .c ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, new_AGEMA_signal_2385, SubCellInst_SboxInst_7_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_XOR8_U1 ( .a ({Ciphertext_s3[29], Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, SubCellInst_SboxInst_7_n3}), .c ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, new_AGEMA_signal_2169, SubCellInst_SboxInst_7_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_U1 ( .a ({Ciphertext_s3[34], Ciphertext_s2[34], Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, SubCellInst_SboxInst_8_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_XOR_i1_U1 ( .a ({Ciphertext_s3[34], Ciphertext_s2[34], Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({Ciphertext_s3[35], Ciphertext_s2[35], Ciphertext_s1[35], Ciphertext_s0[35]}), .c ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, SubCellInst_SboxInst_8_XX_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_XOR_i2_U1 ( .a ({Ciphertext_s3[32], Ciphertext_s2[32], Ciphertext_s1[32], Ciphertext_s0[32]}), .b ({Ciphertext_s3[34], Ciphertext_s2[34], Ciphertext_s1[34], Ciphertext_s0[34]}), .c ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, new_AGEMA_signal_1323, SubCellInst_SboxInst_8_XX_2_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_XOR0_U1 ( .a ({Ciphertext_s3[33], Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, new_AGEMA_signal_1323, SubCellInst_SboxInst_8_XX_2_}), .c ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, new_AGEMA_signal_2175, SubCellInst_SboxInst_8_Q0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_XOR1_U1 ( .a ({Ciphertext_s3[33], Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, SubCellInst_SboxInst_8_XX_1_}), .c ({new_AGEMA_signal_2180, new_AGEMA_signal_2179, new_AGEMA_signal_2178, SubCellInst_SboxInst_8_Q1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_XOR3_U1 ( .a ({Ciphertext_s3[33], Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, SubCellInst_SboxInst_8_n3}), .c ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, new_AGEMA_signal_2181, SubCellInst_SboxInst_8_Q4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_XOR5_U1 ( .a ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, new_AGEMA_signal_1323, SubCellInst_SboxInst_8_XX_2_}), .b ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, SubCellInst_SboxInst_8_n3}), .c ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, new_AGEMA_signal_2184, SubCellInst_SboxInst_8_Q6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_XOR6_U1 ( .a ({new_AGEMA_signal_2180, new_AGEMA_signal_2179, new_AGEMA_signal_2178, SubCellInst_SboxInst_8_Q1}), .b ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, new_AGEMA_signal_2184, SubCellInst_SboxInst_8_Q6}), .c ({new_AGEMA_signal_2396, new_AGEMA_signal_2395, new_AGEMA_signal_2394, SubCellInst_SboxInst_8_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_XOR8_U1 ( .a ({Ciphertext_s3[33], Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, SubCellInst_SboxInst_8_n3}), .c ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, new_AGEMA_signal_2187, SubCellInst_SboxInst_8_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_U1 ( .a ({Ciphertext_s3[38], Ciphertext_s2[38], Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, new_AGEMA_signal_1329, SubCellInst_SboxInst_9_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_XOR_i1_U1 ( .a ({Ciphertext_s3[38], Ciphertext_s2[38], Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({Ciphertext_s3[39], Ciphertext_s2[39], Ciphertext_s1[39], Ciphertext_s0[39]}), .c ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, new_AGEMA_signal_1335, SubCellInst_SboxInst_9_XX_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_XOR_i2_U1 ( .a ({Ciphertext_s3[36], Ciphertext_s2[36], Ciphertext_s1[36], Ciphertext_s0[36]}), .b ({Ciphertext_s3[38], Ciphertext_s2[38], Ciphertext_s1[38], Ciphertext_s0[38]}), .c ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, new_AGEMA_signal_1341, SubCellInst_SboxInst_9_XX_2_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_XOR0_U1 ( .a ({Ciphertext_s3[37], Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, new_AGEMA_signal_1341, SubCellInst_SboxInst_9_XX_2_}), .c ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, new_AGEMA_signal_2193, SubCellInst_SboxInst_9_Q0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_XOR1_U1 ( .a ({Ciphertext_s3[37], Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, new_AGEMA_signal_1335, SubCellInst_SboxInst_9_XX_1_}), .c ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, new_AGEMA_signal_2196, SubCellInst_SboxInst_9_Q1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_XOR3_U1 ( .a ({Ciphertext_s3[37], Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, new_AGEMA_signal_1329, SubCellInst_SboxInst_9_n3}), .c ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, new_AGEMA_signal_2199, SubCellInst_SboxInst_9_Q4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_XOR5_U1 ( .a ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, new_AGEMA_signal_1341, SubCellInst_SboxInst_9_XX_2_}), .b ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, new_AGEMA_signal_1329, SubCellInst_SboxInst_9_n3}), .c ({new_AGEMA_signal_2204, new_AGEMA_signal_2203, new_AGEMA_signal_2202, SubCellInst_SboxInst_9_Q6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_XOR6_U1 ( .a ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, new_AGEMA_signal_2196, SubCellInst_SboxInst_9_Q1}), .b ({new_AGEMA_signal_2204, new_AGEMA_signal_2203, new_AGEMA_signal_2202, SubCellInst_SboxInst_9_Q6}), .c ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, new_AGEMA_signal_2403, SubCellInst_SboxInst_9_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_XOR8_U1 ( .a ({Ciphertext_s3[37], Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, new_AGEMA_signal_1329, SubCellInst_SboxInst_9_n3}), .c ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, new_AGEMA_signal_2205, SubCellInst_SboxInst_9_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_U1 ( .a ({Ciphertext_s3[42], Ciphertext_s2[42], Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, SubCellInst_SboxInst_10_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_XOR_i1_U1 ( .a ({Ciphertext_s3[42], Ciphertext_s2[42], Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({Ciphertext_s3[43], Ciphertext_s2[43], Ciphertext_s1[43], Ciphertext_s0[43]}), .c ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, new_AGEMA_signal_1353, SubCellInst_SboxInst_10_XX_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_XOR_i2_U1 ( .a ({Ciphertext_s3[40], Ciphertext_s2[40], Ciphertext_s1[40], Ciphertext_s0[40]}), .b ({Ciphertext_s3[42], Ciphertext_s2[42], Ciphertext_s1[42], Ciphertext_s0[42]}), .c ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, SubCellInst_SboxInst_10_XX_2_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_XOR0_U1 ( .a ({Ciphertext_s3[41], Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, SubCellInst_SboxInst_10_XX_2_}), .c ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, new_AGEMA_signal_2211, SubCellInst_SboxInst_10_Q0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_XOR1_U1 ( .a ({Ciphertext_s3[41], Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, new_AGEMA_signal_1353, SubCellInst_SboxInst_10_XX_1_}), .c ({new_AGEMA_signal_2216, new_AGEMA_signal_2215, new_AGEMA_signal_2214, SubCellInst_SboxInst_10_Q1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_XOR3_U1 ( .a ({Ciphertext_s3[41], Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, SubCellInst_SboxInst_10_n3}), .c ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, new_AGEMA_signal_2217, SubCellInst_SboxInst_10_Q4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_XOR5_U1 ( .a ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, SubCellInst_SboxInst_10_XX_2_}), .b ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, SubCellInst_SboxInst_10_n3}), .c ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, new_AGEMA_signal_2220, SubCellInst_SboxInst_10_Q6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_XOR6_U1 ( .a ({new_AGEMA_signal_2216, new_AGEMA_signal_2215, new_AGEMA_signal_2214, SubCellInst_SboxInst_10_Q1}), .b ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, new_AGEMA_signal_2220, SubCellInst_SboxInst_10_Q6}), .c ({new_AGEMA_signal_2414, new_AGEMA_signal_2413, new_AGEMA_signal_2412, SubCellInst_SboxInst_10_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_XOR8_U1 ( .a ({Ciphertext_s3[41], Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, SubCellInst_SboxInst_10_n3}), .c ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, new_AGEMA_signal_2223, SubCellInst_SboxInst_10_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_U1 ( .a ({Ciphertext_s3[46], Ciphertext_s2[46], Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, new_AGEMA_signal_1365, SubCellInst_SboxInst_11_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_XOR_i1_U1 ( .a ({Ciphertext_s3[46], Ciphertext_s2[46], Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({Ciphertext_s3[47], Ciphertext_s2[47], Ciphertext_s1[47], Ciphertext_s0[47]}), .c ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, new_AGEMA_signal_1371, SubCellInst_SboxInst_11_XX_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_XOR_i2_U1 ( .a ({Ciphertext_s3[44], Ciphertext_s2[44], Ciphertext_s1[44], Ciphertext_s0[44]}), .b ({Ciphertext_s3[46], Ciphertext_s2[46], Ciphertext_s1[46], Ciphertext_s0[46]}), .c ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, SubCellInst_SboxInst_11_XX_2_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_XOR0_U1 ( .a ({Ciphertext_s3[45], Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, SubCellInst_SboxInst_11_XX_2_}), .c ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, new_AGEMA_signal_2229, SubCellInst_SboxInst_11_Q0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_XOR1_U1 ( .a ({Ciphertext_s3[45], Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, new_AGEMA_signal_1371, SubCellInst_SboxInst_11_XX_1_}), .c ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, new_AGEMA_signal_2232, SubCellInst_SboxInst_11_Q1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_XOR3_U1 ( .a ({Ciphertext_s3[45], Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, new_AGEMA_signal_1365, SubCellInst_SboxInst_11_n3}), .c ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, new_AGEMA_signal_2235, SubCellInst_SboxInst_11_Q4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_XOR5_U1 ( .a ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, SubCellInst_SboxInst_11_XX_2_}), .b ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, new_AGEMA_signal_1365, SubCellInst_SboxInst_11_n3}), .c ({new_AGEMA_signal_2240, new_AGEMA_signal_2239, new_AGEMA_signal_2238, SubCellInst_SboxInst_11_Q6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_XOR6_U1 ( .a ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, new_AGEMA_signal_2232, SubCellInst_SboxInst_11_Q1}), .b ({new_AGEMA_signal_2240, new_AGEMA_signal_2239, new_AGEMA_signal_2238, SubCellInst_SboxInst_11_Q6}), .c ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, new_AGEMA_signal_2421, SubCellInst_SboxInst_11_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_XOR8_U1 ( .a ({Ciphertext_s3[45], Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, new_AGEMA_signal_1365, SubCellInst_SboxInst_11_n3}), .c ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, new_AGEMA_signal_2241, SubCellInst_SboxInst_11_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_U1 ( .a ({Ciphertext_s3[50], Ciphertext_s2[50], Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, SubCellInst_SboxInst_12_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_XOR_i1_U1 ( .a ({Ciphertext_s3[50], Ciphertext_s2[50], Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({Ciphertext_s3[51], Ciphertext_s2[51], Ciphertext_s1[51], Ciphertext_s0[51]}), .c ({new_AGEMA_signal_1391, new_AGEMA_signal_1390, new_AGEMA_signal_1389, SubCellInst_SboxInst_12_XX_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_XOR_i2_U1 ( .a ({Ciphertext_s3[48], Ciphertext_s2[48], Ciphertext_s1[48], Ciphertext_s0[48]}), .b ({Ciphertext_s3[50], Ciphertext_s2[50], Ciphertext_s1[50], Ciphertext_s0[50]}), .c ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, SubCellInst_SboxInst_12_XX_2_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_XOR0_U1 ( .a ({Ciphertext_s3[49], Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, SubCellInst_SboxInst_12_XX_2_}), .c ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, new_AGEMA_signal_2247, SubCellInst_SboxInst_12_Q0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_XOR1_U1 ( .a ({Ciphertext_s3[49], Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1391, new_AGEMA_signal_1390, new_AGEMA_signal_1389, SubCellInst_SboxInst_12_XX_1_}), .c ({new_AGEMA_signal_2252, new_AGEMA_signal_2251, new_AGEMA_signal_2250, SubCellInst_SboxInst_12_Q1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_XOR3_U1 ( .a ({Ciphertext_s3[49], Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, SubCellInst_SboxInst_12_n3}), .c ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, new_AGEMA_signal_2253, SubCellInst_SboxInst_12_Q4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_XOR5_U1 ( .a ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, SubCellInst_SboxInst_12_XX_2_}), .b ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, SubCellInst_SboxInst_12_n3}), .c ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, new_AGEMA_signal_2256, SubCellInst_SboxInst_12_Q6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_XOR6_U1 ( .a ({new_AGEMA_signal_2252, new_AGEMA_signal_2251, new_AGEMA_signal_2250, SubCellInst_SboxInst_12_Q1}), .b ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, new_AGEMA_signal_2256, SubCellInst_SboxInst_12_Q6}), .c ({new_AGEMA_signal_2432, new_AGEMA_signal_2431, new_AGEMA_signal_2430, SubCellInst_SboxInst_12_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_XOR8_U1 ( .a ({Ciphertext_s3[49], Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, SubCellInst_SboxInst_12_n3}), .c ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, new_AGEMA_signal_2259, SubCellInst_SboxInst_12_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_U1 ( .a ({Ciphertext_s3[54], Ciphertext_s2[54], Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, SubCellInst_SboxInst_13_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_XOR_i1_U1 ( .a ({Ciphertext_s3[54], Ciphertext_s2[54], Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({Ciphertext_s3[55], Ciphertext_s2[55], Ciphertext_s1[55], Ciphertext_s0[55]}), .c ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, new_AGEMA_signal_1407, SubCellInst_SboxInst_13_XX_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_XOR_i2_U1 ( .a ({Ciphertext_s3[52], Ciphertext_s2[52], Ciphertext_s1[52], Ciphertext_s0[52]}), .b ({Ciphertext_s3[54], Ciphertext_s2[54], Ciphertext_s1[54], Ciphertext_s0[54]}), .c ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, new_AGEMA_signal_1413, SubCellInst_SboxInst_13_XX_2_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_XOR0_U1 ( .a ({Ciphertext_s3[53], Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, new_AGEMA_signal_1413, SubCellInst_SboxInst_13_XX_2_}), .c ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, new_AGEMA_signal_2265, SubCellInst_SboxInst_13_Q0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_XOR1_U1 ( .a ({Ciphertext_s3[53], Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, new_AGEMA_signal_1407, SubCellInst_SboxInst_13_XX_1_}), .c ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, new_AGEMA_signal_2268, SubCellInst_SboxInst_13_Q1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_XOR3_U1 ( .a ({Ciphertext_s3[53], Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, SubCellInst_SboxInst_13_n3}), .c ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, new_AGEMA_signal_2271, SubCellInst_SboxInst_13_Q4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_XOR5_U1 ( .a ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, new_AGEMA_signal_1413, SubCellInst_SboxInst_13_XX_2_}), .b ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, SubCellInst_SboxInst_13_n3}), .c ({new_AGEMA_signal_2276, new_AGEMA_signal_2275, new_AGEMA_signal_2274, SubCellInst_SboxInst_13_Q6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_XOR6_U1 ( .a ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, new_AGEMA_signal_2268, SubCellInst_SboxInst_13_Q1}), .b ({new_AGEMA_signal_2276, new_AGEMA_signal_2275, new_AGEMA_signal_2274, SubCellInst_SboxInst_13_Q6}), .c ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, new_AGEMA_signal_2439, SubCellInst_SboxInst_13_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_XOR8_U1 ( .a ({Ciphertext_s3[53], Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, SubCellInst_SboxInst_13_n3}), .c ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, new_AGEMA_signal_2277, SubCellInst_SboxInst_13_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_U1 ( .a ({Ciphertext_s3[58], Ciphertext_s2[58], Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, SubCellInst_SboxInst_14_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_XOR_i1_U1 ( .a ({Ciphertext_s3[58], Ciphertext_s2[58], Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({Ciphertext_s3[59], Ciphertext_s2[59], Ciphertext_s1[59], Ciphertext_s0[59]}), .c ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, new_AGEMA_signal_1425, SubCellInst_SboxInst_14_XX_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_XOR_i2_U1 ( .a ({Ciphertext_s3[56], Ciphertext_s2[56], Ciphertext_s1[56], Ciphertext_s0[56]}), .b ({Ciphertext_s3[58], Ciphertext_s2[58], Ciphertext_s1[58], Ciphertext_s0[58]}), .c ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, new_AGEMA_signal_1431, SubCellInst_SboxInst_14_XX_2_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_XOR0_U1 ( .a ({Ciphertext_s3[57], Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, new_AGEMA_signal_1431, SubCellInst_SboxInst_14_XX_2_}), .c ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, new_AGEMA_signal_2283, SubCellInst_SboxInst_14_Q0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_XOR1_U1 ( .a ({Ciphertext_s3[57], Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, new_AGEMA_signal_1425, SubCellInst_SboxInst_14_XX_1_}), .c ({new_AGEMA_signal_2288, new_AGEMA_signal_2287, new_AGEMA_signal_2286, SubCellInst_SboxInst_14_Q1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_XOR3_U1 ( .a ({Ciphertext_s3[57], Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, SubCellInst_SboxInst_14_n3}), .c ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, new_AGEMA_signal_2289, SubCellInst_SboxInst_14_Q4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_XOR5_U1 ( .a ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, new_AGEMA_signal_1431, SubCellInst_SboxInst_14_XX_2_}), .b ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, SubCellInst_SboxInst_14_n3}), .c ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, new_AGEMA_signal_2292, SubCellInst_SboxInst_14_Q6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_XOR6_U1 ( .a ({new_AGEMA_signal_2288, new_AGEMA_signal_2287, new_AGEMA_signal_2286, SubCellInst_SboxInst_14_Q1}), .b ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, new_AGEMA_signal_2292, SubCellInst_SboxInst_14_Q6}), .c ({new_AGEMA_signal_2450, new_AGEMA_signal_2449, new_AGEMA_signal_2448, SubCellInst_SboxInst_14_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_XOR8_U1 ( .a ({Ciphertext_s3[57], Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, SubCellInst_SboxInst_14_n3}), .c ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, new_AGEMA_signal_2295, SubCellInst_SboxInst_14_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_U1 ( .a ({Ciphertext_s3[62], Ciphertext_s2[62], Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, new_AGEMA_signal_1437, SubCellInst_SboxInst_15_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_XOR_i1_U1 ( .a ({Ciphertext_s3[62], Ciphertext_s2[62], Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({Ciphertext_s3[63], Ciphertext_s2[63], Ciphertext_s1[63], Ciphertext_s0[63]}), .c ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, new_AGEMA_signal_1443, SubCellInst_SboxInst_15_XX_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_XOR_i2_U1 ( .a ({Ciphertext_s3[60], Ciphertext_s2[60], Ciphertext_s1[60], Ciphertext_s0[60]}), .b ({Ciphertext_s3[62], Ciphertext_s2[62], Ciphertext_s1[62], Ciphertext_s0[62]}), .c ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, new_AGEMA_signal_1449, SubCellInst_SboxInst_15_XX_2_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_XOR0_U1 ( .a ({Ciphertext_s3[61], Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, new_AGEMA_signal_1449, SubCellInst_SboxInst_15_XX_2_}), .c ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, new_AGEMA_signal_2301, SubCellInst_SboxInst_15_Q0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_XOR1_U1 ( .a ({Ciphertext_s3[61], Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, new_AGEMA_signal_1443, SubCellInst_SboxInst_15_XX_1_}), .c ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, new_AGEMA_signal_2304, SubCellInst_SboxInst_15_Q1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_XOR3_U1 ( .a ({Ciphertext_s3[61], Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, new_AGEMA_signal_1437, SubCellInst_SboxInst_15_n3}), .c ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, new_AGEMA_signal_2307, SubCellInst_SboxInst_15_Q4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_XOR5_U1 ( .a ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, new_AGEMA_signal_1449, SubCellInst_SboxInst_15_XX_2_}), .b ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, new_AGEMA_signal_1437, SubCellInst_SboxInst_15_n3}), .c ({new_AGEMA_signal_2312, new_AGEMA_signal_2311, new_AGEMA_signal_2310, SubCellInst_SboxInst_15_Q6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_XOR6_U1 ( .a ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, new_AGEMA_signal_2304, SubCellInst_SboxInst_15_Q1}), .b ({new_AGEMA_signal_2312, new_AGEMA_signal_2311, new_AGEMA_signal_2310, SubCellInst_SboxInst_15_Q6}), .c ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, new_AGEMA_signal_2457, SubCellInst_SboxInst_15_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_XOR8_U1 ( .a ({Ciphertext_s3[61], Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, new_AGEMA_signal_1437, SubCellInst_SboxInst_15_n3}), .c ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, new_AGEMA_signal_2313, SubCellInst_SboxInst_15_L2}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_0_U1 ( .s (rst), .b ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, new_AGEMA_signal_1452, TweakeyGeneration_key_Feedback[0]}), .a ({Key_s3[0], Key_s2[0], Key_s1[0], Key_s0[0]}), .c ({new_AGEMA_signal_1460, new_AGEMA_signal_1459, new_AGEMA_signal_1458, TweakeyGeneration_StateRegInput[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_1_U1 ( .s (rst), .b ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, new_AGEMA_signal_1461, TweakeyGeneration_key_Feedback[1]}), .a ({Key_s3[1], Key_s2[1], Key_s1[1], Key_s0[1]}), .c ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, new_AGEMA_signal_1467, TweakeyGeneration_StateRegInput[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_2_U1 ( .s (rst), .b ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, new_AGEMA_signal_1470, TweakeyGeneration_key_Feedback[2]}), .a ({Key_s3[2], Key_s2[2], Key_s1[2], Key_s0[2]}), .c ({new_AGEMA_signal_1478, new_AGEMA_signal_1477, new_AGEMA_signal_1476, TweakeyGeneration_StateRegInput[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_3_U1 ( .s (rst), .b ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, new_AGEMA_signal_1479, TweakeyGeneration_key_Feedback[3]}), .a ({Key_s3[3], Key_s2[3], Key_s1[3], Key_s0[3]}), .c ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, new_AGEMA_signal_1485, TweakeyGeneration_StateRegInput[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_4_U1 ( .s (rst), .b ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, new_AGEMA_signal_1488, TweakeyGeneration_key_Feedback[4]}), .a ({Key_s3[4], Key_s2[4], Key_s1[4], Key_s0[4]}), .c ({new_AGEMA_signal_1496, new_AGEMA_signal_1495, new_AGEMA_signal_1494, TweakeyGeneration_StateRegInput[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_5_U1 ( .s (rst), .b ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, new_AGEMA_signal_1497, TweakeyGeneration_key_Feedback[5]}), .a ({Key_s3[5], Key_s2[5], Key_s1[5], Key_s0[5]}), .c ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, new_AGEMA_signal_1503, TweakeyGeneration_StateRegInput[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_6_U1 ( .s (rst), .b ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, new_AGEMA_signal_1506, TweakeyGeneration_key_Feedback[6]}), .a ({Key_s3[6], Key_s2[6], Key_s1[6], Key_s0[6]}), .c ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, new_AGEMA_signal_1512, TweakeyGeneration_StateRegInput[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_7_U1 ( .s (rst), .b ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, TweakeyGeneration_key_Feedback[7]}), .a ({Key_s3[7], Key_s2[7], Key_s1[7], Key_s0[7]}), .c ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, TweakeyGeneration_StateRegInput[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_8_U1 ( .s (rst), .b ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, new_AGEMA_signal_1524, TweakeyGeneration_key_Feedback[8]}), .a ({Key_s3[8], Key_s2[8], Key_s1[8], Key_s0[8]}), .c ({new_AGEMA_signal_1532, new_AGEMA_signal_1531, new_AGEMA_signal_1530, TweakeyGeneration_StateRegInput[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_9_U1 ( .s (rst), .b ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, new_AGEMA_signal_1533, TweakeyGeneration_key_Feedback[9]}), .a ({Key_s3[9], Key_s2[9], Key_s1[9], Key_s0[9]}), .c ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, new_AGEMA_signal_1539, TweakeyGeneration_StateRegInput[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_10_U1 ( .s (rst), .b ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, new_AGEMA_signal_1542, TweakeyGeneration_key_Feedback[10]}), .a ({Key_s3[10], Key_s2[10], Key_s1[10], Key_s0[10]}), .c ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, TweakeyGeneration_StateRegInput[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_11_U1 ( .s (rst), .b ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, new_AGEMA_signal_1551, TweakeyGeneration_key_Feedback[11]}), .a ({Key_s3[11], Key_s2[11], Key_s1[11], Key_s0[11]}), .c ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, new_AGEMA_signal_1557, TweakeyGeneration_StateRegInput[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_12_U1 ( .s (rst), .b ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, TweakeyGeneration_key_Feedback[12]}), .a ({Key_s3[12], Key_s2[12], Key_s1[12], Key_s0[12]}), .c ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, new_AGEMA_signal_1566, TweakeyGeneration_StateRegInput[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_13_U1 ( .s (rst), .b ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, new_AGEMA_signal_1569, TweakeyGeneration_key_Feedback[13]}), .a ({Key_s3[13], Key_s2[13], Key_s1[13], Key_s0[13]}), .c ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, new_AGEMA_signal_1575, TweakeyGeneration_StateRegInput[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_14_U1 ( .s (rst), .b ({new_AGEMA_signal_1580, new_AGEMA_signal_1579, new_AGEMA_signal_1578, TweakeyGeneration_key_Feedback[14]}), .a ({Key_s3[14], Key_s2[14], Key_s1[14], Key_s0[14]}), .c ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, new_AGEMA_signal_1584, TweakeyGeneration_StateRegInput[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_15_U1 ( .s (rst), .b ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, new_AGEMA_signal_1587, TweakeyGeneration_key_Feedback[15]}), .a ({Key_s3[15], Key_s2[15], Key_s1[15], Key_s0[15]}), .c ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, new_AGEMA_signal_1593, TweakeyGeneration_StateRegInput[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_16_U1 ( .s (rst), .b ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, new_AGEMA_signal_1596, TweakeyGeneration_key_Feedback[16]}), .a ({Key_s3[16], Key_s2[16], Key_s1[16], Key_s0[16]}), .c ({new_AGEMA_signal_1604, new_AGEMA_signal_1603, new_AGEMA_signal_1602, TweakeyGeneration_StateRegInput[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_17_U1 ( .s (rst), .b ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, TweakeyGeneration_key_Feedback[17]}), .a ({Key_s3[17], Key_s2[17], Key_s1[17], Key_s0[17]}), .c ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, new_AGEMA_signal_1611, TweakeyGeneration_StateRegInput[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_18_U1 ( .s (rst), .b ({new_AGEMA_signal_1616, new_AGEMA_signal_1615, new_AGEMA_signal_1614, TweakeyGeneration_key_Feedback[18]}), .a ({Key_s3[18], Key_s2[18], Key_s1[18], Key_s0[18]}), .c ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, new_AGEMA_signal_1620, TweakeyGeneration_StateRegInput[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_19_U1 ( .s (rst), .b ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, TweakeyGeneration_key_Feedback[19]}), .a ({Key_s3[19], Key_s2[19], Key_s1[19], Key_s0[19]}), .c ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, new_AGEMA_signal_1629, TweakeyGeneration_StateRegInput[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_20_U1 ( .s (rst), .b ({new_AGEMA_signal_1634, new_AGEMA_signal_1633, new_AGEMA_signal_1632, TweakeyGeneration_key_Feedback[20]}), .a ({Key_s3[20], Key_s2[20], Key_s1[20], Key_s0[20]}), .c ({new_AGEMA_signal_1640, new_AGEMA_signal_1639, new_AGEMA_signal_1638, TweakeyGeneration_StateRegInput[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_21_U1 ( .s (rst), .b ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, TweakeyGeneration_key_Feedback[21]}), .a ({Key_s3[21], Key_s2[21], Key_s1[21], Key_s0[21]}), .c ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, new_AGEMA_signal_1647, TweakeyGeneration_StateRegInput[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_22_U1 ( .s (rst), .b ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, new_AGEMA_signal_1650, TweakeyGeneration_key_Feedback[22]}), .a ({Key_s3[22], Key_s2[22], Key_s1[22], Key_s0[22]}), .c ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, new_AGEMA_signal_1656, TweakeyGeneration_StateRegInput[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_23_U1 ( .s (rst), .b ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, new_AGEMA_signal_1659, TweakeyGeneration_key_Feedback[23]}), .a ({Key_s3[23], Key_s2[23], Key_s1[23], Key_s0[23]}), .c ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, new_AGEMA_signal_1665, TweakeyGeneration_StateRegInput[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_24_U1 ( .s (rst), .b ({new_AGEMA_signal_1670, new_AGEMA_signal_1669, new_AGEMA_signal_1668, TweakeyGeneration_key_Feedback[24]}), .a ({Key_s3[24], Key_s2[24], Key_s1[24], Key_s0[24]}), .c ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, new_AGEMA_signal_1674, TweakeyGeneration_StateRegInput[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_25_U1 ( .s (rst), .b ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, new_AGEMA_signal_1677, TweakeyGeneration_key_Feedback[25]}), .a ({Key_s3[25], Key_s2[25], Key_s1[25], Key_s0[25]}), .c ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1683, TweakeyGeneration_StateRegInput[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_26_U1 ( .s (rst), .b ({new_AGEMA_signal_1688, new_AGEMA_signal_1687, new_AGEMA_signal_1686, TweakeyGeneration_key_Feedback[26]}), .a ({Key_s3[26], Key_s2[26], Key_s1[26], Key_s0[26]}), .c ({new_AGEMA_signal_1694, new_AGEMA_signal_1693, new_AGEMA_signal_1692, TweakeyGeneration_StateRegInput[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_27_U1 ( .s (rst), .b ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, new_AGEMA_signal_1695, TweakeyGeneration_key_Feedback[27]}), .a ({Key_s3[27], Key_s2[27], Key_s1[27], Key_s0[27]}), .c ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, new_AGEMA_signal_1701, TweakeyGeneration_StateRegInput[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_28_U1 ( .s (rst), .b ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, new_AGEMA_signal_1704, TweakeyGeneration_key_Feedback[28]}), .a ({Key_s3[28], Key_s2[28], Key_s1[28], Key_s0[28]}), .c ({new_AGEMA_signal_1712, new_AGEMA_signal_1711, new_AGEMA_signal_1710, TweakeyGeneration_StateRegInput[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_29_U1 ( .s (rst), .b ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, new_AGEMA_signal_1713, TweakeyGeneration_key_Feedback[29]}), .a ({Key_s3[29], Key_s2[29], Key_s1[29], Key_s0[29]}), .c ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, new_AGEMA_signal_1719, TweakeyGeneration_StateRegInput[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_30_U1 ( .s (rst), .b ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, new_AGEMA_signal_1722, TweakeyGeneration_key_Feedback[30]}), .a ({Key_s3[30], Key_s2[30], Key_s1[30], Key_s0[30]}), .c ({new_AGEMA_signal_1730, new_AGEMA_signal_1729, new_AGEMA_signal_1728, TweakeyGeneration_StateRegInput[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_31_U1 ( .s (rst), .b ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, new_AGEMA_signal_1731, TweakeyGeneration_key_Feedback[31]}), .a ({Key_s3[31], Key_s2[31], Key_s1[31], Key_s0[31]}), .c ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, new_AGEMA_signal_1737, TweakeyGeneration_StateRegInput[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_32_U1 ( .s (rst), .b ({new_AGEMA_signal_1742, new_AGEMA_signal_1741, new_AGEMA_signal_1740, TweakeyGeneration_key_Feedback[32]}), .a ({Key_s3[32], Key_s2[32], Key_s1[32], Key_s0[32]}), .c ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, new_AGEMA_signal_1746, TweakeyGeneration_StateRegInput[32]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_33_U1 ( .s (rst), .b ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, new_AGEMA_signal_1749, TweakeyGeneration_key_Feedback[33]}), .a ({Key_s3[33], Key_s2[33], Key_s1[33], Key_s0[33]}), .c ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, new_AGEMA_signal_1755, TweakeyGeneration_StateRegInput[33]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_34_U1 ( .s (rst), .b ({new_AGEMA_signal_1760, new_AGEMA_signal_1759, new_AGEMA_signal_1758, TweakeyGeneration_key_Feedback[34]}), .a ({Key_s3[34], Key_s2[34], Key_s1[34], Key_s0[34]}), .c ({new_AGEMA_signal_1766, new_AGEMA_signal_1765, new_AGEMA_signal_1764, TweakeyGeneration_StateRegInput[34]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_35_U1 ( .s (rst), .b ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, new_AGEMA_signal_1767, TweakeyGeneration_key_Feedback[35]}), .a ({Key_s3[35], Key_s2[35], Key_s1[35], Key_s0[35]}), .c ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, new_AGEMA_signal_1773, TweakeyGeneration_StateRegInput[35]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_36_U1 ( .s (rst), .b ({new_AGEMA_signal_1778, new_AGEMA_signal_1777, new_AGEMA_signal_1776, TweakeyGeneration_key_Feedback[36]}), .a ({Key_s3[36], Key_s2[36], Key_s1[36], Key_s0[36]}), .c ({new_AGEMA_signal_1784, new_AGEMA_signal_1783, new_AGEMA_signal_1782, TweakeyGeneration_StateRegInput[36]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_37_U1 ( .s (rst), .b ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, new_AGEMA_signal_1785, TweakeyGeneration_key_Feedback[37]}), .a ({Key_s3[37], Key_s2[37], Key_s1[37], Key_s0[37]}), .c ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, new_AGEMA_signal_1791, TweakeyGeneration_StateRegInput[37]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_38_U1 ( .s (rst), .b ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, new_AGEMA_signal_1794, TweakeyGeneration_key_Feedback[38]}), .a ({Key_s3[38], Key_s2[38], Key_s1[38], Key_s0[38]}), .c ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, new_AGEMA_signal_1800, TweakeyGeneration_StateRegInput[38]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_39_U1 ( .s (rst), .b ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, new_AGEMA_signal_1803, TweakeyGeneration_key_Feedback[39]}), .a ({Key_s3[39], Key_s2[39], Key_s1[39], Key_s0[39]}), .c ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, new_AGEMA_signal_1809, TweakeyGeneration_StateRegInput[39]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_40_U1 ( .s (rst), .b ({new_AGEMA_signal_1814, new_AGEMA_signal_1813, new_AGEMA_signal_1812, TweakeyGeneration_key_Feedback[40]}), .a ({Key_s3[40], Key_s2[40], Key_s1[40], Key_s0[40]}), .c ({new_AGEMA_signal_1820, new_AGEMA_signal_1819, new_AGEMA_signal_1818, TweakeyGeneration_StateRegInput[40]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_41_U1 ( .s (rst), .b ({new_AGEMA_signal_1823, new_AGEMA_signal_1822, new_AGEMA_signal_1821, TweakeyGeneration_key_Feedback[41]}), .a ({Key_s3[41], Key_s2[41], Key_s1[41], Key_s0[41]}), .c ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, new_AGEMA_signal_1827, TweakeyGeneration_StateRegInput[41]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_42_U1 ( .s (rst), .b ({new_AGEMA_signal_1832, new_AGEMA_signal_1831, new_AGEMA_signal_1830, TweakeyGeneration_key_Feedback[42]}), .a ({Key_s3[42], Key_s2[42], Key_s1[42], Key_s0[42]}), .c ({new_AGEMA_signal_1838, new_AGEMA_signal_1837, new_AGEMA_signal_1836, TweakeyGeneration_StateRegInput[42]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_43_U1 ( .s (rst), .b ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, new_AGEMA_signal_1839, TweakeyGeneration_key_Feedback[43]}), .a ({Key_s3[43], Key_s2[43], Key_s1[43], Key_s0[43]}), .c ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, new_AGEMA_signal_1845, TweakeyGeneration_StateRegInput[43]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_44_U1 ( .s (rst), .b ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, new_AGEMA_signal_1848, TweakeyGeneration_key_Feedback[44]}), .a ({Key_s3[44], Key_s2[44], Key_s1[44], Key_s0[44]}), .c ({new_AGEMA_signal_1856, new_AGEMA_signal_1855, new_AGEMA_signal_1854, TweakeyGeneration_StateRegInput[44]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_45_U1 ( .s (rst), .b ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, new_AGEMA_signal_1857, TweakeyGeneration_key_Feedback[45]}), .a ({Key_s3[45], Key_s2[45], Key_s1[45], Key_s0[45]}), .c ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, new_AGEMA_signal_1863, TweakeyGeneration_StateRegInput[45]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_46_U1 ( .s (rst), .b ({new_AGEMA_signal_1868, new_AGEMA_signal_1867, new_AGEMA_signal_1866, TweakeyGeneration_key_Feedback[46]}), .a ({Key_s3[46], Key_s2[46], Key_s1[46], Key_s0[46]}), .c ({new_AGEMA_signal_1874, new_AGEMA_signal_1873, new_AGEMA_signal_1872, TweakeyGeneration_StateRegInput[46]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_47_U1 ( .s (rst), .b ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, new_AGEMA_signal_1875, TweakeyGeneration_key_Feedback[47]}), .a ({Key_s3[47], Key_s2[47], Key_s1[47], Key_s0[47]}), .c ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, new_AGEMA_signal_1881, TweakeyGeneration_StateRegInput[47]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_48_U1 ( .s (rst), .b ({new_AGEMA_signal_1886, new_AGEMA_signal_1885, new_AGEMA_signal_1884, TweakeyGeneration_key_Feedback[48]}), .a ({Key_s3[48], Key_s2[48], Key_s1[48], Key_s0[48]}), .c ({new_AGEMA_signal_1892, new_AGEMA_signal_1891, new_AGEMA_signal_1890, TweakeyGeneration_StateRegInput[48]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_49_U1 ( .s (rst), .b ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, new_AGEMA_signal_1893, TweakeyGeneration_key_Feedback[49]}), .a ({Key_s3[49], Key_s2[49], Key_s1[49], Key_s0[49]}), .c ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, new_AGEMA_signal_1899, TweakeyGeneration_StateRegInput[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_50_U1 ( .s (rst), .b ({new_AGEMA_signal_1904, new_AGEMA_signal_1903, new_AGEMA_signal_1902, TweakeyGeneration_key_Feedback[50]}), .a ({Key_s3[50], Key_s2[50], Key_s1[50], Key_s0[50]}), .c ({new_AGEMA_signal_1910, new_AGEMA_signal_1909, new_AGEMA_signal_1908, TweakeyGeneration_StateRegInput[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_51_U1 ( .s (rst), .b ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, new_AGEMA_signal_1911, TweakeyGeneration_key_Feedback[51]}), .a ({Key_s3[51], Key_s2[51], Key_s1[51], Key_s0[51]}), .c ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, new_AGEMA_signal_1917, TweakeyGeneration_StateRegInput[51]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_52_U1 ( .s (rst), .b ({new_AGEMA_signal_1922, new_AGEMA_signal_1921, new_AGEMA_signal_1920, TweakeyGeneration_key_Feedback[52]}), .a ({Key_s3[52], Key_s2[52], Key_s1[52], Key_s0[52]}), .c ({new_AGEMA_signal_1928, new_AGEMA_signal_1927, new_AGEMA_signal_1926, TweakeyGeneration_StateRegInput[52]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_53_U1 ( .s (rst), .b ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, new_AGEMA_signal_1929, TweakeyGeneration_key_Feedback[53]}), .a ({Key_s3[53], Key_s2[53], Key_s1[53], Key_s0[53]}), .c ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, new_AGEMA_signal_1935, TweakeyGeneration_StateRegInput[53]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_54_U1 ( .s (rst), .b ({new_AGEMA_signal_1940, new_AGEMA_signal_1939, new_AGEMA_signal_1938, TweakeyGeneration_key_Feedback[54]}), .a ({Key_s3[54], Key_s2[54], Key_s1[54], Key_s0[54]}), .c ({new_AGEMA_signal_1946, new_AGEMA_signal_1945, new_AGEMA_signal_1944, TweakeyGeneration_StateRegInput[54]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_55_U1 ( .s (rst), .b ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, new_AGEMA_signal_1947, TweakeyGeneration_key_Feedback[55]}), .a ({Key_s3[55], Key_s2[55], Key_s1[55], Key_s0[55]}), .c ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, new_AGEMA_signal_1953, TweakeyGeneration_StateRegInput[55]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_56_U1 ( .s (rst), .b ({new_AGEMA_signal_1958, new_AGEMA_signal_1957, new_AGEMA_signal_1956, TweakeyGeneration_key_Feedback[56]}), .a ({Key_s3[56], Key_s2[56], Key_s1[56], Key_s0[56]}), .c ({new_AGEMA_signal_1964, new_AGEMA_signal_1963, new_AGEMA_signal_1962, TweakeyGeneration_StateRegInput[56]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_57_U1 ( .s (rst), .b ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, new_AGEMA_signal_1965, TweakeyGeneration_key_Feedback[57]}), .a ({Key_s3[57], Key_s2[57], Key_s1[57], Key_s0[57]}), .c ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, new_AGEMA_signal_1971, TweakeyGeneration_StateRegInput[57]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_58_U1 ( .s (rst), .b ({new_AGEMA_signal_1976, new_AGEMA_signal_1975, new_AGEMA_signal_1974, TweakeyGeneration_key_Feedback[58]}), .a ({Key_s3[58], Key_s2[58], Key_s1[58], Key_s0[58]}), .c ({new_AGEMA_signal_1982, new_AGEMA_signal_1981, new_AGEMA_signal_1980, TweakeyGeneration_StateRegInput[58]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_59_U1 ( .s (rst), .b ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, new_AGEMA_signal_1983, TweakeyGeneration_key_Feedback[59]}), .a ({Key_s3[59], Key_s2[59], Key_s1[59], Key_s0[59]}), .c ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, new_AGEMA_signal_1989, TweakeyGeneration_StateRegInput[59]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_60_U1 ( .s (rst), .b ({new_AGEMA_signal_1994, new_AGEMA_signal_1993, new_AGEMA_signal_1992, TweakeyGeneration_key_Feedback[60]}), .a ({Key_s3[60], Key_s2[60], Key_s1[60], Key_s0[60]}), .c ({new_AGEMA_signal_2000, new_AGEMA_signal_1999, new_AGEMA_signal_1998, TweakeyGeneration_StateRegInput[60]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_61_U1 ( .s (rst), .b ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, new_AGEMA_signal_2001, TweakeyGeneration_key_Feedback[61]}), .a ({Key_s3[61], Key_s2[61], Key_s1[61], Key_s0[61]}), .c ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, new_AGEMA_signal_2007, TweakeyGeneration_StateRegInput[61]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_62_U1 ( .s (rst), .b ({new_AGEMA_signal_2012, new_AGEMA_signal_2011, new_AGEMA_signal_2010, TweakeyGeneration_key_Feedback[62]}), .a ({Key_s3[62], Key_s2[62], Key_s1[62], Key_s0[62]}), .c ({new_AGEMA_signal_2018, new_AGEMA_signal_2017, new_AGEMA_signal_2016, TweakeyGeneration_StateRegInput[62]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_63_U1 ( .s (rst), .b ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, new_AGEMA_signal_2019, TweakeyGeneration_key_Feedback[63]}), .a ({Key_s3[63], Key_s2[63], Key_s1[63], Key_s0[63]}), .c ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, new_AGEMA_signal_2025, TweakeyGeneration_StateRegInput[63]}) ) ;
    MUX2_X1 FSMMUX_MUXInst_0_U1 ( .S (rst), .A (FSMUpdate[0]), .B (1'b1), .Z (FSMSelected[0]) ) ;
    MUX2_X1 FSMMUX_MUXInst_1_U1 ( .S (rst), .A (FSMUpdate[1]), .B (1'b0), .Z (FSMSelected[1]) ) ;
    MUX2_X1 FSMMUX_MUXInst_2_U1 ( .S (rst), .A (FSMUpdate[2]), .B (1'b0), .Z (FSMSelected[2]) ) ;
    MUX2_X1 FSMMUX_MUXInst_3_U1 ( .S (rst), .A (FSMUpdate[3]), .B (1'b0), .Z (FSMSelected[3]) ) ;
    MUX2_X1 FSMMUX_MUXInst_4_U1 ( .S (rst), .A (FSMUpdate[4]), .B (1'b0), .Z (FSMSelected[4]) ) ;
    MUX2_X1 FSMMUX_MUXInst_5_U1 ( .S (rst), .A (FSMUpdate[5]), .B (1'b0), .Z (FSMSelected[5]) ) ;
    MUX2_X1 FSMUpdateInst_StateUpdateInst_0_U5 ( .S (FSM[4]), .A (FSMUpdateInst_StateUpdateInst_0_n4), .B (FSM[5]), .Z (FSMUpdate[0]) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_0_U4 ( .A1 (FSM[5]), .A2 (FSMUpdateInst_StateUpdateInst_0_n3), .ZN (FSMUpdateInst_StateUpdateInst_0_n4) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_0_U3 ( .A1 (FSMUpdateInst_StateUpdateInst_0_n2), .A2 (FSMUpdateInst_StateUpdateInst_0_n1), .ZN (FSMUpdateInst_StateUpdateInst_0_n3) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_0_U2 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdate[4]), .ZN (FSMUpdateInst_StateUpdateInst_0_n1) ) ;
    AND2_X1 FSMUpdateInst_StateUpdateInst_0_U1 ( .A1 (FSMUpdate[1]), .A2 (FSM[1]), .ZN (FSMUpdateInst_StateUpdateInst_0_n2) ) ;
    AND2_X1 FSMUpdateInst_StateUpdateInst_2_U5 ( .A1 (FSMUpdateInst_StateUpdateInst_2_n4), .A2 (FSM[1]), .ZN (FSMUpdate[2]) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_2_U4 ( .A1 (FSMUpdateInst_StateUpdateInst_2_n3), .A2 (FSM[5]), .ZN (FSMUpdateInst_StateUpdateInst_2_n4) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_2_U3 ( .A1 (FSM[4]), .A2 (FSMUpdateInst_StateUpdateInst_2_n2), .ZN (FSMUpdateInst_StateUpdateInst_2_n3) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_2_U2 ( .A1 (FSMUpdate[1]), .A2 (FSMUpdateInst_StateUpdateInst_2_n1), .ZN (FSMUpdateInst_StateUpdateInst_2_n2) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_2_U1 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdate[4]), .ZN (FSMUpdateInst_StateUpdateInst_2_n1) ) ;
    OR2_X1 FSMUpdateInst_StateUpdateInst_5_U5 ( .A1 (FSM[4]), .A2 (FSMUpdateInst_StateUpdateInst_5_n4), .ZN (FSMUpdate[5]) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_5_U4 ( .A1 (FSMUpdate[4]), .A2 (FSMUpdateInst_StateUpdateInst_5_n3), .ZN (FSMUpdateInst_StateUpdateInst_5_n4) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_5_U3 ( .A1 (FSM[5]), .A2 (FSMUpdateInst_StateUpdateInst_5_n2), .ZN (FSMUpdateInst_StateUpdateInst_5_n3) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_5_U2 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdateInst_StateUpdateInst_5_n1), .ZN (FSMUpdateInst_StateUpdateInst_5_n2) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_5_U1 ( .A1 (FSMUpdate[1]), .A2 (FSM[1]), .ZN (FSMUpdateInst_StateUpdateInst_5_n1) ) ;
    NOR2_X1 FSMSignalsInst_doneInst_U6 ( .A1 (FSMSignalsInst_doneInst_n5), .A2 (FSMSignalsInst_doneInst_n4), .ZN (done) ) ;
    NAND2_X1 FSMSignalsInst_doneInst_U5 ( .A1 (FSM[4]), .A2 (FSM[5]), .ZN (FSMSignalsInst_doneInst_n4) ) ;
    NAND2_X1 FSMSignalsInst_doneInst_U4 ( .A1 (FSMSignalsInst_doneInst_n3), .A2 (FSMSignalsInst_doneInst_n2), .ZN (FSMSignalsInst_doneInst_n5) ) ;
    NOR2_X1 FSMSignalsInst_doneInst_U3 ( .A1 (FSMUpdate[4]), .A2 (FSMSignalsInst_doneInst_n1), .ZN (FSMSignalsInst_doneInst_n2) ) ;
    INV_X1 FSMSignalsInst_doneInst_U2 ( .A (FSMUpdate[1]), .ZN (FSMSignalsInst_doneInst_n1) ) ;
    NOR2_X1 FSMSignalsInst_doneInst_U1 ( .A1 (FSM[1]), .A2 (FSMUpdate[3]), .ZN (FSMSignalsInst_doneInst_n3) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_1000 ( .C (clk), .D (rst), .Q (new_AGEMA_signal_4431) ) ;
    buf_clk new_AGEMA_reg_buffer_1002 ( .C (clk), .D (Plaintext_s0[2]), .Q (new_AGEMA_signal_4433) ) ;
    buf_clk new_AGEMA_reg_buffer_1004 ( .C (clk), .D (Plaintext_s1[2]), .Q (new_AGEMA_signal_4435) ) ;
    buf_clk new_AGEMA_reg_buffer_1006 ( .C (clk), .D (Plaintext_s2[2]), .Q (new_AGEMA_signal_4437) ) ;
    buf_clk new_AGEMA_reg_buffer_1008 ( .C (clk), .D (Plaintext_s3[2]), .Q (new_AGEMA_signal_4439) ) ;
    buf_clk new_AGEMA_reg_buffer_1010 ( .C (clk), .D (Plaintext_s0[3]), .Q (new_AGEMA_signal_4441) ) ;
    buf_clk new_AGEMA_reg_buffer_1012 ( .C (clk), .D (Plaintext_s1[3]), .Q (new_AGEMA_signal_4443) ) ;
    buf_clk new_AGEMA_reg_buffer_1014 ( .C (clk), .D (Plaintext_s2[3]), .Q (new_AGEMA_signal_4445) ) ;
    buf_clk new_AGEMA_reg_buffer_1016 ( .C (clk), .D (Plaintext_s3[3]), .Q (new_AGEMA_signal_4447) ) ;
    buf_clk new_AGEMA_reg_buffer_1018 ( .C (clk), .D (Plaintext_s0[6]), .Q (new_AGEMA_signal_4449) ) ;
    buf_clk new_AGEMA_reg_buffer_1020 ( .C (clk), .D (Plaintext_s1[6]), .Q (new_AGEMA_signal_4451) ) ;
    buf_clk new_AGEMA_reg_buffer_1022 ( .C (clk), .D (Plaintext_s2[6]), .Q (new_AGEMA_signal_4453) ) ;
    buf_clk new_AGEMA_reg_buffer_1024 ( .C (clk), .D (Plaintext_s3[6]), .Q (new_AGEMA_signal_4455) ) ;
    buf_clk new_AGEMA_reg_buffer_1026 ( .C (clk), .D (Plaintext_s0[7]), .Q (new_AGEMA_signal_4457) ) ;
    buf_clk new_AGEMA_reg_buffer_1028 ( .C (clk), .D (Plaintext_s1[7]), .Q (new_AGEMA_signal_4459) ) ;
    buf_clk new_AGEMA_reg_buffer_1030 ( .C (clk), .D (Plaintext_s2[7]), .Q (new_AGEMA_signal_4461) ) ;
    buf_clk new_AGEMA_reg_buffer_1032 ( .C (clk), .D (Plaintext_s3[7]), .Q (new_AGEMA_signal_4463) ) ;
    buf_clk new_AGEMA_reg_buffer_1034 ( .C (clk), .D (Plaintext_s0[10]), .Q (new_AGEMA_signal_4465) ) ;
    buf_clk new_AGEMA_reg_buffer_1036 ( .C (clk), .D (Plaintext_s1[10]), .Q (new_AGEMA_signal_4467) ) ;
    buf_clk new_AGEMA_reg_buffer_1038 ( .C (clk), .D (Plaintext_s2[10]), .Q (new_AGEMA_signal_4469) ) ;
    buf_clk new_AGEMA_reg_buffer_1040 ( .C (clk), .D (Plaintext_s3[10]), .Q (new_AGEMA_signal_4471) ) ;
    buf_clk new_AGEMA_reg_buffer_1042 ( .C (clk), .D (Plaintext_s0[11]), .Q (new_AGEMA_signal_4473) ) ;
    buf_clk new_AGEMA_reg_buffer_1044 ( .C (clk), .D (Plaintext_s1[11]), .Q (new_AGEMA_signal_4475) ) ;
    buf_clk new_AGEMA_reg_buffer_1046 ( .C (clk), .D (Plaintext_s2[11]), .Q (new_AGEMA_signal_4477) ) ;
    buf_clk new_AGEMA_reg_buffer_1048 ( .C (clk), .D (Plaintext_s3[11]), .Q (new_AGEMA_signal_4479) ) ;
    buf_clk new_AGEMA_reg_buffer_1050 ( .C (clk), .D (Plaintext_s0[14]), .Q (new_AGEMA_signal_4481) ) ;
    buf_clk new_AGEMA_reg_buffer_1052 ( .C (clk), .D (Plaintext_s1[14]), .Q (new_AGEMA_signal_4483) ) ;
    buf_clk new_AGEMA_reg_buffer_1054 ( .C (clk), .D (Plaintext_s2[14]), .Q (new_AGEMA_signal_4485) ) ;
    buf_clk new_AGEMA_reg_buffer_1056 ( .C (clk), .D (Plaintext_s3[14]), .Q (new_AGEMA_signal_4487) ) ;
    buf_clk new_AGEMA_reg_buffer_1058 ( .C (clk), .D (Plaintext_s0[15]), .Q (new_AGEMA_signal_4489) ) ;
    buf_clk new_AGEMA_reg_buffer_1060 ( .C (clk), .D (Plaintext_s1[15]), .Q (new_AGEMA_signal_4491) ) ;
    buf_clk new_AGEMA_reg_buffer_1062 ( .C (clk), .D (Plaintext_s2[15]), .Q (new_AGEMA_signal_4493) ) ;
    buf_clk new_AGEMA_reg_buffer_1064 ( .C (clk), .D (Plaintext_s3[15]), .Q (new_AGEMA_signal_4495) ) ;
    buf_clk new_AGEMA_reg_buffer_1066 ( .C (clk), .D (Plaintext_s0[18]), .Q (new_AGEMA_signal_4497) ) ;
    buf_clk new_AGEMA_reg_buffer_1068 ( .C (clk), .D (Plaintext_s1[18]), .Q (new_AGEMA_signal_4499) ) ;
    buf_clk new_AGEMA_reg_buffer_1070 ( .C (clk), .D (Plaintext_s2[18]), .Q (new_AGEMA_signal_4501) ) ;
    buf_clk new_AGEMA_reg_buffer_1072 ( .C (clk), .D (Plaintext_s3[18]), .Q (new_AGEMA_signal_4503) ) ;
    buf_clk new_AGEMA_reg_buffer_1074 ( .C (clk), .D (Plaintext_s0[19]), .Q (new_AGEMA_signal_4505) ) ;
    buf_clk new_AGEMA_reg_buffer_1076 ( .C (clk), .D (Plaintext_s1[19]), .Q (new_AGEMA_signal_4507) ) ;
    buf_clk new_AGEMA_reg_buffer_1078 ( .C (clk), .D (Plaintext_s2[19]), .Q (new_AGEMA_signal_4509) ) ;
    buf_clk new_AGEMA_reg_buffer_1080 ( .C (clk), .D (Plaintext_s3[19]), .Q (new_AGEMA_signal_4511) ) ;
    buf_clk new_AGEMA_reg_buffer_1082 ( .C (clk), .D (Plaintext_s0[22]), .Q (new_AGEMA_signal_4513) ) ;
    buf_clk new_AGEMA_reg_buffer_1084 ( .C (clk), .D (Plaintext_s1[22]), .Q (new_AGEMA_signal_4515) ) ;
    buf_clk new_AGEMA_reg_buffer_1086 ( .C (clk), .D (Plaintext_s2[22]), .Q (new_AGEMA_signal_4517) ) ;
    buf_clk new_AGEMA_reg_buffer_1088 ( .C (clk), .D (Plaintext_s3[22]), .Q (new_AGEMA_signal_4519) ) ;
    buf_clk new_AGEMA_reg_buffer_1090 ( .C (clk), .D (Plaintext_s0[23]), .Q (new_AGEMA_signal_4521) ) ;
    buf_clk new_AGEMA_reg_buffer_1092 ( .C (clk), .D (Plaintext_s1[23]), .Q (new_AGEMA_signal_4523) ) ;
    buf_clk new_AGEMA_reg_buffer_1094 ( .C (clk), .D (Plaintext_s2[23]), .Q (new_AGEMA_signal_4525) ) ;
    buf_clk new_AGEMA_reg_buffer_1096 ( .C (clk), .D (Plaintext_s3[23]), .Q (new_AGEMA_signal_4527) ) ;
    buf_clk new_AGEMA_reg_buffer_1098 ( .C (clk), .D (Plaintext_s0[26]), .Q (new_AGEMA_signal_4529) ) ;
    buf_clk new_AGEMA_reg_buffer_1100 ( .C (clk), .D (Plaintext_s1[26]), .Q (new_AGEMA_signal_4531) ) ;
    buf_clk new_AGEMA_reg_buffer_1102 ( .C (clk), .D (Plaintext_s2[26]), .Q (new_AGEMA_signal_4533) ) ;
    buf_clk new_AGEMA_reg_buffer_1104 ( .C (clk), .D (Plaintext_s3[26]), .Q (new_AGEMA_signal_4535) ) ;
    buf_clk new_AGEMA_reg_buffer_1106 ( .C (clk), .D (Plaintext_s0[27]), .Q (new_AGEMA_signal_4537) ) ;
    buf_clk new_AGEMA_reg_buffer_1108 ( .C (clk), .D (Plaintext_s1[27]), .Q (new_AGEMA_signal_4539) ) ;
    buf_clk new_AGEMA_reg_buffer_1110 ( .C (clk), .D (Plaintext_s2[27]), .Q (new_AGEMA_signal_4541) ) ;
    buf_clk new_AGEMA_reg_buffer_1112 ( .C (clk), .D (Plaintext_s3[27]), .Q (new_AGEMA_signal_4543) ) ;
    buf_clk new_AGEMA_reg_buffer_1114 ( .C (clk), .D (Plaintext_s0[30]), .Q (new_AGEMA_signal_4545) ) ;
    buf_clk new_AGEMA_reg_buffer_1116 ( .C (clk), .D (Plaintext_s1[30]), .Q (new_AGEMA_signal_4547) ) ;
    buf_clk new_AGEMA_reg_buffer_1118 ( .C (clk), .D (Plaintext_s2[30]), .Q (new_AGEMA_signal_4549) ) ;
    buf_clk new_AGEMA_reg_buffer_1120 ( .C (clk), .D (Plaintext_s3[30]), .Q (new_AGEMA_signal_4551) ) ;
    buf_clk new_AGEMA_reg_buffer_1122 ( .C (clk), .D (Plaintext_s0[31]), .Q (new_AGEMA_signal_4553) ) ;
    buf_clk new_AGEMA_reg_buffer_1124 ( .C (clk), .D (Plaintext_s1[31]), .Q (new_AGEMA_signal_4555) ) ;
    buf_clk new_AGEMA_reg_buffer_1126 ( .C (clk), .D (Plaintext_s2[31]), .Q (new_AGEMA_signal_4557) ) ;
    buf_clk new_AGEMA_reg_buffer_1128 ( .C (clk), .D (Plaintext_s3[31]), .Q (new_AGEMA_signal_4559) ) ;
    buf_clk new_AGEMA_reg_buffer_1130 ( .C (clk), .D (Plaintext_s0[34]), .Q (new_AGEMA_signal_4561) ) ;
    buf_clk new_AGEMA_reg_buffer_1132 ( .C (clk), .D (Plaintext_s1[34]), .Q (new_AGEMA_signal_4563) ) ;
    buf_clk new_AGEMA_reg_buffer_1134 ( .C (clk), .D (Plaintext_s2[34]), .Q (new_AGEMA_signal_4565) ) ;
    buf_clk new_AGEMA_reg_buffer_1136 ( .C (clk), .D (Plaintext_s3[34]), .Q (new_AGEMA_signal_4567) ) ;
    buf_clk new_AGEMA_reg_buffer_1138 ( .C (clk), .D (Plaintext_s0[35]), .Q (new_AGEMA_signal_4569) ) ;
    buf_clk new_AGEMA_reg_buffer_1140 ( .C (clk), .D (Plaintext_s1[35]), .Q (new_AGEMA_signal_4571) ) ;
    buf_clk new_AGEMA_reg_buffer_1142 ( .C (clk), .D (Plaintext_s2[35]), .Q (new_AGEMA_signal_4573) ) ;
    buf_clk new_AGEMA_reg_buffer_1144 ( .C (clk), .D (Plaintext_s3[35]), .Q (new_AGEMA_signal_4575) ) ;
    buf_clk new_AGEMA_reg_buffer_1146 ( .C (clk), .D (Plaintext_s0[38]), .Q (new_AGEMA_signal_4577) ) ;
    buf_clk new_AGEMA_reg_buffer_1148 ( .C (clk), .D (Plaintext_s1[38]), .Q (new_AGEMA_signal_4579) ) ;
    buf_clk new_AGEMA_reg_buffer_1150 ( .C (clk), .D (Plaintext_s2[38]), .Q (new_AGEMA_signal_4581) ) ;
    buf_clk new_AGEMA_reg_buffer_1152 ( .C (clk), .D (Plaintext_s3[38]), .Q (new_AGEMA_signal_4583) ) ;
    buf_clk new_AGEMA_reg_buffer_1154 ( .C (clk), .D (Plaintext_s0[39]), .Q (new_AGEMA_signal_4585) ) ;
    buf_clk new_AGEMA_reg_buffer_1156 ( .C (clk), .D (Plaintext_s1[39]), .Q (new_AGEMA_signal_4587) ) ;
    buf_clk new_AGEMA_reg_buffer_1158 ( .C (clk), .D (Plaintext_s2[39]), .Q (new_AGEMA_signal_4589) ) ;
    buf_clk new_AGEMA_reg_buffer_1160 ( .C (clk), .D (Plaintext_s3[39]), .Q (new_AGEMA_signal_4591) ) ;
    buf_clk new_AGEMA_reg_buffer_1162 ( .C (clk), .D (Plaintext_s0[42]), .Q (new_AGEMA_signal_4593) ) ;
    buf_clk new_AGEMA_reg_buffer_1164 ( .C (clk), .D (Plaintext_s1[42]), .Q (new_AGEMA_signal_4595) ) ;
    buf_clk new_AGEMA_reg_buffer_1166 ( .C (clk), .D (Plaintext_s2[42]), .Q (new_AGEMA_signal_4597) ) ;
    buf_clk new_AGEMA_reg_buffer_1168 ( .C (clk), .D (Plaintext_s3[42]), .Q (new_AGEMA_signal_4599) ) ;
    buf_clk new_AGEMA_reg_buffer_1170 ( .C (clk), .D (Plaintext_s0[43]), .Q (new_AGEMA_signal_4601) ) ;
    buf_clk new_AGEMA_reg_buffer_1172 ( .C (clk), .D (Plaintext_s1[43]), .Q (new_AGEMA_signal_4603) ) ;
    buf_clk new_AGEMA_reg_buffer_1174 ( .C (clk), .D (Plaintext_s2[43]), .Q (new_AGEMA_signal_4605) ) ;
    buf_clk new_AGEMA_reg_buffer_1176 ( .C (clk), .D (Plaintext_s3[43]), .Q (new_AGEMA_signal_4607) ) ;
    buf_clk new_AGEMA_reg_buffer_1178 ( .C (clk), .D (Plaintext_s0[46]), .Q (new_AGEMA_signal_4609) ) ;
    buf_clk new_AGEMA_reg_buffer_1180 ( .C (clk), .D (Plaintext_s1[46]), .Q (new_AGEMA_signal_4611) ) ;
    buf_clk new_AGEMA_reg_buffer_1182 ( .C (clk), .D (Plaintext_s2[46]), .Q (new_AGEMA_signal_4613) ) ;
    buf_clk new_AGEMA_reg_buffer_1184 ( .C (clk), .D (Plaintext_s3[46]), .Q (new_AGEMA_signal_4615) ) ;
    buf_clk new_AGEMA_reg_buffer_1186 ( .C (clk), .D (Plaintext_s0[47]), .Q (new_AGEMA_signal_4617) ) ;
    buf_clk new_AGEMA_reg_buffer_1188 ( .C (clk), .D (Plaintext_s1[47]), .Q (new_AGEMA_signal_4619) ) ;
    buf_clk new_AGEMA_reg_buffer_1190 ( .C (clk), .D (Plaintext_s2[47]), .Q (new_AGEMA_signal_4621) ) ;
    buf_clk new_AGEMA_reg_buffer_1192 ( .C (clk), .D (Plaintext_s3[47]), .Q (new_AGEMA_signal_4623) ) ;
    buf_clk new_AGEMA_reg_buffer_1194 ( .C (clk), .D (Plaintext_s0[50]), .Q (new_AGEMA_signal_4625) ) ;
    buf_clk new_AGEMA_reg_buffer_1196 ( .C (clk), .D (Plaintext_s1[50]), .Q (new_AGEMA_signal_4627) ) ;
    buf_clk new_AGEMA_reg_buffer_1198 ( .C (clk), .D (Plaintext_s2[50]), .Q (new_AGEMA_signal_4629) ) ;
    buf_clk new_AGEMA_reg_buffer_1200 ( .C (clk), .D (Plaintext_s3[50]), .Q (new_AGEMA_signal_4631) ) ;
    buf_clk new_AGEMA_reg_buffer_1202 ( .C (clk), .D (Plaintext_s0[51]), .Q (new_AGEMA_signal_4633) ) ;
    buf_clk new_AGEMA_reg_buffer_1204 ( .C (clk), .D (Plaintext_s1[51]), .Q (new_AGEMA_signal_4635) ) ;
    buf_clk new_AGEMA_reg_buffer_1206 ( .C (clk), .D (Plaintext_s2[51]), .Q (new_AGEMA_signal_4637) ) ;
    buf_clk new_AGEMA_reg_buffer_1208 ( .C (clk), .D (Plaintext_s3[51]), .Q (new_AGEMA_signal_4639) ) ;
    buf_clk new_AGEMA_reg_buffer_1210 ( .C (clk), .D (Plaintext_s0[54]), .Q (new_AGEMA_signal_4641) ) ;
    buf_clk new_AGEMA_reg_buffer_1212 ( .C (clk), .D (Plaintext_s1[54]), .Q (new_AGEMA_signal_4643) ) ;
    buf_clk new_AGEMA_reg_buffer_1214 ( .C (clk), .D (Plaintext_s2[54]), .Q (new_AGEMA_signal_4645) ) ;
    buf_clk new_AGEMA_reg_buffer_1216 ( .C (clk), .D (Plaintext_s3[54]), .Q (new_AGEMA_signal_4647) ) ;
    buf_clk new_AGEMA_reg_buffer_1218 ( .C (clk), .D (Plaintext_s0[55]), .Q (new_AGEMA_signal_4649) ) ;
    buf_clk new_AGEMA_reg_buffer_1220 ( .C (clk), .D (Plaintext_s1[55]), .Q (new_AGEMA_signal_4651) ) ;
    buf_clk new_AGEMA_reg_buffer_1222 ( .C (clk), .D (Plaintext_s2[55]), .Q (new_AGEMA_signal_4653) ) ;
    buf_clk new_AGEMA_reg_buffer_1224 ( .C (clk), .D (Plaintext_s3[55]), .Q (new_AGEMA_signal_4655) ) ;
    buf_clk new_AGEMA_reg_buffer_1226 ( .C (clk), .D (Plaintext_s0[58]), .Q (new_AGEMA_signal_4657) ) ;
    buf_clk new_AGEMA_reg_buffer_1228 ( .C (clk), .D (Plaintext_s1[58]), .Q (new_AGEMA_signal_4659) ) ;
    buf_clk new_AGEMA_reg_buffer_1230 ( .C (clk), .D (Plaintext_s2[58]), .Q (new_AGEMA_signal_4661) ) ;
    buf_clk new_AGEMA_reg_buffer_1232 ( .C (clk), .D (Plaintext_s3[58]), .Q (new_AGEMA_signal_4663) ) ;
    buf_clk new_AGEMA_reg_buffer_1234 ( .C (clk), .D (Plaintext_s0[59]), .Q (new_AGEMA_signal_4665) ) ;
    buf_clk new_AGEMA_reg_buffer_1236 ( .C (clk), .D (Plaintext_s1[59]), .Q (new_AGEMA_signal_4667) ) ;
    buf_clk new_AGEMA_reg_buffer_1238 ( .C (clk), .D (Plaintext_s2[59]), .Q (new_AGEMA_signal_4669) ) ;
    buf_clk new_AGEMA_reg_buffer_1240 ( .C (clk), .D (Plaintext_s3[59]), .Q (new_AGEMA_signal_4671) ) ;
    buf_clk new_AGEMA_reg_buffer_1242 ( .C (clk), .D (Plaintext_s0[62]), .Q (new_AGEMA_signal_4673) ) ;
    buf_clk new_AGEMA_reg_buffer_1244 ( .C (clk), .D (Plaintext_s1[62]), .Q (new_AGEMA_signal_4675) ) ;
    buf_clk new_AGEMA_reg_buffer_1246 ( .C (clk), .D (Plaintext_s2[62]), .Q (new_AGEMA_signal_4677) ) ;
    buf_clk new_AGEMA_reg_buffer_1248 ( .C (clk), .D (Plaintext_s3[62]), .Q (new_AGEMA_signal_4679) ) ;
    buf_clk new_AGEMA_reg_buffer_1250 ( .C (clk), .D (Plaintext_s0[63]), .Q (new_AGEMA_signal_4681) ) ;
    buf_clk new_AGEMA_reg_buffer_1252 ( .C (clk), .D (Plaintext_s1[63]), .Q (new_AGEMA_signal_4683) ) ;
    buf_clk new_AGEMA_reg_buffer_1254 ( .C (clk), .D (Plaintext_s2[63]), .Q (new_AGEMA_signal_4685) ) ;
    buf_clk new_AGEMA_reg_buffer_1256 ( .C (clk), .D (Plaintext_s3[63]), .Q (new_AGEMA_signal_4687) ) ;
    buf_clk new_AGEMA_reg_buffer_1258 ( .C (clk), .D (SubCellInst_SboxInst_0_Q0), .Q (new_AGEMA_signal_4689) ) ;
    buf_clk new_AGEMA_reg_buffer_1260 ( .C (clk), .D (new_AGEMA_signal_2031), .Q (new_AGEMA_signal_4691) ) ;
    buf_clk new_AGEMA_reg_buffer_1262 ( .C (clk), .D (new_AGEMA_signal_2032), .Q (new_AGEMA_signal_4693) ) ;
    buf_clk new_AGEMA_reg_buffer_1264 ( .C (clk), .D (new_AGEMA_signal_2033), .Q (new_AGEMA_signal_4695) ) ;
    buf_clk new_AGEMA_reg_buffer_1266 ( .C (clk), .D (SubCellInst_SboxInst_0_L1), .Q (new_AGEMA_signal_4697) ) ;
    buf_clk new_AGEMA_reg_buffer_1268 ( .C (clk), .D (new_AGEMA_signal_2322), .Q (new_AGEMA_signal_4699) ) ;
    buf_clk new_AGEMA_reg_buffer_1270 ( .C (clk), .D (new_AGEMA_signal_2323), .Q (new_AGEMA_signal_4701) ) ;
    buf_clk new_AGEMA_reg_buffer_1272 ( .C (clk), .D (new_AGEMA_signal_2324), .Q (new_AGEMA_signal_4703) ) ;
    buf_clk new_AGEMA_reg_buffer_1274 ( .C (clk), .D (SubCellInst_SboxInst_0_XX_2_), .Q (new_AGEMA_signal_4705) ) ;
    buf_clk new_AGEMA_reg_buffer_1276 ( .C (clk), .D (new_AGEMA_signal_1179), .Q (new_AGEMA_signal_4707) ) ;
    buf_clk new_AGEMA_reg_buffer_1278 ( .C (clk), .D (new_AGEMA_signal_1180), .Q (new_AGEMA_signal_4709) ) ;
    buf_clk new_AGEMA_reg_buffer_1280 ( .C (clk), .D (new_AGEMA_signal_1181), .Q (new_AGEMA_signal_4711) ) ;
    buf_clk new_AGEMA_reg_buffer_1282 ( .C (clk), .D (SubCellInst_SboxInst_0_XX_1_), .Q (new_AGEMA_signal_4713) ) ;
    buf_clk new_AGEMA_reg_buffer_1284 ( .C (clk), .D (new_AGEMA_signal_1173), .Q (new_AGEMA_signal_4715) ) ;
    buf_clk new_AGEMA_reg_buffer_1286 ( .C (clk), .D (new_AGEMA_signal_1174), .Q (new_AGEMA_signal_4717) ) ;
    buf_clk new_AGEMA_reg_buffer_1288 ( .C (clk), .D (new_AGEMA_signal_1175), .Q (new_AGEMA_signal_4719) ) ;
    buf_clk new_AGEMA_reg_buffer_1290 ( .C (clk), .D (SubCellInst_SboxInst_1_Q0), .Q (new_AGEMA_signal_4721) ) ;
    buf_clk new_AGEMA_reg_buffer_1292 ( .C (clk), .D (new_AGEMA_signal_2049), .Q (new_AGEMA_signal_4723) ) ;
    buf_clk new_AGEMA_reg_buffer_1294 ( .C (clk), .D (new_AGEMA_signal_2050), .Q (new_AGEMA_signal_4725) ) ;
    buf_clk new_AGEMA_reg_buffer_1296 ( .C (clk), .D (new_AGEMA_signal_2051), .Q (new_AGEMA_signal_4727) ) ;
    buf_clk new_AGEMA_reg_buffer_1298 ( .C (clk), .D (SubCellInst_SboxInst_1_L1), .Q (new_AGEMA_signal_4729) ) ;
    buf_clk new_AGEMA_reg_buffer_1300 ( .C (clk), .D (new_AGEMA_signal_2331), .Q (new_AGEMA_signal_4731) ) ;
    buf_clk new_AGEMA_reg_buffer_1302 ( .C (clk), .D (new_AGEMA_signal_2332), .Q (new_AGEMA_signal_4733) ) ;
    buf_clk new_AGEMA_reg_buffer_1304 ( .C (clk), .D (new_AGEMA_signal_2333), .Q (new_AGEMA_signal_4735) ) ;
    buf_clk new_AGEMA_reg_buffer_1306 ( .C (clk), .D (SubCellInst_SboxInst_1_XX_2_), .Q (new_AGEMA_signal_4737) ) ;
    buf_clk new_AGEMA_reg_buffer_1308 ( .C (clk), .D (new_AGEMA_signal_1197), .Q (new_AGEMA_signal_4739) ) ;
    buf_clk new_AGEMA_reg_buffer_1310 ( .C (clk), .D (new_AGEMA_signal_1198), .Q (new_AGEMA_signal_4741) ) ;
    buf_clk new_AGEMA_reg_buffer_1312 ( .C (clk), .D (new_AGEMA_signal_1199), .Q (new_AGEMA_signal_4743) ) ;
    buf_clk new_AGEMA_reg_buffer_1314 ( .C (clk), .D (SubCellInst_SboxInst_1_XX_1_), .Q (new_AGEMA_signal_4745) ) ;
    buf_clk new_AGEMA_reg_buffer_1316 ( .C (clk), .D (new_AGEMA_signal_1191), .Q (new_AGEMA_signal_4747) ) ;
    buf_clk new_AGEMA_reg_buffer_1318 ( .C (clk), .D (new_AGEMA_signal_1192), .Q (new_AGEMA_signal_4749) ) ;
    buf_clk new_AGEMA_reg_buffer_1320 ( .C (clk), .D (new_AGEMA_signal_1193), .Q (new_AGEMA_signal_4751) ) ;
    buf_clk new_AGEMA_reg_buffer_1322 ( .C (clk), .D (SubCellInst_SboxInst_2_Q0), .Q (new_AGEMA_signal_4753) ) ;
    buf_clk new_AGEMA_reg_buffer_1324 ( .C (clk), .D (new_AGEMA_signal_2067), .Q (new_AGEMA_signal_4755) ) ;
    buf_clk new_AGEMA_reg_buffer_1326 ( .C (clk), .D (new_AGEMA_signal_2068), .Q (new_AGEMA_signal_4757) ) ;
    buf_clk new_AGEMA_reg_buffer_1328 ( .C (clk), .D (new_AGEMA_signal_2069), .Q (new_AGEMA_signal_4759) ) ;
    buf_clk new_AGEMA_reg_buffer_1330 ( .C (clk), .D (SubCellInst_SboxInst_2_L1), .Q (new_AGEMA_signal_4761) ) ;
    buf_clk new_AGEMA_reg_buffer_1332 ( .C (clk), .D (new_AGEMA_signal_2340), .Q (new_AGEMA_signal_4763) ) ;
    buf_clk new_AGEMA_reg_buffer_1334 ( .C (clk), .D (new_AGEMA_signal_2341), .Q (new_AGEMA_signal_4765) ) ;
    buf_clk new_AGEMA_reg_buffer_1336 ( .C (clk), .D (new_AGEMA_signal_2342), .Q (new_AGEMA_signal_4767) ) ;
    buf_clk new_AGEMA_reg_buffer_1338 ( .C (clk), .D (SubCellInst_SboxInst_2_XX_2_), .Q (new_AGEMA_signal_4769) ) ;
    buf_clk new_AGEMA_reg_buffer_1340 ( .C (clk), .D (new_AGEMA_signal_1215), .Q (new_AGEMA_signal_4771) ) ;
    buf_clk new_AGEMA_reg_buffer_1342 ( .C (clk), .D (new_AGEMA_signal_1216), .Q (new_AGEMA_signal_4773) ) ;
    buf_clk new_AGEMA_reg_buffer_1344 ( .C (clk), .D (new_AGEMA_signal_1217), .Q (new_AGEMA_signal_4775) ) ;
    buf_clk new_AGEMA_reg_buffer_1346 ( .C (clk), .D (SubCellInst_SboxInst_2_XX_1_), .Q (new_AGEMA_signal_4777) ) ;
    buf_clk new_AGEMA_reg_buffer_1348 ( .C (clk), .D (new_AGEMA_signal_1209), .Q (new_AGEMA_signal_4779) ) ;
    buf_clk new_AGEMA_reg_buffer_1350 ( .C (clk), .D (new_AGEMA_signal_1210), .Q (new_AGEMA_signal_4781) ) ;
    buf_clk new_AGEMA_reg_buffer_1352 ( .C (clk), .D (new_AGEMA_signal_1211), .Q (new_AGEMA_signal_4783) ) ;
    buf_clk new_AGEMA_reg_buffer_1354 ( .C (clk), .D (SubCellInst_SboxInst_3_Q0), .Q (new_AGEMA_signal_4785) ) ;
    buf_clk new_AGEMA_reg_buffer_1356 ( .C (clk), .D (new_AGEMA_signal_2085), .Q (new_AGEMA_signal_4787) ) ;
    buf_clk new_AGEMA_reg_buffer_1358 ( .C (clk), .D (new_AGEMA_signal_2086), .Q (new_AGEMA_signal_4789) ) ;
    buf_clk new_AGEMA_reg_buffer_1360 ( .C (clk), .D (new_AGEMA_signal_2087), .Q (new_AGEMA_signal_4791) ) ;
    buf_clk new_AGEMA_reg_buffer_1362 ( .C (clk), .D (SubCellInst_SboxInst_3_L1), .Q (new_AGEMA_signal_4793) ) ;
    buf_clk new_AGEMA_reg_buffer_1364 ( .C (clk), .D (new_AGEMA_signal_2349), .Q (new_AGEMA_signal_4795) ) ;
    buf_clk new_AGEMA_reg_buffer_1366 ( .C (clk), .D (new_AGEMA_signal_2350), .Q (new_AGEMA_signal_4797) ) ;
    buf_clk new_AGEMA_reg_buffer_1368 ( .C (clk), .D (new_AGEMA_signal_2351), .Q (new_AGEMA_signal_4799) ) ;
    buf_clk new_AGEMA_reg_buffer_1370 ( .C (clk), .D (SubCellInst_SboxInst_3_XX_2_), .Q (new_AGEMA_signal_4801) ) ;
    buf_clk new_AGEMA_reg_buffer_1372 ( .C (clk), .D (new_AGEMA_signal_1233), .Q (new_AGEMA_signal_4803) ) ;
    buf_clk new_AGEMA_reg_buffer_1374 ( .C (clk), .D (new_AGEMA_signal_1234), .Q (new_AGEMA_signal_4805) ) ;
    buf_clk new_AGEMA_reg_buffer_1376 ( .C (clk), .D (new_AGEMA_signal_1235), .Q (new_AGEMA_signal_4807) ) ;
    buf_clk new_AGEMA_reg_buffer_1378 ( .C (clk), .D (SubCellInst_SboxInst_3_XX_1_), .Q (new_AGEMA_signal_4809) ) ;
    buf_clk new_AGEMA_reg_buffer_1380 ( .C (clk), .D (new_AGEMA_signal_1227), .Q (new_AGEMA_signal_4811) ) ;
    buf_clk new_AGEMA_reg_buffer_1382 ( .C (clk), .D (new_AGEMA_signal_1228), .Q (new_AGEMA_signal_4813) ) ;
    buf_clk new_AGEMA_reg_buffer_1384 ( .C (clk), .D (new_AGEMA_signal_1229), .Q (new_AGEMA_signal_4815) ) ;
    buf_clk new_AGEMA_reg_buffer_1386 ( .C (clk), .D (SubCellInst_SboxInst_4_Q0), .Q (new_AGEMA_signal_4817) ) ;
    buf_clk new_AGEMA_reg_buffer_1388 ( .C (clk), .D (new_AGEMA_signal_2103), .Q (new_AGEMA_signal_4819) ) ;
    buf_clk new_AGEMA_reg_buffer_1390 ( .C (clk), .D (new_AGEMA_signal_2104), .Q (new_AGEMA_signal_4821) ) ;
    buf_clk new_AGEMA_reg_buffer_1392 ( .C (clk), .D (new_AGEMA_signal_2105), .Q (new_AGEMA_signal_4823) ) ;
    buf_clk new_AGEMA_reg_buffer_1394 ( .C (clk), .D (SubCellInst_SboxInst_4_L1), .Q (new_AGEMA_signal_4825) ) ;
    buf_clk new_AGEMA_reg_buffer_1396 ( .C (clk), .D (new_AGEMA_signal_2358), .Q (new_AGEMA_signal_4827) ) ;
    buf_clk new_AGEMA_reg_buffer_1398 ( .C (clk), .D (new_AGEMA_signal_2359), .Q (new_AGEMA_signal_4829) ) ;
    buf_clk new_AGEMA_reg_buffer_1400 ( .C (clk), .D (new_AGEMA_signal_2360), .Q (new_AGEMA_signal_4831) ) ;
    buf_clk new_AGEMA_reg_buffer_1402 ( .C (clk), .D (SubCellInst_SboxInst_4_XX_2_), .Q (new_AGEMA_signal_4833) ) ;
    buf_clk new_AGEMA_reg_buffer_1404 ( .C (clk), .D (new_AGEMA_signal_1251), .Q (new_AGEMA_signal_4835) ) ;
    buf_clk new_AGEMA_reg_buffer_1406 ( .C (clk), .D (new_AGEMA_signal_1252), .Q (new_AGEMA_signal_4837) ) ;
    buf_clk new_AGEMA_reg_buffer_1408 ( .C (clk), .D (new_AGEMA_signal_1253), .Q (new_AGEMA_signal_4839) ) ;
    buf_clk new_AGEMA_reg_buffer_1410 ( .C (clk), .D (SubCellInst_SboxInst_4_XX_1_), .Q (new_AGEMA_signal_4841) ) ;
    buf_clk new_AGEMA_reg_buffer_1412 ( .C (clk), .D (new_AGEMA_signal_1245), .Q (new_AGEMA_signal_4843) ) ;
    buf_clk new_AGEMA_reg_buffer_1414 ( .C (clk), .D (new_AGEMA_signal_1246), .Q (new_AGEMA_signal_4845) ) ;
    buf_clk new_AGEMA_reg_buffer_1416 ( .C (clk), .D (new_AGEMA_signal_1247), .Q (new_AGEMA_signal_4847) ) ;
    buf_clk new_AGEMA_reg_buffer_1418 ( .C (clk), .D (SubCellInst_SboxInst_5_Q0), .Q (new_AGEMA_signal_4849) ) ;
    buf_clk new_AGEMA_reg_buffer_1420 ( .C (clk), .D (new_AGEMA_signal_2121), .Q (new_AGEMA_signal_4851) ) ;
    buf_clk new_AGEMA_reg_buffer_1422 ( .C (clk), .D (new_AGEMA_signal_2122), .Q (new_AGEMA_signal_4853) ) ;
    buf_clk new_AGEMA_reg_buffer_1424 ( .C (clk), .D (new_AGEMA_signal_2123), .Q (new_AGEMA_signal_4855) ) ;
    buf_clk new_AGEMA_reg_buffer_1426 ( .C (clk), .D (SubCellInst_SboxInst_5_L1), .Q (new_AGEMA_signal_4857) ) ;
    buf_clk new_AGEMA_reg_buffer_1428 ( .C (clk), .D (new_AGEMA_signal_2367), .Q (new_AGEMA_signal_4859) ) ;
    buf_clk new_AGEMA_reg_buffer_1430 ( .C (clk), .D (new_AGEMA_signal_2368), .Q (new_AGEMA_signal_4861) ) ;
    buf_clk new_AGEMA_reg_buffer_1432 ( .C (clk), .D (new_AGEMA_signal_2369), .Q (new_AGEMA_signal_4863) ) ;
    buf_clk new_AGEMA_reg_buffer_1434 ( .C (clk), .D (SubCellInst_SboxInst_5_XX_2_), .Q (new_AGEMA_signal_4865) ) ;
    buf_clk new_AGEMA_reg_buffer_1436 ( .C (clk), .D (new_AGEMA_signal_1269), .Q (new_AGEMA_signal_4867) ) ;
    buf_clk new_AGEMA_reg_buffer_1438 ( .C (clk), .D (new_AGEMA_signal_1270), .Q (new_AGEMA_signal_4869) ) ;
    buf_clk new_AGEMA_reg_buffer_1440 ( .C (clk), .D (new_AGEMA_signal_1271), .Q (new_AGEMA_signal_4871) ) ;
    buf_clk new_AGEMA_reg_buffer_1442 ( .C (clk), .D (SubCellInst_SboxInst_5_XX_1_), .Q (new_AGEMA_signal_4873) ) ;
    buf_clk new_AGEMA_reg_buffer_1444 ( .C (clk), .D (new_AGEMA_signal_1263), .Q (new_AGEMA_signal_4875) ) ;
    buf_clk new_AGEMA_reg_buffer_1446 ( .C (clk), .D (new_AGEMA_signal_1264), .Q (new_AGEMA_signal_4877) ) ;
    buf_clk new_AGEMA_reg_buffer_1448 ( .C (clk), .D (new_AGEMA_signal_1265), .Q (new_AGEMA_signal_4879) ) ;
    buf_clk new_AGEMA_reg_buffer_1450 ( .C (clk), .D (SubCellInst_SboxInst_6_Q0), .Q (new_AGEMA_signal_4881) ) ;
    buf_clk new_AGEMA_reg_buffer_1452 ( .C (clk), .D (new_AGEMA_signal_2139), .Q (new_AGEMA_signal_4883) ) ;
    buf_clk new_AGEMA_reg_buffer_1454 ( .C (clk), .D (new_AGEMA_signal_2140), .Q (new_AGEMA_signal_4885) ) ;
    buf_clk new_AGEMA_reg_buffer_1456 ( .C (clk), .D (new_AGEMA_signal_2141), .Q (new_AGEMA_signal_4887) ) ;
    buf_clk new_AGEMA_reg_buffer_1458 ( .C (clk), .D (SubCellInst_SboxInst_6_L1), .Q (new_AGEMA_signal_4889) ) ;
    buf_clk new_AGEMA_reg_buffer_1460 ( .C (clk), .D (new_AGEMA_signal_2376), .Q (new_AGEMA_signal_4891) ) ;
    buf_clk new_AGEMA_reg_buffer_1462 ( .C (clk), .D (new_AGEMA_signal_2377), .Q (new_AGEMA_signal_4893) ) ;
    buf_clk new_AGEMA_reg_buffer_1464 ( .C (clk), .D (new_AGEMA_signal_2378), .Q (new_AGEMA_signal_4895) ) ;
    buf_clk new_AGEMA_reg_buffer_1466 ( .C (clk), .D (SubCellInst_SboxInst_6_XX_2_), .Q (new_AGEMA_signal_4897) ) ;
    buf_clk new_AGEMA_reg_buffer_1468 ( .C (clk), .D (new_AGEMA_signal_1287), .Q (new_AGEMA_signal_4899) ) ;
    buf_clk new_AGEMA_reg_buffer_1470 ( .C (clk), .D (new_AGEMA_signal_1288), .Q (new_AGEMA_signal_4901) ) ;
    buf_clk new_AGEMA_reg_buffer_1472 ( .C (clk), .D (new_AGEMA_signal_1289), .Q (new_AGEMA_signal_4903) ) ;
    buf_clk new_AGEMA_reg_buffer_1474 ( .C (clk), .D (SubCellInst_SboxInst_6_XX_1_), .Q (new_AGEMA_signal_4905) ) ;
    buf_clk new_AGEMA_reg_buffer_1476 ( .C (clk), .D (new_AGEMA_signal_1281), .Q (new_AGEMA_signal_4907) ) ;
    buf_clk new_AGEMA_reg_buffer_1478 ( .C (clk), .D (new_AGEMA_signal_1282), .Q (new_AGEMA_signal_4909) ) ;
    buf_clk new_AGEMA_reg_buffer_1480 ( .C (clk), .D (new_AGEMA_signal_1283), .Q (new_AGEMA_signal_4911) ) ;
    buf_clk new_AGEMA_reg_buffer_1482 ( .C (clk), .D (SubCellInst_SboxInst_7_Q0), .Q (new_AGEMA_signal_4913) ) ;
    buf_clk new_AGEMA_reg_buffer_1484 ( .C (clk), .D (new_AGEMA_signal_2157), .Q (new_AGEMA_signal_4915) ) ;
    buf_clk new_AGEMA_reg_buffer_1486 ( .C (clk), .D (new_AGEMA_signal_2158), .Q (new_AGEMA_signal_4917) ) ;
    buf_clk new_AGEMA_reg_buffer_1488 ( .C (clk), .D (new_AGEMA_signal_2159), .Q (new_AGEMA_signal_4919) ) ;
    buf_clk new_AGEMA_reg_buffer_1490 ( .C (clk), .D (SubCellInst_SboxInst_7_L1), .Q (new_AGEMA_signal_4921) ) ;
    buf_clk new_AGEMA_reg_buffer_1492 ( .C (clk), .D (new_AGEMA_signal_2385), .Q (new_AGEMA_signal_4923) ) ;
    buf_clk new_AGEMA_reg_buffer_1494 ( .C (clk), .D (new_AGEMA_signal_2386), .Q (new_AGEMA_signal_4925) ) ;
    buf_clk new_AGEMA_reg_buffer_1496 ( .C (clk), .D (new_AGEMA_signal_2387), .Q (new_AGEMA_signal_4927) ) ;
    buf_clk new_AGEMA_reg_buffer_1498 ( .C (clk), .D (SubCellInst_SboxInst_7_XX_2_), .Q (new_AGEMA_signal_4929) ) ;
    buf_clk new_AGEMA_reg_buffer_1500 ( .C (clk), .D (new_AGEMA_signal_1305), .Q (new_AGEMA_signal_4931) ) ;
    buf_clk new_AGEMA_reg_buffer_1502 ( .C (clk), .D (new_AGEMA_signal_1306), .Q (new_AGEMA_signal_4933) ) ;
    buf_clk new_AGEMA_reg_buffer_1504 ( .C (clk), .D (new_AGEMA_signal_1307), .Q (new_AGEMA_signal_4935) ) ;
    buf_clk new_AGEMA_reg_buffer_1506 ( .C (clk), .D (SubCellInst_SboxInst_7_XX_1_), .Q (new_AGEMA_signal_4937) ) ;
    buf_clk new_AGEMA_reg_buffer_1508 ( .C (clk), .D (new_AGEMA_signal_1299), .Q (new_AGEMA_signal_4939) ) ;
    buf_clk new_AGEMA_reg_buffer_1510 ( .C (clk), .D (new_AGEMA_signal_1300), .Q (new_AGEMA_signal_4941) ) ;
    buf_clk new_AGEMA_reg_buffer_1512 ( .C (clk), .D (new_AGEMA_signal_1301), .Q (new_AGEMA_signal_4943) ) ;
    buf_clk new_AGEMA_reg_buffer_1514 ( .C (clk), .D (SubCellInst_SboxInst_8_Q0), .Q (new_AGEMA_signal_4945) ) ;
    buf_clk new_AGEMA_reg_buffer_1516 ( .C (clk), .D (new_AGEMA_signal_2175), .Q (new_AGEMA_signal_4947) ) ;
    buf_clk new_AGEMA_reg_buffer_1518 ( .C (clk), .D (new_AGEMA_signal_2176), .Q (new_AGEMA_signal_4949) ) ;
    buf_clk new_AGEMA_reg_buffer_1520 ( .C (clk), .D (new_AGEMA_signal_2177), .Q (new_AGEMA_signal_4951) ) ;
    buf_clk new_AGEMA_reg_buffer_1522 ( .C (clk), .D (SubCellInst_SboxInst_8_L1), .Q (new_AGEMA_signal_4953) ) ;
    buf_clk new_AGEMA_reg_buffer_1524 ( .C (clk), .D (new_AGEMA_signal_2394), .Q (new_AGEMA_signal_4955) ) ;
    buf_clk new_AGEMA_reg_buffer_1526 ( .C (clk), .D (new_AGEMA_signal_2395), .Q (new_AGEMA_signal_4957) ) ;
    buf_clk new_AGEMA_reg_buffer_1528 ( .C (clk), .D (new_AGEMA_signal_2396), .Q (new_AGEMA_signal_4959) ) ;
    buf_clk new_AGEMA_reg_buffer_1530 ( .C (clk), .D (SubCellInst_SboxInst_8_XX_2_), .Q (new_AGEMA_signal_4961) ) ;
    buf_clk new_AGEMA_reg_buffer_1532 ( .C (clk), .D (new_AGEMA_signal_1323), .Q (new_AGEMA_signal_4963) ) ;
    buf_clk new_AGEMA_reg_buffer_1534 ( .C (clk), .D (new_AGEMA_signal_1324), .Q (new_AGEMA_signal_4965) ) ;
    buf_clk new_AGEMA_reg_buffer_1536 ( .C (clk), .D (new_AGEMA_signal_1325), .Q (new_AGEMA_signal_4967) ) ;
    buf_clk new_AGEMA_reg_buffer_1538 ( .C (clk), .D (SubCellInst_SboxInst_8_XX_1_), .Q (new_AGEMA_signal_4969) ) ;
    buf_clk new_AGEMA_reg_buffer_1540 ( .C (clk), .D (new_AGEMA_signal_1317), .Q (new_AGEMA_signal_4971) ) ;
    buf_clk new_AGEMA_reg_buffer_1542 ( .C (clk), .D (new_AGEMA_signal_1318), .Q (new_AGEMA_signal_4973) ) ;
    buf_clk new_AGEMA_reg_buffer_1544 ( .C (clk), .D (new_AGEMA_signal_1319), .Q (new_AGEMA_signal_4975) ) ;
    buf_clk new_AGEMA_reg_buffer_1546 ( .C (clk), .D (SubCellInst_SboxInst_9_Q0), .Q (new_AGEMA_signal_4977) ) ;
    buf_clk new_AGEMA_reg_buffer_1548 ( .C (clk), .D (new_AGEMA_signal_2193), .Q (new_AGEMA_signal_4979) ) ;
    buf_clk new_AGEMA_reg_buffer_1550 ( .C (clk), .D (new_AGEMA_signal_2194), .Q (new_AGEMA_signal_4981) ) ;
    buf_clk new_AGEMA_reg_buffer_1552 ( .C (clk), .D (new_AGEMA_signal_2195), .Q (new_AGEMA_signal_4983) ) ;
    buf_clk new_AGEMA_reg_buffer_1554 ( .C (clk), .D (SubCellInst_SboxInst_9_L1), .Q (new_AGEMA_signal_4985) ) ;
    buf_clk new_AGEMA_reg_buffer_1556 ( .C (clk), .D (new_AGEMA_signal_2403), .Q (new_AGEMA_signal_4987) ) ;
    buf_clk new_AGEMA_reg_buffer_1558 ( .C (clk), .D (new_AGEMA_signal_2404), .Q (new_AGEMA_signal_4989) ) ;
    buf_clk new_AGEMA_reg_buffer_1560 ( .C (clk), .D (new_AGEMA_signal_2405), .Q (new_AGEMA_signal_4991) ) ;
    buf_clk new_AGEMA_reg_buffer_1562 ( .C (clk), .D (SubCellInst_SboxInst_9_XX_2_), .Q (new_AGEMA_signal_4993) ) ;
    buf_clk new_AGEMA_reg_buffer_1564 ( .C (clk), .D (new_AGEMA_signal_1341), .Q (new_AGEMA_signal_4995) ) ;
    buf_clk new_AGEMA_reg_buffer_1566 ( .C (clk), .D (new_AGEMA_signal_1342), .Q (new_AGEMA_signal_4997) ) ;
    buf_clk new_AGEMA_reg_buffer_1568 ( .C (clk), .D (new_AGEMA_signal_1343), .Q (new_AGEMA_signal_4999) ) ;
    buf_clk new_AGEMA_reg_buffer_1570 ( .C (clk), .D (SubCellInst_SboxInst_9_XX_1_), .Q (new_AGEMA_signal_5001) ) ;
    buf_clk new_AGEMA_reg_buffer_1572 ( .C (clk), .D (new_AGEMA_signal_1335), .Q (new_AGEMA_signal_5003) ) ;
    buf_clk new_AGEMA_reg_buffer_1574 ( .C (clk), .D (new_AGEMA_signal_1336), .Q (new_AGEMA_signal_5005) ) ;
    buf_clk new_AGEMA_reg_buffer_1576 ( .C (clk), .D (new_AGEMA_signal_1337), .Q (new_AGEMA_signal_5007) ) ;
    buf_clk new_AGEMA_reg_buffer_1578 ( .C (clk), .D (SubCellInst_SboxInst_10_Q0), .Q (new_AGEMA_signal_5009) ) ;
    buf_clk new_AGEMA_reg_buffer_1580 ( .C (clk), .D (new_AGEMA_signal_2211), .Q (new_AGEMA_signal_5011) ) ;
    buf_clk new_AGEMA_reg_buffer_1582 ( .C (clk), .D (new_AGEMA_signal_2212), .Q (new_AGEMA_signal_5013) ) ;
    buf_clk new_AGEMA_reg_buffer_1584 ( .C (clk), .D (new_AGEMA_signal_2213), .Q (new_AGEMA_signal_5015) ) ;
    buf_clk new_AGEMA_reg_buffer_1586 ( .C (clk), .D (SubCellInst_SboxInst_10_L1), .Q (new_AGEMA_signal_5017) ) ;
    buf_clk new_AGEMA_reg_buffer_1588 ( .C (clk), .D (new_AGEMA_signal_2412), .Q (new_AGEMA_signal_5019) ) ;
    buf_clk new_AGEMA_reg_buffer_1590 ( .C (clk), .D (new_AGEMA_signal_2413), .Q (new_AGEMA_signal_5021) ) ;
    buf_clk new_AGEMA_reg_buffer_1592 ( .C (clk), .D (new_AGEMA_signal_2414), .Q (new_AGEMA_signal_5023) ) ;
    buf_clk new_AGEMA_reg_buffer_1594 ( .C (clk), .D (SubCellInst_SboxInst_10_XX_2_), .Q (new_AGEMA_signal_5025) ) ;
    buf_clk new_AGEMA_reg_buffer_1596 ( .C (clk), .D (new_AGEMA_signal_1359), .Q (new_AGEMA_signal_5027) ) ;
    buf_clk new_AGEMA_reg_buffer_1598 ( .C (clk), .D (new_AGEMA_signal_1360), .Q (new_AGEMA_signal_5029) ) ;
    buf_clk new_AGEMA_reg_buffer_1600 ( .C (clk), .D (new_AGEMA_signal_1361), .Q (new_AGEMA_signal_5031) ) ;
    buf_clk new_AGEMA_reg_buffer_1602 ( .C (clk), .D (SubCellInst_SboxInst_10_XX_1_), .Q (new_AGEMA_signal_5033) ) ;
    buf_clk new_AGEMA_reg_buffer_1604 ( .C (clk), .D (new_AGEMA_signal_1353), .Q (new_AGEMA_signal_5035) ) ;
    buf_clk new_AGEMA_reg_buffer_1606 ( .C (clk), .D (new_AGEMA_signal_1354), .Q (new_AGEMA_signal_5037) ) ;
    buf_clk new_AGEMA_reg_buffer_1608 ( .C (clk), .D (new_AGEMA_signal_1355), .Q (new_AGEMA_signal_5039) ) ;
    buf_clk new_AGEMA_reg_buffer_1610 ( .C (clk), .D (SubCellInst_SboxInst_11_Q0), .Q (new_AGEMA_signal_5041) ) ;
    buf_clk new_AGEMA_reg_buffer_1612 ( .C (clk), .D (new_AGEMA_signal_2229), .Q (new_AGEMA_signal_5043) ) ;
    buf_clk new_AGEMA_reg_buffer_1614 ( .C (clk), .D (new_AGEMA_signal_2230), .Q (new_AGEMA_signal_5045) ) ;
    buf_clk new_AGEMA_reg_buffer_1616 ( .C (clk), .D (new_AGEMA_signal_2231), .Q (new_AGEMA_signal_5047) ) ;
    buf_clk new_AGEMA_reg_buffer_1618 ( .C (clk), .D (SubCellInst_SboxInst_11_L1), .Q (new_AGEMA_signal_5049) ) ;
    buf_clk new_AGEMA_reg_buffer_1620 ( .C (clk), .D (new_AGEMA_signal_2421), .Q (new_AGEMA_signal_5051) ) ;
    buf_clk new_AGEMA_reg_buffer_1622 ( .C (clk), .D (new_AGEMA_signal_2422), .Q (new_AGEMA_signal_5053) ) ;
    buf_clk new_AGEMA_reg_buffer_1624 ( .C (clk), .D (new_AGEMA_signal_2423), .Q (new_AGEMA_signal_5055) ) ;
    buf_clk new_AGEMA_reg_buffer_1626 ( .C (clk), .D (SubCellInst_SboxInst_11_XX_2_), .Q (new_AGEMA_signal_5057) ) ;
    buf_clk new_AGEMA_reg_buffer_1628 ( .C (clk), .D (new_AGEMA_signal_1377), .Q (new_AGEMA_signal_5059) ) ;
    buf_clk new_AGEMA_reg_buffer_1630 ( .C (clk), .D (new_AGEMA_signal_1378), .Q (new_AGEMA_signal_5061) ) ;
    buf_clk new_AGEMA_reg_buffer_1632 ( .C (clk), .D (new_AGEMA_signal_1379), .Q (new_AGEMA_signal_5063) ) ;
    buf_clk new_AGEMA_reg_buffer_1634 ( .C (clk), .D (SubCellInst_SboxInst_11_XX_1_), .Q (new_AGEMA_signal_5065) ) ;
    buf_clk new_AGEMA_reg_buffer_1636 ( .C (clk), .D (new_AGEMA_signal_1371), .Q (new_AGEMA_signal_5067) ) ;
    buf_clk new_AGEMA_reg_buffer_1638 ( .C (clk), .D (new_AGEMA_signal_1372), .Q (new_AGEMA_signal_5069) ) ;
    buf_clk new_AGEMA_reg_buffer_1640 ( .C (clk), .D (new_AGEMA_signal_1373), .Q (new_AGEMA_signal_5071) ) ;
    buf_clk new_AGEMA_reg_buffer_1642 ( .C (clk), .D (SubCellInst_SboxInst_12_Q0), .Q (new_AGEMA_signal_5073) ) ;
    buf_clk new_AGEMA_reg_buffer_1644 ( .C (clk), .D (new_AGEMA_signal_2247), .Q (new_AGEMA_signal_5075) ) ;
    buf_clk new_AGEMA_reg_buffer_1646 ( .C (clk), .D (new_AGEMA_signal_2248), .Q (new_AGEMA_signal_5077) ) ;
    buf_clk new_AGEMA_reg_buffer_1648 ( .C (clk), .D (new_AGEMA_signal_2249), .Q (new_AGEMA_signal_5079) ) ;
    buf_clk new_AGEMA_reg_buffer_1650 ( .C (clk), .D (SubCellInst_SboxInst_12_L1), .Q (new_AGEMA_signal_5081) ) ;
    buf_clk new_AGEMA_reg_buffer_1652 ( .C (clk), .D (new_AGEMA_signal_2430), .Q (new_AGEMA_signal_5083) ) ;
    buf_clk new_AGEMA_reg_buffer_1654 ( .C (clk), .D (new_AGEMA_signal_2431), .Q (new_AGEMA_signal_5085) ) ;
    buf_clk new_AGEMA_reg_buffer_1656 ( .C (clk), .D (new_AGEMA_signal_2432), .Q (new_AGEMA_signal_5087) ) ;
    buf_clk new_AGEMA_reg_buffer_1658 ( .C (clk), .D (SubCellInst_SboxInst_12_XX_2_), .Q (new_AGEMA_signal_5089) ) ;
    buf_clk new_AGEMA_reg_buffer_1660 ( .C (clk), .D (new_AGEMA_signal_1395), .Q (new_AGEMA_signal_5091) ) ;
    buf_clk new_AGEMA_reg_buffer_1662 ( .C (clk), .D (new_AGEMA_signal_1396), .Q (new_AGEMA_signal_5093) ) ;
    buf_clk new_AGEMA_reg_buffer_1664 ( .C (clk), .D (new_AGEMA_signal_1397), .Q (new_AGEMA_signal_5095) ) ;
    buf_clk new_AGEMA_reg_buffer_1666 ( .C (clk), .D (SubCellInst_SboxInst_12_XX_1_), .Q (new_AGEMA_signal_5097) ) ;
    buf_clk new_AGEMA_reg_buffer_1668 ( .C (clk), .D (new_AGEMA_signal_1389), .Q (new_AGEMA_signal_5099) ) ;
    buf_clk new_AGEMA_reg_buffer_1670 ( .C (clk), .D (new_AGEMA_signal_1390), .Q (new_AGEMA_signal_5101) ) ;
    buf_clk new_AGEMA_reg_buffer_1672 ( .C (clk), .D (new_AGEMA_signal_1391), .Q (new_AGEMA_signal_5103) ) ;
    buf_clk new_AGEMA_reg_buffer_1674 ( .C (clk), .D (SubCellInst_SboxInst_13_Q0), .Q (new_AGEMA_signal_5105) ) ;
    buf_clk new_AGEMA_reg_buffer_1676 ( .C (clk), .D (new_AGEMA_signal_2265), .Q (new_AGEMA_signal_5107) ) ;
    buf_clk new_AGEMA_reg_buffer_1678 ( .C (clk), .D (new_AGEMA_signal_2266), .Q (new_AGEMA_signal_5109) ) ;
    buf_clk new_AGEMA_reg_buffer_1680 ( .C (clk), .D (new_AGEMA_signal_2267), .Q (new_AGEMA_signal_5111) ) ;
    buf_clk new_AGEMA_reg_buffer_1682 ( .C (clk), .D (SubCellInst_SboxInst_13_L1), .Q (new_AGEMA_signal_5113) ) ;
    buf_clk new_AGEMA_reg_buffer_1684 ( .C (clk), .D (new_AGEMA_signal_2439), .Q (new_AGEMA_signal_5115) ) ;
    buf_clk new_AGEMA_reg_buffer_1686 ( .C (clk), .D (new_AGEMA_signal_2440), .Q (new_AGEMA_signal_5117) ) ;
    buf_clk new_AGEMA_reg_buffer_1688 ( .C (clk), .D (new_AGEMA_signal_2441), .Q (new_AGEMA_signal_5119) ) ;
    buf_clk new_AGEMA_reg_buffer_1690 ( .C (clk), .D (SubCellInst_SboxInst_13_XX_2_), .Q (new_AGEMA_signal_5121) ) ;
    buf_clk new_AGEMA_reg_buffer_1692 ( .C (clk), .D (new_AGEMA_signal_1413), .Q (new_AGEMA_signal_5123) ) ;
    buf_clk new_AGEMA_reg_buffer_1694 ( .C (clk), .D (new_AGEMA_signal_1414), .Q (new_AGEMA_signal_5125) ) ;
    buf_clk new_AGEMA_reg_buffer_1696 ( .C (clk), .D (new_AGEMA_signal_1415), .Q (new_AGEMA_signal_5127) ) ;
    buf_clk new_AGEMA_reg_buffer_1698 ( .C (clk), .D (SubCellInst_SboxInst_13_XX_1_), .Q (new_AGEMA_signal_5129) ) ;
    buf_clk new_AGEMA_reg_buffer_1700 ( .C (clk), .D (new_AGEMA_signal_1407), .Q (new_AGEMA_signal_5131) ) ;
    buf_clk new_AGEMA_reg_buffer_1702 ( .C (clk), .D (new_AGEMA_signal_1408), .Q (new_AGEMA_signal_5133) ) ;
    buf_clk new_AGEMA_reg_buffer_1704 ( .C (clk), .D (new_AGEMA_signal_1409), .Q (new_AGEMA_signal_5135) ) ;
    buf_clk new_AGEMA_reg_buffer_1706 ( .C (clk), .D (SubCellInst_SboxInst_14_Q0), .Q (new_AGEMA_signal_5137) ) ;
    buf_clk new_AGEMA_reg_buffer_1708 ( .C (clk), .D (new_AGEMA_signal_2283), .Q (new_AGEMA_signal_5139) ) ;
    buf_clk new_AGEMA_reg_buffer_1710 ( .C (clk), .D (new_AGEMA_signal_2284), .Q (new_AGEMA_signal_5141) ) ;
    buf_clk new_AGEMA_reg_buffer_1712 ( .C (clk), .D (new_AGEMA_signal_2285), .Q (new_AGEMA_signal_5143) ) ;
    buf_clk new_AGEMA_reg_buffer_1714 ( .C (clk), .D (SubCellInst_SboxInst_14_L1), .Q (new_AGEMA_signal_5145) ) ;
    buf_clk new_AGEMA_reg_buffer_1716 ( .C (clk), .D (new_AGEMA_signal_2448), .Q (new_AGEMA_signal_5147) ) ;
    buf_clk new_AGEMA_reg_buffer_1718 ( .C (clk), .D (new_AGEMA_signal_2449), .Q (new_AGEMA_signal_5149) ) ;
    buf_clk new_AGEMA_reg_buffer_1720 ( .C (clk), .D (new_AGEMA_signal_2450), .Q (new_AGEMA_signal_5151) ) ;
    buf_clk new_AGEMA_reg_buffer_1722 ( .C (clk), .D (SubCellInst_SboxInst_14_XX_2_), .Q (new_AGEMA_signal_5153) ) ;
    buf_clk new_AGEMA_reg_buffer_1724 ( .C (clk), .D (new_AGEMA_signal_1431), .Q (new_AGEMA_signal_5155) ) ;
    buf_clk new_AGEMA_reg_buffer_1726 ( .C (clk), .D (new_AGEMA_signal_1432), .Q (new_AGEMA_signal_5157) ) ;
    buf_clk new_AGEMA_reg_buffer_1728 ( .C (clk), .D (new_AGEMA_signal_1433), .Q (new_AGEMA_signal_5159) ) ;
    buf_clk new_AGEMA_reg_buffer_1730 ( .C (clk), .D (SubCellInst_SboxInst_14_XX_1_), .Q (new_AGEMA_signal_5161) ) ;
    buf_clk new_AGEMA_reg_buffer_1732 ( .C (clk), .D (new_AGEMA_signal_1425), .Q (new_AGEMA_signal_5163) ) ;
    buf_clk new_AGEMA_reg_buffer_1734 ( .C (clk), .D (new_AGEMA_signal_1426), .Q (new_AGEMA_signal_5165) ) ;
    buf_clk new_AGEMA_reg_buffer_1736 ( .C (clk), .D (new_AGEMA_signal_1427), .Q (new_AGEMA_signal_5167) ) ;
    buf_clk new_AGEMA_reg_buffer_1738 ( .C (clk), .D (SubCellInst_SboxInst_15_Q0), .Q (new_AGEMA_signal_5169) ) ;
    buf_clk new_AGEMA_reg_buffer_1740 ( .C (clk), .D (new_AGEMA_signal_2301), .Q (new_AGEMA_signal_5171) ) ;
    buf_clk new_AGEMA_reg_buffer_1742 ( .C (clk), .D (new_AGEMA_signal_2302), .Q (new_AGEMA_signal_5173) ) ;
    buf_clk new_AGEMA_reg_buffer_1744 ( .C (clk), .D (new_AGEMA_signal_2303), .Q (new_AGEMA_signal_5175) ) ;
    buf_clk new_AGEMA_reg_buffer_1746 ( .C (clk), .D (SubCellInst_SboxInst_15_L1), .Q (new_AGEMA_signal_5177) ) ;
    buf_clk new_AGEMA_reg_buffer_1748 ( .C (clk), .D (new_AGEMA_signal_2457), .Q (new_AGEMA_signal_5179) ) ;
    buf_clk new_AGEMA_reg_buffer_1750 ( .C (clk), .D (new_AGEMA_signal_2458), .Q (new_AGEMA_signal_5181) ) ;
    buf_clk new_AGEMA_reg_buffer_1752 ( .C (clk), .D (new_AGEMA_signal_2459), .Q (new_AGEMA_signal_5183) ) ;
    buf_clk new_AGEMA_reg_buffer_1754 ( .C (clk), .D (SubCellInst_SboxInst_15_XX_2_), .Q (new_AGEMA_signal_5185) ) ;
    buf_clk new_AGEMA_reg_buffer_1756 ( .C (clk), .D (new_AGEMA_signal_1449), .Q (new_AGEMA_signal_5187) ) ;
    buf_clk new_AGEMA_reg_buffer_1758 ( .C (clk), .D (new_AGEMA_signal_1450), .Q (new_AGEMA_signal_5189) ) ;
    buf_clk new_AGEMA_reg_buffer_1760 ( .C (clk), .D (new_AGEMA_signal_1451), .Q (new_AGEMA_signal_5191) ) ;
    buf_clk new_AGEMA_reg_buffer_1762 ( .C (clk), .D (SubCellInst_SboxInst_15_XX_1_), .Q (new_AGEMA_signal_5193) ) ;
    buf_clk new_AGEMA_reg_buffer_1764 ( .C (clk), .D (new_AGEMA_signal_1443), .Q (new_AGEMA_signal_5195) ) ;
    buf_clk new_AGEMA_reg_buffer_1766 ( .C (clk), .D (new_AGEMA_signal_1444), .Q (new_AGEMA_signal_5197) ) ;
    buf_clk new_AGEMA_reg_buffer_1768 ( .C (clk), .D (new_AGEMA_signal_1445), .Q (new_AGEMA_signal_5199) ) ;
    buf_clk new_AGEMA_reg_buffer_1770 ( .C (clk), .D (FSMUpdate[3]), .Q (new_AGEMA_signal_5201) ) ;
    buf_clk new_AGEMA_reg_buffer_1772 ( .C (clk), .D (FSMUpdate[4]), .Q (new_AGEMA_signal_5203) ) ;
    buf_clk new_AGEMA_reg_buffer_1774 ( .C (clk), .D (TweakeyGeneration_key_Feedback[2]), .Q (new_AGEMA_signal_5205) ) ;
    buf_clk new_AGEMA_reg_buffer_1776 ( .C (clk), .D (new_AGEMA_signal_1470), .Q (new_AGEMA_signal_5207) ) ;
    buf_clk new_AGEMA_reg_buffer_1778 ( .C (clk), .D (new_AGEMA_signal_1471), .Q (new_AGEMA_signal_5209) ) ;
    buf_clk new_AGEMA_reg_buffer_1780 ( .C (clk), .D (new_AGEMA_signal_1472), .Q (new_AGEMA_signal_5211) ) ;
    buf_clk new_AGEMA_reg_buffer_1782 ( .C (clk), .D (TweakeyGeneration_key_Feedback[3]), .Q (new_AGEMA_signal_5213) ) ;
    buf_clk new_AGEMA_reg_buffer_1784 ( .C (clk), .D (new_AGEMA_signal_1479), .Q (new_AGEMA_signal_5215) ) ;
    buf_clk new_AGEMA_reg_buffer_1786 ( .C (clk), .D (new_AGEMA_signal_1480), .Q (new_AGEMA_signal_5217) ) ;
    buf_clk new_AGEMA_reg_buffer_1788 ( .C (clk), .D (new_AGEMA_signal_1481), .Q (new_AGEMA_signal_5219) ) ;
    buf_clk new_AGEMA_reg_buffer_1790 ( .C (clk), .D (TweakeyGeneration_key_Feedback[6]), .Q (new_AGEMA_signal_5221) ) ;
    buf_clk new_AGEMA_reg_buffer_1792 ( .C (clk), .D (new_AGEMA_signal_1506), .Q (new_AGEMA_signal_5223) ) ;
    buf_clk new_AGEMA_reg_buffer_1794 ( .C (clk), .D (new_AGEMA_signal_1507), .Q (new_AGEMA_signal_5225) ) ;
    buf_clk new_AGEMA_reg_buffer_1796 ( .C (clk), .D (new_AGEMA_signal_1508), .Q (new_AGEMA_signal_5227) ) ;
    buf_clk new_AGEMA_reg_buffer_1798 ( .C (clk), .D (TweakeyGeneration_key_Feedback[7]), .Q (new_AGEMA_signal_5229) ) ;
    buf_clk new_AGEMA_reg_buffer_1800 ( .C (clk), .D (new_AGEMA_signal_1515), .Q (new_AGEMA_signal_5231) ) ;
    buf_clk new_AGEMA_reg_buffer_1802 ( .C (clk), .D (new_AGEMA_signal_1516), .Q (new_AGEMA_signal_5233) ) ;
    buf_clk new_AGEMA_reg_buffer_1804 ( .C (clk), .D (new_AGEMA_signal_1517), .Q (new_AGEMA_signal_5235) ) ;
    buf_clk new_AGEMA_reg_buffer_1806 ( .C (clk), .D (TweakeyGeneration_key_Feedback[10]), .Q (new_AGEMA_signal_5237) ) ;
    buf_clk new_AGEMA_reg_buffer_1808 ( .C (clk), .D (new_AGEMA_signal_1542), .Q (new_AGEMA_signal_5239) ) ;
    buf_clk new_AGEMA_reg_buffer_1810 ( .C (clk), .D (new_AGEMA_signal_1543), .Q (new_AGEMA_signal_5241) ) ;
    buf_clk new_AGEMA_reg_buffer_1812 ( .C (clk), .D (new_AGEMA_signal_1544), .Q (new_AGEMA_signal_5243) ) ;
    buf_clk new_AGEMA_reg_buffer_1814 ( .C (clk), .D (TweakeyGeneration_key_Feedback[11]), .Q (new_AGEMA_signal_5245) ) ;
    buf_clk new_AGEMA_reg_buffer_1816 ( .C (clk), .D (new_AGEMA_signal_1551), .Q (new_AGEMA_signal_5247) ) ;
    buf_clk new_AGEMA_reg_buffer_1818 ( .C (clk), .D (new_AGEMA_signal_1552), .Q (new_AGEMA_signal_5249) ) ;
    buf_clk new_AGEMA_reg_buffer_1820 ( .C (clk), .D (new_AGEMA_signal_1553), .Q (new_AGEMA_signal_5251) ) ;
    buf_clk new_AGEMA_reg_buffer_1822 ( .C (clk), .D (TweakeyGeneration_key_Feedback[14]), .Q (new_AGEMA_signal_5253) ) ;
    buf_clk new_AGEMA_reg_buffer_1824 ( .C (clk), .D (new_AGEMA_signal_1578), .Q (new_AGEMA_signal_5255) ) ;
    buf_clk new_AGEMA_reg_buffer_1826 ( .C (clk), .D (new_AGEMA_signal_1579), .Q (new_AGEMA_signal_5257) ) ;
    buf_clk new_AGEMA_reg_buffer_1828 ( .C (clk), .D (new_AGEMA_signal_1580), .Q (new_AGEMA_signal_5259) ) ;
    buf_clk new_AGEMA_reg_buffer_1830 ( .C (clk), .D (TweakeyGeneration_key_Feedback[15]), .Q (new_AGEMA_signal_5261) ) ;
    buf_clk new_AGEMA_reg_buffer_1832 ( .C (clk), .D (new_AGEMA_signal_1587), .Q (new_AGEMA_signal_5263) ) ;
    buf_clk new_AGEMA_reg_buffer_1834 ( .C (clk), .D (new_AGEMA_signal_1588), .Q (new_AGEMA_signal_5265) ) ;
    buf_clk new_AGEMA_reg_buffer_1836 ( .C (clk), .D (new_AGEMA_signal_1589), .Q (new_AGEMA_signal_5267) ) ;
    buf_clk new_AGEMA_reg_buffer_1838 ( .C (clk), .D (TweakeyGeneration_key_Feedback[18]), .Q (new_AGEMA_signal_5269) ) ;
    buf_clk new_AGEMA_reg_buffer_1840 ( .C (clk), .D (new_AGEMA_signal_1614), .Q (new_AGEMA_signal_5271) ) ;
    buf_clk new_AGEMA_reg_buffer_1842 ( .C (clk), .D (new_AGEMA_signal_1615), .Q (new_AGEMA_signal_5273) ) ;
    buf_clk new_AGEMA_reg_buffer_1844 ( .C (clk), .D (new_AGEMA_signal_1616), .Q (new_AGEMA_signal_5275) ) ;
    buf_clk new_AGEMA_reg_buffer_1846 ( .C (clk), .D (TweakeyGeneration_key_Feedback[19]), .Q (new_AGEMA_signal_5277) ) ;
    buf_clk new_AGEMA_reg_buffer_1848 ( .C (clk), .D (new_AGEMA_signal_1623), .Q (new_AGEMA_signal_5279) ) ;
    buf_clk new_AGEMA_reg_buffer_1850 ( .C (clk), .D (new_AGEMA_signal_1624), .Q (new_AGEMA_signal_5281) ) ;
    buf_clk new_AGEMA_reg_buffer_1852 ( .C (clk), .D (new_AGEMA_signal_1625), .Q (new_AGEMA_signal_5283) ) ;
    buf_clk new_AGEMA_reg_buffer_1854 ( .C (clk), .D (TweakeyGeneration_key_Feedback[22]), .Q (new_AGEMA_signal_5285) ) ;
    buf_clk new_AGEMA_reg_buffer_1856 ( .C (clk), .D (new_AGEMA_signal_1650), .Q (new_AGEMA_signal_5287) ) ;
    buf_clk new_AGEMA_reg_buffer_1858 ( .C (clk), .D (new_AGEMA_signal_1651), .Q (new_AGEMA_signal_5289) ) ;
    buf_clk new_AGEMA_reg_buffer_1860 ( .C (clk), .D (new_AGEMA_signal_1652), .Q (new_AGEMA_signal_5291) ) ;
    buf_clk new_AGEMA_reg_buffer_1862 ( .C (clk), .D (TweakeyGeneration_key_Feedback[23]), .Q (new_AGEMA_signal_5293) ) ;
    buf_clk new_AGEMA_reg_buffer_1864 ( .C (clk), .D (new_AGEMA_signal_1659), .Q (new_AGEMA_signal_5295) ) ;
    buf_clk new_AGEMA_reg_buffer_1866 ( .C (clk), .D (new_AGEMA_signal_1660), .Q (new_AGEMA_signal_5297) ) ;
    buf_clk new_AGEMA_reg_buffer_1868 ( .C (clk), .D (new_AGEMA_signal_1661), .Q (new_AGEMA_signal_5299) ) ;
    buf_clk new_AGEMA_reg_buffer_1870 ( .C (clk), .D (TweakeyGeneration_key_Feedback[26]), .Q (new_AGEMA_signal_5301) ) ;
    buf_clk new_AGEMA_reg_buffer_1872 ( .C (clk), .D (new_AGEMA_signal_1686), .Q (new_AGEMA_signal_5303) ) ;
    buf_clk new_AGEMA_reg_buffer_1874 ( .C (clk), .D (new_AGEMA_signal_1687), .Q (new_AGEMA_signal_5305) ) ;
    buf_clk new_AGEMA_reg_buffer_1876 ( .C (clk), .D (new_AGEMA_signal_1688), .Q (new_AGEMA_signal_5307) ) ;
    buf_clk new_AGEMA_reg_buffer_1878 ( .C (clk), .D (TweakeyGeneration_key_Feedback[27]), .Q (new_AGEMA_signal_5309) ) ;
    buf_clk new_AGEMA_reg_buffer_1880 ( .C (clk), .D (new_AGEMA_signal_1695), .Q (new_AGEMA_signal_5311) ) ;
    buf_clk new_AGEMA_reg_buffer_1882 ( .C (clk), .D (new_AGEMA_signal_1696), .Q (new_AGEMA_signal_5313) ) ;
    buf_clk new_AGEMA_reg_buffer_1884 ( .C (clk), .D (new_AGEMA_signal_1697), .Q (new_AGEMA_signal_5315) ) ;
    buf_clk new_AGEMA_reg_buffer_1886 ( .C (clk), .D (TweakeyGeneration_key_Feedback[30]), .Q (new_AGEMA_signal_5317) ) ;
    buf_clk new_AGEMA_reg_buffer_1888 ( .C (clk), .D (new_AGEMA_signal_1722), .Q (new_AGEMA_signal_5319) ) ;
    buf_clk new_AGEMA_reg_buffer_1890 ( .C (clk), .D (new_AGEMA_signal_1723), .Q (new_AGEMA_signal_5321) ) ;
    buf_clk new_AGEMA_reg_buffer_1892 ( .C (clk), .D (new_AGEMA_signal_1724), .Q (new_AGEMA_signal_5323) ) ;
    buf_clk new_AGEMA_reg_buffer_1894 ( .C (clk), .D (TweakeyGeneration_key_Feedback[31]), .Q (new_AGEMA_signal_5325) ) ;
    buf_clk new_AGEMA_reg_buffer_1896 ( .C (clk), .D (new_AGEMA_signal_1731), .Q (new_AGEMA_signal_5327) ) ;
    buf_clk new_AGEMA_reg_buffer_1898 ( .C (clk), .D (new_AGEMA_signal_1732), .Q (new_AGEMA_signal_5329) ) ;
    buf_clk new_AGEMA_reg_buffer_1900 ( .C (clk), .D (new_AGEMA_signal_1733), .Q (new_AGEMA_signal_5331) ) ;
    buf_clk new_AGEMA_reg_buffer_1904 ( .C (clk), .D (Plaintext_s0[0]), .Q (new_AGEMA_signal_5335) ) ;
    buf_clk new_AGEMA_reg_buffer_1908 ( .C (clk), .D (Plaintext_s1[0]), .Q (new_AGEMA_signal_5339) ) ;
    buf_clk new_AGEMA_reg_buffer_1912 ( .C (clk), .D (Plaintext_s2[0]), .Q (new_AGEMA_signal_5343) ) ;
    buf_clk new_AGEMA_reg_buffer_1916 ( .C (clk), .D (Plaintext_s3[0]), .Q (new_AGEMA_signal_5347) ) ;
    buf_clk new_AGEMA_reg_buffer_1920 ( .C (clk), .D (Plaintext_s0[1]), .Q (new_AGEMA_signal_5351) ) ;
    buf_clk new_AGEMA_reg_buffer_1924 ( .C (clk), .D (Plaintext_s1[1]), .Q (new_AGEMA_signal_5355) ) ;
    buf_clk new_AGEMA_reg_buffer_1928 ( .C (clk), .D (Plaintext_s2[1]), .Q (new_AGEMA_signal_5359) ) ;
    buf_clk new_AGEMA_reg_buffer_1932 ( .C (clk), .D (Plaintext_s3[1]), .Q (new_AGEMA_signal_5363) ) ;
    buf_clk new_AGEMA_reg_buffer_1936 ( .C (clk), .D (Plaintext_s0[4]), .Q (new_AGEMA_signal_5367) ) ;
    buf_clk new_AGEMA_reg_buffer_1940 ( .C (clk), .D (Plaintext_s1[4]), .Q (new_AGEMA_signal_5371) ) ;
    buf_clk new_AGEMA_reg_buffer_1944 ( .C (clk), .D (Plaintext_s2[4]), .Q (new_AGEMA_signal_5375) ) ;
    buf_clk new_AGEMA_reg_buffer_1948 ( .C (clk), .D (Plaintext_s3[4]), .Q (new_AGEMA_signal_5379) ) ;
    buf_clk new_AGEMA_reg_buffer_1952 ( .C (clk), .D (Plaintext_s0[5]), .Q (new_AGEMA_signal_5383) ) ;
    buf_clk new_AGEMA_reg_buffer_1956 ( .C (clk), .D (Plaintext_s1[5]), .Q (new_AGEMA_signal_5387) ) ;
    buf_clk new_AGEMA_reg_buffer_1960 ( .C (clk), .D (Plaintext_s2[5]), .Q (new_AGEMA_signal_5391) ) ;
    buf_clk new_AGEMA_reg_buffer_1964 ( .C (clk), .D (Plaintext_s3[5]), .Q (new_AGEMA_signal_5395) ) ;
    buf_clk new_AGEMA_reg_buffer_1968 ( .C (clk), .D (Plaintext_s0[8]), .Q (new_AGEMA_signal_5399) ) ;
    buf_clk new_AGEMA_reg_buffer_1972 ( .C (clk), .D (Plaintext_s1[8]), .Q (new_AGEMA_signal_5403) ) ;
    buf_clk new_AGEMA_reg_buffer_1976 ( .C (clk), .D (Plaintext_s2[8]), .Q (new_AGEMA_signal_5407) ) ;
    buf_clk new_AGEMA_reg_buffer_1980 ( .C (clk), .D (Plaintext_s3[8]), .Q (new_AGEMA_signal_5411) ) ;
    buf_clk new_AGEMA_reg_buffer_1984 ( .C (clk), .D (Plaintext_s0[9]), .Q (new_AGEMA_signal_5415) ) ;
    buf_clk new_AGEMA_reg_buffer_1988 ( .C (clk), .D (Plaintext_s1[9]), .Q (new_AGEMA_signal_5419) ) ;
    buf_clk new_AGEMA_reg_buffer_1992 ( .C (clk), .D (Plaintext_s2[9]), .Q (new_AGEMA_signal_5423) ) ;
    buf_clk new_AGEMA_reg_buffer_1996 ( .C (clk), .D (Plaintext_s3[9]), .Q (new_AGEMA_signal_5427) ) ;
    buf_clk new_AGEMA_reg_buffer_2000 ( .C (clk), .D (Plaintext_s0[12]), .Q (new_AGEMA_signal_5431) ) ;
    buf_clk new_AGEMA_reg_buffer_2004 ( .C (clk), .D (Plaintext_s1[12]), .Q (new_AGEMA_signal_5435) ) ;
    buf_clk new_AGEMA_reg_buffer_2008 ( .C (clk), .D (Plaintext_s2[12]), .Q (new_AGEMA_signal_5439) ) ;
    buf_clk new_AGEMA_reg_buffer_2012 ( .C (clk), .D (Plaintext_s3[12]), .Q (new_AGEMA_signal_5443) ) ;
    buf_clk new_AGEMA_reg_buffer_2016 ( .C (clk), .D (Plaintext_s0[13]), .Q (new_AGEMA_signal_5447) ) ;
    buf_clk new_AGEMA_reg_buffer_2020 ( .C (clk), .D (Plaintext_s1[13]), .Q (new_AGEMA_signal_5451) ) ;
    buf_clk new_AGEMA_reg_buffer_2024 ( .C (clk), .D (Plaintext_s2[13]), .Q (new_AGEMA_signal_5455) ) ;
    buf_clk new_AGEMA_reg_buffer_2028 ( .C (clk), .D (Plaintext_s3[13]), .Q (new_AGEMA_signal_5459) ) ;
    buf_clk new_AGEMA_reg_buffer_2032 ( .C (clk), .D (Plaintext_s0[16]), .Q (new_AGEMA_signal_5463) ) ;
    buf_clk new_AGEMA_reg_buffer_2036 ( .C (clk), .D (Plaintext_s1[16]), .Q (new_AGEMA_signal_5467) ) ;
    buf_clk new_AGEMA_reg_buffer_2040 ( .C (clk), .D (Plaintext_s2[16]), .Q (new_AGEMA_signal_5471) ) ;
    buf_clk new_AGEMA_reg_buffer_2044 ( .C (clk), .D (Plaintext_s3[16]), .Q (new_AGEMA_signal_5475) ) ;
    buf_clk new_AGEMA_reg_buffer_2048 ( .C (clk), .D (Plaintext_s0[17]), .Q (new_AGEMA_signal_5479) ) ;
    buf_clk new_AGEMA_reg_buffer_2052 ( .C (clk), .D (Plaintext_s1[17]), .Q (new_AGEMA_signal_5483) ) ;
    buf_clk new_AGEMA_reg_buffer_2056 ( .C (clk), .D (Plaintext_s2[17]), .Q (new_AGEMA_signal_5487) ) ;
    buf_clk new_AGEMA_reg_buffer_2060 ( .C (clk), .D (Plaintext_s3[17]), .Q (new_AGEMA_signal_5491) ) ;
    buf_clk new_AGEMA_reg_buffer_2064 ( .C (clk), .D (Plaintext_s0[20]), .Q (new_AGEMA_signal_5495) ) ;
    buf_clk new_AGEMA_reg_buffer_2068 ( .C (clk), .D (Plaintext_s1[20]), .Q (new_AGEMA_signal_5499) ) ;
    buf_clk new_AGEMA_reg_buffer_2072 ( .C (clk), .D (Plaintext_s2[20]), .Q (new_AGEMA_signal_5503) ) ;
    buf_clk new_AGEMA_reg_buffer_2076 ( .C (clk), .D (Plaintext_s3[20]), .Q (new_AGEMA_signal_5507) ) ;
    buf_clk new_AGEMA_reg_buffer_2080 ( .C (clk), .D (Plaintext_s0[21]), .Q (new_AGEMA_signal_5511) ) ;
    buf_clk new_AGEMA_reg_buffer_2084 ( .C (clk), .D (Plaintext_s1[21]), .Q (new_AGEMA_signal_5515) ) ;
    buf_clk new_AGEMA_reg_buffer_2088 ( .C (clk), .D (Plaintext_s2[21]), .Q (new_AGEMA_signal_5519) ) ;
    buf_clk new_AGEMA_reg_buffer_2092 ( .C (clk), .D (Plaintext_s3[21]), .Q (new_AGEMA_signal_5523) ) ;
    buf_clk new_AGEMA_reg_buffer_2096 ( .C (clk), .D (Plaintext_s0[24]), .Q (new_AGEMA_signal_5527) ) ;
    buf_clk new_AGEMA_reg_buffer_2100 ( .C (clk), .D (Plaintext_s1[24]), .Q (new_AGEMA_signal_5531) ) ;
    buf_clk new_AGEMA_reg_buffer_2104 ( .C (clk), .D (Plaintext_s2[24]), .Q (new_AGEMA_signal_5535) ) ;
    buf_clk new_AGEMA_reg_buffer_2108 ( .C (clk), .D (Plaintext_s3[24]), .Q (new_AGEMA_signal_5539) ) ;
    buf_clk new_AGEMA_reg_buffer_2112 ( .C (clk), .D (Plaintext_s0[25]), .Q (new_AGEMA_signal_5543) ) ;
    buf_clk new_AGEMA_reg_buffer_2116 ( .C (clk), .D (Plaintext_s1[25]), .Q (new_AGEMA_signal_5547) ) ;
    buf_clk new_AGEMA_reg_buffer_2120 ( .C (clk), .D (Plaintext_s2[25]), .Q (new_AGEMA_signal_5551) ) ;
    buf_clk new_AGEMA_reg_buffer_2124 ( .C (clk), .D (Plaintext_s3[25]), .Q (new_AGEMA_signal_5555) ) ;
    buf_clk new_AGEMA_reg_buffer_2128 ( .C (clk), .D (Plaintext_s0[28]), .Q (new_AGEMA_signal_5559) ) ;
    buf_clk new_AGEMA_reg_buffer_2132 ( .C (clk), .D (Plaintext_s1[28]), .Q (new_AGEMA_signal_5563) ) ;
    buf_clk new_AGEMA_reg_buffer_2136 ( .C (clk), .D (Plaintext_s2[28]), .Q (new_AGEMA_signal_5567) ) ;
    buf_clk new_AGEMA_reg_buffer_2140 ( .C (clk), .D (Plaintext_s3[28]), .Q (new_AGEMA_signal_5571) ) ;
    buf_clk new_AGEMA_reg_buffer_2144 ( .C (clk), .D (Plaintext_s0[29]), .Q (new_AGEMA_signal_5575) ) ;
    buf_clk new_AGEMA_reg_buffer_2148 ( .C (clk), .D (Plaintext_s1[29]), .Q (new_AGEMA_signal_5579) ) ;
    buf_clk new_AGEMA_reg_buffer_2152 ( .C (clk), .D (Plaintext_s2[29]), .Q (new_AGEMA_signal_5583) ) ;
    buf_clk new_AGEMA_reg_buffer_2156 ( .C (clk), .D (Plaintext_s3[29]), .Q (new_AGEMA_signal_5587) ) ;
    buf_clk new_AGEMA_reg_buffer_2160 ( .C (clk), .D (Plaintext_s0[32]), .Q (new_AGEMA_signal_5591) ) ;
    buf_clk new_AGEMA_reg_buffer_2164 ( .C (clk), .D (Plaintext_s1[32]), .Q (new_AGEMA_signal_5595) ) ;
    buf_clk new_AGEMA_reg_buffer_2168 ( .C (clk), .D (Plaintext_s2[32]), .Q (new_AGEMA_signal_5599) ) ;
    buf_clk new_AGEMA_reg_buffer_2172 ( .C (clk), .D (Plaintext_s3[32]), .Q (new_AGEMA_signal_5603) ) ;
    buf_clk new_AGEMA_reg_buffer_2176 ( .C (clk), .D (Plaintext_s0[33]), .Q (new_AGEMA_signal_5607) ) ;
    buf_clk new_AGEMA_reg_buffer_2180 ( .C (clk), .D (Plaintext_s1[33]), .Q (new_AGEMA_signal_5611) ) ;
    buf_clk new_AGEMA_reg_buffer_2184 ( .C (clk), .D (Plaintext_s2[33]), .Q (new_AGEMA_signal_5615) ) ;
    buf_clk new_AGEMA_reg_buffer_2188 ( .C (clk), .D (Plaintext_s3[33]), .Q (new_AGEMA_signal_5619) ) ;
    buf_clk new_AGEMA_reg_buffer_2192 ( .C (clk), .D (Plaintext_s0[36]), .Q (new_AGEMA_signal_5623) ) ;
    buf_clk new_AGEMA_reg_buffer_2196 ( .C (clk), .D (Plaintext_s1[36]), .Q (new_AGEMA_signal_5627) ) ;
    buf_clk new_AGEMA_reg_buffer_2200 ( .C (clk), .D (Plaintext_s2[36]), .Q (new_AGEMA_signal_5631) ) ;
    buf_clk new_AGEMA_reg_buffer_2204 ( .C (clk), .D (Plaintext_s3[36]), .Q (new_AGEMA_signal_5635) ) ;
    buf_clk new_AGEMA_reg_buffer_2208 ( .C (clk), .D (Plaintext_s0[37]), .Q (new_AGEMA_signal_5639) ) ;
    buf_clk new_AGEMA_reg_buffer_2212 ( .C (clk), .D (Plaintext_s1[37]), .Q (new_AGEMA_signal_5643) ) ;
    buf_clk new_AGEMA_reg_buffer_2216 ( .C (clk), .D (Plaintext_s2[37]), .Q (new_AGEMA_signal_5647) ) ;
    buf_clk new_AGEMA_reg_buffer_2220 ( .C (clk), .D (Plaintext_s3[37]), .Q (new_AGEMA_signal_5651) ) ;
    buf_clk new_AGEMA_reg_buffer_2224 ( .C (clk), .D (Plaintext_s0[40]), .Q (new_AGEMA_signal_5655) ) ;
    buf_clk new_AGEMA_reg_buffer_2228 ( .C (clk), .D (Plaintext_s1[40]), .Q (new_AGEMA_signal_5659) ) ;
    buf_clk new_AGEMA_reg_buffer_2232 ( .C (clk), .D (Plaintext_s2[40]), .Q (new_AGEMA_signal_5663) ) ;
    buf_clk new_AGEMA_reg_buffer_2236 ( .C (clk), .D (Plaintext_s3[40]), .Q (new_AGEMA_signal_5667) ) ;
    buf_clk new_AGEMA_reg_buffer_2240 ( .C (clk), .D (Plaintext_s0[41]), .Q (new_AGEMA_signal_5671) ) ;
    buf_clk new_AGEMA_reg_buffer_2244 ( .C (clk), .D (Plaintext_s1[41]), .Q (new_AGEMA_signal_5675) ) ;
    buf_clk new_AGEMA_reg_buffer_2248 ( .C (clk), .D (Plaintext_s2[41]), .Q (new_AGEMA_signal_5679) ) ;
    buf_clk new_AGEMA_reg_buffer_2252 ( .C (clk), .D (Plaintext_s3[41]), .Q (new_AGEMA_signal_5683) ) ;
    buf_clk new_AGEMA_reg_buffer_2256 ( .C (clk), .D (Plaintext_s0[44]), .Q (new_AGEMA_signal_5687) ) ;
    buf_clk new_AGEMA_reg_buffer_2260 ( .C (clk), .D (Plaintext_s1[44]), .Q (new_AGEMA_signal_5691) ) ;
    buf_clk new_AGEMA_reg_buffer_2264 ( .C (clk), .D (Plaintext_s2[44]), .Q (new_AGEMA_signal_5695) ) ;
    buf_clk new_AGEMA_reg_buffer_2268 ( .C (clk), .D (Plaintext_s3[44]), .Q (new_AGEMA_signal_5699) ) ;
    buf_clk new_AGEMA_reg_buffer_2272 ( .C (clk), .D (Plaintext_s0[45]), .Q (new_AGEMA_signal_5703) ) ;
    buf_clk new_AGEMA_reg_buffer_2276 ( .C (clk), .D (Plaintext_s1[45]), .Q (new_AGEMA_signal_5707) ) ;
    buf_clk new_AGEMA_reg_buffer_2280 ( .C (clk), .D (Plaintext_s2[45]), .Q (new_AGEMA_signal_5711) ) ;
    buf_clk new_AGEMA_reg_buffer_2284 ( .C (clk), .D (Plaintext_s3[45]), .Q (new_AGEMA_signal_5715) ) ;
    buf_clk new_AGEMA_reg_buffer_2288 ( .C (clk), .D (Plaintext_s0[48]), .Q (new_AGEMA_signal_5719) ) ;
    buf_clk new_AGEMA_reg_buffer_2292 ( .C (clk), .D (Plaintext_s1[48]), .Q (new_AGEMA_signal_5723) ) ;
    buf_clk new_AGEMA_reg_buffer_2296 ( .C (clk), .D (Plaintext_s2[48]), .Q (new_AGEMA_signal_5727) ) ;
    buf_clk new_AGEMA_reg_buffer_2300 ( .C (clk), .D (Plaintext_s3[48]), .Q (new_AGEMA_signal_5731) ) ;
    buf_clk new_AGEMA_reg_buffer_2304 ( .C (clk), .D (Plaintext_s0[49]), .Q (new_AGEMA_signal_5735) ) ;
    buf_clk new_AGEMA_reg_buffer_2308 ( .C (clk), .D (Plaintext_s1[49]), .Q (new_AGEMA_signal_5739) ) ;
    buf_clk new_AGEMA_reg_buffer_2312 ( .C (clk), .D (Plaintext_s2[49]), .Q (new_AGEMA_signal_5743) ) ;
    buf_clk new_AGEMA_reg_buffer_2316 ( .C (clk), .D (Plaintext_s3[49]), .Q (new_AGEMA_signal_5747) ) ;
    buf_clk new_AGEMA_reg_buffer_2320 ( .C (clk), .D (Plaintext_s0[52]), .Q (new_AGEMA_signal_5751) ) ;
    buf_clk new_AGEMA_reg_buffer_2324 ( .C (clk), .D (Plaintext_s1[52]), .Q (new_AGEMA_signal_5755) ) ;
    buf_clk new_AGEMA_reg_buffer_2328 ( .C (clk), .D (Plaintext_s2[52]), .Q (new_AGEMA_signal_5759) ) ;
    buf_clk new_AGEMA_reg_buffer_2332 ( .C (clk), .D (Plaintext_s3[52]), .Q (new_AGEMA_signal_5763) ) ;
    buf_clk new_AGEMA_reg_buffer_2336 ( .C (clk), .D (Plaintext_s0[53]), .Q (new_AGEMA_signal_5767) ) ;
    buf_clk new_AGEMA_reg_buffer_2340 ( .C (clk), .D (Plaintext_s1[53]), .Q (new_AGEMA_signal_5771) ) ;
    buf_clk new_AGEMA_reg_buffer_2344 ( .C (clk), .D (Plaintext_s2[53]), .Q (new_AGEMA_signal_5775) ) ;
    buf_clk new_AGEMA_reg_buffer_2348 ( .C (clk), .D (Plaintext_s3[53]), .Q (new_AGEMA_signal_5779) ) ;
    buf_clk new_AGEMA_reg_buffer_2352 ( .C (clk), .D (Plaintext_s0[56]), .Q (new_AGEMA_signal_5783) ) ;
    buf_clk new_AGEMA_reg_buffer_2356 ( .C (clk), .D (Plaintext_s1[56]), .Q (new_AGEMA_signal_5787) ) ;
    buf_clk new_AGEMA_reg_buffer_2360 ( .C (clk), .D (Plaintext_s2[56]), .Q (new_AGEMA_signal_5791) ) ;
    buf_clk new_AGEMA_reg_buffer_2364 ( .C (clk), .D (Plaintext_s3[56]), .Q (new_AGEMA_signal_5795) ) ;
    buf_clk new_AGEMA_reg_buffer_2368 ( .C (clk), .D (Plaintext_s0[57]), .Q (new_AGEMA_signal_5799) ) ;
    buf_clk new_AGEMA_reg_buffer_2372 ( .C (clk), .D (Plaintext_s1[57]), .Q (new_AGEMA_signal_5803) ) ;
    buf_clk new_AGEMA_reg_buffer_2376 ( .C (clk), .D (Plaintext_s2[57]), .Q (new_AGEMA_signal_5807) ) ;
    buf_clk new_AGEMA_reg_buffer_2380 ( .C (clk), .D (Plaintext_s3[57]), .Q (new_AGEMA_signal_5811) ) ;
    buf_clk new_AGEMA_reg_buffer_2384 ( .C (clk), .D (Plaintext_s0[60]), .Q (new_AGEMA_signal_5815) ) ;
    buf_clk new_AGEMA_reg_buffer_2388 ( .C (clk), .D (Plaintext_s1[60]), .Q (new_AGEMA_signal_5819) ) ;
    buf_clk new_AGEMA_reg_buffer_2392 ( .C (clk), .D (Plaintext_s2[60]), .Q (new_AGEMA_signal_5823) ) ;
    buf_clk new_AGEMA_reg_buffer_2396 ( .C (clk), .D (Plaintext_s3[60]), .Q (new_AGEMA_signal_5827) ) ;
    buf_clk new_AGEMA_reg_buffer_2400 ( .C (clk), .D (Plaintext_s0[61]), .Q (new_AGEMA_signal_5831) ) ;
    buf_clk new_AGEMA_reg_buffer_2404 ( .C (clk), .D (Plaintext_s1[61]), .Q (new_AGEMA_signal_5835) ) ;
    buf_clk new_AGEMA_reg_buffer_2408 ( .C (clk), .D (Plaintext_s2[61]), .Q (new_AGEMA_signal_5839) ) ;
    buf_clk new_AGEMA_reg_buffer_2412 ( .C (clk), .D (Plaintext_s3[61]), .Q (new_AGEMA_signal_5843) ) ;
    buf_clk new_AGEMA_reg_buffer_2416 ( .C (clk), .D (Ciphertext_s0[1]), .Q (new_AGEMA_signal_5847) ) ;
    buf_clk new_AGEMA_reg_buffer_2418 ( .C (clk), .D (Ciphertext_s1[1]), .Q (new_AGEMA_signal_5849) ) ;
    buf_clk new_AGEMA_reg_buffer_2420 ( .C (clk), .D (Ciphertext_s2[1]), .Q (new_AGEMA_signal_5851) ) ;
    buf_clk new_AGEMA_reg_buffer_2422 ( .C (clk), .D (Ciphertext_s3[1]), .Q (new_AGEMA_signal_5853) ) ;
    buf_clk new_AGEMA_reg_buffer_2432 ( .C (clk), .D (SubCellInst_SboxInst_0_Q6), .Q (new_AGEMA_signal_5863) ) ;
    buf_clk new_AGEMA_reg_buffer_2434 ( .C (clk), .D (new_AGEMA_signal_2040), .Q (new_AGEMA_signal_5865) ) ;
    buf_clk new_AGEMA_reg_buffer_2436 ( .C (clk), .D (new_AGEMA_signal_2041), .Q (new_AGEMA_signal_5867) ) ;
    buf_clk new_AGEMA_reg_buffer_2438 ( .C (clk), .D (new_AGEMA_signal_2042), .Q (new_AGEMA_signal_5869) ) ;
    buf_clk new_AGEMA_reg_buffer_2440 ( .C (clk), .D (SubCellInst_SboxInst_0_L2), .Q (new_AGEMA_signal_5871) ) ;
    buf_clk new_AGEMA_reg_buffer_2444 ( .C (clk), .D (new_AGEMA_signal_2043), .Q (new_AGEMA_signal_5875) ) ;
    buf_clk new_AGEMA_reg_buffer_2448 ( .C (clk), .D (new_AGEMA_signal_2044), .Q (new_AGEMA_signal_5879) ) ;
    buf_clk new_AGEMA_reg_buffer_2452 ( .C (clk), .D (new_AGEMA_signal_2045), .Q (new_AGEMA_signal_5883) ) ;
    buf_clk new_AGEMA_reg_buffer_2464 ( .C (clk), .D (Ciphertext_s0[5]), .Q (new_AGEMA_signal_5895) ) ;
    buf_clk new_AGEMA_reg_buffer_2466 ( .C (clk), .D (Ciphertext_s1[5]), .Q (new_AGEMA_signal_5897) ) ;
    buf_clk new_AGEMA_reg_buffer_2468 ( .C (clk), .D (Ciphertext_s2[5]), .Q (new_AGEMA_signal_5899) ) ;
    buf_clk new_AGEMA_reg_buffer_2470 ( .C (clk), .D (Ciphertext_s3[5]), .Q (new_AGEMA_signal_5901) ) ;
    buf_clk new_AGEMA_reg_buffer_2480 ( .C (clk), .D (SubCellInst_SboxInst_1_Q6), .Q (new_AGEMA_signal_5911) ) ;
    buf_clk new_AGEMA_reg_buffer_2482 ( .C (clk), .D (new_AGEMA_signal_2058), .Q (new_AGEMA_signal_5913) ) ;
    buf_clk new_AGEMA_reg_buffer_2484 ( .C (clk), .D (new_AGEMA_signal_2059), .Q (new_AGEMA_signal_5915) ) ;
    buf_clk new_AGEMA_reg_buffer_2486 ( .C (clk), .D (new_AGEMA_signal_2060), .Q (new_AGEMA_signal_5917) ) ;
    buf_clk new_AGEMA_reg_buffer_2488 ( .C (clk), .D (SubCellInst_SboxInst_1_L2), .Q (new_AGEMA_signal_5919) ) ;
    buf_clk new_AGEMA_reg_buffer_2492 ( .C (clk), .D (new_AGEMA_signal_2061), .Q (new_AGEMA_signal_5923) ) ;
    buf_clk new_AGEMA_reg_buffer_2496 ( .C (clk), .D (new_AGEMA_signal_2062), .Q (new_AGEMA_signal_5927) ) ;
    buf_clk new_AGEMA_reg_buffer_2500 ( .C (clk), .D (new_AGEMA_signal_2063), .Q (new_AGEMA_signal_5931) ) ;
    buf_clk new_AGEMA_reg_buffer_2512 ( .C (clk), .D (Ciphertext_s0[9]), .Q (new_AGEMA_signal_5943) ) ;
    buf_clk new_AGEMA_reg_buffer_2514 ( .C (clk), .D (Ciphertext_s1[9]), .Q (new_AGEMA_signal_5945) ) ;
    buf_clk new_AGEMA_reg_buffer_2516 ( .C (clk), .D (Ciphertext_s2[9]), .Q (new_AGEMA_signal_5947) ) ;
    buf_clk new_AGEMA_reg_buffer_2518 ( .C (clk), .D (Ciphertext_s3[9]), .Q (new_AGEMA_signal_5949) ) ;
    buf_clk new_AGEMA_reg_buffer_2528 ( .C (clk), .D (SubCellInst_SboxInst_2_Q6), .Q (new_AGEMA_signal_5959) ) ;
    buf_clk new_AGEMA_reg_buffer_2530 ( .C (clk), .D (new_AGEMA_signal_2076), .Q (new_AGEMA_signal_5961) ) ;
    buf_clk new_AGEMA_reg_buffer_2532 ( .C (clk), .D (new_AGEMA_signal_2077), .Q (new_AGEMA_signal_5963) ) ;
    buf_clk new_AGEMA_reg_buffer_2534 ( .C (clk), .D (new_AGEMA_signal_2078), .Q (new_AGEMA_signal_5965) ) ;
    buf_clk new_AGEMA_reg_buffer_2536 ( .C (clk), .D (SubCellInst_SboxInst_2_L2), .Q (new_AGEMA_signal_5967) ) ;
    buf_clk new_AGEMA_reg_buffer_2540 ( .C (clk), .D (new_AGEMA_signal_2079), .Q (new_AGEMA_signal_5971) ) ;
    buf_clk new_AGEMA_reg_buffer_2544 ( .C (clk), .D (new_AGEMA_signal_2080), .Q (new_AGEMA_signal_5975) ) ;
    buf_clk new_AGEMA_reg_buffer_2548 ( .C (clk), .D (new_AGEMA_signal_2081), .Q (new_AGEMA_signal_5979) ) ;
    buf_clk new_AGEMA_reg_buffer_2560 ( .C (clk), .D (Ciphertext_s0[13]), .Q (new_AGEMA_signal_5991) ) ;
    buf_clk new_AGEMA_reg_buffer_2562 ( .C (clk), .D (Ciphertext_s1[13]), .Q (new_AGEMA_signal_5993) ) ;
    buf_clk new_AGEMA_reg_buffer_2564 ( .C (clk), .D (Ciphertext_s2[13]), .Q (new_AGEMA_signal_5995) ) ;
    buf_clk new_AGEMA_reg_buffer_2566 ( .C (clk), .D (Ciphertext_s3[13]), .Q (new_AGEMA_signal_5997) ) ;
    buf_clk new_AGEMA_reg_buffer_2576 ( .C (clk), .D (SubCellInst_SboxInst_3_Q6), .Q (new_AGEMA_signal_6007) ) ;
    buf_clk new_AGEMA_reg_buffer_2578 ( .C (clk), .D (new_AGEMA_signal_2094), .Q (new_AGEMA_signal_6009) ) ;
    buf_clk new_AGEMA_reg_buffer_2580 ( .C (clk), .D (new_AGEMA_signal_2095), .Q (new_AGEMA_signal_6011) ) ;
    buf_clk new_AGEMA_reg_buffer_2582 ( .C (clk), .D (new_AGEMA_signal_2096), .Q (new_AGEMA_signal_6013) ) ;
    buf_clk new_AGEMA_reg_buffer_2584 ( .C (clk), .D (SubCellInst_SboxInst_3_L2), .Q (new_AGEMA_signal_6015) ) ;
    buf_clk new_AGEMA_reg_buffer_2588 ( .C (clk), .D (new_AGEMA_signal_2097), .Q (new_AGEMA_signal_6019) ) ;
    buf_clk new_AGEMA_reg_buffer_2592 ( .C (clk), .D (new_AGEMA_signal_2098), .Q (new_AGEMA_signal_6023) ) ;
    buf_clk new_AGEMA_reg_buffer_2596 ( .C (clk), .D (new_AGEMA_signal_2099), .Q (new_AGEMA_signal_6027) ) ;
    buf_clk new_AGEMA_reg_buffer_2608 ( .C (clk), .D (Ciphertext_s0[17]), .Q (new_AGEMA_signal_6039) ) ;
    buf_clk new_AGEMA_reg_buffer_2610 ( .C (clk), .D (Ciphertext_s1[17]), .Q (new_AGEMA_signal_6041) ) ;
    buf_clk new_AGEMA_reg_buffer_2612 ( .C (clk), .D (Ciphertext_s2[17]), .Q (new_AGEMA_signal_6043) ) ;
    buf_clk new_AGEMA_reg_buffer_2614 ( .C (clk), .D (Ciphertext_s3[17]), .Q (new_AGEMA_signal_6045) ) ;
    buf_clk new_AGEMA_reg_buffer_2624 ( .C (clk), .D (SubCellInst_SboxInst_4_Q6), .Q (new_AGEMA_signal_6055) ) ;
    buf_clk new_AGEMA_reg_buffer_2626 ( .C (clk), .D (new_AGEMA_signal_2112), .Q (new_AGEMA_signal_6057) ) ;
    buf_clk new_AGEMA_reg_buffer_2628 ( .C (clk), .D (new_AGEMA_signal_2113), .Q (new_AGEMA_signal_6059) ) ;
    buf_clk new_AGEMA_reg_buffer_2630 ( .C (clk), .D (new_AGEMA_signal_2114), .Q (new_AGEMA_signal_6061) ) ;
    buf_clk new_AGEMA_reg_buffer_2632 ( .C (clk), .D (SubCellInst_SboxInst_4_L2), .Q (new_AGEMA_signal_6063) ) ;
    buf_clk new_AGEMA_reg_buffer_2636 ( .C (clk), .D (new_AGEMA_signal_2115), .Q (new_AGEMA_signal_6067) ) ;
    buf_clk new_AGEMA_reg_buffer_2640 ( .C (clk), .D (new_AGEMA_signal_2116), .Q (new_AGEMA_signal_6071) ) ;
    buf_clk new_AGEMA_reg_buffer_2644 ( .C (clk), .D (new_AGEMA_signal_2117), .Q (new_AGEMA_signal_6075) ) ;
    buf_clk new_AGEMA_reg_buffer_2656 ( .C (clk), .D (Ciphertext_s0[21]), .Q (new_AGEMA_signal_6087) ) ;
    buf_clk new_AGEMA_reg_buffer_2658 ( .C (clk), .D (Ciphertext_s1[21]), .Q (new_AGEMA_signal_6089) ) ;
    buf_clk new_AGEMA_reg_buffer_2660 ( .C (clk), .D (Ciphertext_s2[21]), .Q (new_AGEMA_signal_6091) ) ;
    buf_clk new_AGEMA_reg_buffer_2662 ( .C (clk), .D (Ciphertext_s3[21]), .Q (new_AGEMA_signal_6093) ) ;
    buf_clk new_AGEMA_reg_buffer_2672 ( .C (clk), .D (SubCellInst_SboxInst_5_Q6), .Q (new_AGEMA_signal_6103) ) ;
    buf_clk new_AGEMA_reg_buffer_2674 ( .C (clk), .D (new_AGEMA_signal_2130), .Q (new_AGEMA_signal_6105) ) ;
    buf_clk new_AGEMA_reg_buffer_2676 ( .C (clk), .D (new_AGEMA_signal_2131), .Q (new_AGEMA_signal_6107) ) ;
    buf_clk new_AGEMA_reg_buffer_2678 ( .C (clk), .D (new_AGEMA_signal_2132), .Q (new_AGEMA_signal_6109) ) ;
    buf_clk new_AGEMA_reg_buffer_2680 ( .C (clk), .D (SubCellInst_SboxInst_5_L2), .Q (new_AGEMA_signal_6111) ) ;
    buf_clk new_AGEMA_reg_buffer_2684 ( .C (clk), .D (new_AGEMA_signal_2133), .Q (new_AGEMA_signal_6115) ) ;
    buf_clk new_AGEMA_reg_buffer_2688 ( .C (clk), .D (new_AGEMA_signal_2134), .Q (new_AGEMA_signal_6119) ) ;
    buf_clk new_AGEMA_reg_buffer_2692 ( .C (clk), .D (new_AGEMA_signal_2135), .Q (new_AGEMA_signal_6123) ) ;
    buf_clk new_AGEMA_reg_buffer_2704 ( .C (clk), .D (Ciphertext_s0[25]), .Q (new_AGEMA_signal_6135) ) ;
    buf_clk new_AGEMA_reg_buffer_2706 ( .C (clk), .D (Ciphertext_s1[25]), .Q (new_AGEMA_signal_6137) ) ;
    buf_clk new_AGEMA_reg_buffer_2708 ( .C (clk), .D (Ciphertext_s2[25]), .Q (new_AGEMA_signal_6139) ) ;
    buf_clk new_AGEMA_reg_buffer_2710 ( .C (clk), .D (Ciphertext_s3[25]), .Q (new_AGEMA_signal_6141) ) ;
    buf_clk new_AGEMA_reg_buffer_2720 ( .C (clk), .D (SubCellInst_SboxInst_6_Q6), .Q (new_AGEMA_signal_6151) ) ;
    buf_clk new_AGEMA_reg_buffer_2722 ( .C (clk), .D (new_AGEMA_signal_2148), .Q (new_AGEMA_signal_6153) ) ;
    buf_clk new_AGEMA_reg_buffer_2724 ( .C (clk), .D (new_AGEMA_signal_2149), .Q (new_AGEMA_signal_6155) ) ;
    buf_clk new_AGEMA_reg_buffer_2726 ( .C (clk), .D (new_AGEMA_signal_2150), .Q (new_AGEMA_signal_6157) ) ;
    buf_clk new_AGEMA_reg_buffer_2728 ( .C (clk), .D (SubCellInst_SboxInst_6_L2), .Q (new_AGEMA_signal_6159) ) ;
    buf_clk new_AGEMA_reg_buffer_2732 ( .C (clk), .D (new_AGEMA_signal_2151), .Q (new_AGEMA_signal_6163) ) ;
    buf_clk new_AGEMA_reg_buffer_2736 ( .C (clk), .D (new_AGEMA_signal_2152), .Q (new_AGEMA_signal_6167) ) ;
    buf_clk new_AGEMA_reg_buffer_2740 ( .C (clk), .D (new_AGEMA_signal_2153), .Q (new_AGEMA_signal_6171) ) ;
    buf_clk new_AGEMA_reg_buffer_2752 ( .C (clk), .D (Ciphertext_s0[29]), .Q (new_AGEMA_signal_6183) ) ;
    buf_clk new_AGEMA_reg_buffer_2754 ( .C (clk), .D (Ciphertext_s1[29]), .Q (new_AGEMA_signal_6185) ) ;
    buf_clk new_AGEMA_reg_buffer_2756 ( .C (clk), .D (Ciphertext_s2[29]), .Q (new_AGEMA_signal_6187) ) ;
    buf_clk new_AGEMA_reg_buffer_2758 ( .C (clk), .D (Ciphertext_s3[29]), .Q (new_AGEMA_signal_6189) ) ;
    buf_clk new_AGEMA_reg_buffer_2768 ( .C (clk), .D (SubCellInst_SboxInst_7_Q6), .Q (new_AGEMA_signal_6199) ) ;
    buf_clk new_AGEMA_reg_buffer_2770 ( .C (clk), .D (new_AGEMA_signal_2166), .Q (new_AGEMA_signal_6201) ) ;
    buf_clk new_AGEMA_reg_buffer_2772 ( .C (clk), .D (new_AGEMA_signal_2167), .Q (new_AGEMA_signal_6203) ) ;
    buf_clk new_AGEMA_reg_buffer_2774 ( .C (clk), .D (new_AGEMA_signal_2168), .Q (new_AGEMA_signal_6205) ) ;
    buf_clk new_AGEMA_reg_buffer_2776 ( .C (clk), .D (SubCellInst_SboxInst_7_L2), .Q (new_AGEMA_signal_6207) ) ;
    buf_clk new_AGEMA_reg_buffer_2780 ( .C (clk), .D (new_AGEMA_signal_2169), .Q (new_AGEMA_signal_6211) ) ;
    buf_clk new_AGEMA_reg_buffer_2784 ( .C (clk), .D (new_AGEMA_signal_2170), .Q (new_AGEMA_signal_6215) ) ;
    buf_clk new_AGEMA_reg_buffer_2788 ( .C (clk), .D (new_AGEMA_signal_2171), .Q (new_AGEMA_signal_6219) ) ;
    buf_clk new_AGEMA_reg_buffer_2800 ( .C (clk), .D (Ciphertext_s0[33]), .Q (new_AGEMA_signal_6231) ) ;
    buf_clk new_AGEMA_reg_buffer_2802 ( .C (clk), .D (Ciphertext_s1[33]), .Q (new_AGEMA_signal_6233) ) ;
    buf_clk new_AGEMA_reg_buffer_2804 ( .C (clk), .D (Ciphertext_s2[33]), .Q (new_AGEMA_signal_6235) ) ;
    buf_clk new_AGEMA_reg_buffer_2806 ( .C (clk), .D (Ciphertext_s3[33]), .Q (new_AGEMA_signal_6237) ) ;
    buf_clk new_AGEMA_reg_buffer_2816 ( .C (clk), .D (SubCellInst_SboxInst_8_Q6), .Q (new_AGEMA_signal_6247) ) ;
    buf_clk new_AGEMA_reg_buffer_2818 ( .C (clk), .D (new_AGEMA_signal_2184), .Q (new_AGEMA_signal_6249) ) ;
    buf_clk new_AGEMA_reg_buffer_2820 ( .C (clk), .D (new_AGEMA_signal_2185), .Q (new_AGEMA_signal_6251) ) ;
    buf_clk new_AGEMA_reg_buffer_2822 ( .C (clk), .D (new_AGEMA_signal_2186), .Q (new_AGEMA_signal_6253) ) ;
    buf_clk new_AGEMA_reg_buffer_2824 ( .C (clk), .D (SubCellInst_SboxInst_8_L2), .Q (new_AGEMA_signal_6255) ) ;
    buf_clk new_AGEMA_reg_buffer_2828 ( .C (clk), .D (new_AGEMA_signal_2187), .Q (new_AGEMA_signal_6259) ) ;
    buf_clk new_AGEMA_reg_buffer_2832 ( .C (clk), .D (new_AGEMA_signal_2188), .Q (new_AGEMA_signal_6263) ) ;
    buf_clk new_AGEMA_reg_buffer_2836 ( .C (clk), .D (new_AGEMA_signal_2189), .Q (new_AGEMA_signal_6267) ) ;
    buf_clk new_AGEMA_reg_buffer_2848 ( .C (clk), .D (Ciphertext_s0[37]), .Q (new_AGEMA_signal_6279) ) ;
    buf_clk new_AGEMA_reg_buffer_2850 ( .C (clk), .D (Ciphertext_s1[37]), .Q (new_AGEMA_signal_6281) ) ;
    buf_clk new_AGEMA_reg_buffer_2852 ( .C (clk), .D (Ciphertext_s2[37]), .Q (new_AGEMA_signal_6283) ) ;
    buf_clk new_AGEMA_reg_buffer_2854 ( .C (clk), .D (Ciphertext_s3[37]), .Q (new_AGEMA_signal_6285) ) ;
    buf_clk new_AGEMA_reg_buffer_2864 ( .C (clk), .D (SubCellInst_SboxInst_9_Q6), .Q (new_AGEMA_signal_6295) ) ;
    buf_clk new_AGEMA_reg_buffer_2866 ( .C (clk), .D (new_AGEMA_signal_2202), .Q (new_AGEMA_signal_6297) ) ;
    buf_clk new_AGEMA_reg_buffer_2868 ( .C (clk), .D (new_AGEMA_signal_2203), .Q (new_AGEMA_signal_6299) ) ;
    buf_clk new_AGEMA_reg_buffer_2870 ( .C (clk), .D (new_AGEMA_signal_2204), .Q (new_AGEMA_signal_6301) ) ;
    buf_clk new_AGEMA_reg_buffer_2872 ( .C (clk), .D (SubCellInst_SboxInst_9_L2), .Q (new_AGEMA_signal_6303) ) ;
    buf_clk new_AGEMA_reg_buffer_2876 ( .C (clk), .D (new_AGEMA_signal_2205), .Q (new_AGEMA_signal_6307) ) ;
    buf_clk new_AGEMA_reg_buffer_2880 ( .C (clk), .D (new_AGEMA_signal_2206), .Q (new_AGEMA_signal_6311) ) ;
    buf_clk new_AGEMA_reg_buffer_2884 ( .C (clk), .D (new_AGEMA_signal_2207), .Q (new_AGEMA_signal_6315) ) ;
    buf_clk new_AGEMA_reg_buffer_2896 ( .C (clk), .D (Ciphertext_s0[41]), .Q (new_AGEMA_signal_6327) ) ;
    buf_clk new_AGEMA_reg_buffer_2898 ( .C (clk), .D (Ciphertext_s1[41]), .Q (new_AGEMA_signal_6329) ) ;
    buf_clk new_AGEMA_reg_buffer_2900 ( .C (clk), .D (Ciphertext_s2[41]), .Q (new_AGEMA_signal_6331) ) ;
    buf_clk new_AGEMA_reg_buffer_2902 ( .C (clk), .D (Ciphertext_s3[41]), .Q (new_AGEMA_signal_6333) ) ;
    buf_clk new_AGEMA_reg_buffer_2912 ( .C (clk), .D (SubCellInst_SboxInst_10_Q6), .Q (new_AGEMA_signal_6343) ) ;
    buf_clk new_AGEMA_reg_buffer_2914 ( .C (clk), .D (new_AGEMA_signal_2220), .Q (new_AGEMA_signal_6345) ) ;
    buf_clk new_AGEMA_reg_buffer_2916 ( .C (clk), .D (new_AGEMA_signal_2221), .Q (new_AGEMA_signal_6347) ) ;
    buf_clk new_AGEMA_reg_buffer_2918 ( .C (clk), .D (new_AGEMA_signal_2222), .Q (new_AGEMA_signal_6349) ) ;
    buf_clk new_AGEMA_reg_buffer_2920 ( .C (clk), .D (SubCellInst_SboxInst_10_L2), .Q (new_AGEMA_signal_6351) ) ;
    buf_clk new_AGEMA_reg_buffer_2924 ( .C (clk), .D (new_AGEMA_signal_2223), .Q (new_AGEMA_signal_6355) ) ;
    buf_clk new_AGEMA_reg_buffer_2928 ( .C (clk), .D (new_AGEMA_signal_2224), .Q (new_AGEMA_signal_6359) ) ;
    buf_clk new_AGEMA_reg_buffer_2932 ( .C (clk), .D (new_AGEMA_signal_2225), .Q (new_AGEMA_signal_6363) ) ;
    buf_clk new_AGEMA_reg_buffer_2944 ( .C (clk), .D (Ciphertext_s0[45]), .Q (new_AGEMA_signal_6375) ) ;
    buf_clk new_AGEMA_reg_buffer_2946 ( .C (clk), .D (Ciphertext_s1[45]), .Q (new_AGEMA_signal_6377) ) ;
    buf_clk new_AGEMA_reg_buffer_2948 ( .C (clk), .D (Ciphertext_s2[45]), .Q (new_AGEMA_signal_6379) ) ;
    buf_clk new_AGEMA_reg_buffer_2950 ( .C (clk), .D (Ciphertext_s3[45]), .Q (new_AGEMA_signal_6381) ) ;
    buf_clk new_AGEMA_reg_buffer_2960 ( .C (clk), .D (SubCellInst_SboxInst_11_Q6), .Q (new_AGEMA_signal_6391) ) ;
    buf_clk new_AGEMA_reg_buffer_2962 ( .C (clk), .D (new_AGEMA_signal_2238), .Q (new_AGEMA_signal_6393) ) ;
    buf_clk new_AGEMA_reg_buffer_2964 ( .C (clk), .D (new_AGEMA_signal_2239), .Q (new_AGEMA_signal_6395) ) ;
    buf_clk new_AGEMA_reg_buffer_2966 ( .C (clk), .D (new_AGEMA_signal_2240), .Q (new_AGEMA_signal_6397) ) ;
    buf_clk new_AGEMA_reg_buffer_2968 ( .C (clk), .D (SubCellInst_SboxInst_11_L2), .Q (new_AGEMA_signal_6399) ) ;
    buf_clk new_AGEMA_reg_buffer_2972 ( .C (clk), .D (new_AGEMA_signal_2241), .Q (new_AGEMA_signal_6403) ) ;
    buf_clk new_AGEMA_reg_buffer_2976 ( .C (clk), .D (new_AGEMA_signal_2242), .Q (new_AGEMA_signal_6407) ) ;
    buf_clk new_AGEMA_reg_buffer_2980 ( .C (clk), .D (new_AGEMA_signal_2243), .Q (new_AGEMA_signal_6411) ) ;
    buf_clk new_AGEMA_reg_buffer_2992 ( .C (clk), .D (Ciphertext_s0[49]), .Q (new_AGEMA_signal_6423) ) ;
    buf_clk new_AGEMA_reg_buffer_2994 ( .C (clk), .D (Ciphertext_s1[49]), .Q (new_AGEMA_signal_6425) ) ;
    buf_clk new_AGEMA_reg_buffer_2996 ( .C (clk), .D (Ciphertext_s2[49]), .Q (new_AGEMA_signal_6427) ) ;
    buf_clk new_AGEMA_reg_buffer_2998 ( .C (clk), .D (Ciphertext_s3[49]), .Q (new_AGEMA_signal_6429) ) ;
    buf_clk new_AGEMA_reg_buffer_3008 ( .C (clk), .D (SubCellInst_SboxInst_12_Q6), .Q (new_AGEMA_signal_6439) ) ;
    buf_clk new_AGEMA_reg_buffer_3010 ( .C (clk), .D (new_AGEMA_signal_2256), .Q (new_AGEMA_signal_6441) ) ;
    buf_clk new_AGEMA_reg_buffer_3012 ( .C (clk), .D (new_AGEMA_signal_2257), .Q (new_AGEMA_signal_6443) ) ;
    buf_clk new_AGEMA_reg_buffer_3014 ( .C (clk), .D (new_AGEMA_signal_2258), .Q (new_AGEMA_signal_6445) ) ;
    buf_clk new_AGEMA_reg_buffer_3016 ( .C (clk), .D (SubCellInst_SboxInst_12_L2), .Q (new_AGEMA_signal_6447) ) ;
    buf_clk new_AGEMA_reg_buffer_3020 ( .C (clk), .D (new_AGEMA_signal_2259), .Q (new_AGEMA_signal_6451) ) ;
    buf_clk new_AGEMA_reg_buffer_3024 ( .C (clk), .D (new_AGEMA_signal_2260), .Q (new_AGEMA_signal_6455) ) ;
    buf_clk new_AGEMA_reg_buffer_3028 ( .C (clk), .D (new_AGEMA_signal_2261), .Q (new_AGEMA_signal_6459) ) ;
    buf_clk new_AGEMA_reg_buffer_3040 ( .C (clk), .D (Ciphertext_s0[53]), .Q (new_AGEMA_signal_6471) ) ;
    buf_clk new_AGEMA_reg_buffer_3042 ( .C (clk), .D (Ciphertext_s1[53]), .Q (new_AGEMA_signal_6473) ) ;
    buf_clk new_AGEMA_reg_buffer_3044 ( .C (clk), .D (Ciphertext_s2[53]), .Q (new_AGEMA_signal_6475) ) ;
    buf_clk new_AGEMA_reg_buffer_3046 ( .C (clk), .D (Ciphertext_s3[53]), .Q (new_AGEMA_signal_6477) ) ;
    buf_clk new_AGEMA_reg_buffer_3056 ( .C (clk), .D (SubCellInst_SboxInst_13_Q6), .Q (new_AGEMA_signal_6487) ) ;
    buf_clk new_AGEMA_reg_buffer_3058 ( .C (clk), .D (new_AGEMA_signal_2274), .Q (new_AGEMA_signal_6489) ) ;
    buf_clk new_AGEMA_reg_buffer_3060 ( .C (clk), .D (new_AGEMA_signal_2275), .Q (new_AGEMA_signal_6491) ) ;
    buf_clk new_AGEMA_reg_buffer_3062 ( .C (clk), .D (new_AGEMA_signal_2276), .Q (new_AGEMA_signal_6493) ) ;
    buf_clk new_AGEMA_reg_buffer_3064 ( .C (clk), .D (SubCellInst_SboxInst_13_L2), .Q (new_AGEMA_signal_6495) ) ;
    buf_clk new_AGEMA_reg_buffer_3068 ( .C (clk), .D (new_AGEMA_signal_2277), .Q (new_AGEMA_signal_6499) ) ;
    buf_clk new_AGEMA_reg_buffer_3072 ( .C (clk), .D (new_AGEMA_signal_2278), .Q (new_AGEMA_signal_6503) ) ;
    buf_clk new_AGEMA_reg_buffer_3076 ( .C (clk), .D (new_AGEMA_signal_2279), .Q (new_AGEMA_signal_6507) ) ;
    buf_clk new_AGEMA_reg_buffer_3088 ( .C (clk), .D (Ciphertext_s0[57]), .Q (new_AGEMA_signal_6519) ) ;
    buf_clk new_AGEMA_reg_buffer_3090 ( .C (clk), .D (Ciphertext_s1[57]), .Q (new_AGEMA_signal_6521) ) ;
    buf_clk new_AGEMA_reg_buffer_3092 ( .C (clk), .D (Ciphertext_s2[57]), .Q (new_AGEMA_signal_6523) ) ;
    buf_clk new_AGEMA_reg_buffer_3094 ( .C (clk), .D (Ciphertext_s3[57]), .Q (new_AGEMA_signal_6525) ) ;
    buf_clk new_AGEMA_reg_buffer_3104 ( .C (clk), .D (SubCellInst_SboxInst_14_Q6), .Q (new_AGEMA_signal_6535) ) ;
    buf_clk new_AGEMA_reg_buffer_3106 ( .C (clk), .D (new_AGEMA_signal_2292), .Q (new_AGEMA_signal_6537) ) ;
    buf_clk new_AGEMA_reg_buffer_3108 ( .C (clk), .D (new_AGEMA_signal_2293), .Q (new_AGEMA_signal_6539) ) ;
    buf_clk new_AGEMA_reg_buffer_3110 ( .C (clk), .D (new_AGEMA_signal_2294), .Q (new_AGEMA_signal_6541) ) ;
    buf_clk new_AGEMA_reg_buffer_3112 ( .C (clk), .D (SubCellInst_SboxInst_14_L2), .Q (new_AGEMA_signal_6543) ) ;
    buf_clk new_AGEMA_reg_buffer_3116 ( .C (clk), .D (new_AGEMA_signal_2295), .Q (new_AGEMA_signal_6547) ) ;
    buf_clk new_AGEMA_reg_buffer_3120 ( .C (clk), .D (new_AGEMA_signal_2296), .Q (new_AGEMA_signal_6551) ) ;
    buf_clk new_AGEMA_reg_buffer_3124 ( .C (clk), .D (new_AGEMA_signal_2297), .Q (new_AGEMA_signal_6555) ) ;
    buf_clk new_AGEMA_reg_buffer_3136 ( .C (clk), .D (Ciphertext_s0[61]), .Q (new_AGEMA_signal_6567) ) ;
    buf_clk new_AGEMA_reg_buffer_3138 ( .C (clk), .D (Ciphertext_s1[61]), .Q (new_AGEMA_signal_6569) ) ;
    buf_clk new_AGEMA_reg_buffer_3140 ( .C (clk), .D (Ciphertext_s2[61]), .Q (new_AGEMA_signal_6571) ) ;
    buf_clk new_AGEMA_reg_buffer_3142 ( .C (clk), .D (Ciphertext_s3[61]), .Q (new_AGEMA_signal_6573) ) ;
    buf_clk new_AGEMA_reg_buffer_3152 ( .C (clk), .D (SubCellInst_SboxInst_15_Q6), .Q (new_AGEMA_signal_6583) ) ;
    buf_clk new_AGEMA_reg_buffer_3154 ( .C (clk), .D (new_AGEMA_signal_2310), .Q (new_AGEMA_signal_6585) ) ;
    buf_clk new_AGEMA_reg_buffer_3156 ( .C (clk), .D (new_AGEMA_signal_2311), .Q (new_AGEMA_signal_6587) ) ;
    buf_clk new_AGEMA_reg_buffer_3158 ( .C (clk), .D (new_AGEMA_signal_2312), .Q (new_AGEMA_signal_6589) ) ;
    buf_clk new_AGEMA_reg_buffer_3160 ( .C (clk), .D (SubCellInst_SboxInst_15_L2), .Q (new_AGEMA_signal_6591) ) ;
    buf_clk new_AGEMA_reg_buffer_3164 ( .C (clk), .D (new_AGEMA_signal_2313), .Q (new_AGEMA_signal_6595) ) ;
    buf_clk new_AGEMA_reg_buffer_3168 ( .C (clk), .D (new_AGEMA_signal_2314), .Q (new_AGEMA_signal_6599) ) ;
    buf_clk new_AGEMA_reg_buffer_3172 ( .C (clk), .D (new_AGEMA_signal_2315), .Q (new_AGEMA_signal_6603) ) ;
    buf_clk new_AGEMA_reg_buffer_3184 ( .C (clk), .D (FSMUpdate[1]), .Q (new_AGEMA_signal_6615) ) ;
    buf_clk new_AGEMA_reg_buffer_3188 ( .C (clk), .D (FSM[1]), .Q (new_AGEMA_signal_6619) ) ;
    buf_clk new_AGEMA_reg_buffer_3192 ( .C (clk), .D (FSM[4]), .Q (new_AGEMA_signal_6623) ) ;
    buf_clk new_AGEMA_reg_buffer_3196 ( .C (clk), .D (FSM[5]), .Q (new_AGEMA_signal_6627) ) ;
    buf_clk new_AGEMA_reg_buffer_3200 ( .C (clk), .D (TweakeyGeneration_key_Feedback[0]), .Q (new_AGEMA_signal_6631) ) ;
    buf_clk new_AGEMA_reg_buffer_3204 ( .C (clk), .D (new_AGEMA_signal_1452), .Q (new_AGEMA_signal_6635) ) ;
    buf_clk new_AGEMA_reg_buffer_3208 ( .C (clk), .D (new_AGEMA_signal_1453), .Q (new_AGEMA_signal_6639) ) ;
    buf_clk new_AGEMA_reg_buffer_3212 ( .C (clk), .D (new_AGEMA_signal_1454), .Q (new_AGEMA_signal_6643) ) ;
    buf_clk new_AGEMA_reg_buffer_3216 ( .C (clk), .D (TweakeyGeneration_key_Feedback[1]), .Q (new_AGEMA_signal_6647) ) ;
    buf_clk new_AGEMA_reg_buffer_3220 ( .C (clk), .D (new_AGEMA_signal_1461), .Q (new_AGEMA_signal_6651) ) ;
    buf_clk new_AGEMA_reg_buffer_3224 ( .C (clk), .D (new_AGEMA_signal_1462), .Q (new_AGEMA_signal_6655) ) ;
    buf_clk new_AGEMA_reg_buffer_3228 ( .C (clk), .D (new_AGEMA_signal_1463), .Q (new_AGEMA_signal_6659) ) ;
    buf_clk new_AGEMA_reg_buffer_3232 ( .C (clk), .D (TweakeyGeneration_key_Feedback[4]), .Q (new_AGEMA_signal_6663) ) ;
    buf_clk new_AGEMA_reg_buffer_3236 ( .C (clk), .D (new_AGEMA_signal_1488), .Q (new_AGEMA_signal_6667) ) ;
    buf_clk new_AGEMA_reg_buffer_3240 ( .C (clk), .D (new_AGEMA_signal_1489), .Q (new_AGEMA_signal_6671) ) ;
    buf_clk new_AGEMA_reg_buffer_3244 ( .C (clk), .D (new_AGEMA_signal_1490), .Q (new_AGEMA_signal_6675) ) ;
    buf_clk new_AGEMA_reg_buffer_3248 ( .C (clk), .D (TweakeyGeneration_key_Feedback[5]), .Q (new_AGEMA_signal_6679) ) ;
    buf_clk new_AGEMA_reg_buffer_3252 ( .C (clk), .D (new_AGEMA_signal_1497), .Q (new_AGEMA_signal_6683) ) ;
    buf_clk new_AGEMA_reg_buffer_3256 ( .C (clk), .D (new_AGEMA_signal_1498), .Q (new_AGEMA_signal_6687) ) ;
    buf_clk new_AGEMA_reg_buffer_3260 ( .C (clk), .D (new_AGEMA_signal_1499), .Q (new_AGEMA_signal_6691) ) ;
    buf_clk new_AGEMA_reg_buffer_3264 ( .C (clk), .D (TweakeyGeneration_key_Feedback[8]), .Q (new_AGEMA_signal_6695) ) ;
    buf_clk new_AGEMA_reg_buffer_3268 ( .C (clk), .D (new_AGEMA_signal_1524), .Q (new_AGEMA_signal_6699) ) ;
    buf_clk new_AGEMA_reg_buffer_3272 ( .C (clk), .D (new_AGEMA_signal_1525), .Q (new_AGEMA_signal_6703) ) ;
    buf_clk new_AGEMA_reg_buffer_3276 ( .C (clk), .D (new_AGEMA_signal_1526), .Q (new_AGEMA_signal_6707) ) ;
    buf_clk new_AGEMA_reg_buffer_3280 ( .C (clk), .D (TweakeyGeneration_key_Feedback[9]), .Q (new_AGEMA_signal_6711) ) ;
    buf_clk new_AGEMA_reg_buffer_3284 ( .C (clk), .D (new_AGEMA_signal_1533), .Q (new_AGEMA_signal_6715) ) ;
    buf_clk new_AGEMA_reg_buffer_3288 ( .C (clk), .D (new_AGEMA_signal_1534), .Q (new_AGEMA_signal_6719) ) ;
    buf_clk new_AGEMA_reg_buffer_3292 ( .C (clk), .D (new_AGEMA_signal_1535), .Q (new_AGEMA_signal_6723) ) ;
    buf_clk new_AGEMA_reg_buffer_3296 ( .C (clk), .D (TweakeyGeneration_key_Feedback[12]), .Q (new_AGEMA_signal_6727) ) ;
    buf_clk new_AGEMA_reg_buffer_3300 ( .C (clk), .D (new_AGEMA_signal_1560), .Q (new_AGEMA_signal_6731) ) ;
    buf_clk new_AGEMA_reg_buffer_3304 ( .C (clk), .D (new_AGEMA_signal_1561), .Q (new_AGEMA_signal_6735) ) ;
    buf_clk new_AGEMA_reg_buffer_3308 ( .C (clk), .D (new_AGEMA_signal_1562), .Q (new_AGEMA_signal_6739) ) ;
    buf_clk new_AGEMA_reg_buffer_3312 ( .C (clk), .D (TweakeyGeneration_key_Feedback[13]), .Q (new_AGEMA_signal_6743) ) ;
    buf_clk new_AGEMA_reg_buffer_3316 ( .C (clk), .D (new_AGEMA_signal_1569), .Q (new_AGEMA_signal_6747) ) ;
    buf_clk new_AGEMA_reg_buffer_3320 ( .C (clk), .D (new_AGEMA_signal_1570), .Q (new_AGEMA_signal_6751) ) ;
    buf_clk new_AGEMA_reg_buffer_3324 ( .C (clk), .D (new_AGEMA_signal_1571), .Q (new_AGEMA_signal_6755) ) ;
    buf_clk new_AGEMA_reg_buffer_3328 ( .C (clk), .D (TweakeyGeneration_key_Feedback[16]), .Q (new_AGEMA_signal_6759) ) ;
    buf_clk new_AGEMA_reg_buffer_3332 ( .C (clk), .D (new_AGEMA_signal_1596), .Q (new_AGEMA_signal_6763) ) ;
    buf_clk new_AGEMA_reg_buffer_3336 ( .C (clk), .D (new_AGEMA_signal_1597), .Q (new_AGEMA_signal_6767) ) ;
    buf_clk new_AGEMA_reg_buffer_3340 ( .C (clk), .D (new_AGEMA_signal_1598), .Q (new_AGEMA_signal_6771) ) ;
    buf_clk new_AGEMA_reg_buffer_3344 ( .C (clk), .D (TweakeyGeneration_key_Feedback[17]), .Q (new_AGEMA_signal_6775) ) ;
    buf_clk new_AGEMA_reg_buffer_3348 ( .C (clk), .D (new_AGEMA_signal_1605), .Q (new_AGEMA_signal_6779) ) ;
    buf_clk new_AGEMA_reg_buffer_3352 ( .C (clk), .D (new_AGEMA_signal_1606), .Q (new_AGEMA_signal_6783) ) ;
    buf_clk new_AGEMA_reg_buffer_3356 ( .C (clk), .D (new_AGEMA_signal_1607), .Q (new_AGEMA_signal_6787) ) ;
    buf_clk new_AGEMA_reg_buffer_3360 ( .C (clk), .D (TweakeyGeneration_key_Feedback[20]), .Q (new_AGEMA_signal_6791) ) ;
    buf_clk new_AGEMA_reg_buffer_3364 ( .C (clk), .D (new_AGEMA_signal_1632), .Q (new_AGEMA_signal_6795) ) ;
    buf_clk new_AGEMA_reg_buffer_3368 ( .C (clk), .D (new_AGEMA_signal_1633), .Q (new_AGEMA_signal_6799) ) ;
    buf_clk new_AGEMA_reg_buffer_3372 ( .C (clk), .D (new_AGEMA_signal_1634), .Q (new_AGEMA_signal_6803) ) ;
    buf_clk new_AGEMA_reg_buffer_3376 ( .C (clk), .D (TweakeyGeneration_key_Feedback[21]), .Q (new_AGEMA_signal_6807) ) ;
    buf_clk new_AGEMA_reg_buffer_3380 ( .C (clk), .D (new_AGEMA_signal_1641), .Q (new_AGEMA_signal_6811) ) ;
    buf_clk new_AGEMA_reg_buffer_3384 ( .C (clk), .D (new_AGEMA_signal_1642), .Q (new_AGEMA_signal_6815) ) ;
    buf_clk new_AGEMA_reg_buffer_3388 ( .C (clk), .D (new_AGEMA_signal_1643), .Q (new_AGEMA_signal_6819) ) ;
    buf_clk new_AGEMA_reg_buffer_3392 ( .C (clk), .D (TweakeyGeneration_key_Feedback[24]), .Q (new_AGEMA_signal_6823) ) ;
    buf_clk new_AGEMA_reg_buffer_3396 ( .C (clk), .D (new_AGEMA_signal_1668), .Q (new_AGEMA_signal_6827) ) ;
    buf_clk new_AGEMA_reg_buffer_3400 ( .C (clk), .D (new_AGEMA_signal_1669), .Q (new_AGEMA_signal_6831) ) ;
    buf_clk new_AGEMA_reg_buffer_3404 ( .C (clk), .D (new_AGEMA_signal_1670), .Q (new_AGEMA_signal_6835) ) ;
    buf_clk new_AGEMA_reg_buffer_3408 ( .C (clk), .D (TweakeyGeneration_key_Feedback[25]), .Q (new_AGEMA_signal_6839) ) ;
    buf_clk new_AGEMA_reg_buffer_3412 ( .C (clk), .D (new_AGEMA_signal_1677), .Q (new_AGEMA_signal_6843) ) ;
    buf_clk new_AGEMA_reg_buffer_3416 ( .C (clk), .D (new_AGEMA_signal_1678), .Q (new_AGEMA_signal_6847) ) ;
    buf_clk new_AGEMA_reg_buffer_3420 ( .C (clk), .D (new_AGEMA_signal_1679), .Q (new_AGEMA_signal_6851) ) ;
    buf_clk new_AGEMA_reg_buffer_3424 ( .C (clk), .D (TweakeyGeneration_key_Feedback[28]), .Q (new_AGEMA_signal_6855) ) ;
    buf_clk new_AGEMA_reg_buffer_3428 ( .C (clk), .D (new_AGEMA_signal_1704), .Q (new_AGEMA_signal_6859) ) ;
    buf_clk new_AGEMA_reg_buffer_3432 ( .C (clk), .D (new_AGEMA_signal_1705), .Q (new_AGEMA_signal_6863) ) ;
    buf_clk new_AGEMA_reg_buffer_3436 ( .C (clk), .D (new_AGEMA_signal_1706), .Q (new_AGEMA_signal_6867) ) ;
    buf_clk new_AGEMA_reg_buffer_3440 ( .C (clk), .D (TweakeyGeneration_key_Feedback[29]), .Q (new_AGEMA_signal_6871) ) ;
    buf_clk new_AGEMA_reg_buffer_3444 ( .C (clk), .D (new_AGEMA_signal_1713), .Q (new_AGEMA_signal_6875) ) ;
    buf_clk new_AGEMA_reg_buffer_3448 ( .C (clk), .D (new_AGEMA_signal_1714), .Q (new_AGEMA_signal_6879) ) ;
    buf_clk new_AGEMA_reg_buffer_3452 ( .C (clk), .D (new_AGEMA_signal_1715), .Q (new_AGEMA_signal_6883) ) ;
    buf_clk new_AGEMA_reg_buffer_3712 ( .C (clk), .D (TweakeyGeneration_StateRegInput[63]), .Q (new_AGEMA_signal_7143) ) ;
    buf_clk new_AGEMA_reg_buffer_3716 ( .C (clk), .D (new_AGEMA_signal_2025), .Q (new_AGEMA_signal_7147) ) ;
    buf_clk new_AGEMA_reg_buffer_3720 ( .C (clk), .D (new_AGEMA_signal_2026), .Q (new_AGEMA_signal_7151) ) ;
    buf_clk new_AGEMA_reg_buffer_3724 ( .C (clk), .D (new_AGEMA_signal_2027), .Q (new_AGEMA_signal_7155) ) ;
    buf_clk new_AGEMA_reg_buffer_3728 ( .C (clk), .D (TweakeyGeneration_StateRegInput[62]), .Q (new_AGEMA_signal_7159) ) ;
    buf_clk new_AGEMA_reg_buffer_3732 ( .C (clk), .D (new_AGEMA_signal_2016), .Q (new_AGEMA_signal_7163) ) ;
    buf_clk new_AGEMA_reg_buffer_3736 ( .C (clk), .D (new_AGEMA_signal_2017), .Q (new_AGEMA_signal_7167) ) ;
    buf_clk new_AGEMA_reg_buffer_3740 ( .C (clk), .D (new_AGEMA_signal_2018), .Q (new_AGEMA_signal_7171) ) ;
    buf_clk new_AGEMA_reg_buffer_3744 ( .C (clk), .D (TweakeyGeneration_StateRegInput[61]), .Q (new_AGEMA_signal_7175) ) ;
    buf_clk new_AGEMA_reg_buffer_3748 ( .C (clk), .D (new_AGEMA_signal_2007), .Q (new_AGEMA_signal_7179) ) ;
    buf_clk new_AGEMA_reg_buffer_3752 ( .C (clk), .D (new_AGEMA_signal_2008), .Q (new_AGEMA_signal_7183) ) ;
    buf_clk new_AGEMA_reg_buffer_3756 ( .C (clk), .D (new_AGEMA_signal_2009), .Q (new_AGEMA_signal_7187) ) ;
    buf_clk new_AGEMA_reg_buffer_3760 ( .C (clk), .D (TweakeyGeneration_StateRegInput[60]), .Q (new_AGEMA_signal_7191) ) ;
    buf_clk new_AGEMA_reg_buffer_3764 ( .C (clk), .D (new_AGEMA_signal_1998), .Q (new_AGEMA_signal_7195) ) ;
    buf_clk new_AGEMA_reg_buffer_3768 ( .C (clk), .D (new_AGEMA_signal_1999), .Q (new_AGEMA_signal_7199) ) ;
    buf_clk new_AGEMA_reg_buffer_3772 ( .C (clk), .D (new_AGEMA_signal_2000), .Q (new_AGEMA_signal_7203) ) ;
    buf_clk new_AGEMA_reg_buffer_3776 ( .C (clk), .D (TweakeyGeneration_StateRegInput[59]), .Q (new_AGEMA_signal_7207) ) ;
    buf_clk new_AGEMA_reg_buffer_3780 ( .C (clk), .D (new_AGEMA_signal_1989), .Q (new_AGEMA_signal_7211) ) ;
    buf_clk new_AGEMA_reg_buffer_3784 ( .C (clk), .D (new_AGEMA_signal_1990), .Q (new_AGEMA_signal_7215) ) ;
    buf_clk new_AGEMA_reg_buffer_3788 ( .C (clk), .D (new_AGEMA_signal_1991), .Q (new_AGEMA_signal_7219) ) ;
    buf_clk new_AGEMA_reg_buffer_3792 ( .C (clk), .D (TweakeyGeneration_StateRegInput[58]), .Q (new_AGEMA_signal_7223) ) ;
    buf_clk new_AGEMA_reg_buffer_3796 ( .C (clk), .D (new_AGEMA_signal_1980), .Q (new_AGEMA_signal_7227) ) ;
    buf_clk new_AGEMA_reg_buffer_3800 ( .C (clk), .D (new_AGEMA_signal_1981), .Q (new_AGEMA_signal_7231) ) ;
    buf_clk new_AGEMA_reg_buffer_3804 ( .C (clk), .D (new_AGEMA_signal_1982), .Q (new_AGEMA_signal_7235) ) ;
    buf_clk new_AGEMA_reg_buffer_3808 ( .C (clk), .D (TweakeyGeneration_StateRegInput[57]), .Q (new_AGEMA_signal_7239) ) ;
    buf_clk new_AGEMA_reg_buffer_3812 ( .C (clk), .D (new_AGEMA_signal_1971), .Q (new_AGEMA_signal_7243) ) ;
    buf_clk new_AGEMA_reg_buffer_3816 ( .C (clk), .D (new_AGEMA_signal_1972), .Q (new_AGEMA_signal_7247) ) ;
    buf_clk new_AGEMA_reg_buffer_3820 ( .C (clk), .D (new_AGEMA_signal_1973), .Q (new_AGEMA_signal_7251) ) ;
    buf_clk new_AGEMA_reg_buffer_3824 ( .C (clk), .D (TweakeyGeneration_StateRegInput[56]), .Q (new_AGEMA_signal_7255) ) ;
    buf_clk new_AGEMA_reg_buffer_3828 ( .C (clk), .D (new_AGEMA_signal_1962), .Q (new_AGEMA_signal_7259) ) ;
    buf_clk new_AGEMA_reg_buffer_3832 ( .C (clk), .D (new_AGEMA_signal_1963), .Q (new_AGEMA_signal_7263) ) ;
    buf_clk new_AGEMA_reg_buffer_3836 ( .C (clk), .D (new_AGEMA_signal_1964), .Q (new_AGEMA_signal_7267) ) ;
    buf_clk new_AGEMA_reg_buffer_3840 ( .C (clk), .D (TweakeyGeneration_StateRegInput[55]), .Q (new_AGEMA_signal_7271) ) ;
    buf_clk new_AGEMA_reg_buffer_3844 ( .C (clk), .D (new_AGEMA_signal_1953), .Q (new_AGEMA_signal_7275) ) ;
    buf_clk new_AGEMA_reg_buffer_3848 ( .C (clk), .D (new_AGEMA_signal_1954), .Q (new_AGEMA_signal_7279) ) ;
    buf_clk new_AGEMA_reg_buffer_3852 ( .C (clk), .D (new_AGEMA_signal_1955), .Q (new_AGEMA_signal_7283) ) ;
    buf_clk new_AGEMA_reg_buffer_3856 ( .C (clk), .D (TweakeyGeneration_StateRegInput[54]), .Q (new_AGEMA_signal_7287) ) ;
    buf_clk new_AGEMA_reg_buffer_3860 ( .C (clk), .D (new_AGEMA_signal_1944), .Q (new_AGEMA_signal_7291) ) ;
    buf_clk new_AGEMA_reg_buffer_3864 ( .C (clk), .D (new_AGEMA_signal_1945), .Q (new_AGEMA_signal_7295) ) ;
    buf_clk new_AGEMA_reg_buffer_3868 ( .C (clk), .D (new_AGEMA_signal_1946), .Q (new_AGEMA_signal_7299) ) ;
    buf_clk new_AGEMA_reg_buffer_3872 ( .C (clk), .D (TweakeyGeneration_StateRegInput[53]), .Q (new_AGEMA_signal_7303) ) ;
    buf_clk new_AGEMA_reg_buffer_3876 ( .C (clk), .D (new_AGEMA_signal_1935), .Q (new_AGEMA_signal_7307) ) ;
    buf_clk new_AGEMA_reg_buffer_3880 ( .C (clk), .D (new_AGEMA_signal_1936), .Q (new_AGEMA_signal_7311) ) ;
    buf_clk new_AGEMA_reg_buffer_3884 ( .C (clk), .D (new_AGEMA_signal_1937), .Q (new_AGEMA_signal_7315) ) ;
    buf_clk new_AGEMA_reg_buffer_3888 ( .C (clk), .D (TweakeyGeneration_StateRegInput[52]), .Q (new_AGEMA_signal_7319) ) ;
    buf_clk new_AGEMA_reg_buffer_3892 ( .C (clk), .D (new_AGEMA_signal_1926), .Q (new_AGEMA_signal_7323) ) ;
    buf_clk new_AGEMA_reg_buffer_3896 ( .C (clk), .D (new_AGEMA_signal_1927), .Q (new_AGEMA_signal_7327) ) ;
    buf_clk new_AGEMA_reg_buffer_3900 ( .C (clk), .D (new_AGEMA_signal_1928), .Q (new_AGEMA_signal_7331) ) ;
    buf_clk new_AGEMA_reg_buffer_3904 ( .C (clk), .D (TweakeyGeneration_StateRegInput[51]), .Q (new_AGEMA_signal_7335) ) ;
    buf_clk new_AGEMA_reg_buffer_3908 ( .C (clk), .D (new_AGEMA_signal_1917), .Q (new_AGEMA_signal_7339) ) ;
    buf_clk new_AGEMA_reg_buffer_3912 ( .C (clk), .D (new_AGEMA_signal_1918), .Q (new_AGEMA_signal_7343) ) ;
    buf_clk new_AGEMA_reg_buffer_3916 ( .C (clk), .D (new_AGEMA_signal_1919), .Q (new_AGEMA_signal_7347) ) ;
    buf_clk new_AGEMA_reg_buffer_3920 ( .C (clk), .D (TweakeyGeneration_StateRegInput[50]), .Q (new_AGEMA_signal_7351) ) ;
    buf_clk new_AGEMA_reg_buffer_3924 ( .C (clk), .D (new_AGEMA_signal_1908), .Q (new_AGEMA_signal_7355) ) ;
    buf_clk new_AGEMA_reg_buffer_3928 ( .C (clk), .D (new_AGEMA_signal_1909), .Q (new_AGEMA_signal_7359) ) ;
    buf_clk new_AGEMA_reg_buffer_3932 ( .C (clk), .D (new_AGEMA_signal_1910), .Q (new_AGEMA_signal_7363) ) ;
    buf_clk new_AGEMA_reg_buffer_3936 ( .C (clk), .D (TweakeyGeneration_StateRegInput[49]), .Q (new_AGEMA_signal_7367) ) ;
    buf_clk new_AGEMA_reg_buffer_3940 ( .C (clk), .D (new_AGEMA_signal_1899), .Q (new_AGEMA_signal_7371) ) ;
    buf_clk new_AGEMA_reg_buffer_3944 ( .C (clk), .D (new_AGEMA_signal_1900), .Q (new_AGEMA_signal_7375) ) ;
    buf_clk new_AGEMA_reg_buffer_3948 ( .C (clk), .D (new_AGEMA_signal_1901), .Q (new_AGEMA_signal_7379) ) ;
    buf_clk new_AGEMA_reg_buffer_3952 ( .C (clk), .D (TweakeyGeneration_StateRegInput[48]), .Q (new_AGEMA_signal_7383) ) ;
    buf_clk new_AGEMA_reg_buffer_3956 ( .C (clk), .D (new_AGEMA_signal_1890), .Q (new_AGEMA_signal_7387) ) ;
    buf_clk new_AGEMA_reg_buffer_3960 ( .C (clk), .D (new_AGEMA_signal_1891), .Q (new_AGEMA_signal_7391) ) ;
    buf_clk new_AGEMA_reg_buffer_3964 ( .C (clk), .D (new_AGEMA_signal_1892), .Q (new_AGEMA_signal_7395) ) ;
    buf_clk new_AGEMA_reg_buffer_3968 ( .C (clk), .D (TweakeyGeneration_StateRegInput[47]), .Q (new_AGEMA_signal_7399) ) ;
    buf_clk new_AGEMA_reg_buffer_3972 ( .C (clk), .D (new_AGEMA_signal_1881), .Q (new_AGEMA_signal_7403) ) ;
    buf_clk new_AGEMA_reg_buffer_3976 ( .C (clk), .D (new_AGEMA_signal_1882), .Q (new_AGEMA_signal_7407) ) ;
    buf_clk new_AGEMA_reg_buffer_3980 ( .C (clk), .D (new_AGEMA_signal_1883), .Q (new_AGEMA_signal_7411) ) ;
    buf_clk new_AGEMA_reg_buffer_3984 ( .C (clk), .D (TweakeyGeneration_StateRegInput[46]), .Q (new_AGEMA_signal_7415) ) ;
    buf_clk new_AGEMA_reg_buffer_3988 ( .C (clk), .D (new_AGEMA_signal_1872), .Q (new_AGEMA_signal_7419) ) ;
    buf_clk new_AGEMA_reg_buffer_3992 ( .C (clk), .D (new_AGEMA_signal_1873), .Q (new_AGEMA_signal_7423) ) ;
    buf_clk new_AGEMA_reg_buffer_3996 ( .C (clk), .D (new_AGEMA_signal_1874), .Q (new_AGEMA_signal_7427) ) ;
    buf_clk new_AGEMA_reg_buffer_4000 ( .C (clk), .D (TweakeyGeneration_StateRegInput[45]), .Q (new_AGEMA_signal_7431) ) ;
    buf_clk new_AGEMA_reg_buffer_4004 ( .C (clk), .D (new_AGEMA_signal_1863), .Q (new_AGEMA_signal_7435) ) ;
    buf_clk new_AGEMA_reg_buffer_4008 ( .C (clk), .D (new_AGEMA_signal_1864), .Q (new_AGEMA_signal_7439) ) ;
    buf_clk new_AGEMA_reg_buffer_4012 ( .C (clk), .D (new_AGEMA_signal_1865), .Q (new_AGEMA_signal_7443) ) ;
    buf_clk new_AGEMA_reg_buffer_4016 ( .C (clk), .D (TweakeyGeneration_StateRegInput[44]), .Q (new_AGEMA_signal_7447) ) ;
    buf_clk new_AGEMA_reg_buffer_4020 ( .C (clk), .D (new_AGEMA_signal_1854), .Q (new_AGEMA_signal_7451) ) ;
    buf_clk new_AGEMA_reg_buffer_4024 ( .C (clk), .D (new_AGEMA_signal_1855), .Q (new_AGEMA_signal_7455) ) ;
    buf_clk new_AGEMA_reg_buffer_4028 ( .C (clk), .D (new_AGEMA_signal_1856), .Q (new_AGEMA_signal_7459) ) ;
    buf_clk new_AGEMA_reg_buffer_4032 ( .C (clk), .D (TweakeyGeneration_StateRegInput[43]), .Q (new_AGEMA_signal_7463) ) ;
    buf_clk new_AGEMA_reg_buffer_4036 ( .C (clk), .D (new_AGEMA_signal_1845), .Q (new_AGEMA_signal_7467) ) ;
    buf_clk new_AGEMA_reg_buffer_4040 ( .C (clk), .D (new_AGEMA_signal_1846), .Q (new_AGEMA_signal_7471) ) ;
    buf_clk new_AGEMA_reg_buffer_4044 ( .C (clk), .D (new_AGEMA_signal_1847), .Q (new_AGEMA_signal_7475) ) ;
    buf_clk new_AGEMA_reg_buffer_4048 ( .C (clk), .D (TweakeyGeneration_StateRegInput[42]), .Q (new_AGEMA_signal_7479) ) ;
    buf_clk new_AGEMA_reg_buffer_4052 ( .C (clk), .D (new_AGEMA_signal_1836), .Q (new_AGEMA_signal_7483) ) ;
    buf_clk new_AGEMA_reg_buffer_4056 ( .C (clk), .D (new_AGEMA_signal_1837), .Q (new_AGEMA_signal_7487) ) ;
    buf_clk new_AGEMA_reg_buffer_4060 ( .C (clk), .D (new_AGEMA_signal_1838), .Q (new_AGEMA_signal_7491) ) ;
    buf_clk new_AGEMA_reg_buffer_4064 ( .C (clk), .D (TweakeyGeneration_StateRegInput[41]), .Q (new_AGEMA_signal_7495) ) ;
    buf_clk new_AGEMA_reg_buffer_4068 ( .C (clk), .D (new_AGEMA_signal_1827), .Q (new_AGEMA_signal_7499) ) ;
    buf_clk new_AGEMA_reg_buffer_4072 ( .C (clk), .D (new_AGEMA_signal_1828), .Q (new_AGEMA_signal_7503) ) ;
    buf_clk new_AGEMA_reg_buffer_4076 ( .C (clk), .D (new_AGEMA_signal_1829), .Q (new_AGEMA_signal_7507) ) ;
    buf_clk new_AGEMA_reg_buffer_4080 ( .C (clk), .D (TweakeyGeneration_StateRegInput[40]), .Q (new_AGEMA_signal_7511) ) ;
    buf_clk new_AGEMA_reg_buffer_4084 ( .C (clk), .D (new_AGEMA_signal_1818), .Q (new_AGEMA_signal_7515) ) ;
    buf_clk new_AGEMA_reg_buffer_4088 ( .C (clk), .D (new_AGEMA_signal_1819), .Q (new_AGEMA_signal_7519) ) ;
    buf_clk new_AGEMA_reg_buffer_4092 ( .C (clk), .D (new_AGEMA_signal_1820), .Q (new_AGEMA_signal_7523) ) ;
    buf_clk new_AGEMA_reg_buffer_4096 ( .C (clk), .D (TweakeyGeneration_StateRegInput[39]), .Q (new_AGEMA_signal_7527) ) ;
    buf_clk new_AGEMA_reg_buffer_4100 ( .C (clk), .D (new_AGEMA_signal_1809), .Q (new_AGEMA_signal_7531) ) ;
    buf_clk new_AGEMA_reg_buffer_4104 ( .C (clk), .D (new_AGEMA_signal_1810), .Q (new_AGEMA_signal_7535) ) ;
    buf_clk new_AGEMA_reg_buffer_4108 ( .C (clk), .D (new_AGEMA_signal_1811), .Q (new_AGEMA_signal_7539) ) ;
    buf_clk new_AGEMA_reg_buffer_4112 ( .C (clk), .D (TweakeyGeneration_StateRegInput[38]), .Q (new_AGEMA_signal_7543) ) ;
    buf_clk new_AGEMA_reg_buffer_4116 ( .C (clk), .D (new_AGEMA_signal_1800), .Q (new_AGEMA_signal_7547) ) ;
    buf_clk new_AGEMA_reg_buffer_4120 ( .C (clk), .D (new_AGEMA_signal_1801), .Q (new_AGEMA_signal_7551) ) ;
    buf_clk new_AGEMA_reg_buffer_4124 ( .C (clk), .D (new_AGEMA_signal_1802), .Q (new_AGEMA_signal_7555) ) ;
    buf_clk new_AGEMA_reg_buffer_4128 ( .C (clk), .D (TweakeyGeneration_StateRegInput[37]), .Q (new_AGEMA_signal_7559) ) ;
    buf_clk new_AGEMA_reg_buffer_4132 ( .C (clk), .D (new_AGEMA_signal_1791), .Q (new_AGEMA_signal_7563) ) ;
    buf_clk new_AGEMA_reg_buffer_4136 ( .C (clk), .D (new_AGEMA_signal_1792), .Q (new_AGEMA_signal_7567) ) ;
    buf_clk new_AGEMA_reg_buffer_4140 ( .C (clk), .D (new_AGEMA_signal_1793), .Q (new_AGEMA_signal_7571) ) ;
    buf_clk new_AGEMA_reg_buffer_4144 ( .C (clk), .D (TweakeyGeneration_StateRegInput[36]), .Q (new_AGEMA_signal_7575) ) ;
    buf_clk new_AGEMA_reg_buffer_4148 ( .C (clk), .D (new_AGEMA_signal_1782), .Q (new_AGEMA_signal_7579) ) ;
    buf_clk new_AGEMA_reg_buffer_4152 ( .C (clk), .D (new_AGEMA_signal_1783), .Q (new_AGEMA_signal_7583) ) ;
    buf_clk new_AGEMA_reg_buffer_4156 ( .C (clk), .D (new_AGEMA_signal_1784), .Q (new_AGEMA_signal_7587) ) ;
    buf_clk new_AGEMA_reg_buffer_4160 ( .C (clk), .D (TweakeyGeneration_StateRegInput[35]), .Q (new_AGEMA_signal_7591) ) ;
    buf_clk new_AGEMA_reg_buffer_4164 ( .C (clk), .D (new_AGEMA_signal_1773), .Q (new_AGEMA_signal_7595) ) ;
    buf_clk new_AGEMA_reg_buffer_4168 ( .C (clk), .D (new_AGEMA_signal_1774), .Q (new_AGEMA_signal_7599) ) ;
    buf_clk new_AGEMA_reg_buffer_4172 ( .C (clk), .D (new_AGEMA_signal_1775), .Q (new_AGEMA_signal_7603) ) ;
    buf_clk new_AGEMA_reg_buffer_4176 ( .C (clk), .D (TweakeyGeneration_StateRegInput[34]), .Q (new_AGEMA_signal_7607) ) ;
    buf_clk new_AGEMA_reg_buffer_4180 ( .C (clk), .D (new_AGEMA_signal_1764), .Q (new_AGEMA_signal_7611) ) ;
    buf_clk new_AGEMA_reg_buffer_4184 ( .C (clk), .D (new_AGEMA_signal_1765), .Q (new_AGEMA_signal_7615) ) ;
    buf_clk new_AGEMA_reg_buffer_4188 ( .C (clk), .D (new_AGEMA_signal_1766), .Q (new_AGEMA_signal_7619) ) ;
    buf_clk new_AGEMA_reg_buffer_4192 ( .C (clk), .D (TweakeyGeneration_StateRegInput[33]), .Q (new_AGEMA_signal_7623) ) ;
    buf_clk new_AGEMA_reg_buffer_4196 ( .C (clk), .D (new_AGEMA_signal_1755), .Q (new_AGEMA_signal_7627) ) ;
    buf_clk new_AGEMA_reg_buffer_4200 ( .C (clk), .D (new_AGEMA_signal_1756), .Q (new_AGEMA_signal_7631) ) ;
    buf_clk new_AGEMA_reg_buffer_4204 ( .C (clk), .D (new_AGEMA_signal_1757), .Q (new_AGEMA_signal_7635) ) ;
    buf_clk new_AGEMA_reg_buffer_4208 ( .C (clk), .D (TweakeyGeneration_StateRegInput[32]), .Q (new_AGEMA_signal_7639) ) ;
    buf_clk new_AGEMA_reg_buffer_4212 ( .C (clk), .D (new_AGEMA_signal_1746), .Q (new_AGEMA_signal_7643) ) ;
    buf_clk new_AGEMA_reg_buffer_4216 ( .C (clk), .D (new_AGEMA_signal_1747), .Q (new_AGEMA_signal_7647) ) ;
    buf_clk new_AGEMA_reg_buffer_4220 ( .C (clk), .D (new_AGEMA_signal_1748), .Q (new_AGEMA_signal_7651) ) ;
    buf_clk new_AGEMA_reg_buffer_4224 ( .C (clk), .D (TweakeyGeneration_StateRegInput[31]), .Q (new_AGEMA_signal_7655) ) ;
    buf_clk new_AGEMA_reg_buffer_4228 ( .C (clk), .D (new_AGEMA_signal_1737), .Q (new_AGEMA_signal_7659) ) ;
    buf_clk new_AGEMA_reg_buffer_4232 ( .C (clk), .D (new_AGEMA_signal_1738), .Q (new_AGEMA_signal_7663) ) ;
    buf_clk new_AGEMA_reg_buffer_4236 ( .C (clk), .D (new_AGEMA_signal_1739), .Q (new_AGEMA_signal_7667) ) ;
    buf_clk new_AGEMA_reg_buffer_4240 ( .C (clk), .D (TweakeyGeneration_StateRegInput[30]), .Q (new_AGEMA_signal_7671) ) ;
    buf_clk new_AGEMA_reg_buffer_4244 ( .C (clk), .D (new_AGEMA_signal_1728), .Q (new_AGEMA_signal_7675) ) ;
    buf_clk new_AGEMA_reg_buffer_4248 ( .C (clk), .D (new_AGEMA_signal_1729), .Q (new_AGEMA_signal_7679) ) ;
    buf_clk new_AGEMA_reg_buffer_4252 ( .C (clk), .D (new_AGEMA_signal_1730), .Q (new_AGEMA_signal_7683) ) ;
    buf_clk new_AGEMA_reg_buffer_4256 ( .C (clk), .D (TweakeyGeneration_StateRegInput[29]), .Q (new_AGEMA_signal_7687) ) ;
    buf_clk new_AGEMA_reg_buffer_4260 ( .C (clk), .D (new_AGEMA_signal_1719), .Q (new_AGEMA_signal_7691) ) ;
    buf_clk new_AGEMA_reg_buffer_4264 ( .C (clk), .D (new_AGEMA_signal_1720), .Q (new_AGEMA_signal_7695) ) ;
    buf_clk new_AGEMA_reg_buffer_4268 ( .C (clk), .D (new_AGEMA_signal_1721), .Q (new_AGEMA_signal_7699) ) ;
    buf_clk new_AGEMA_reg_buffer_4272 ( .C (clk), .D (TweakeyGeneration_StateRegInput[28]), .Q (new_AGEMA_signal_7703) ) ;
    buf_clk new_AGEMA_reg_buffer_4276 ( .C (clk), .D (new_AGEMA_signal_1710), .Q (new_AGEMA_signal_7707) ) ;
    buf_clk new_AGEMA_reg_buffer_4280 ( .C (clk), .D (new_AGEMA_signal_1711), .Q (new_AGEMA_signal_7711) ) ;
    buf_clk new_AGEMA_reg_buffer_4284 ( .C (clk), .D (new_AGEMA_signal_1712), .Q (new_AGEMA_signal_7715) ) ;
    buf_clk new_AGEMA_reg_buffer_4288 ( .C (clk), .D (TweakeyGeneration_StateRegInput[27]), .Q (new_AGEMA_signal_7719) ) ;
    buf_clk new_AGEMA_reg_buffer_4292 ( .C (clk), .D (new_AGEMA_signal_1701), .Q (new_AGEMA_signal_7723) ) ;
    buf_clk new_AGEMA_reg_buffer_4296 ( .C (clk), .D (new_AGEMA_signal_1702), .Q (new_AGEMA_signal_7727) ) ;
    buf_clk new_AGEMA_reg_buffer_4300 ( .C (clk), .D (new_AGEMA_signal_1703), .Q (new_AGEMA_signal_7731) ) ;
    buf_clk new_AGEMA_reg_buffer_4304 ( .C (clk), .D (TweakeyGeneration_StateRegInput[26]), .Q (new_AGEMA_signal_7735) ) ;
    buf_clk new_AGEMA_reg_buffer_4308 ( .C (clk), .D (new_AGEMA_signal_1692), .Q (new_AGEMA_signal_7739) ) ;
    buf_clk new_AGEMA_reg_buffer_4312 ( .C (clk), .D (new_AGEMA_signal_1693), .Q (new_AGEMA_signal_7743) ) ;
    buf_clk new_AGEMA_reg_buffer_4316 ( .C (clk), .D (new_AGEMA_signal_1694), .Q (new_AGEMA_signal_7747) ) ;
    buf_clk new_AGEMA_reg_buffer_4320 ( .C (clk), .D (TweakeyGeneration_StateRegInput[25]), .Q (new_AGEMA_signal_7751) ) ;
    buf_clk new_AGEMA_reg_buffer_4324 ( .C (clk), .D (new_AGEMA_signal_1683), .Q (new_AGEMA_signal_7755) ) ;
    buf_clk new_AGEMA_reg_buffer_4328 ( .C (clk), .D (new_AGEMA_signal_1684), .Q (new_AGEMA_signal_7759) ) ;
    buf_clk new_AGEMA_reg_buffer_4332 ( .C (clk), .D (new_AGEMA_signal_1685), .Q (new_AGEMA_signal_7763) ) ;
    buf_clk new_AGEMA_reg_buffer_4336 ( .C (clk), .D (TweakeyGeneration_StateRegInput[24]), .Q (new_AGEMA_signal_7767) ) ;
    buf_clk new_AGEMA_reg_buffer_4340 ( .C (clk), .D (new_AGEMA_signal_1674), .Q (new_AGEMA_signal_7771) ) ;
    buf_clk new_AGEMA_reg_buffer_4344 ( .C (clk), .D (new_AGEMA_signal_1675), .Q (new_AGEMA_signal_7775) ) ;
    buf_clk new_AGEMA_reg_buffer_4348 ( .C (clk), .D (new_AGEMA_signal_1676), .Q (new_AGEMA_signal_7779) ) ;
    buf_clk new_AGEMA_reg_buffer_4352 ( .C (clk), .D (TweakeyGeneration_StateRegInput[23]), .Q (new_AGEMA_signal_7783) ) ;
    buf_clk new_AGEMA_reg_buffer_4356 ( .C (clk), .D (new_AGEMA_signal_1665), .Q (new_AGEMA_signal_7787) ) ;
    buf_clk new_AGEMA_reg_buffer_4360 ( .C (clk), .D (new_AGEMA_signal_1666), .Q (new_AGEMA_signal_7791) ) ;
    buf_clk new_AGEMA_reg_buffer_4364 ( .C (clk), .D (new_AGEMA_signal_1667), .Q (new_AGEMA_signal_7795) ) ;
    buf_clk new_AGEMA_reg_buffer_4368 ( .C (clk), .D (TweakeyGeneration_StateRegInput[22]), .Q (new_AGEMA_signal_7799) ) ;
    buf_clk new_AGEMA_reg_buffer_4372 ( .C (clk), .D (new_AGEMA_signal_1656), .Q (new_AGEMA_signal_7803) ) ;
    buf_clk new_AGEMA_reg_buffer_4376 ( .C (clk), .D (new_AGEMA_signal_1657), .Q (new_AGEMA_signal_7807) ) ;
    buf_clk new_AGEMA_reg_buffer_4380 ( .C (clk), .D (new_AGEMA_signal_1658), .Q (new_AGEMA_signal_7811) ) ;
    buf_clk new_AGEMA_reg_buffer_4384 ( .C (clk), .D (TweakeyGeneration_StateRegInput[21]), .Q (new_AGEMA_signal_7815) ) ;
    buf_clk new_AGEMA_reg_buffer_4388 ( .C (clk), .D (new_AGEMA_signal_1647), .Q (new_AGEMA_signal_7819) ) ;
    buf_clk new_AGEMA_reg_buffer_4392 ( .C (clk), .D (new_AGEMA_signal_1648), .Q (new_AGEMA_signal_7823) ) ;
    buf_clk new_AGEMA_reg_buffer_4396 ( .C (clk), .D (new_AGEMA_signal_1649), .Q (new_AGEMA_signal_7827) ) ;
    buf_clk new_AGEMA_reg_buffer_4400 ( .C (clk), .D (TweakeyGeneration_StateRegInput[20]), .Q (new_AGEMA_signal_7831) ) ;
    buf_clk new_AGEMA_reg_buffer_4404 ( .C (clk), .D (new_AGEMA_signal_1638), .Q (new_AGEMA_signal_7835) ) ;
    buf_clk new_AGEMA_reg_buffer_4408 ( .C (clk), .D (new_AGEMA_signal_1639), .Q (new_AGEMA_signal_7839) ) ;
    buf_clk new_AGEMA_reg_buffer_4412 ( .C (clk), .D (new_AGEMA_signal_1640), .Q (new_AGEMA_signal_7843) ) ;
    buf_clk new_AGEMA_reg_buffer_4416 ( .C (clk), .D (TweakeyGeneration_StateRegInput[19]), .Q (new_AGEMA_signal_7847) ) ;
    buf_clk new_AGEMA_reg_buffer_4420 ( .C (clk), .D (new_AGEMA_signal_1629), .Q (new_AGEMA_signal_7851) ) ;
    buf_clk new_AGEMA_reg_buffer_4424 ( .C (clk), .D (new_AGEMA_signal_1630), .Q (new_AGEMA_signal_7855) ) ;
    buf_clk new_AGEMA_reg_buffer_4428 ( .C (clk), .D (new_AGEMA_signal_1631), .Q (new_AGEMA_signal_7859) ) ;
    buf_clk new_AGEMA_reg_buffer_4432 ( .C (clk), .D (TweakeyGeneration_StateRegInput[18]), .Q (new_AGEMA_signal_7863) ) ;
    buf_clk new_AGEMA_reg_buffer_4436 ( .C (clk), .D (new_AGEMA_signal_1620), .Q (new_AGEMA_signal_7867) ) ;
    buf_clk new_AGEMA_reg_buffer_4440 ( .C (clk), .D (new_AGEMA_signal_1621), .Q (new_AGEMA_signal_7871) ) ;
    buf_clk new_AGEMA_reg_buffer_4444 ( .C (clk), .D (new_AGEMA_signal_1622), .Q (new_AGEMA_signal_7875) ) ;
    buf_clk new_AGEMA_reg_buffer_4448 ( .C (clk), .D (TweakeyGeneration_StateRegInput[17]), .Q (new_AGEMA_signal_7879) ) ;
    buf_clk new_AGEMA_reg_buffer_4452 ( .C (clk), .D (new_AGEMA_signal_1611), .Q (new_AGEMA_signal_7883) ) ;
    buf_clk new_AGEMA_reg_buffer_4456 ( .C (clk), .D (new_AGEMA_signal_1612), .Q (new_AGEMA_signal_7887) ) ;
    buf_clk new_AGEMA_reg_buffer_4460 ( .C (clk), .D (new_AGEMA_signal_1613), .Q (new_AGEMA_signal_7891) ) ;
    buf_clk new_AGEMA_reg_buffer_4464 ( .C (clk), .D (TweakeyGeneration_StateRegInput[16]), .Q (new_AGEMA_signal_7895) ) ;
    buf_clk new_AGEMA_reg_buffer_4468 ( .C (clk), .D (new_AGEMA_signal_1602), .Q (new_AGEMA_signal_7899) ) ;
    buf_clk new_AGEMA_reg_buffer_4472 ( .C (clk), .D (new_AGEMA_signal_1603), .Q (new_AGEMA_signal_7903) ) ;
    buf_clk new_AGEMA_reg_buffer_4476 ( .C (clk), .D (new_AGEMA_signal_1604), .Q (new_AGEMA_signal_7907) ) ;
    buf_clk new_AGEMA_reg_buffer_4480 ( .C (clk), .D (TweakeyGeneration_StateRegInput[15]), .Q (new_AGEMA_signal_7911) ) ;
    buf_clk new_AGEMA_reg_buffer_4484 ( .C (clk), .D (new_AGEMA_signal_1593), .Q (new_AGEMA_signal_7915) ) ;
    buf_clk new_AGEMA_reg_buffer_4488 ( .C (clk), .D (new_AGEMA_signal_1594), .Q (new_AGEMA_signal_7919) ) ;
    buf_clk new_AGEMA_reg_buffer_4492 ( .C (clk), .D (new_AGEMA_signal_1595), .Q (new_AGEMA_signal_7923) ) ;
    buf_clk new_AGEMA_reg_buffer_4496 ( .C (clk), .D (TweakeyGeneration_StateRegInput[14]), .Q (new_AGEMA_signal_7927) ) ;
    buf_clk new_AGEMA_reg_buffer_4500 ( .C (clk), .D (new_AGEMA_signal_1584), .Q (new_AGEMA_signal_7931) ) ;
    buf_clk new_AGEMA_reg_buffer_4504 ( .C (clk), .D (new_AGEMA_signal_1585), .Q (new_AGEMA_signal_7935) ) ;
    buf_clk new_AGEMA_reg_buffer_4508 ( .C (clk), .D (new_AGEMA_signal_1586), .Q (new_AGEMA_signal_7939) ) ;
    buf_clk new_AGEMA_reg_buffer_4512 ( .C (clk), .D (TweakeyGeneration_StateRegInput[13]), .Q (new_AGEMA_signal_7943) ) ;
    buf_clk new_AGEMA_reg_buffer_4516 ( .C (clk), .D (new_AGEMA_signal_1575), .Q (new_AGEMA_signal_7947) ) ;
    buf_clk new_AGEMA_reg_buffer_4520 ( .C (clk), .D (new_AGEMA_signal_1576), .Q (new_AGEMA_signal_7951) ) ;
    buf_clk new_AGEMA_reg_buffer_4524 ( .C (clk), .D (new_AGEMA_signal_1577), .Q (new_AGEMA_signal_7955) ) ;
    buf_clk new_AGEMA_reg_buffer_4528 ( .C (clk), .D (TweakeyGeneration_StateRegInput[12]), .Q (new_AGEMA_signal_7959) ) ;
    buf_clk new_AGEMA_reg_buffer_4532 ( .C (clk), .D (new_AGEMA_signal_1566), .Q (new_AGEMA_signal_7963) ) ;
    buf_clk new_AGEMA_reg_buffer_4536 ( .C (clk), .D (new_AGEMA_signal_1567), .Q (new_AGEMA_signal_7967) ) ;
    buf_clk new_AGEMA_reg_buffer_4540 ( .C (clk), .D (new_AGEMA_signal_1568), .Q (new_AGEMA_signal_7971) ) ;
    buf_clk new_AGEMA_reg_buffer_4544 ( .C (clk), .D (TweakeyGeneration_StateRegInput[11]), .Q (new_AGEMA_signal_7975) ) ;
    buf_clk new_AGEMA_reg_buffer_4548 ( .C (clk), .D (new_AGEMA_signal_1557), .Q (new_AGEMA_signal_7979) ) ;
    buf_clk new_AGEMA_reg_buffer_4552 ( .C (clk), .D (new_AGEMA_signal_1558), .Q (new_AGEMA_signal_7983) ) ;
    buf_clk new_AGEMA_reg_buffer_4556 ( .C (clk), .D (new_AGEMA_signal_1559), .Q (new_AGEMA_signal_7987) ) ;
    buf_clk new_AGEMA_reg_buffer_4560 ( .C (clk), .D (TweakeyGeneration_StateRegInput[10]), .Q (new_AGEMA_signal_7991) ) ;
    buf_clk new_AGEMA_reg_buffer_4564 ( .C (clk), .D (new_AGEMA_signal_1548), .Q (new_AGEMA_signal_7995) ) ;
    buf_clk new_AGEMA_reg_buffer_4568 ( .C (clk), .D (new_AGEMA_signal_1549), .Q (new_AGEMA_signal_7999) ) ;
    buf_clk new_AGEMA_reg_buffer_4572 ( .C (clk), .D (new_AGEMA_signal_1550), .Q (new_AGEMA_signal_8003) ) ;
    buf_clk new_AGEMA_reg_buffer_4576 ( .C (clk), .D (TweakeyGeneration_StateRegInput[9]), .Q (new_AGEMA_signal_8007) ) ;
    buf_clk new_AGEMA_reg_buffer_4580 ( .C (clk), .D (new_AGEMA_signal_1539), .Q (new_AGEMA_signal_8011) ) ;
    buf_clk new_AGEMA_reg_buffer_4584 ( .C (clk), .D (new_AGEMA_signal_1540), .Q (new_AGEMA_signal_8015) ) ;
    buf_clk new_AGEMA_reg_buffer_4588 ( .C (clk), .D (new_AGEMA_signal_1541), .Q (new_AGEMA_signal_8019) ) ;
    buf_clk new_AGEMA_reg_buffer_4592 ( .C (clk), .D (TweakeyGeneration_StateRegInput[8]), .Q (new_AGEMA_signal_8023) ) ;
    buf_clk new_AGEMA_reg_buffer_4596 ( .C (clk), .D (new_AGEMA_signal_1530), .Q (new_AGEMA_signal_8027) ) ;
    buf_clk new_AGEMA_reg_buffer_4600 ( .C (clk), .D (new_AGEMA_signal_1531), .Q (new_AGEMA_signal_8031) ) ;
    buf_clk new_AGEMA_reg_buffer_4604 ( .C (clk), .D (new_AGEMA_signal_1532), .Q (new_AGEMA_signal_8035) ) ;
    buf_clk new_AGEMA_reg_buffer_4608 ( .C (clk), .D (TweakeyGeneration_StateRegInput[7]), .Q (new_AGEMA_signal_8039) ) ;
    buf_clk new_AGEMA_reg_buffer_4612 ( .C (clk), .D (new_AGEMA_signal_1521), .Q (new_AGEMA_signal_8043) ) ;
    buf_clk new_AGEMA_reg_buffer_4616 ( .C (clk), .D (new_AGEMA_signal_1522), .Q (new_AGEMA_signal_8047) ) ;
    buf_clk new_AGEMA_reg_buffer_4620 ( .C (clk), .D (new_AGEMA_signal_1523), .Q (new_AGEMA_signal_8051) ) ;
    buf_clk new_AGEMA_reg_buffer_4624 ( .C (clk), .D (TweakeyGeneration_StateRegInput[6]), .Q (new_AGEMA_signal_8055) ) ;
    buf_clk new_AGEMA_reg_buffer_4628 ( .C (clk), .D (new_AGEMA_signal_1512), .Q (new_AGEMA_signal_8059) ) ;
    buf_clk new_AGEMA_reg_buffer_4632 ( .C (clk), .D (new_AGEMA_signal_1513), .Q (new_AGEMA_signal_8063) ) ;
    buf_clk new_AGEMA_reg_buffer_4636 ( .C (clk), .D (new_AGEMA_signal_1514), .Q (new_AGEMA_signal_8067) ) ;
    buf_clk new_AGEMA_reg_buffer_4640 ( .C (clk), .D (TweakeyGeneration_StateRegInput[5]), .Q (new_AGEMA_signal_8071) ) ;
    buf_clk new_AGEMA_reg_buffer_4644 ( .C (clk), .D (new_AGEMA_signal_1503), .Q (new_AGEMA_signal_8075) ) ;
    buf_clk new_AGEMA_reg_buffer_4648 ( .C (clk), .D (new_AGEMA_signal_1504), .Q (new_AGEMA_signal_8079) ) ;
    buf_clk new_AGEMA_reg_buffer_4652 ( .C (clk), .D (new_AGEMA_signal_1505), .Q (new_AGEMA_signal_8083) ) ;
    buf_clk new_AGEMA_reg_buffer_4656 ( .C (clk), .D (TweakeyGeneration_StateRegInput[4]), .Q (new_AGEMA_signal_8087) ) ;
    buf_clk new_AGEMA_reg_buffer_4660 ( .C (clk), .D (new_AGEMA_signal_1494), .Q (new_AGEMA_signal_8091) ) ;
    buf_clk new_AGEMA_reg_buffer_4664 ( .C (clk), .D (new_AGEMA_signal_1495), .Q (new_AGEMA_signal_8095) ) ;
    buf_clk new_AGEMA_reg_buffer_4668 ( .C (clk), .D (new_AGEMA_signal_1496), .Q (new_AGEMA_signal_8099) ) ;
    buf_clk new_AGEMA_reg_buffer_4672 ( .C (clk), .D (TweakeyGeneration_StateRegInput[3]), .Q (new_AGEMA_signal_8103) ) ;
    buf_clk new_AGEMA_reg_buffer_4676 ( .C (clk), .D (new_AGEMA_signal_1485), .Q (new_AGEMA_signal_8107) ) ;
    buf_clk new_AGEMA_reg_buffer_4680 ( .C (clk), .D (new_AGEMA_signal_1486), .Q (new_AGEMA_signal_8111) ) ;
    buf_clk new_AGEMA_reg_buffer_4684 ( .C (clk), .D (new_AGEMA_signal_1487), .Q (new_AGEMA_signal_8115) ) ;
    buf_clk new_AGEMA_reg_buffer_4688 ( .C (clk), .D (TweakeyGeneration_StateRegInput[2]), .Q (new_AGEMA_signal_8119) ) ;
    buf_clk new_AGEMA_reg_buffer_4692 ( .C (clk), .D (new_AGEMA_signal_1476), .Q (new_AGEMA_signal_8123) ) ;
    buf_clk new_AGEMA_reg_buffer_4696 ( .C (clk), .D (new_AGEMA_signal_1477), .Q (new_AGEMA_signal_8127) ) ;
    buf_clk new_AGEMA_reg_buffer_4700 ( .C (clk), .D (new_AGEMA_signal_1478), .Q (new_AGEMA_signal_8131) ) ;
    buf_clk new_AGEMA_reg_buffer_4704 ( .C (clk), .D (TweakeyGeneration_StateRegInput[1]), .Q (new_AGEMA_signal_8135) ) ;
    buf_clk new_AGEMA_reg_buffer_4708 ( .C (clk), .D (new_AGEMA_signal_1467), .Q (new_AGEMA_signal_8139) ) ;
    buf_clk new_AGEMA_reg_buffer_4712 ( .C (clk), .D (new_AGEMA_signal_1468), .Q (new_AGEMA_signal_8143) ) ;
    buf_clk new_AGEMA_reg_buffer_4716 ( .C (clk), .D (new_AGEMA_signal_1469), .Q (new_AGEMA_signal_8147) ) ;
    buf_clk new_AGEMA_reg_buffer_4720 ( .C (clk), .D (TweakeyGeneration_StateRegInput[0]), .Q (new_AGEMA_signal_8151) ) ;
    buf_clk new_AGEMA_reg_buffer_4724 ( .C (clk), .D (new_AGEMA_signal_1458), .Q (new_AGEMA_signal_8155) ) ;
    buf_clk new_AGEMA_reg_buffer_4728 ( .C (clk), .D (new_AGEMA_signal_1459), .Q (new_AGEMA_signal_8159) ) ;
    buf_clk new_AGEMA_reg_buffer_4732 ( .C (clk), .D (new_AGEMA_signal_1460), .Q (new_AGEMA_signal_8163) ) ;
    buf_clk new_AGEMA_reg_buffer_4736 ( .C (clk), .D (FSMSelected[5]), .Q (new_AGEMA_signal_8167) ) ;
    buf_clk new_AGEMA_reg_buffer_4740 ( .C (clk), .D (FSMSelected[4]), .Q (new_AGEMA_signal_8171) ) ;
    buf_clk new_AGEMA_reg_buffer_4744 ( .C (clk), .D (FSMSelected[3]), .Q (new_AGEMA_signal_8175) ) ;
    buf_clk new_AGEMA_reg_buffer_4748 ( .C (clk), .D (FSMSelected[2]), .Q (new_AGEMA_signal_8179) ) ;
    buf_clk new_AGEMA_reg_buffer_4752 ( .C (clk), .D (FSMSelected[1]), .Q (new_AGEMA_signal_8183) ) ;
    buf_clk new_AGEMA_reg_buffer_4756 ( .C (clk), .D (FSMSelected[0]), .Q (new_AGEMA_signal_8187) ) ;

    /* cells in depth 2 */
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_2_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, new_AGEMA_signal_3417, MCOutput[2]}), .a ({new_AGEMA_signal_4440, new_AGEMA_signal_4438, new_AGEMA_signal_4436, new_AGEMA_signal_4434}), .c ({new_AGEMA_signal_3440, new_AGEMA_signal_3439, new_AGEMA_signal_3438, StateRegInput[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_3_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, new_AGEMA_signal_3597, MCOutput[3]}), .a ({new_AGEMA_signal_4448, new_AGEMA_signal_4446, new_AGEMA_signal_4444, new_AGEMA_signal_4442}), .c ({new_AGEMA_signal_3620, new_AGEMA_signal_3619, new_AGEMA_signal_3618, StateRegInput[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_6_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, new_AGEMA_signal_3423, MCOutput[6]}), .a ({new_AGEMA_signal_4456, new_AGEMA_signal_4454, new_AGEMA_signal_4452, new_AGEMA_signal_4450}), .c ({new_AGEMA_signal_3446, new_AGEMA_signal_3445, new_AGEMA_signal_3444, StateRegInput[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_7_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, new_AGEMA_signal_3603, MCOutput[7]}), .a ({new_AGEMA_signal_4464, new_AGEMA_signal_4462, new_AGEMA_signal_4460, new_AGEMA_signal_4458}), .c ({new_AGEMA_signal_3626, new_AGEMA_signal_3625, new_AGEMA_signal_3624, StateRegInput[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_10_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, new_AGEMA_signal_3429, MCOutput[10]}), .a ({new_AGEMA_signal_4472, new_AGEMA_signal_4470, new_AGEMA_signal_4468, new_AGEMA_signal_4466}), .c ({new_AGEMA_signal_3452, new_AGEMA_signal_3451, new_AGEMA_signal_3450, StateRegInput[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_11_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, new_AGEMA_signal_3609, MCOutput[11]}), .a ({new_AGEMA_signal_4480, new_AGEMA_signal_4478, new_AGEMA_signal_4476, new_AGEMA_signal_4474}), .c ({new_AGEMA_signal_3632, new_AGEMA_signal_3631, new_AGEMA_signal_3630, StateRegInput[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_14_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, new_AGEMA_signal_3771, MCOutput[14]}), .a ({new_AGEMA_signal_4488, new_AGEMA_signal_4486, new_AGEMA_signal_4484, new_AGEMA_signal_4482}), .c ({new_AGEMA_signal_3800, new_AGEMA_signal_3799, new_AGEMA_signal_3798, StateRegInput[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_15_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, new_AGEMA_signal_3903, MCOutput[15]}), .a ({new_AGEMA_signal_4496, new_AGEMA_signal_4494, new_AGEMA_signal_4492, new_AGEMA_signal_4490}), .c ({new_AGEMA_signal_3929, new_AGEMA_signal_3928, new_AGEMA_signal_3927, StateRegInput[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_18_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, new_AGEMA_signal_3399, MCOutput[18]}), .a ({new_AGEMA_signal_4504, new_AGEMA_signal_4502, new_AGEMA_signal_4500, new_AGEMA_signal_4498}), .c ({new_AGEMA_signal_3458, new_AGEMA_signal_3457, new_AGEMA_signal_3456, StateRegInput[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_19_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3578, new_AGEMA_signal_3577, new_AGEMA_signal_3576, MCOutput[19]}), .a ({new_AGEMA_signal_4512, new_AGEMA_signal_4510, new_AGEMA_signal_4508, new_AGEMA_signal_4506}), .c ({new_AGEMA_signal_3638, new_AGEMA_signal_3637, new_AGEMA_signal_3636, StateRegInput[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_22_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, new_AGEMA_signal_3405, MCOutput[22]}), .a ({new_AGEMA_signal_4520, new_AGEMA_signal_4518, new_AGEMA_signal_4516, new_AGEMA_signal_4514}), .c ({new_AGEMA_signal_3464, new_AGEMA_signal_3463, new_AGEMA_signal_3462, StateRegInput[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_23_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3584, new_AGEMA_signal_3583, new_AGEMA_signal_3582, MCOutput[23]}), .a ({new_AGEMA_signal_4528, new_AGEMA_signal_4526, new_AGEMA_signal_4524, new_AGEMA_signal_4522}), .c ({new_AGEMA_signal_3644, new_AGEMA_signal_3643, new_AGEMA_signal_3642, StateRegInput[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_26_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3743, new_AGEMA_signal_3742, new_AGEMA_signal_3741, MCOutput[26]}), .a ({new_AGEMA_signal_4536, new_AGEMA_signal_4534, new_AGEMA_signal_4532, new_AGEMA_signal_4530}), .c ({new_AGEMA_signal_3818, new_AGEMA_signal_3817, new_AGEMA_signal_3816, StateRegInput[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_27_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3887, new_AGEMA_signal_3886, new_AGEMA_signal_3885, MCOutput[27]}), .a ({new_AGEMA_signal_4544, new_AGEMA_signal_4542, new_AGEMA_signal_4540, new_AGEMA_signal_4538}), .c ({new_AGEMA_signal_3947, new_AGEMA_signal_3946, new_AGEMA_signal_3945, StateRegInput[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_30_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, new_AGEMA_signal_3411, MCOutput[30]}), .a ({new_AGEMA_signal_4552, new_AGEMA_signal_4550, new_AGEMA_signal_4548, new_AGEMA_signal_4546}), .c ({new_AGEMA_signal_3470, new_AGEMA_signal_3469, new_AGEMA_signal_3468, StateRegInput[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_31_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, new_AGEMA_signal_3591, MCOutput[31]}), .a ({new_AGEMA_signal_4560, new_AGEMA_signal_4558, new_AGEMA_signal_4556, new_AGEMA_signal_4554}), .c ({new_AGEMA_signal_3650, new_AGEMA_signal_3649, new_AGEMA_signal_3648, StateRegInput[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_34_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3104, new_AGEMA_signal_3103, new_AGEMA_signal_3102, MCOutput[34]}), .a ({new_AGEMA_signal_4568, new_AGEMA_signal_4566, new_AGEMA_signal_4564, new_AGEMA_signal_4562}), .c ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, new_AGEMA_signal_3135, StateRegInput[34]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_35_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3236, new_AGEMA_signal_3235, new_AGEMA_signal_3234, MCOutput[35]}), .a ({new_AGEMA_signal_4576, new_AGEMA_signal_4574, new_AGEMA_signal_4572, new_AGEMA_signal_4570}), .c ({new_AGEMA_signal_3296, new_AGEMA_signal_3295, new_AGEMA_signal_3294, StateRegInput[35]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_38_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3110, new_AGEMA_signal_3109, new_AGEMA_signal_3108, MCOutput[38]}), .a ({new_AGEMA_signal_4584, new_AGEMA_signal_4582, new_AGEMA_signal_4580, new_AGEMA_signal_4578}), .c ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, new_AGEMA_signal_3141, StateRegInput[38]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_39_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3242, new_AGEMA_signal_3241, new_AGEMA_signal_3240, MCOutput[39]}), .a ({new_AGEMA_signal_4592, new_AGEMA_signal_4590, new_AGEMA_signal_4588, new_AGEMA_signal_4586}), .c ({new_AGEMA_signal_3302, new_AGEMA_signal_3301, new_AGEMA_signal_3300, StateRegInput[39]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_42_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3116, new_AGEMA_signal_3115, new_AGEMA_signal_3114, MCOutput[42]}), .a ({new_AGEMA_signal_4600, new_AGEMA_signal_4598, new_AGEMA_signal_4596, new_AGEMA_signal_4594}), .c ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, new_AGEMA_signal_3147, StateRegInput[42]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_43_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3248, new_AGEMA_signal_3247, new_AGEMA_signal_3246, MCOutput[43]}), .a ({new_AGEMA_signal_4608, new_AGEMA_signal_4606, new_AGEMA_signal_4604, new_AGEMA_signal_4602}), .c ({new_AGEMA_signal_3308, new_AGEMA_signal_3307, new_AGEMA_signal_3306, StateRegInput[43]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_46_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3368, new_AGEMA_signal_3367, new_AGEMA_signal_3366, MCOutput[46]}), .a ({new_AGEMA_signal_4616, new_AGEMA_signal_4614, new_AGEMA_signal_4612, new_AGEMA_signal_4610}), .c ({new_AGEMA_signal_3494, new_AGEMA_signal_3493, new_AGEMA_signal_3492, StateRegInput[46]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_47_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3548, new_AGEMA_signal_3547, new_AGEMA_signal_3546, MCOutput[47]}), .a ({new_AGEMA_signal_4624, new_AGEMA_signal_4622, new_AGEMA_signal_4620, new_AGEMA_signal_4618}), .c ({new_AGEMA_signal_3674, new_AGEMA_signal_3673, new_AGEMA_signal_3672, StateRegInput[47]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_50_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, new_AGEMA_signal_3375, MCOutput[50]}), .a ({new_AGEMA_signal_4632, new_AGEMA_signal_4630, new_AGEMA_signal_4628, new_AGEMA_signal_4626}), .c ({new_AGEMA_signal_3500, new_AGEMA_signal_3499, new_AGEMA_signal_3498, StateRegInput[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_51_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3554, new_AGEMA_signal_3553, new_AGEMA_signal_3552, MCOutput[51]}), .a ({new_AGEMA_signal_4640, new_AGEMA_signal_4638, new_AGEMA_signal_4636, new_AGEMA_signal_4634}), .c ({new_AGEMA_signal_3680, new_AGEMA_signal_3679, new_AGEMA_signal_3678, StateRegInput[51]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_54_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, new_AGEMA_signal_3381, MCOutput[54]}), .a ({new_AGEMA_signal_4648, new_AGEMA_signal_4646, new_AGEMA_signal_4644, new_AGEMA_signal_4642}), .c ({new_AGEMA_signal_3506, new_AGEMA_signal_3505, new_AGEMA_signal_3504, StateRegInput[54]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_55_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, new_AGEMA_signal_3561, MCOutput[55]}), .a ({new_AGEMA_signal_4656, new_AGEMA_signal_4654, new_AGEMA_signal_4652, new_AGEMA_signal_4650}), .c ({new_AGEMA_signal_3686, new_AGEMA_signal_3685, new_AGEMA_signal_3684, StateRegInput[55]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_58_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3392, new_AGEMA_signal_3391, new_AGEMA_signal_3390, MCOutput[58]}), .a ({new_AGEMA_signal_4664, new_AGEMA_signal_4662, new_AGEMA_signal_4660, new_AGEMA_signal_4658}), .c ({new_AGEMA_signal_3512, new_AGEMA_signal_3511, new_AGEMA_signal_3510, StateRegInput[58]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_59_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, new_AGEMA_signal_3567, MCOutput[59]}), .a ({new_AGEMA_signal_4672, new_AGEMA_signal_4670, new_AGEMA_signal_4668, new_AGEMA_signal_4666}), .c ({new_AGEMA_signal_3692, new_AGEMA_signal_3691, new_AGEMA_signal_3690, StateRegInput[59]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_62_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, new_AGEMA_signal_3723, MCOutput[62]}), .a ({new_AGEMA_signal_4680, new_AGEMA_signal_4678, new_AGEMA_signal_4676, new_AGEMA_signal_4674}), .c ({new_AGEMA_signal_3854, new_AGEMA_signal_3853, new_AGEMA_signal_3852, StateRegInput[62]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_63_U1 ( .s (new_AGEMA_signal_4432), .b ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, new_AGEMA_signal_3873, MCOutput[63]}), .a ({new_AGEMA_signal_4688, new_AGEMA_signal_4686, new_AGEMA_signal_4684, new_AGEMA_signal_4682}), .c ({new_AGEMA_signal_3983, new_AGEMA_signal_3982, new_AGEMA_signal_3981, StateRegInput[63]}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_U3 ( .a ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, new_AGEMA_signal_2661, SubCellInst_SboxInst_0_YY_1_}), .b ({new_AGEMA_signal_2846, new_AGEMA_signal_2845, new_AGEMA_signal_2844, ShiftRowsOutput[7]}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_U2 ( .a ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, new_AGEMA_signal_2469, SubCellInst_SboxInst_0_YY_0_}), .b ({new_AGEMA_signal_2654, new_AGEMA_signal_2653, new_AGEMA_signal_2652, ShiftRowsOutput[6]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_AND1_U1 ( .a ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, SubCellInst_SboxInst_0_n3}), .b ({new_AGEMA_signal_2036, new_AGEMA_signal_2035, new_AGEMA_signal_2034, SubCellInst_SboxInst_0_Q1}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_2318, new_AGEMA_signal_2317, new_AGEMA_signal_2316, SubCellInst_SboxInst_0_T0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_XOR2_U1 ( .a ({new_AGEMA_signal_4696, new_AGEMA_signal_4694, new_AGEMA_signal_4692, new_AGEMA_signal_4690}), .b ({new_AGEMA_signal_2318, new_AGEMA_signal_2317, new_AGEMA_signal_2316, SubCellInst_SboxInst_0_T0}), .c ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, new_AGEMA_signal_2460, SubCellInst_SboxInst_0_Q2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_AND3_U1 ( .a ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, SubCellInst_SboxInst_0_n3}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, new_AGEMA_signal_2037, SubCellInst_SboxInst_0_Q4}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, new_AGEMA_signal_2319, SubCellInst_SboxInst_0_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_XOR7_U1 ( .a ({new_AGEMA_signal_4704, new_AGEMA_signal_4702, new_AGEMA_signal_4700, new_AGEMA_signal_4698}), .b ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, new_AGEMA_signal_2319, SubCellInst_SboxInst_0_T2}), .c ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, new_AGEMA_signal_2463, SubCellInst_SboxInst_0_Q7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_XOR11_U1 ( .a ({new_AGEMA_signal_4712, new_AGEMA_signal_4710, new_AGEMA_signal_4708, new_AGEMA_signal_4706}), .b ({new_AGEMA_signal_2318, new_AGEMA_signal_2317, new_AGEMA_signal_2316, SubCellInst_SboxInst_0_T0}), .c ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, new_AGEMA_signal_2466, SubCellInst_SboxInst_0_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_XOR12_U1 ( .a ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, new_AGEMA_signal_2466, SubCellInst_SboxInst_0_L3}), .b ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, new_AGEMA_signal_2319, SubCellInst_SboxInst_0_T2}), .c ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, new_AGEMA_signal_2661, SubCellInst_SboxInst_0_YY_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_XOR13_U1 ( .a ({new_AGEMA_signal_4720, new_AGEMA_signal_4718, new_AGEMA_signal_4716, new_AGEMA_signal_4714}), .b ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, new_AGEMA_signal_2319, SubCellInst_SboxInst_0_T2}), .c ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, new_AGEMA_signal_2469, SubCellInst_SboxInst_0_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_U3 ( .a ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, new_AGEMA_signal_2673, SubCellInst_SboxInst_1_YY_1_}), .b ({new_AGEMA_signal_2852, new_AGEMA_signal_2851, new_AGEMA_signal_2850, ShiftRowsOutput[11]}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_U2 ( .a ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, new_AGEMA_signal_2481, SubCellInst_SboxInst_1_YY_0_}), .b ({new_AGEMA_signal_2666, new_AGEMA_signal_2665, new_AGEMA_signal_2664, ShiftRowsOutput[10]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_AND1_U1 ( .a ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, SubCellInst_SboxInst_1_n3}), .b ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, new_AGEMA_signal_2052, SubCellInst_SboxInst_1_Q1}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, new_AGEMA_signal_2325, SubCellInst_SboxInst_1_T0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_XOR2_U1 ( .a ({new_AGEMA_signal_4728, new_AGEMA_signal_4726, new_AGEMA_signal_4724, new_AGEMA_signal_4722}), .b ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, new_AGEMA_signal_2325, SubCellInst_SboxInst_1_T0}), .c ({new_AGEMA_signal_2474, new_AGEMA_signal_2473, new_AGEMA_signal_2472, SubCellInst_SboxInst_1_Q2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_AND3_U1 ( .a ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, SubCellInst_SboxInst_1_n3}), .b ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, new_AGEMA_signal_2055, SubCellInst_SboxInst_1_Q4}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, new_AGEMA_signal_2328, SubCellInst_SboxInst_1_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_XOR7_U1 ( .a ({new_AGEMA_signal_4736, new_AGEMA_signal_4734, new_AGEMA_signal_4732, new_AGEMA_signal_4730}), .b ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, new_AGEMA_signal_2328, SubCellInst_SboxInst_1_T2}), .c ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, new_AGEMA_signal_2475, SubCellInst_SboxInst_1_Q7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_XOR11_U1 ( .a ({new_AGEMA_signal_4744, new_AGEMA_signal_4742, new_AGEMA_signal_4740, new_AGEMA_signal_4738}), .b ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, new_AGEMA_signal_2325, SubCellInst_SboxInst_1_T0}), .c ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, new_AGEMA_signal_2478, SubCellInst_SboxInst_1_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_XOR12_U1 ( .a ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, new_AGEMA_signal_2478, SubCellInst_SboxInst_1_L3}), .b ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, new_AGEMA_signal_2328, SubCellInst_SboxInst_1_T2}), .c ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, new_AGEMA_signal_2673, SubCellInst_SboxInst_1_YY_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_XOR13_U1 ( .a ({new_AGEMA_signal_4752, new_AGEMA_signal_4750, new_AGEMA_signal_4748, new_AGEMA_signal_4746}), .b ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, new_AGEMA_signal_2328, SubCellInst_SboxInst_1_T2}), .c ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, new_AGEMA_signal_2481, SubCellInst_SboxInst_1_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_U3 ( .a ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, new_AGEMA_signal_2685, SubCellInst_SboxInst_2_YY_1_}), .b ({new_AGEMA_signal_2858, new_AGEMA_signal_2857, new_AGEMA_signal_2856, ShiftRowsOutput[15]}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_U2 ( .a ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, new_AGEMA_signal_2493, SubCellInst_SboxInst_2_YY_0_}), .b ({new_AGEMA_signal_2678, new_AGEMA_signal_2677, new_AGEMA_signal_2676, ShiftRowsOutput[14]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_AND1_U1 ( .a ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, SubCellInst_SboxInst_2_n3}), .b ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, new_AGEMA_signal_2070, SubCellInst_SboxInst_2_Q1}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_2336, new_AGEMA_signal_2335, new_AGEMA_signal_2334, SubCellInst_SboxInst_2_T0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_XOR2_U1 ( .a ({new_AGEMA_signal_4760, new_AGEMA_signal_4758, new_AGEMA_signal_4756, new_AGEMA_signal_4754}), .b ({new_AGEMA_signal_2336, new_AGEMA_signal_2335, new_AGEMA_signal_2334, SubCellInst_SboxInst_2_T0}), .c ({new_AGEMA_signal_2486, new_AGEMA_signal_2485, new_AGEMA_signal_2484, SubCellInst_SboxInst_2_Q2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_AND3_U1 ( .a ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, SubCellInst_SboxInst_2_n3}), .b ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, new_AGEMA_signal_2073, SubCellInst_SboxInst_2_Q4}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, new_AGEMA_signal_2337, SubCellInst_SboxInst_2_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_XOR7_U1 ( .a ({new_AGEMA_signal_4768, new_AGEMA_signal_4766, new_AGEMA_signal_4764, new_AGEMA_signal_4762}), .b ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, new_AGEMA_signal_2337, SubCellInst_SboxInst_2_T2}), .c ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, new_AGEMA_signal_2487, SubCellInst_SboxInst_2_Q7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_XOR11_U1 ( .a ({new_AGEMA_signal_4776, new_AGEMA_signal_4774, new_AGEMA_signal_4772, new_AGEMA_signal_4770}), .b ({new_AGEMA_signal_2336, new_AGEMA_signal_2335, new_AGEMA_signal_2334, SubCellInst_SboxInst_2_T0}), .c ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, new_AGEMA_signal_2490, SubCellInst_SboxInst_2_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_XOR12_U1 ( .a ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, new_AGEMA_signal_2490, SubCellInst_SboxInst_2_L3}), .b ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, new_AGEMA_signal_2337, SubCellInst_SboxInst_2_T2}), .c ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, new_AGEMA_signal_2685, SubCellInst_SboxInst_2_YY_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_XOR13_U1 ( .a ({new_AGEMA_signal_4784, new_AGEMA_signal_4782, new_AGEMA_signal_4780, new_AGEMA_signal_4778}), .b ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, new_AGEMA_signal_2337, SubCellInst_SboxInst_2_T2}), .c ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, new_AGEMA_signal_2493, SubCellInst_SboxInst_2_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_U3 ( .a ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, new_AGEMA_signal_2697, SubCellInst_SboxInst_3_YY_1_}), .b ({new_AGEMA_signal_2864, new_AGEMA_signal_2863, new_AGEMA_signal_2862, ShiftRowsOutput[3]}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_U2 ( .a ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, new_AGEMA_signal_2505, SubCellInst_SboxInst_3_YY_0_}), .b ({new_AGEMA_signal_2690, new_AGEMA_signal_2689, new_AGEMA_signal_2688, ShiftRowsOutput[2]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_AND1_U1 ( .a ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, SubCellInst_SboxInst_3_n3}), .b ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, SubCellInst_SboxInst_3_Q1}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, new_AGEMA_signal_2343, SubCellInst_SboxInst_3_T0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_XOR2_U1 ( .a ({new_AGEMA_signal_4792, new_AGEMA_signal_4790, new_AGEMA_signal_4788, new_AGEMA_signal_4786}), .b ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, new_AGEMA_signal_2343, SubCellInst_SboxInst_3_T0}), .c ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, new_AGEMA_signal_2496, SubCellInst_SboxInst_3_Q2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_AND3_U1 ( .a ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, SubCellInst_SboxInst_3_n3}), .b ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, new_AGEMA_signal_2091, SubCellInst_SboxInst_3_Q4}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_2348, new_AGEMA_signal_2347, new_AGEMA_signal_2346, SubCellInst_SboxInst_3_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_XOR7_U1 ( .a ({new_AGEMA_signal_4800, new_AGEMA_signal_4798, new_AGEMA_signal_4796, new_AGEMA_signal_4794}), .b ({new_AGEMA_signal_2348, new_AGEMA_signal_2347, new_AGEMA_signal_2346, SubCellInst_SboxInst_3_T2}), .c ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, new_AGEMA_signal_2499, SubCellInst_SboxInst_3_Q7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_XOR11_U1 ( .a ({new_AGEMA_signal_4808, new_AGEMA_signal_4806, new_AGEMA_signal_4804, new_AGEMA_signal_4802}), .b ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, new_AGEMA_signal_2343, SubCellInst_SboxInst_3_T0}), .c ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, new_AGEMA_signal_2502, SubCellInst_SboxInst_3_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_XOR12_U1 ( .a ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, new_AGEMA_signal_2502, SubCellInst_SboxInst_3_L3}), .b ({new_AGEMA_signal_2348, new_AGEMA_signal_2347, new_AGEMA_signal_2346, SubCellInst_SboxInst_3_T2}), .c ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, new_AGEMA_signal_2697, SubCellInst_SboxInst_3_YY_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_XOR13_U1 ( .a ({new_AGEMA_signal_4816, new_AGEMA_signal_4814, new_AGEMA_signal_4812, new_AGEMA_signal_4810}), .b ({new_AGEMA_signal_2348, new_AGEMA_signal_2347, new_AGEMA_signal_2346, SubCellInst_SboxInst_3_T2}), .c ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, new_AGEMA_signal_2505, SubCellInst_SboxInst_3_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_U3 ( .a ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, new_AGEMA_signal_2709, SubCellInst_SboxInst_4_YY_1_}), .b ({new_AGEMA_signal_2870, new_AGEMA_signal_2869, new_AGEMA_signal_2868, ShiftRowsOutput[27]}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_U2 ( .a ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, new_AGEMA_signal_2517, SubCellInst_SboxInst_4_YY_0_}), .b ({new_AGEMA_signal_2702, new_AGEMA_signal_2701, new_AGEMA_signal_2700, ShiftRowsOutput[26]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_AND1_U1 ( .a ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_4_n3}), .b ({new_AGEMA_signal_2108, new_AGEMA_signal_2107, new_AGEMA_signal_2106, SubCellInst_SboxInst_4_Q1}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, new_AGEMA_signal_2352, SubCellInst_SboxInst_4_T0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_XOR2_U1 ( .a ({new_AGEMA_signal_4824, new_AGEMA_signal_4822, new_AGEMA_signal_4820, new_AGEMA_signal_4818}), .b ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, new_AGEMA_signal_2352, SubCellInst_SboxInst_4_T0}), .c ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, new_AGEMA_signal_2508, SubCellInst_SboxInst_4_Q2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_AND3_U1 ( .a ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_4_n3}), .b ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, new_AGEMA_signal_2109, SubCellInst_SboxInst_4_Q4}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, new_AGEMA_signal_2355, SubCellInst_SboxInst_4_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_XOR7_U1 ( .a ({new_AGEMA_signal_4832, new_AGEMA_signal_4830, new_AGEMA_signal_4828, new_AGEMA_signal_4826}), .b ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, new_AGEMA_signal_2355, SubCellInst_SboxInst_4_T2}), .c ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, new_AGEMA_signal_2511, SubCellInst_SboxInst_4_Q7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_XOR11_U1 ( .a ({new_AGEMA_signal_4840, new_AGEMA_signal_4838, new_AGEMA_signal_4836, new_AGEMA_signal_4834}), .b ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, new_AGEMA_signal_2352, SubCellInst_SboxInst_4_T0}), .c ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, new_AGEMA_signal_2514, SubCellInst_SboxInst_4_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_XOR12_U1 ( .a ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, new_AGEMA_signal_2514, SubCellInst_SboxInst_4_L3}), .b ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, new_AGEMA_signal_2355, SubCellInst_SboxInst_4_T2}), .c ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, new_AGEMA_signal_2709, SubCellInst_SboxInst_4_YY_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_XOR13_U1 ( .a ({new_AGEMA_signal_4848, new_AGEMA_signal_4846, new_AGEMA_signal_4844, new_AGEMA_signal_4842}), .b ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, new_AGEMA_signal_2355, SubCellInst_SboxInst_4_T2}), .c ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, new_AGEMA_signal_2517, SubCellInst_SboxInst_4_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_U3 ( .a ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, new_AGEMA_signal_2721, SubCellInst_SboxInst_5_YY_1_}), .b ({new_AGEMA_signal_2876, new_AGEMA_signal_2875, new_AGEMA_signal_2874, ShiftRowsOutput[31]}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_U2 ( .a ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, new_AGEMA_signal_2529, SubCellInst_SboxInst_5_YY_0_}), .b ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, new_AGEMA_signal_2712, ShiftRowsOutput[30]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_AND1_U1 ( .a ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_5_n3}), .b ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, new_AGEMA_signal_2124, SubCellInst_SboxInst_5_Q1}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, new_AGEMA_signal_2361, SubCellInst_SboxInst_5_T0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_XOR2_U1 ( .a ({new_AGEMA_signal_4856, new_AGEMA_signal_4854, new_AGEMA_signal_4852, new_AGEMA_signal_4850}), .b ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, new_AGEMA_signal_2361, SubCellInst_SboxInst_5_T0}), .c ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, new_AGEMA_signal_2520, SubCellInst_SboxInst_5_Q2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_AND3_U1 ( .a ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_5_n3}), .b ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, new_AGEMA_signal_2127, SubCellInst_SboxInst_5_Q4}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, new_AGEMA_signal_2364, SubCellInst_SboxInst_5_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_XOR7_U1 ( .a ({new_AGEMA_signal_4864, new_AGEMA_signal_4862, new_AGEMA_signal_4860, new_AGEMA_signal_4858}), .b ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, new_AGEMA_signal_2364, SubCellInst_SboxInst_5_T2}), .c ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, new_AGEMA_signal_2523, SubCellInst_SboxInst_5_Q7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_XOR11_U1 ( .a ({new_AGEMA_signal_4872, new_AGEMA_signal_4870, new_AGEMA_signal_4868, new_AGEMA_signal_4866}), .b ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, new_AGEMA_signal_2361, SubCellInst_SboxInst_5_T0}), .c ({new_AGEMA_signal_2528, new_AGEMA_signal_2527, new_AGEMA_signal_2526, SubCellInst_SboxInst_5_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_XOR12_U1 ( .a ({new_AGEMA_signal_2528, new_AGEMA_signal_2527, new_AGEMA_signal_2526, SubCellInst_SboxInst_5_L3}), .b ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, new_AGEMA_signal_2364, SubCellInst_SboxInst_5_T2}), .c ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, new_AGEMA_signal_2721, SubCellInst_SboxInst_5_YY_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_XOR13_U1 ( .a ({new_AGEMA_signal_4880, new_AGEMA_signal_4878, new_AGEMA_signal_4876, new_AGEMA_signal_4874}), .b ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, new_AGEMA_signal_2364, SubCellInst_SboxInst_5_T2}), .c ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, new_AGEMA_signal_2529, SubCellInst_SboxInst_5_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_U3 ( .a ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, new_AGEMA_signal_2733, SubCellInst_SboxInst_6_YY_1_}), .b ({new_AGEMA_signal_2882, new_AGEMA_signal_2881, new_AGEMA_signal_2880, ShiftRowsOutput[19]}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_U2 ( .a ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, new_AGEMA_signal_2541, SubCellInst_SboxInst_6_YY_0_}), .b ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, new_AGEMA_signal_2724, ShiftRowsOutput[18]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_AND1_U1 ( .a ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_6_n3}), .b ({new_AGEMA_signal_2144, new_AGEMA_signal_2143, new_AGEMA_signal_2142, SubCellInst_SboxInst_6_Q1}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_2372, new_AGEMA_signal_2371, new_AGEMA_signal_2370, SubCellInst_SboxInst_6_T0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_XOR2_U1 ( .a ({new_AGEMA_signal_4888, new_AGEMA_signal_4886, new_AGEMA_signal_4884, new_AGEMA_signal_4882}), .b ({new_AGEMA_signal_2372, new_AGEMA_signal_2371, new_AGEMA_signal_2370, SubCellInst_SboxInst_6_T0}), .c ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, new_AGEMA_signal_2532, SubCellInst_SboxInst_6_Q2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_AND3_U1 ( .a ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_6_n3}), .b ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, new_AGEMA_signal_2145, SubCellInst_SboxInst_6_Q4}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, new_AGEMA_signal_2373, SubCellInst_SboxInst_6_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_XOR7_U1 ( .a ({new_AGEMA_signal_4896, new_AGEMA_signal_4894, new_AGEMA_signal_4892, new_AGEMA_signal_4890}), .b ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, new_AGEMA_signal_2373, SubCellInst_SboxInst_6_T2}), .c ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, new_AGEMA_signal_2535, SubCellInst_SboxInst_6_Q7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_XOR11_U1 ( .a ({new_AGEMA_signal_4904, new_AGEMA_signal_4902, new_AGEMA_signal_4900, new_AGEMA_signal_4898}), .b ({new_AGEMA_signal_2372, new_AGEMA_signal_2371, new_AGEMA_signal_2370, SubCellInst_SboxInst_6_T0}), .c ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, new_AGEMA_signal_2538, SubCellInst_SboxInst_6_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_XOR12_U1 ( .a ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, new_AGEMA_signal_2538, SubCellInst_SboxInst_6_L3}), .b ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, new_AGEMA_signal_2373, SubCellInst_SboxInst_6_T2}), .c ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, new_AGEMA_signal_2733, SubCellInst_SboxInst_6_YY_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_XOR13_U1 ( .a ({new_AGEMA_signal_4912, new_AGEMA_signal_4910, new_AGEMA_signal_4908, new_AGEMA_signal_4906}), .b ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, new_AGEMA_signal_2373, SubCellInst_SboxInst_6_T2}), .c ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, new_AGEMA_signal_2541, SubCellInst_SboxInst_6_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_U3 ( .a ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, new_AGEMA_signal_2745, SubCellInst_SboxInst_7_YY_1_}), .b ({new_AGEMA_signal_2888, new_AGEMA_signal_2887, new_AGEMA_signal_2886, ShiftRowsOutput[23]}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_U2 ( .a ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, new_AGEMA_signal_2553, SubCellInst_SboxInst_7_YY_0_}), .b ({new_AGEMA_signal_2738, new_AGEMA_signal_2737, new_AGEMA_signal_2736, ShiftRowsOutput[22]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_AND1_U1 ( .a ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, SubCellInst_SboxInst_7_n3}), .b ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, new_AGEMA_signal_2160, SubCellInst_SboxInst_7_Q1}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, new_AGEMA_signal_2379, SubCellInst_SboxInst_7_T0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_XOR2_U1 ( .a ({new_AGEMA_signal_4920, new_AGEMA_signal_4918, new_AGEMA_signal_4916, new_AGEMA_signal_4914}), .b ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, new_AGEMA_signal_2379, SubCellInst_SboxInst_7_T0}), .c ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, new_AGEMA_signal_2544, SubCellInst_SboxInst_7_Q2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_AND3_U1 ( .a ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, SubCellInst_SboxInst_7_n3}), .b ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, new_AGEMA_signal_2163, SubCellInst_SboxInst_7_Q4}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_2384, new_AGEMA_signal_2383, new_AGEMA_signal_2382, SubCellInst_SboxInst_7_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_XOR7_U1 ( .a ({new_AGEMA_signal_4928, new_AGEMA_signal_4926, new_AGEMA_signal_4924, new_AGEMA_signal_4922}), .b ({new_AGEMA_signal_2384, new_AGEMA_signal_2383, new_AGEMA_signal_2382, SubCellInst_SboxInst_7_T2}), .c ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, new_AGEMA_signal_2547, SubCellInst_SboxInst_7_Q7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_XOR11_U1 ( .a ({new_AGEMA_signal_4936, new_AGEMA_signal_4934, new_AGEMA_signal_4932, new_AGEMA_signal_4930}), .b ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, new_AGEMA_signal_2379, SubCellInst_SboxInst_7_T0}), .c ({new_AGEMA_signal_2552, new_AGEMA_signal_2551, new_AGEMA_signal_2550, SubCellInst_SboxInst_7_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_XOR12_U1 ( .a ({new_AGEMA_signal_2552, new_AGEMA_signal_2551, new_AGEMA_signal_2550, SubCellInst_SboxInst_7_L3}), .b ({new_AGEMA_signal_2384, new_AGEMA_signal_2383, new_AGEMA_signal_2382, SubCellInst_SboxInst_7_T2}), .c ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, new_AGEMA_signal_2745, SubCellInst_SboxInst_7_YY_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_XOR13_U1 ( .a ({new_AGEMA_signal_4944, new_AGEMA_signal_4942, new_AGEMA_signal_4940, new_AGEMA_signal_4938}), .b ({new_AGEMA_signal_2384, new_AGEMA_signal_2383, new_AGEMA_signal_2382, SubCellInst_SboxInst_7_T2}), .c ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, new_AGEMA_signal_2553, SubCellInst_SboxInst_7_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_U3 ( .a ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, new_AGEMA_signal_2757, SubCellInst_SboxInst_8_YY_1_}), .b ({new_AGEMA_signal_2894, new_AGEMA_signal_2893, new_AGEMA_signal_2892, AddRoundConstantOutput[35]}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_U2 ( .a ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, new_AGEMA_signal_2565, SubCellInst_SboxInst_8_YY_0_}), .b ({new_AGEMA_signal_2750, new_AGEMA_signal_2749, new_AGEMA_signal_2748, AddRoundConstantOutput[34]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_AND1_U1 ( .a ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, SubCellInst_SboxInst_8_n3}), .b ({new_AGEMA_signal_2180, new_AGEMA_signal_2179, new_AGEMA_signal_2178, SubCellInst_SboxInst_8_Q1}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, new_AGEMA_signal_2388, SubCellInst_SboxInst_8_T0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_XOR2_U1 ( .a ({new_AGEMA_signal_4952, new_AGEMA_signal_4950, new_AGEMA_signal_4948, new_AGEMA_signal_4946}), .b ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, new_AGEMA_signal_2388, SubCellInst_SboxInst_8_T0}), .c ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, new_AGEMA_signal_2556, SubCellInst_SboxInst_8_Q2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_AND3_U1 ( .a ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, SubCellInst_SboxInst_8_n3}), .b ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, new_AGEMA_signal_2181, SubCellInst_SboxInst_8_Q4}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, new_AGEMA_signal_2391, SubCellInst_SboxInst_8_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_XOR7_U1 ( .a ({new_AGEMA_signal_4960, new_AGEMA_signal_4958, new_AGEMA_signal_4956, new_AGEMA_signal_4954}), .b ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, new_AGEMA_signal_2391, SubCellInst_SboxInst_8_T2}), .c ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, new_AGEMA_signal_2559, SubCellInst_SboxInst_8_Q7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_XOR11_U1 ( .a ({new_AGEMA_signal_4968, new_AGEMA_signal_4966, new_AGEMA_signal_4964, new_AGEMA_signal_4962}), .b ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, new_AGEMA_signal_2388, SubCellInst_SboxInst_8_T0}), .c ({new_AGEMA_signal_2564, new_AGEMA_signal_2563, new_AGEMA_signal_2562, SubCellInst_SboxInst_8_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_XOR12_U1 ( .a ({new_AGEMA_signal_2564, new_AGEMA_signal_2563, new_AGEMA_signal_2562, SubCellInst_SboxInst_8_L3}), .b ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, new_AGEMA_signal_2391, SubCellInst_SboxInst_8_T2}), .c ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, new_AGEMA_signal_2757, SubCellInst_SboxInst_8_YY_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_XOR13_U1 ( .a ({new_AGEMA_signal_4976, new_AGEMA_signal_4974, new_AGEMA_signal_4972, new_AGEMA_signal_4970}), .b ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, new_AGEMA_signal_2391, SubCellInst_SboxInst_8_T2}), .c ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, new_AGEMA_signal_2565, SubCellInst_SboxInst_8_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_U3 ( .a ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, new_AGEMA_signal_2769, SubCellInst_SboxInst_9_YY_1_}), .b ({new_AGEMA_signal_2900, new_AGEMA_signal_2899, new_AGEMA_signal_2898, AddRoundConstantOutput[39]}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_U2 ( .a ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, new_AGEMA_signal_2577, SubCellInst_SboxInst_9_YY_0_}), .b ({new_AGEMA_signal_2762, new_AGEMA_signal_2761, new_AGEMA_signal_2760, AddRoundConstantOutput[38]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_AND1_U1 ( .a ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, new_AGEMA_signal_1329, SubCellInst_SboxInst_9_n3}), .b ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, new_AGEMA_signal_2196, SubCellInst_SboxInst_9_Q1}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, new_AGEMA_signal_2397, SubCellInst_SboxInst_9_T0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_XOR2_U1 ( .a ({new_AGEMA_signal_4984, new_AGEMA_signal_4982, new_AGEMA_signal_4980, new_AGEMA_signal_4978}), .b ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, new_AGEMA_signal_2397, SubCellInst_SboxInst_9_T0}), .c ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, new_AGEMA_signal_2568, SubCellInst_SboxInst_9_Q2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_AND3_U1 ( .a ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, new_AGEMA_signal_1329, SubCellInst_SboxInst_9_n3}), .b ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, new_AGEMA_signal_2199, SubCellInst_SboxInst_9_Q4}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, new_AGEMA_signal_2400, SubCellInst_SboxInst_9_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_XOR7_U1 ( .a ({new_AGEMA_signal_4992, new_AGEMA_signal_4990, new_AGEMA_signal_4988, new_AGEMA_signal_4986}), .b ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, new_AGEMA_signal_2400, SubCellInst_SboxInst_9_T2}), .c ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, new_AGEMA_signal_2571, SubCellInst_SboxInst_9_Q7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_XOR11_U1 ( .a ({new_AGEMA_signal_5000, new_AGEMA_signal_4998, new_AGEMA_signal_4996, new_AGEMA_signal_4994}), .b ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, new_AGEMA_signal_2397, SubCellInst_SboxInst_9_T0}), .c ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, new_AGEMA_signal_2574, SubCellInst_SboxInst_9_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_XOR12_U1 ( .a ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, new_AGEMA_signal_2574, SubCellInst_SboxInst_9_L3}), .b ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, new_AGEMA_signal_2400, SubCellInst_SboxInst_9_T2}), .c ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, new_AGEMA_signal_2769, SubCellInst_SboxInst_9_YY_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_XOR13_U1 ( .a ({new_AGEMA_signal_5008, new_AGEMA_signal_5006, new_AGEMA_signal_5004, new_AGEMA_signal_5002}), .b ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, new_AGEMA_signal_2400, SubCellInst_SboxInst_9_T2}), .c ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, new_AGEMA_signal_2577, SubCellInst_SboxInst_9_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_U3 ( .a ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, new_AGEMA_signal_2781, SubCellInst_SboxInst_10_YY_1_}), .b ({new_AGEMA_signal_2906, new_AGEMA_signal_2905, new_AGEMA_signal_2904, AddRoundConstantOutput[43]}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_U2 ( .a ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, new_AGEMA_signal_2589, SubCellInst_SboxInst_10_YY_0_}), .b ({new_AGEMA_signal_2774, new_AGEMA_signal_2773, new_AGEMA_signal_2772, AddRoundConstantOutput[42]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_AND1_U1 ( .a ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, SubCellInst_SboxInst_10_n3}), .b ({new_AGEMA_signal_2216, new_AGEMA_signal_2215, new_AGEMA_signal_2214, SubCellInst_SboxInst_10_Q1}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, new_AGEMA_signal_2406, SubCellInst_SboxInst_10_T0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_XOR2_U1 ( .a ({new_AGEMA_signal_5016, new_AGEMA_signal_5014, new_AGEMA_signal_5012, new_AGEMA_signal_5010}), .b ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, new_AGEMA_signal_2406, SubCellInst_SboxInst_10_T0}), .c ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, new_AGEMA_signal_2580, SubCellInst_SboxInst_10_Q2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_AND3_U1 ( .a ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, SubCellInst_SboxInst_10_n3}), .b ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, new_AGEMA_signal_2217, SubCellInst_SboxInst_10_Q4}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, new_AGEMA_signal_2409, SubCellInst_SboxInst_10_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_XOR7_U1 ( .a ({new_AGEMA_signal_5024, new_AGEMA_signal_5022, new_AGEMA_signal_5020, new_AGEMA_signal_5018}), .b ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, new_AGEMA_signal_2409, SubCellInst_SboxInst_10_T2}), .c ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, new_AGEMA_signal_2583, SubCellInst_SboxInst_10_Q7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_XOR11_U1 ( .a ({new_AGEMA_signal_5032, new_AGEMA_signal_5030, new_AGEMA_signal_5028, new_AGEMA_signal_5026}), .b ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, new_AGEMA_signal_2406, SubCellInst_SboxInst_10_T0}), .c ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, new_AGEMA_signal_2586, SubCellInst_SboxInst_10_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_XOR12_U1 ( .a ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, new_AGEMA_signal_2586, SubCellInst_SboxInst_10_L3}), .b ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, new_AGEMA_signal_2409, SubCellInst_SboxInst_10_T2}), .c ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, new_AGEMA_signal_2781, SubCellInst_SboxInst_10_YY_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_XOR13_U1 ( .a ({new_AGEMA_signal_5040, new_AGEMA_signal_5038, new_AGEMA_signal_5036, new_AGEMA_signal_5034}), .b ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, new_AGEMA_signal_2409, SubCellInst_SboxInst_10_T2}), .c ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, new_AGEMA_signal_2589, SubCellInst_SboxInst_10_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_U3 ( .a ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, new_AGEMA_signal_2793, SubCellInst_SboxInst_11_YY_1_}), .b ({new_AGEMA_signal_2912, new_AGEMA_signal_2911, new_AGEMA_signal_2910, SubCellOutput[47]}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_U2 ( .a ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, new_AGEMA_signal_2601, SubCellInst_SboxInst_11_YY_0_}), .b ({new_AGEMA_signal_2786, new_AGEMA_signal_2785, new_AGEMA_signal_2784, SubCellOutput[46]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_AND1_U1 ( .a ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, new_AGEMA_signal_1365, SubCellInst_SboxInst_11_n3}), .b ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, new_AGEMA_signal_2232, SubCellInst_SboxInst_11_Q1}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, new_AGEMA_signal_2415, SubCellInst_SboxInst_11_T0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_XOR2_U1 ( .a ({new_AGEMA_signal_5048, new_AGEMA_signal_5046, new_AGEMA_signal_5044, new_AGEMA_signal_5042}), .b ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, new_AGEMA_signal_2415, SubCellInst_SboxInst_11_T0}), .c ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, new_AGEMA_signal_2592, SubCellInst_SboxInst_11_Q2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_AND3_U1 ( .a ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, new_AGEMA_signal_1365, SubCellInst_SboxInst_11_n3}), .b ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, new_AGEMA_signal_2235, SubCellInst_SboxInst_11_Q4}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, new_AGEMA_signal_2418, SubCellInst_SboxInst_11_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_XOR7_U1 ( .a ({new_AGEMA_signal_5056, new_AGEMA_signal_5054, new_AGEMA_signal_5052, new_AGEMA_signal_5050}), .b ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, new_AGEMA_signal_2418, SubCellInst_SboxInst_11_T2}), .c ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, new_AGEMA_signal_2595, SubCellInst_SboxInst_11_Q7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_XOR11_U1 ( .a ({new_AGEMA_signal_5064, new_AGEMA_signal_5062, new_AGEMA_signal_5060, new_AGEMA_signal_5058}), .b ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, new_AGEMA_signal_2415, SubCellInst_SboxInst_11_T0}), .c ({new_AGEMA_signal_2600, new_AGEMA_signal_2599, new_AGEMA_signal_2598, SubCellInst_SboxInst_11_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_XOR12_U1 ( .a ({new_AGEMA_signal_2600, new_AGEMA_signal_2599, new_AGEMA_signal_2598, SubCellInst_SboxInst_11_L3}), .b ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, new_AGEMA_signal_2418, SubCellInst_SboxInst_11_T2}), .c ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, new_AGEMA_signal_2793, SubCellInst_SboxInst_11_YY_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_XOR13_U1 ( .a ({new_AGEMA_signal_5072, new_AGEMA_signal_5070, new_AGEMA_signal_5068, new_AGEMA_signal_5066}), .b ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, new_AGEMA_signal_2418, SubCellInst_SboxInst_11_T2}), .c ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, new_AGEMA_signal_2601, SubCellInst_SboxInst_11_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_U3 ( .a ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, new_AGEMA_signal_2805, SubCellInst_SboxInst_12_YY_1_}), .b ({new_AGEMA_signal_2918, new_AGEMA_signal_2917, new_AGEMA_signal_2916, AddRoundConstantOutput[51]}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_U2 ( .a ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, new_AGEMA_signal_2613, SubCellInst_SboxInst_12_YY_0_}), .b ({new_AGEMA_signal_2798, new_AGEMA_signal_2797, new_AGEMA_signal_2796, AddRoundConstantOutput[50]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_AND1_U1 ( .a ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, SubCellInst_SboxInst_12_n3}), .b ({new_AGEMA_signal_2252, new_AGEMA_signal_2251, new_AGEMA_signal_2250, SubCellInst_SboxInst_12_Q1}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, new_AGEMA_signal_2424, SubCellInst_SboxInst_12_T0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_XOR2_U1 ( .a ({new_AGEMA_signal_5080, new_AGEMA_signal_5078, new_AGEMA_signal_5076, new_AGEMA_signal_5074}), .b ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, new_AGEMA_signal_2424, SubCellInst_SboxInst_12_T0}), .c ({new_AGEMA_signal_2606, new_AGEMA_signal_2605, new_AGEMA_signal_2604, SubCellInst_SboxInst_12_Q2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_AND3_U1 ( .a ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, SubCellInst_SboxInst_12_n3}), .b ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, new_AGEMA_signal_2253, SubCellInst_SboxInst_12_Q4}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, new_AGEMA_signal_2427, SubCellInst_SboxInst_12_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_XOR7_U1 ( .a ({new_AGEMA_signal_5088, new_AGEMA_signal_5086, new_AGEMA_signal_5084, new_AGEMA_signal_5082}), .b ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, new_AGEMA_signal_2427, SubCellInst_SboxInst_12_T2}), .c ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, new_AGEMA_signal_2607, SubCellInst_SboxInst_12_Q7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_XOR11_U1 ( .a ({new_AGEMA_signal_5096, new_AGEMA_signal_5094, new_AGEMA_signal_5092, new_AGEMA_signal_5090}), .b ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, new_AGEMA_signal_2424, SubCellInst_SboxInst_12_T0}), .c ({new_AGEMA_signal_2612, new_AGEMA_signal_2611, new_AGEMA_signal_2610, SubCellInst_SboxInst_12_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_XOR12_U1 ( .a ({new_AGEMA_signal_2612, new_AGEMA_signal_2611, new_AGEMA_signal_2610, SubCellInst_SboxInst_12_L3}), .b ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, new_AGEMA_signal_2427, SubCellInst_SboxInst_12_T2}), .c ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, new_AGEMA_signal_2805, SubCellInst_SboxInst_12_YY_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_XOR13_U1 ( .a ({new_AGEMA_signal_5104, new_AGEMA_signal_5102, new_AGEMA_signal_5100, new_AGEMA_signal_5098}), .b ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, new_AGEMA_signal_2427, SubCellInst_SboxInst_12_T2}), .c ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, new_AGEMA_signal_2613, SubCellInst_SboxInst_12_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_U3 ( .a ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, new_AGEMA_signal_2817, SubCellInst_SboxInst_13_YY_1_}), .b ({new_AGEMA_signal_2924, new_AGEMA_signal_2923, new_AGEMA_signal_2922, AddRoundConstantOutput[55]}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_U2 ( .a ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, new_AGEMA_signal_2625, SubCellInst_SboxInst_13_YY_0_}), .b ({new_AGEMA_signal_2810, new_AGEMA_signal_2809, new_AGEMA_signal_2808, AddRoundConstantOutput[54]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_AND1_U1 ( .a ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, SubCellInst_SboxInst_13_n3}), .b ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, new_AGEMA_signal_2268, SubCellInst_SboxInst_13_Q1}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, new_AGEMA_signal_2433, SubCellInst_SboxInst_13_T0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_XOR2_U1 ( .a ({new_AGEMA_signal_5112, new_AGEMA_signal_5110, new_AGEMA_signal_5108, new_AGEMA_signal_5106}), .b ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, new_AGEMA_signal_2433, SubCellInst_SboxInst_13_T0}), .c ({new_AGEMA_signal_2618, new_AGEMA_signal_2617, new_AGEMA_signal_2616, SubCellInst_SboxInst_13_Q2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_AND3_U1 ( .a ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, SubCellInst_SboxInst_13_n3}), .b ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, new_AGEMA_signal_2271, SubCellInst_SboxInst_13_Q4}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, new_AGEMA_signal_2436, SubCellInst_SboxInst_13_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_XOR7_U1 ( .a ({new_AGEMA_signal_5120, new_AGEMA_signal_5118, new_AGEMA_signal_5116, new_AGEMA_signal_5114}), .b ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, new_AGEMA_signal_2436, SubCellInst_SboxInst_13_T2}), .c ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, new_AGEMA_signal_2619, SubCellInst_SboxInst_13_Q7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_XOR11_U1 ( .a ({new_AGEMA_signal_5128, new_AGEMA_signal_5126, new_AGEMA_signal_5124, new_AGEMA_signal_5122}), .b ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, new_AGEMA_signal_2433, SubCellInst_SboxInst_13_T0}), .c ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, new_AGEMA_signal_2622, SubCellInst_SboxInst_13_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_XOR12_U1 ( .a ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, new_AGEMA_signal_2622, SubCellInst_SboxInst_13_L3}), .b ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, new_AGEMA_signal_2436, SubCellInst_SboxInst_13_T2}), .c ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, new_AGEMA_signal_2817, SubCellInst_SboxInst_13_YY_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_XOR13_U1 ( .a ({new_AGEMA_signal_5136, new_AGEMA_signal_5134, new_AGEMA_signal_5132, new_AGEMA_signal_5130}), .b ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, new_AGEMA_signal_2436, SubCellInst_SboxInst_13_T2}), .c ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, new_AGEMA_signal_2625, SubCellInst_SboxInst_13_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_U3 ( .a ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, new_AGEMA_signal_2829, SubCellInst_SboxInst_14_YY_1_}), .b ({new_AGEMA_signal_2930, new_AGEMA_signal_2929, new_AGEMA_signal_2928, AddRoundConstantOutput[59]}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_U2 ( .a ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, new_AGEMA_signal_2637, SubCellInst_SboxInst_14_YY_0_}), .b ({new_AGEMA_signal_2822, new_AGEMA_signal_2821, new_AGEMA_signal_2820, AddRoundConstantOutput[58]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_AND1_U1 ( .a ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, SubCellInst_SboxInst_14_n3}), .b ({new_AGEMA_signal_2288, new_AGEMA_signal_2287, new_AGEMA_signal_2286, SubCellInst_SboxInst_14_Q1}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, new_AGEMA_signal_2442, SubCellInst_SboxInst_14_T0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_XOR2_U1 ( .a ({new_AGEMA_signal_5144, new_AGEMA_signal_5142, new_AGEMA_signal_5140, new_AGEMA_signal_5138}), .b ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, new_AGEMA_signal_2442, SubCellInst_SboxInst_14_T0}), .c ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, new_AGEMA_signal_2628, SubCellInst_SboxInst_14_Q2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_AND3_U1 ( .a ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, SubCellInst_SboxInst_14_n3}), .b ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, new_AGEMA_signal_2289, SubCellInst_SboxInst_14_Q4}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, new_AGEMA_signal_2445, SubCellInst_SboxInst_14_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_XOR7_U1 ( .a ({new_AGEMA_signal_5152, new_AGEMA_signal_5150, new_AGEMA_signal_5148, new_AGEMA_signal_5146}), .b ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, new_AGEMA_signal_2445, SubCellInst_SboxInst_14_T2}), .c ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, new_AGEMA_signal_2631, SubCellInst_SboxInst_14_Q7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_XOR11_U1 ( .a ({new_AGEMA_signal_5160, new_AGEMA_signal_5158, new_AGEMA_signal_5156, new_AGEMA_signal_5154}), .b ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, new_AGEMA_signal_2442, SubCellInst_SboxInst_14_T0}), .c ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, new_AGEMA_signal_2634, SubCellInst_SboxInst_14_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_XOR12_U1 ( .a ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, new_AGEMA_signal_2634, SubCellInst_SboxInst_14_L3}), .b ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, new_AGEMA_signal_2445, SubCellInst_SboxInst_14_T2}), .c ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, new_AGEMA_signal_2829, SubCellInst_SboxInst_14_YY_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_XOR13_U1 ( .a ({new_AGEMA_signal_5168, new_AGEMA_signal_5166, new_AGEMA_signal_5164, new_AGEMA_signal_5162}), .b ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, new_AGEMA_signal_2445, SubCellInst_SboxInst_14_T2}), .c ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, new_AGEMA_signal_2637, SubCellInst_SboxInst_14_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_U3 ( .a ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, new_AGEMA_signal_2841, SubCellInst_SboxInst_15_YY_1_}), .b ({new_AGEMA_signal_2936, new_AGEMA_signal_2935, new_AGEMA_signal_2934, SubCellOutput[63]}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_U2 ( .a ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, new_AGEMA_signal_2649, SubCellInst_SboxInst_15_YY_0_}), .b ({new_AGEMA_signal_2834, new_AGEMA_signal_2833, new_AGEMA_signal_2832, SubCellOutput[62]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_AND1_U1 ( .a ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, new_AGEMA_signal_1437, SubCellInst_SboxInst_15_n3}), .b ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, new_AGEMA_signal_2304, SubCellInst_SboxInst_15_Q1}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, new_AGEMA_signal_2451, SubCellInst_SboxInst_15_T0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_XOR2_U1 ( .a ({new_AGEMA_signal_5176, new_AGEMA_signal_5174, new_AGEMA_signal_5172, new_AGEMA_signal_5170}), .b ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, new_AGEMA_signal_2451, SubCellInst_SboxInst_15_T0}), .c ({new_AGEMA_signal_2642, new_AGEMA_signal_2641, new_AGEMA_signal_2640, SubCellInst_SboxInst_15_Q2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_AND3_U1 ( .a ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, new_AGEMA_signal_1437, SubCellInst_SboxInst_15_n3}), .b ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, new_AGEMA_signal_2307, SubCellInst_SboxInst_15_Q4}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, new_AGEMA_signal_2454, SubCellInst_SboxInst_15_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_XOR7_U1 ( .a ({new_AGEMA_signal_5184, new_AGEMA_signal_5182, new_AGEMA_signal_5180, new_AGEMA_signal_5178}), .b ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, new_AGEMA_signal_2454, SubCellInst_SboxInst_15_T2}), .c ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, new_AGEMA_signal_2643, SubCellInst_SboxInst_15_Q7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_XOR11_U1 ( .a ({new_AGEMA_signal_5192, new_AGEMA_signal_5190, new_AGEMA_signal_5188, new_AGEMA_signal_5186}), .b ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, new_AGEMA_signal_2451, SubCellInst_SboxInst_15_T0}), .c ({new_AGEMA_signal_2648, new_AGEMA_signal_2647, new_AGEMA_signal_2646, SubCellInst_SboxInst_15_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_XOR12_U1 ( .a ({new_AGEMA_signal_2648, new_AGEMA_signal_2647, new_AGEMA_signal_2646, SubCellInst_SboxInst_15_L3}), .b ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, new_AGEMA_signal_2454, SubCellInst_SboxInst_15_T2}), .c ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, new_AGEMA_signal_2841, SubCellInst_SboxInst_15_YY_1_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_XOR13_U1 ( .a ({new_AGEMA_signal_5200, new_AGEMA_signal_5198, new_AGEMA_signal_5196, new_AGEMA_signal_5194}), .b ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, new_AGEMA_signal_2454, SubCellInst_SboxInst_15_T2}), .c ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, new_AGEMA_signal_2649, SubCellInst_SboxInst_15_YY_0_}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2942, new_AGEMA_signal_2941, new_AGEMA_signal_2940, AddConstXOR_AddConstXOR_XORInst_0_2_n1}), .b ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_5202}), .c ({new_AGEMA_signal_3074, new_AGEMA_signal_3073, new_AGEMA_signal_3072, AddRoundConstantOutput[62]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2834, new_AGEMA_signal_2833, new_AGEMA_signal_2832, SubCellOutput[62]}), .c ({new_AGEMA_signal_2942, new_AGEMA_signal_2941, new_AGEMA_signal_2940, AddConstXOR_AddConstXOR_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, new_AGEMA_signal_3075, AddConstXOR_AddConstXOR_XORInst_0_3_n1}), .b ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_5204}), .c ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, new_AGEMA_signal_3201, AddRoundConstantOutput[63]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2936, new_AGEMA_signal_2935, new_AGEMA_signal_2934, SubCellOutput[63]}), .c ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, new_AGEMA_signal_3075, AddConstXOR_AddConstXOR_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, new_AGEMA_signal_2943, AddConstXOR_AddConstXOR_XORInst_1_2_n1}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .c ({new_AGEMA_signal_3080, new_AGEMA_signal_3079, new_AGEMA_signal_3078, AddRoundConstantOutput[46]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2786, new_AGEMA_signal_2785, new_AGEMA_signal_2784, SubCellOutput[46]}), .c ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, new_AGEMA_signal_2943, AddConstXOR_AddConstXOR_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_3083, new_AGEMA_signal_3082, new_AGEMA_signal_3081, AddConstXOR_AddConstXOR_XORInst_1_3_n1}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .c ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, new_AGEMA_signal_3207, AddRoundConstantOutput[47]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2912, new_AGEMA_signal_2911, new_AGEMA_signal_2910, SubCellOutput[47]}), .c ({new_AGEMA_signal_3083, new_AGEMA_signal_3082, new_AGEMA_signal_3081, AddConstXOR_AddConstXOR_XORInst_1_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2948, new_AGEMA_signal_2947, new_AGEMA_signal_2946, AddRoundTweakeyXOR_XORInst_0_2_n1}), .b ({new_AGEMA_signal_5212, new_AGEMA_signal_5210, new_AGEMA_signal_5208, new_AGEMA_signal_5206}), .c ({new_AGEMA_signal_3086, new_AGEMA_signal_3085, new_AGEMA_signal_3084, ShiftRowsOutput[46]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2750, new_AGEMA_signal_2749, new_AGEMA_signal_2748, AddRoundConstantOutput[34]}), .c ({new_AGEMA_signal_2948, new_AGEMA_signal_2947, new_AGEMA_signal_2946, AddRoundTweakeyXOR_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, new_AGEMA_signal_3087, AddRoundTweakeyXOR_XORInst_0_3_n1}), .b ({new_AGEMA_signal_5220, new_AGEMA_signal_5218, new_AGEMA_signal_5216, new_AGEMA_signal_5214}), .c ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, new_AGEMA_signal_3213, ShiftRowsOutput[47]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2894, new_AGEMA_signal_2893, new_AGEMA_signal_2892, AddRoundConstantOutput[35]}), .c ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, new_AGEMA_signal_3087, AddRoundTweakeyXOR_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, new_AGEMA_signal_2949, AddRoundTweakeyXOR_XORInst_1_2_n1}), .b ({new_AGEMA_signal_5228, new_AGEMA_signal_5226, new_AGEMA_signal_5224, new_AGEMA_signal_5222}), .c ({new_AGEMA_signal_3092, new_AGEMA_signal_3091, new_AGEMA_signal_3090, ShiftRowsOutput[34]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2762, new_AGEMA_signal_2761, new_AGEMA_signal_2760, AddRoundConstantOutput[38]}), .c ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, new_AGEMA_signal_2949, AddRoundTweakeyXOR_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, new_AGEMA_signal_3093, AddRoundTweakeyXOR_XORInst_1_3_n1}), .b ({new_AGEMA_signal_5236, new_AGEMA_signal_5234, new_AGEMA_signal_5232, new_AGEMA_signal_5230}), .c ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, new_AGEMA_signal_3219, ShiftRowsOutput[35]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2900, new_AGEMA_signal_2899, new_AGEMA_signal_2898, AddRoundConstantOutput[39]}), .c ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, new_AGEMA_signal_3093, AddRoundTweakeyXOR_XORInst_1_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_2954, new_AGEMA_signal_2953, new_AGEMA_signal_2952, AddRoundTweakeyXOR_XORInst_2_2_n1}), .b ({new_AGEMA_signal_5244, new_AGEMA_signal_5242, new_AGEMA_signal_5240, new_AGEMA_signal_5238}), .c ({new_AGEMA_signal_3098, new_AGEMA_signal_3097, new_AGEMA_signal_3096, ShiftRowsOutput[38]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2774, new_AGEMA_signal_2773, new_AGEMA_signal_2772, AddRoundConstantOutput[42]}), .c ({new_AGEMA_signal_2954, new_AGEMA_signal_2953, new_AGEMA_signal_2952, AddRoundTweakeyXOR_XORInst_2_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, new_AGEMA_signal_3099, AddRoundTweakeyXOR_XORInst_2_3_n1}), .b ({new_AGEMA_signal_5252, new_AGEMA_signal_5250, new_AGEMA_signal_5248, new_AGEMA_signal_5246}), .c ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, new_AGEMA_signal_3225, ShiftRowsOutput[39]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2906, new_AGEMA_signal_2905, new_AGEMA_signal_2904, AddRoundConstantOutput[43]}), .c ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, new_AGEMA_signal_3099, AddRoundTweakeyXOR_XORInst_2_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_3230, new_AGEMA_signal_3229, new_AGEMA_signal_3228, AddRoundTweakeyXOR_XORInst_3_2_n1}), .b ({new_AGEMA_signal_5260, new_AGEMA_signal_5258, new_AGEMA_signal_5256, new_AGEMA_signal_5254}), .c ({new_AGEMA_signal_3344, new_AGEMA_signal_3343, new_AGEMA_signal_3342, ShiftRowsOutput[42]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3080, new_AGEMA_signal_3079, new_AGEMA_signal_3078, AddRoundConstantOutput[46]}), .c ({new_AGEMA_signal_3230, new_AGEMA_signal_3229, new_AGEMA_signal_3228, AddRoundTweakeyXOR_XORInst_3_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, new_AGEMA_signal_3345, AddRoundTweakeyXOR_XORInst_3_3_n1}), .b ({new_AGEMA_signal_5268, new_AGEMA_signal_5266, new_AGEMA_signal_5264, new_AGEMA_signal_5262}), .c ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, new_AGEMA_signal_3531, ShiftRowsOutput[43]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, new_AGEMA_signal_3207, AddRoundConstantOutput[47]}), .c ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, new_AGEMA_signal_3345, AddRoundTweakeyXOR_XORInst_3_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_4_2_U2 ( .a ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, new_AGEMA_signal_2955, AddRoundTweakeyXOR_XORInst_4_2_n1}), .b ({new_AGEMA_signal_5276, new_AGEMA_signal_5274, new_AGEMA_signal_5272, new_AGEMA_signal_5270}), .c ({new_AGEMA_signal_3104, new_AGEMA_signal_3103, new_AGEMA_signal_3102, MCOutput[34]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_4_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2798, new_AGEMA_signal_2797, new_AGEMA_signal_2796, AddRoundConstantOutput[50]}), .c ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, new_AGEMA_signal_2955, AddRoundTweakeyXOR_XORInst_4_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_4_3_U2 ( .a ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, new_AGEMA_signal_3105, AddRoundTweakeyXOR_XORInst_4_3_n1}), .b ({new_AGEMA_signal_5284, new_AGEMA_signal_5282, new_AGEMA_signal_5280, new_AGEMA_signal_5278}), .c ({new_AGEMA_signal_3236, new_AGEMA_signal_3235, new_AGEMA_signal_3234, MCOutput[35]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_4_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2918, new_AGEMA_signal_2917, new_AGEMA_signal_2916, AddRoundConstantOutput[51]}), .c ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, new_AGEMA_signal_3105, AddRoundTweakeyXOR_XORInst_4_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_5_2_U2 ( .a ({new_AGEMA_signal_2960, new_AGEMA_signal_2959, new_AGEMA_signal_2958, AddRoundTweakeyXOR_XORInst_5_2_n1}), .b ({new_AGEMA_signal_5292, new_AGEMA_signal_5290, new_AGEMA_signal_5288, new_AGEMA_signal_5286}), .c ({new_AGEMA_signal_3110, new_AGEMA_signal_3109, new_AGEMA_signal_3108, MCOutput[38]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_5_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2810, new_AGEMA_signal_2809, new_AGEMA_signal_2808, AddRoundConstantOutput[54]}), .c ({new_AGEMA_signal_2960, new_AGEMA_signal_2959, new_AGEMA_signal_2958, AddRoundTweakeyXOR_XORInst_5_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_5_3_U2 ( .a ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, new_AGEMA_signal_3111, AddRoundTweakeyXOR_XORInst_5_3_n1}), .b ({new_AGEMA_signal_5300, new_AGEMA_signal_5298, new_AGEMA_signal_5296, new_AGEMA_signal_5294}), .c ({new_AGEMA_signal_3242, new_AGEMA_signal_3241, new_AGEMA_signal_3240, MCOutput[39]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_5_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2924, new_AGEMA_signal_2923, new_AGEMA_signal_2922, AddRoundConstantOutput[55]}), .c ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, new_AGEMA_signal_3111, AddRoundTweakeyXOR_XORInst_5_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_6_2_U2 ( .a ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, new_AGEMA_signal_2961, AddRoundTweakeyXOR_XORInst_6_2_n1}), .b ({new_AGEMA_signal_5308, new_AGEMA_signal_5306, new_AGEMA_signal_5304, new_AGEMA_signal_5302}), .c ({new_AGEMA_signal_3116, new_AGEMA_signal_3115, new_AGEMA_signal_3114, MCOutput[42]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_6_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2822, new_AGEMA_signal_2821, new_AGEMA_signal_2820, AddRoundConstantOutput[58]}), .c ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, new_AGEMA_signal_2961, AddRoundTweakeyXOR_XORInst_6_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_6_3_U2 ( .a ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, new_AGEMA_signal_3117, AddRoundTweakeyXOR_XORInst_6_3_n1}), .b ({new_AGEMA_signal_5316, new_AGEMA_signal_5314, new_AGEMA_signal_5312, new_AGEMA_signal_5310}), .c ({new_AGEMA_signal_3248, new_AGEMA_signal_3247, new_AGEMA_signal_3246, MCOutput[43]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_6_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2930, new_AGEMA_signal_2929, new_AGEMA_signal_2928, AddRoundConstantOutput[59]}), .c ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, new_AGEMA_signal_3117, AddRoundTweakeyXOR_XORInst_6_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_7_2_U2 ( .a ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, new_AGEMA_signal_3249, AddRoundTweakeyXOR_XORInst_7_2_n1}), .b ({new_AGEMA_signal_5324, new_AGEMA_signal_5322, new_AGEMA_signal_5320, new_AGEMA_signal_5318}), .c ({new_AGEMA_signal_3368, new_AGEMA_signal_3367, new_AGEMA_signal_3366, MCOutput[46]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_7_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3074, new_AGEMA_signal_3073, new_AGEMA_signal_3072, AddRoundConstantOutput[62]}), .c ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, new_AGEMA_signal_3249, AddRoundTweakeyXOR_XORInst_7_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_7_3_U2 ( .a ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, new_AGEMA_signal_3369, AddRoundTweakeyXOR_XORInst_7_3_n1}), .b ({new_AGEMA_signal_5332, new_AGEMA_signal_5330, new_AGEMA_signal_5328, new_AGEMA_signal_5326}), .c ({new_AGEMA_signal_3548, new_AGEMA_signal_3547, new_AGEMA_signal_3546, MCOutput[47]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_7_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, new_AGEMA_signal_3201, AddRoundConstantOutput[63]}), .c ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, new_AGEMA_signal_3369, AddRoundTweakeyXOR_XORInst_7_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_0_2_U3 ( .a ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, new_AGEMA_signal_3255, MCInst_MCR0_XORInst_0_2_n2}), .b ({new_AGEMA_signal_2966, new_AGEMA_signal_2965, new_AGEMA_signal_2964, MCInst_MCR0_XORInst_0_2_n1}), .c ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, new_AGEMA_signal_3375, MCOutput[50]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, new_AGEMA_signal_2724, ShiftRowsOutput[18]}), .b ({new_AGEMA_signal_2690, new_AGEMA_signal_2689, new_AGEMA_signal_2688, ShiftRowsOutput[2]}), .c ({new_AGEMA_signal_2966, new_AGEMA_signal_2965, new_AGEMA_signal_2964, MCInst_MCR0_XORInst_0_2_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3104, new_AGEMA_signal_3103, new_AGEMA_signal_3102, MCOutput[34]}), .c ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, new_AGEMA_signal_3255, MCInst_MCR0_XORInst_0_2_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_0_3_U3 ( .a ({new_AGEMA_signal_3380, new_AGEMA_signal_3379, new_AGEMA_signal_3378, MCInst_MCR0_XORInst_0_3_n2}), .b ({new_AGEMA_signal_3122, new_AGEMA_signal_3121, new_AGEMA_signal_3120, MCInst_MCR0_XORInst_0_3_n1}), .c ({new_AGEMA_signal_3554, new_AGEMA_signal_3553, new_AGEMA_signal_3552, MCOutput[51]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2882, new_AGEMA_signal_2881, new_AGEMA_signal_2880, ShiftRowsOutput[19]}), .b ({new_AGEMA_signal_2864, new_AGEMA_signal_2863, new_AGEMA_signal_2862, ShiftRowsOutput[3]}), .c ({new_AGEMA_signal_3122, new_AGEMA_signal_3121, new_AGEMA_signal_3120, MCInst_MCR0_XORInst_0_3_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3236, new_AGEMA_signal_3235, new_AGEMA_signal_3234, MCOutput[35]}), .c ({new_AGEMA_signal_3380, new_AGEMA_signal_3379, new_AGEMA_signal_3378, MCInst_MCR0_XORInst_0_3_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_1_2_U3 ( .a ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, new_AGEMA_signal_3261, MCInst_MCR0_XORInst_1_2_n2}), .b ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, new_AGEMA_signal_2967, MCInst_MCR0_XORInst_1_2_n1}), .c ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, new_AGEMA_signal_3381, MCOutput[54]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2738, new_AGEMA_signal_2737, new_AGEMA_signal_2736, ShiftRowsOutput[22]}), .b ({new_AGEMA_signal_2654, new_AGEMA_signal_2653, new_AGEMA_signal_2652, ShiftRowsOutput[6]}), .c ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, new_AGEMA_signal_2967, MCInst_MCR0_XORInst_1_2_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3110, new_AGEMA_signal_3109, new_AGEMA_signal_3108, MCOutput[38]}), .c ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, new_AGEMA_signal_3261, MCInst_MCR0_XORInst_1_2_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_1_3_U3 ( .a ({new_AGEMA_signal_3386, new_AGEMA_signal_3385, new_AGEMA_signal_3384, MCInst_MCR0_XORInst_1_3_n2}), .b ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, new_AGEMA_signal_3123, MCInst_MCR0_XORInst_1_3_n1}), .c ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, new_AGEMA_signal_3561, MCOutput[55]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2888, new_AGEMA_signal_2887, new_AGEMA_signal_2886, ShiftRowsOutput[23]}), .b ({new_AGEMA_signal_2846, new_AGEMA_signal_2845, new_AGEMA_signal_2844, ShiftRowsOutput[7]}), .c ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, new_AGEMA_signal_3123, MCInst_MCR0_XORInst_1_3_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3242, new_AGEMA_signal_3241, new_AGEMA_signal_3240, MCOutput[39]}), .c ({new_AGEMA_signal_3386, new_AGEMA_signal_3385, new_AGEMA_signal_3384, MCInst_MCR0_XORInst_1_3_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_2_2_U3 ( .a ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, new_AGEMA_signal_3267, MCInst_MCR0_XORInst_2_2_n2}), .b ({new_AGEMA_signal_2972, new_AGEMA_signal_2971, new_AGEMA_signal_2970, MCInst_MCR0_XORInst_2_2_n1}), .c ({new_AGEMA_signal_3392, new_AGEMA_signal_3391, new_AGEMA_signal_3390, MCOutput[58]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_2702, new_AGEMA_signal_2701, new_AGEMA_signal_2700, ShiftRowsOutput[26]}), .b ({new_AGEMA_signal_2666, new_AGEMA_signal_2665, new_AGEMA_signal_2664, ShiftRowsOutput[10]}), .c ({new_AGEMA_signal_2972, new_AGEMA_signal_2971, new_AGEMA_signal_2970, MCInst_MCR0_XORInst_2_2_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3116, new_AGEMA_signal_3115, new_AGEMA_signal_3114, MCOutput[42]}), .c ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, new_AGEMA_signal_3267, MCInst_MCR0_XORInst_2_2_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_2_3_U3 ( .a ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, new_AGEMA_signal_3393, MCInst_MCR0_XORInst_2_3_n2}), .b ({new_AGEMA_signal_3128, new_AGEMA_signal_3127, new_AGEMA_signal_3126, MCInst_MCR0_XORInst_2_3_n1}), .c ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, new_AGEMA_signal_3567, MCOutput[59]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_2870, new_AGEMA_signal_2869, new_AGEMA_signal_2868, ShiftRowsOutput[27]}), .b ({new_AGEMA_signal_2852, new_AGEMA_signal_2851, new_AGEMA_signal_2850, ShiftRowsOutput[11]}), .c ({new_AGEMA_signal_3128, new_AGEMA_signal_3127, new_AGEMA_signal_3126, MCInst_MCR0_XORInst_2_3_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3248, new_AGEMA_signal_3247, new_AGEMA_signal_3246, MCOutput[43]}), .c ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, new_AGEMA_signal_3393, MCInst_MCR0_XORInst_2_3_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_3_2_U3 ( .a ({new_AGEMA_signal_3572, new_AGEMA_signal_3571, new_AGEMA_signal_3570, MCInst_MCR0_XORInst_3_2_n2}), .b ({new_AGEMA_signal_2975, new_AGEMA_signal_2974, new_AGEMA_signal_2973, MCInst_MCR0_XORInst_3_2_n1}), .c ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, new_AGEMA_signal_3723, MCOutput[62]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, new_AGEMA_signal_2712, ShiftRowsOutput[30]}), .b ({new_AGEMA_signal_2678, new_AGEMA_signal_2677, new_AGEMA_signal_2676, ShiftRowsOutput[14]}), .c ({new_AGEMA_signal_2975, new_AGEMA_signal_2974, new_AGEMA_signal_2973, MCInst_MCR0_XORInst_3_2_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3368, new_AGEMA_signal_3367, new_AGEMA_signal_3366, MCOutput[46]}), .c ({new_AGEMA_signal_3572, new_AGEMA_signal_3571, new_AGEMA_signal_3570, MCInst_MCR0_XORInst_3_2_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_3_3_U3 ( .a ({new_AGEMA_signal_3728, new_AGEMA_signal_3727, new_AGEMA_signal_3726, MCInst_MCR0_XORInst_3_3_n2}), .b ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, new_AGEMA_signal_3129, MCInst_MCR0_XORInst_3_3_n1}), .c ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, new_AGEMA_signal_3873, MCOutput[63]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_2876, new_AGEMA_signal_2875, new_AGEMA_signal_2874, ShiftRowsOutput[31]}), .b ({new_AGEMA_signal_2858, new_AGEMA_signal_2857, new_AGEMA_signal_2856, ShiftRowsOutput[15]}), .c ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, new_AGEMA_signal_3129, MCInst_MCR0_XORInst_3_3_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3548, new_AGEMA_signal_3547, new_AGEMA_signal_3546, MCOutput[47]}), .c ({new_AGEMA_signal_3728, new_AGEMA_signal_3727, new_AGEMA_signal_3726, MCInst_MCR0_XORInst_3_3_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, new_AGEMA_signal_3273, MCInst_MCR2_XORInst_0_2_n1}), .b ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, new_AGEMA_signal_2724, ShiftRowsOutput[18]}), .c ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, new_AGEMA_signal_3399, MCOutput[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3092, new_AGEMA_signal_3091, new_AGEMA_signal_3090, ShiftRowsOutput[34]}), .c ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, new_AGEMA_signal_3273, MCInst_MCR2_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_3404, new_AGEMA_signal_3403, new_AGEMA_signal_3402, MCInst_MCR2_XORInst_0_3_n1}), .b ({new_AGEMA_signal_2882, new_AGEMA_signal_2881, new_AGEMA_signal_2880, ShiftRowsOutput[19]}), .c ({new_AGEMA_signal_3578, new_AGEMA_signal_3577, new_AGEMA_signal_3576, MCOutput[19]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, new_AGEMA_signal_3219, ShiftRowsOutput[35]}), .c ({new_AGEMA_signal_3404, new_AGEMA_signal_3403, new_AGEMA_signal_3402, MCInst_MCR2_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_3278, new_AGEMA_signal_3277, new_AGEMA_signal_3276, MCInst_MCR2_XORInst_1_2_n1}), .b ({new_AGEMA_signal_2738, new_AGEMA_signal_2737, new_AGEMA_signal_2736, ShiftRowsOutput[22]}), .c ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, new_AGEMA_signal_3405, MCOutput[22]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3098, new_AGEMA_signal_3097, new_AGEMA_signal_3096, ShiftRowsOutput[38]}), .c ({new_AGEMA_signal_3278, new_AGEMA_signal_3277, new_AGEMA_signal_3276, MCInst_MCR2_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_3410, new_AGEMA_signal_3409, new_AGEMA_signal_3408, MCInst_MCR2_XORInst_1_3_n1}), .b ({new_AGEMA_signal_2888, new_AGEMA_signal_2887, new_AGEMA_signal_2886, ShiftRowsOutput[23]}), .c ({new_AGEMA_signal_3584, new_AGEMA_signal_3583, new_AGEMA_signal_3582, MCOutput[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, new_AGEMA_signal_3225, ShiftRowsOutput[39]}), .c ({new_AGEMA_signal_3410, new_AGEMA_signal_3409, new_AGEMA_signal_3408, MCInst_MCR2_XORInst_1_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, new_AGEMA_signal_3585, MCInst_MCR2_XORInst_2_2_n1}), .b ({new_AGEMA_signal_2702, new_AGEMA_signal_2701, new_AGEMA_signal_2700, ShiftRowsOutput[26]}), .c ({new_AGEMA_signal_3743, new_AGEMA_signal_3742, new_AGEMA_signal_3741, MCOutput[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3344, new_AGEMA_signal_3343, new_AGEMA_signal_3342, ShiftRowsOutput[42]}), .c ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, new_AGEMA_signal_3585, MCInst_MCR2_XORInst_2_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_3746, new_AGEMA_signal_3745, new_AGEMA_signal_3744, MCInst_MCR2_XORInst_2_3_n1}), .b ({new_AGEMA_signal_2870, new_AGEMA_signal_2869, new_AGEMA_signal_2868, ShiftRowsOutput[27]}), .c ({new_AGEMA_signal_3887, new_AGEMA_signal_3886, new_AGEMA_signal_3885, MCOutput[27]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, new_AGEMA_signal_3531, ShiftRowsOutput[43]}), .c ({new_AGEMA_signal_3746, new_AGEMA_signal_3745, new_AGEMA_signal_3744, MCInst_MCR2_XORInst_2_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, new_AGEMA_signal_3279, MCInst_MCR2_XORInst_3_2_n1}), .b ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, new_AGEMA_signal_2712, ShiftRowsOutput[30]}), .c ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, new_AGEMA_signal_3411, MCOutput[30]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3086, new_AGEMA_signal_3085, new_AGEMA_signal_3084, ShiftRowsOutput[46]}), .c ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, new_AGEMA_signal_3279, MCInst_MCR2_XORInst_3_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_3416, new_AGEMA_signal_3415, new_AGEMA_signal_3414, MCInst_MCR2_XORInst_3_3_n1}), .b ({new_AGEMA_signal_2876, new_AGEMA_signal_2875, new_AGEMA_signal_2874, ShiftRowsOutput[31]}), .c ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, new_AGEMA_signal_3591, MCOutput[31]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, new_AGEMA_signal_3213, ShiftRowsOutput[47]}), .c ({new_AGEMA_signal_3416, new_AGEMA_signal_3415, new_AGEMA_signal_3414, MCInst_MCR2_XORInst_3_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_3284, new_AGEMA_signal_3283, new_AGEMA_signal_3282, MCInst_MCR3_XORInst_0_2_n1}), .b ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, new_AGEMA_signal_2724, ShiftRowsOutput[18]}), .c ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, new_AGEMA_signal_3417, MCOutput[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3104, new_AGEMA_signal_3103, new_AGEMA_signal_3102, MCOutput[34]}), .c ({new_AGEMA_signal_3284, new_AGEMA_signal_3283, new_AGEMA_signal_3282, MCInst_MCR3_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_3422, new_AGEMA_signal_3421, new_AGEMA_signal_3420, MCInst_MCR3_XORInst_0_3_n1}), .b ({new_AGEMA_signal_2882, new_AGEMA_signal_2881, new_AGEMA_signal_2880, ShiftRowsOutput[19]}), .c ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, new_AGEMA_signal_3597, MCOutput[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3236, new_AGEMA_signal_3235, new_AGEMA_signal_3234, MCOutput[35]}), .c ({new_AGEMA_signal_3422, new_AGEMA_signal_3421, new_AGEMA_signal_3420, MCInst_MCR3_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, new_AGEMA_signal_3285, MCInst_MCR3_XORInst_1_2_n1}), .b ({new_AGEMA_signal_2738, new_AGEMA_signal_2737, new_AGEMA_signal_2736, ShiftRowsOutput[22]}), .c ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, new_AGEMA_signal_3423, MCOutput[6]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3110, new_AGEMA_signal_3109, new_AGEMA_signal_3108, MCOutput[38]}), .c ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, new_AGEMA_signal_3285, MCInst_MCR3_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_3428, new_AGEMA_signal_3427, new_AGEMA_signal_3426, MCInst_MCR3_XORInst_1_3_n1}), .b ({new_AGEMA_signal_2888, new_AGEMA_signal_2887, new_AGEMA_signal_2886, ShiftRowsOutput[23]}), .c ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, new_AGEMA_signal_3603, MCOutput[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3242, new_AGEMA_signal_3241, new_AGEMA_signal_3240, MCOutput[39]}), .c ({new_AGEMA_signal_3428, new_AGEMA_signal_3427, new_AGEMA_signal_3426, MCInst_MCR3_XORInst_1_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_3290, new_AGEMA_signal_3289, new_AGEMA_signal_3288, MCInst_MCR3_XORInst_2_2_n1}), .b ({new_AGEMA_signal_2702, new_AGEMA_signal_2701, new_AGEMA_signal_2700, ShiftRowsOutput[26]}), .c ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, new_AGEMA_signal_3429, MCOutput[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3116, new_AGEMA_signal_3115, new_AGEMA_signal_3114, MCOutput[42]}), .c ({new_AGEMA_signal_3290, new_AGEMA_signal_3289, new_AGEMA_signal_3288, MCInst_MCR3_XORInst_2_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_3434, new_AGEMA_signal_3433, new_AGEMA_signal_3432, MCInst_MCR3_XORInst_2_3_n1}), .b ({new_AGEMA_signal_2870, new_AGEMA_signal_2869, new_AGEMA_signal_2868, ShiftRowsOutput[27]}), .c ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, new_AGEMA_signal_3609, MCOutput[11]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3248, new_AGEMA_signal_3247, new_AGEMA_signal_3246, MCOutput[43]}), .c ({new_AGEMA_signal_3434, new_AGEMA_signal_3433, new_AGEMA_signal_3432, MCInst_MCR3_XORInst_2_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_3614, new_AGEMA_signal_3613, new_AGEMA_signal_3612, MCInst_MCR3_XORInst_3_2_n1}), .b ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, new_AGEMA_signal_2712, ShiftRowsOutput[30]}), .c ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, new_AGEMA_signal_3771, MCOutput[14]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3368, new_AGEMA_signal_3367, new_AGEMA_signal_3366, MCOutput[46]}), .c ({new_AGEMA_signal_3614, new_AGEMA_signal_3613, new_AGEMA_signal_3612, MCInst_MCR3_XORInst_3_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_3776, new_AGEMA_signal_3775, new_AGEMA_signal_3774, MCInst_MCR3_XORInst_3_3_n1}), .b ({new_AGEMA_signal_2876, new_AGEMA_signal_2875, new_AGEMA_signal_2874, ShiftRowsOutput[31]}), .c ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, new_AGEMA_signal_3903, MCOutput[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3548, new_AGEMA_signal_3547, new_AGEMA_signal_3546, MCOutput[47]}), .c ({new_AGEMA_signal_3776, new_AGEMA_signal_3775, new_AGEMA_signal_3774, MCInst_MCR3_XORInst_3_3_n1}) ) ;
    buf_clk new_AGEMA_reg_buffer_1001 ( .C (clk), .D (new_AGEMA_signal_4431), .Q (new_AGEMA_signal_4432) ) ;
    buf_clk new_AGEMA_reg_buffer_1003 ( .C (clk), .D (new_AGEMA_signal_4433), .Q (new_AGEMA_signal_4434) ) ;
    buf_clk new_AGEMA_reg_buffer_1005 ( .C (clk), .D (new_AGEMA_signal_4435), .Q (new_AGEMA_signal_4436) ) ;
    buf_clk new_AGEMA_reg_buffer_1007 ( .C (clk), .D (new_AGEMA_signal_4437), .Q (new_AGEMA_signal_4438) ) ;
    buf_clk new_AGEMA_reg_buffer_1009 ( .C (clk), .D (new_AGEMA_signal_4439), .Q (new_AGEMA_signal_4440) ) ;
    buf_clk new_AGEMA_reg_buffer_1011 ( .C (clk), .D (new_AGEMA_signal_4441), .Q (new_AGEMA_signal_4442) ) ;
    buf_clk new_AGEMA_reg_buffer_1013 ( .C (clk), .D (new_AGEMA_signal_4443), .Q (new_AGEMA_signal_4444) ) ;
    buf_clk new_AGEMA_reg_buffer_1015 ( .C (clk), .D (new_AGEMA_signal_4445), .Q (new_AGEMA_signal_4446) ) ;
    buf_clk new_AGEMA_reg_buffer_1017 ( .C (clk), .D (new_AGEMA_signal_4447), .Q (new_AGEMA_signal_4448) ) ;
    buf_clk new_AGEMA_reg_buffer_1019 ( .C (clk), .D (new_AGEMA_signal_4449), .Q (new_AGEMA_signal_4450) ) ;
    buf_clk new_AGEMA_reg_buffer_1021 ( .C (clk), .D (new_AGEMA_signal_4451), .Q (new_AGEMA_signal_4452) ) ;
    buf_clk new_AGEMA_reg_buffer_1023 ( .C (clk), .D (new_AGEMA_signal_4453), .Q (new_AGEMA_signal_4454) ) ;
    buf_clk new_AGEMA_reg_buffer_1025 ( .C (clk), .D (new_AGEMA_signal_4455), .Q (new_AGEMA_signal_4456) ) ;
    buf_clk new_AGEMA_reg_buffer_1027 ( .C (clk), .D (new_AGEMA_signal_4457), .Q (new_AGEMA_signal_4458) ) ;
    buf_clk new_AGEMA_reg_buffer_1029 ( .C (clk), .D (new_AGEMA_signal_4459), .Q (new_AGEMA_signal_4460) ) ;
    buf_clk new_AGEMA_reg_buffer_1031 ( .C (clk), .D (new_AGEMA_signal_4461), .Q (new_AGEMA_signal_4462) ) ;
    buf_clk new_AGEMA_reg_buffer_1033 ( .C (clk), .D (new_AGEMA_signal_4463), .Q (new_AGEMA_signal_4464) ) ;
    buf_clk new_AGEMA_reg_buffer_1035 ( .C (clk), .D (new_AGEMA_signal_4465), .Q (new_AGEMA_signal_4466) ) ;
    buf_clk new_AGEMA_reg_buffer_1037 ( .C (clk), .D (new_AGEMA_signal_4467), .Q (new_AGEMA_signal_4468) ) ;
    buf_clk new_AGEMA_reg_buffer_1039 ( .C (clk), .D (new_AGEMA_signal_4469), .Q (new_AGEMA_signal_4470) ) ;
    buf_clk new_AGEMA_reg_buffer_1041 ( .C (clk), .D (new_AGEMA_signal_4471), .Q (new_AGEMA_signal_4472) ) ;
    buf_clk new_AGEMA_reg_buffer_1043 ( .C (clk), .D (new_AGEMA_signal_4473), .Q (new_AGEMA_signal_4474) ) ;
    buf_clk new_AGEMA_reg_buffer_1045 ( .C (clk), .D (new_AGEMA_signal_4475), .Q (new_AGEMA_signal_4476) ) ;
    buf_clk new_AGEMA_reg_buffer_1047 ( .C (clk), .D (new_AGEMA_signal_4477), .Q (new_AGEMA_signal_4478) ) ;
    buf_clk new_AGEMA_reg_buffer_1049 ( .C (clk), .D (new_AGEMA_signal_4479), .Q (new_AGEMA_signal_4480) ) ;
    buf_clk new_AGEMA_reg_buffer_1051 ( .C (clk), .D (new_AGEMA_signal_4481), .Q (new_AGEMA_signal_4482) ) ;
    buf_clk new_AGEMA_reg_buffer_1053 ( .C (clk), .D (new_AGEMA_signal_4483), .Q (new_AGEMA_signal_4484) ) ;
    buf_clk new_AGEMA_reg_buffer_1055 ( .C (clk), .D (new_AGEMA_signal_4485), .Q (new_AGEMA_signal_4486) ) ;
    buf_clk new_AGEMA_reg_buffer_1057 ( .C (clk), .D (new_AGEMA_signal_4487), .Q (new_AGEMA_signal_4488) ) ;
    buf_clk new_AGEMA_reg_buffer_1059 ( .C (clk), .D (new_AGEMA_signal_4489), .Q (new_AGEMA_signal_4490) ) ;
    buf_clk new_AGEMA_reg_buffer_1061 ( .C (clk), .D (new_AGEMA_signal_4491), .Q (new_AGEMA_signal_4492) ) ;
    buf_clk new_AGEMA_reg_buffer_1063 ( .C (clk), .D (new_AGEMA_signal_4493), .Q (new_AGEMA_signal_4494) ) ;
    buf_clk new_AGEMA_reg_buffer_1065 ( .C (clk), .D (new_AGEMA_signal_4495), .Q (new_AGEMA_signal_4496) ) ;
    buf_clk new_AGEMA_reg_buffer_1067 ( .C (clk), .D (new_AGEMA_signal_4497), .Q (new_AGEMA_signal_4498) ) ;
    buf_clk new_AGEMA_reg_buffer_1069 ( .C (clk), .D (new_AGEMA_signal_4499), .Q (new_AGEMA_signal_4500) ) ;
    buf_clk new_AGEMA_reg_buffer_1071 ( .C (clk), .D (new_AGEMA_signal_4501), .Q (new_AGEMA_signal_4502) ) ;
    buf_clk new_AGEMA_reg_buffer_1073 ( .C (clk), .D (new_AGEMA_signal_4503), .Q (new_AGEMA_signal_4504) ) ;
    buf_clk new_AGEMA_reg_buffer_1075 ( .C (clk), .D (new_AGEMA_signal_4505), .Q (new_AGEMA_signal_4506) ) ;
    buf_clk new_AGEMA_reg_buffer_1077 ( .C (clk), .D (new_AGEMA_signal_4507), .Q (new_AGEMA_signal_4508) ) ;
    buf_clk new_AGEMA_reg_buffer_1079 ( .C (clk), .D (new_AGEMA_signal_4509), .Q (new_AGEMA_signal_4510) ) ;
    buf_clk new_AGEMA_reg_buffer_1081 ( .C (clk), .D (new_AGEMA_signal_4511), .Q (new_AGEMA_signal_4512) ) ;
    buf_clk new_AGEMA_reg_buffer_1083 ( .C (clk), .D (new_AGEMA_signal_4513), .Q (new_AGEMA_signal_4514) ) ;
    buf_clk new_AGEMA_reg_buffer_1085 ( .C (clk), .D (new_AGEMA_signal_4515), .Q (new_AGEMA_signal_4516) ) ;
    buf_clk new_AGEMA_reg_buffer_1087 ( .C (clk), .D (new_AGEMA_signal_4517), .Q (new_AGEMA_signal_4518) ) ;
    buf_clk new_AGEMA_reg_buffer_1089 ( .C (clk), .D (new_AGEMA_signal_4519), .Q (new_AGEMA_signal_4520) ) ;
    buf_clk new_AGEMA_reg_buffer_1091 ( .C (clk), .D (new_AGEMA_signal_4521), .Q (new_AGEMA_signal_4522) ) ;
    buf_clk new_AGEMA_reg_buffer_1093 ( .C (clk), .D (new_AGEMA_signal_4523), .Q (new_AGEMA_signal_4524) ) ;
    buf_clk new_AGEMA_reg_buffer_1095 ( .C (clk), .D (new_AGEMA_signal_4525), .Q (new_AGEMA_signal_4526) ) ;
    buf_clk new_AGEMA_reg_buffer_1097 ( .C (clk), .D (new_AGEMA_signal_4527), .Q (new_AGEMA_signal_4528) ) ;
    buf_clk new_AGEMA_reg_buffer_1099 ( .C (clk), .D (new_AGEMA_signal_4529), .Q (new_AGEMA_signal_4530) ) ;
    buf_clk new_AGEMA_reg_buffer_1101 ( .C (clk), .D (new_AGEMA_signal_4531), .Q (new_AGEMA_signal_4532) ) ;
    buf_clk new_AGEMA_reg_buffer_1103 ( .C (clk), .D (new_AGEMA_signal_4533), .Q (new_AGEMA_signal_4534) ) ;
    buf_clk new_AGEMA_reg_buffer_1105 ( .C (clk), .D (new_AGEMA_signal_4535), .Q (new_AGEMA_signal_4536) ) ;
    buf_clk new_AGEMA_reg_buffer_1107 ( .C (clk), .D (new_AGEMA_signal_4537), .Q (new_AGEMA_signal_4538) ) ;
    buf_clk new_AGEMA_reg_buffer_1109 ( .C (clk), .D (new_AGEMA_signal_4539), .Q (new_AGEMA_signal_4540) ) ;
    buf_clk new_AGEMA_reg_buffer_1111 ( .C (clk), .D (new_AGEMA_signal_4541), .Q (new_AGEMA_signal_4542) ) ;
    buf_clk new_AGEMA_reg_buffer_1113 ( .C (clk), .D (new_AGEMA_signal_4543), .Q (new_AGEMA_signal_4544) ) ;
    buf_clk new_AGEMA_reg_buffer_1115 ( .C (clk), .D (new_AGEMA_signal_4545), .Q (new_AGEMA_signal_4546) ) ;
    buf_clk new_AGEMA_reg_buffer_1117 ( .C (clk), .D (new_AGEMA_signal_4547), .Q (new_AGEMA_signal_4548) ) ;
    buf_clk new_AGEMA_reg_buffer_1119 ( .C (clk), .D (new_AGEMA_signal_4549), .Q (new_AGEMA_signal_4550) ) ;
    buf_clk new_AGEMA_reg_buffer_1121 ( .C (clk), .D (new_AGEMA_signal_4551), .Q (new_AGEMA_signal_4552) ) ;
    buf_clk new_AGEMA_reg_buffer_1123 ( .C (clk), .D (new_AGEMA_signal_4553), .Q (new_AGEMA_signal_4554) ) ;
    buf_clk new_AGEMA_reg_buffer_1125 ( .C (clk), .D (new_AGEMA_signal_4555), .Q (new_AGEMA_signal_4556) ) ;
    buf_clk new_AGEMA_reg_buffer_1127 ( .C (clk), .D (new_AGEMA_signal_4557), .Q (new_AGEMA_signal_4558) ) ;
    buf_clk new_AGEMA_reg_buffer_1129 ( .C (clk), .D (new_AGEMA_signal_4559), .Q (new_AGEMA_signal_4560) ) ;
    buf_clk new_AGEMA_reg_buffer_1131 ( .C (clk), .D (new_AGEMA_signal_4561), .Q (new_AGEMA_signal_4562) ) ;
    buf_clk new_AGEMA_reg_buffer_1133 ( .C (clk), .D (new_AGEMA_signal_4563), .Q (new_AGEMA_signal_4564) ) ;
    buf_clk new_AGEMA_reg_buffer_1135 ( .C (clk), .D (new_AGEMA_signal_4565), .Q (new_AGEMA_signal_4566) ) ;
    buf_clk new_AGEMA_reg_buffer_1137 ( .C (clk), .D (new_AGEMA_signal_4567), .Q (new_AGEMA_signal_4568) ) ;
    buf_clk new_AGEMA_reg_buffer_1139 ( .C (clk), .D (new_AGEMA_signal_4569), .Q (new_AGEMA_signal_4570) ) ;
    buf_clk new_AGEMA_reg_buffer_1141 ( .C (clk), .D (new_AGEMA_signal_4571), .Q (new_AGEMA_signal_4572) ) ;
    buf_clk new_AGEMA_reg_buffer_1143 ( .C (clk), .D (new_AGEMA_signal_4573), .Q (new_AGEMA_signal_4574) ) ;
    buf_clk new_AGEMA_reg_buffer_1145 ( .C (clk), .D (new_AGEMA_signal_4575), .Q (new_AGEMA_signal_4576) ) ;
    buf_clk new_AGEMA_reg_buffer_1147 ( .C (clk), .D (new_AGEMA_signal_4577), .Q (new_AGEMA_signal_4578) ) ;
    buf_clk new_AGEMA_reg_buffer_1149 ( .C (clk), .D (new_AGEMA_signal_4579), .Q (new_AGEMA_signal_4580) ) ;
    buf_clk new_AGEMA_reg_buffer_1151 ( .C (clk), .D (new_AGEMA_signal_4581), .Q (new_AGEMA_signal_4582) ) ;
    buf_clk new_AGEMA_reg_buffer_1153 ( .C (clk), .D (new_AGEMA_signal_4583), .Q (new_AGEMA_signal_4584) ) ;
    buf_clk new_AGEMA_reg_buffer_1155 ( .C (clk), .D (new_AGEMA_signal_4585), .Q (new_AGEMA_signal_4586) ) ;
    buf_clk new_AGEMA_reg_buffer_1157 ( .C (clk), .D (new_AGEMA_signal_4587), .Q (new_AGEMA_signal_4588) ) ;
    buf_clk new_AGEMA_reg_buffer_1159 ( .C (clk), .D (new_AGEMA_signal_4589), .Q (new_AGEMA_signal_4590) ) ;
    buf_clk new_AGEMA_reg_buffer_1161 ( .C (clk), .D (new_AGEMA_signal_4591), .Q (new_AGEMA_signal_4592) ) ;
    buf_clk new_AGEMA_reg_buffer_1163 ( .C (clk), .D (new_AGEMA_signal_4593), .Q (new_AGEMA_signal_4594) ) ;
    buf_clk new_AGEMA_reg_buffer_1165 ( .C (clk), .D (new_AGEMA_signal_4595), .Q (new_AGEMA_signal_4596) ) ;
    buf_clk new_AGEMA_reg_buffer_1167 ( .C (clk), .D (new_AGEMA_signal_4597), .Q (new_AGEMA_signal_4598) ) ;
    buf_clk new_AGEMA_reg_buffer_1169 ( .C (clk), .D (new_AGEMA_signal_4599), .Q (new_AGEMA_signal_4600) ) ;
    buf_clk new_AGEMA_reg_buffer_1171 ( .C (clk), .D (new_AGEMA_signal_4601), .Q (new_AGEMA_signal_4602) ) ;
    buf_clk new_AGEMA_reg_buffer_1173 ( .C (clk), .D (new_AGEMA_signal_4603), .Q (new_AGEMA_signal_4604) ) ;
    buf_clk new_AGEMA_reg_buffer_1175 ( .C (clk), .D (new_AGEMA_signal_4605), .Q (new_AGEMA_signal_4606) ) ;
    buf_clk new_AGEMA_reg_buffer_1177 ( .C (clk), .D (new_AGEMA_signal_4607), .Q (new_AGEMA_signal_4608) ) ;
    buf_clk new_AGEMA_reg_buffer_1179 ( .C (clk), .D (new_AGEMA_signal_4609), .Q (new_AGEMA_signal_4610) ) ;
    buf_clk new_AGEMA_reg_buffer_1181 ( .C (clk), .D (new_AGEMA_signal_4611), .Q (new_AGEMA_signal_4612) ) ;
    buf_clk new_AGEMA_reg_buffer_1183 ( .C (clk), .D (new_AGEMA_signal_4613), .Q (new_AGEMA_signal_4614) ) ;
    buf_clk new_AGEMA_reg_buffer_1185 ( .C (clk), .D (new_AGEMA_signal_4615), .Q (new_AGEMA_signal_4616) ) ;
    buf_clk new_AGEMA_reg_buffer_1187 ( .C (clk), .D (new_AGEMA_signal_4617), .Q (new_AGEMA_signal_4618) ) ;
    buf_clk new_AGEMA_reg_buffer_1189 ( .C (clk), .D (new_AGEMA_signal_4619), .Q (new_AGEMA_signal_4620) ) ;
    buf_clk new_AGEMA_reg_buffer_1191 ( .C (clk), .D (new_AGEMA_signal_4621), .Q (new_AGEMA_signal_4622) ) ;
    buf_clk new_AGEMA_reg_buffer_1193 ( .C (clk), .D (new_AGEMA_signal_4623), .Q (new_AGEMA_signal_4624) ) ;
    buf_clk new_AGEMA_reg_buffer_1195 ( .C (clk), .D (new_AGEMA_signal_4625), .Q (new_AGEMA_signal_4626) ) ;
    buf_clk new_AGEMA_reg_buffer_1197 ( .C (clk), .D (new_AGEMA_signal_4627), .Q (new_AGEMA_signal_4628) ) ;
    buf_clk new_AGEMA_reg_buffer_1199 ( .C (clk), .D (new_AGEMA_signal_4629), .Q (new_AGEMA_signal_4630) ) ;
    buf_clk new_AGEMA_reg_buffer_1201 ( .C (clk), .D (new_AGEMA_signal_4631), .Q (new_AGEMA_signal_4632) ) ;
    buf_clk new_AGEMA_reg_buffer_1203 ( .C (clk), .D (new_AGEMA_signal_4633), .Q (new_AGEMA_signal_4634) ) ;
    buf_clk new_AGEMA_reg_buffer_1205 ( .C (clk), .D (new_AGEMA_signal_4635), .Q (new_AGEMA_signal_4636) ) ;
    buf_clk new_AGEMA_reg_buffer_1207 ( .C (clk), .D (new_AGEMA_signal_4637), .Q (new_AGEMA_signal_4638) ) ;
    buf_clk new_AGEMA_reg_buffer_1209 ( .C (clk), .D (new_AGEMA_signal_4639), .Q (new_AGEMA_signal_4640) ) ;
    buf_clk new_AGEMA_reg_buffer_1211 ( .C (clk), .D (new_AGEMA_signal_4641), .Q (new_AGEMA_signal_4642) ) ;
    buf_clk new_AGEMA_reg_buffer_1213 ( .C (clk), .D (new_AGEMA_signal_4643), .Q (new_AGEMA_signal_4644) ) ;
    buf_clk new_AGEMA_reg_buffer_1215 ( .C (clk), .D (new_AGEMA_signal_4645), .Q (new_AGEMA_signal_4646) ) ;
    buf_clk new_AGEMA_reg_buffer_1217 ( .C (clk), .D (new_AGEMA_signal_4647), .Q (new_AGEMA_signal_4648) ) ;
    buf_clk new_AGEMA_reg_buffer_1219 ( .C (clk), .D (new_AGEMA_signal_4649), .Q (new_AGEMA_signal_4650) ) ;
    buf_clk new_AGEMA_reg_buffer_1221 ( .C (clk), .D (new_AGEMA_signal_4651), .Q (new_AGEMA_signal_4652) ) ;
    buf_clk new_AGEMA_reg_buffer_1223 ( .C (clk), .D (new_AGEMA_signal_4653), .Q (new_AGEMA_signal_4654) ) ;
    buf_clk new_AGEMA_reg_buffer_1225 ( .C (clk), .D (new_AGEMA_signal_4655), .Q (new_AGEMA_signal_4656) ) ;
    buf_clk new_AGEMA_reg_buffer_1227 ( .C (clk), .D (new_AGEMA_signal_4657), .Q (new_AGEMA_signal_4658) ) ;
    buf_clk new_AGEMA_reg_buffer_1229 ( .C (clk), .D (new_AGEMA_signal_4659), .Q (new_AGEMA_signal_4660) ) ;
    buf_clk new_AGEMA_reg_buffer_1231 ( .C (clk), .D (new_AGEMA_signal_4661), .Q (new_AGEMA_signal_4662) ) ;
    buf_clk new_AGEMA_reg_buffer_1233 ( .C (clk), .D (new_AGEMA_signal_4663), .Q (new_AGEMA_signal_4664) ) ;
    buf_clk new_AGEMA_reg_buffer_1235 ( .C (clk), .D (new_AGEMA_signal_4665), .Q (new_AGEMA_signal_4666) ) ;
    buf_clk new_AGEMA_reg_buffer_1237 ( .C (clk), .D (new_AGEMA_signal_4667), .Q (new_AGEMA_signal_4668) ) ;
    buf_clk new_AGEMA_reg_buffer_1239 ( .C (clk), .D (new_AGEMA_signal_4669), .Q (new_AGEMA_signal_4670) ) ;
    buf_clk new_AGEMA_reg_buffer_1241 ( .C (clk), .D (new_AGEMA_signal_4671), .Q (new_AGEMA_signal_4672) ) ;
    buf_clk new_AGEMA_reg_buffer_1243 ( .C (clk), .D (new_AGEMA_signal_4673), .Q (new_AGEMA_signal_4674) ) ;
    buf_clk new_AGEMA_reg_buffer_1245 ( .C (clk), .D (new_AGEMA_signal_4675), .Q (new_AGEMA_signal_4676) ) ;
    buf_clk new_AGEMA_reg_buffer_1247 ( .C (clk), .D (new_AGEMA_signal_4677), .Q (new_AGEMA_signal_4678) ) ;
    buf_clk new_AGEMA_reg_buffer_1249 ( .C (clk), .D (new_AGEMA_signal_4679), .Q (new_AGEMA_signal_4680) ) ;
    buf_clk new_AGEMA_reg_buffer_1251 ( .C (clk), .D (new_AGEMA_signal_4681), .Q (new_AGEMA_signal_4682) ) ;
    buf_clk new_AGEMA_reg_buffer_1253 ( .C (clk), .D (new_AGEMA_signal_4683), .Q (new_AGEMA_signal_4684) ) ;
    buf_clk new_AGEMA_reg_buffer_1255 ( .C (clk), .D (new_AGEMA_signal_4685), .Q (new_AGEMA_signal_4686) ) ;
    buf_clk new_AGEMA_reg_buffer_1257 ( .C (clk), .D (new_AGEMA_signal_4687), .Q (new_AGEMA_signal_4688) ) ;
    buf_clk new_AGEMA_reg_buffer_1259 ( .C (clk), .D (new_AGEMA_signal_4689), .Q (new_AGEMA_signal_4690) ) ;
    buf_clk new_AGEMA_reg_buffer_1261 ( .C (clk), .D (new_AGEMA_signal_4691), .Q (new_AGEMA_signal_4692) ) ;
    buf_clk new_AGEMA_reg_buffer_1263 ( .C (clk), .D (new_AGEMA_signal_4693), .Q (new_AGEMA_signal_4694) ) ;
    buf_clk new_AGEMA_reg_buffer_1265 ( .C (clk), .D (new_AGEMA_signal_4695), .Q (new_AGEMA_signal_4696) ) ;
    buf_clk new_AGEMA_reg_buffer_1267 ( .C (clk), .D (new_AGEMA_signal_4697), .Q (new_AGEMA_signal_4698) ) ;
    buf_clk new_AGEMA_reg_buffer_1269 ( .C (clk), .D (new_AGEMA_signal_4699), .Q (new_AGEMA_signal_4700) ) ;
    buf_clk new_AGEMA_reg_buffer_1271 ( .C (clk), .D (new_AGEMA_signal_4701), .Q (new_AGEMA_signal_4702) ) ;
    buf_clk new_AGEMA_reg_buffer_1273 ( .C (clk), .D (new_AGEMA_signal_4703), .Q (new_AGEMA_signal_4704) ) ;
    buf_clk new_AGEMA_reg_buffer_1275 ( .C (clk), .D (new_AGEMA_signal_4705), .Q (new_AGEMA_signal_4706) ) ;
    buf_clk new_AGEMA_reg_buffer_1277 ( .C (clk), .D (new_AGEMA_signal_4707), .Q (new_AGEMA_signal_4708) ) ;
    buf_clk new_AGEMA_reg_buffer_1279 ( .C (clk), .D (new_AGEMA_signal_4709), .Q (new_AGEMA_signal_4710) ) ;
    buf_clk new_AGEMA_reg_buffer_1281 ( .C (clk), .D (new_AGEMA_signal_4711), .Q (new_AGEMA_signal_4712) ) ;
    buf_clk new_AGEMA_reg_buffer_1283 ( .C (clk), .D (new_AGEMA_signal_4713), .Q (new_AGEMA_signal_4714) ) ;
    buf_clk new_AGEMA_reg_buffer_1285 ( .C (clk), .D (new_AGEMA_signal_4715), .Q (new_AGEMA_signal_4716) ) ;
    buf_clk new_AGEMA_reg_buffer_1287 ( .C (clk), .D (new_AGEMA_signal_4717), .Q (new_AGEMA_signal_4718) ) ;
    buf_clk new_AGEMA_reg_buffer_1289 ( .C (clk), .D (new_AGEMA_signal_4719), .Q (new_AGEMA_signal_4720) ) ;
    buf_clk new_AGEMA_reg_buffer_1291 ( .C (clk), .D (new_AGEMA_signal_4721), .Q (new_AGEMA_signal_4722) ) ;
    buf_clk new_AGEMA_reg_buffer_1293 ( .C (clk), .D (new_AGEMA_signal_4723), .Q (new_AGEMA_signal_4724) ) ;
    buf_clk new_AGEMA_reg_buffer_1295 ( .C (clk), .D (new_AGEMA_signal_4725), .Q (new_AGEMA_signal_4726) ) ;
    buf_clk new_AGEMA_reg_buffer_1297 ( .C (clk), .D (new_AGEMA_signal_4727), .Q (new_AGEMA_signal_4728) ) ;
    buf_clk new_AGEMA_reg_buffer_1299 ( .C (clk), .D (new_AGEMA_signal_4729), .Q (new_AGEMA_signal_4730) ) ;
    buf_clk new_AGEMA_reg_buffer_1301 ( .C (clk), .D (new_AGEMA_signal_4731), .Q (new_AGEMA_signal_4732) ) ;
    buf_clk new_AGEMA_reg_buffer_1303 ( .C (clk), .D (new_AGEMA_signal_4733), .Q (new_AGEMA_signal_4734) ) ;
    buf_clk new_AGEMA_reg_buffer_1305 ( .C (clk), .D (new_AGEMA_signal_4735), .Q (new_AGEMA_signal_4736) ) ;
    buf_clk new_AGEMA_reg_buffer_1307 ( .C (clk), .D (new_AGEMA_signal_4737), .Q (new_AGEMA_signal_4738) ) ;
    buf_clk new_AGEMA_reg_buffer_1309 ( .C (clk), .D (new_AGEMA_signal_4739), .Q (new_AGEMA_signal_4740) ) ;
    buf_clk new_AGEMA_reg_buffer_1311 ( .C (clk), .D (new_AGEMA_signal_4741), .Q (new_AGEMA_signal_4742) ) ;
    buf_clk new_AGEMA_reg_buffer_1313 ( .C (clk), .D (new_AGEMA_signal_4743), .Q (new_AGEMA_signal_4744) ) ;
    buf_clk new_AGEMA_reg_buffer_1315 ( .C (clk), .D (new_AGEMA_signal_4745), .Q (new_AGEMA_signal_4746) ) ;
    buf_clk new_AGEMA_reg_buffer_1317 ( .C (clk), .D (new_AGEMA_signal_4747), .Q (new_AGEMA_signal_4748) ) ;
    buf_clk new_AGEMA_reg_buffer_1319 ( .C (clk), .D (new_AGEMA_signal_4749), .Q (new_AGEMA_signal_4750) ) ;
    buf_clk new_AGEMA_reg_buffer_1321 ( .C (clk), .D (new_AGEMA_signal_4751), .Q (new_AGEMA_signal_4752) ) ;
    buf_clk new_AGEMA_reg_buffer_1323 ( .C (clk), .D (new_AGEMA_signal_4753), .Q (new_AGEMA_signal_4754) ) ;
    buf_clk new_AGEMA_reg_buffer_1325 ( .C (clk), .D (new_AGEMA_signal_4755), .Q (new_AGEMA_signal_4756) ) ;
    buf_clk new_AGEMA_reg_buffer_1327 ( .C (clk), .D (new_AGEMA_signal_4757), .Q (new_AGEMA_signal_4758) ) ;
    buf_clk new_AGEMA_reg_buffer_1329 ( .C (clk), .D (new_AGEMA_signal_4759), .Q (new_AGEMA_signal_4760) ) ;
    buf_clk new_AGEMA_reg_buffer_1331 ( .C (clk), .D (new_AGEMA_signal_4761), .Q (new_AGEMA_signal_4762) ) ;
    buf_clk new_AGEMA_reg_buffer_1333 ( .C (clk), .D (new_AGEMA_signal_4763), .Q (new_AGEMA_signal_4764) ) ;
    buf_clk new_AGEMA_reg_buffer_1335 ( .C (clk), .D (new_AGEMA_signal_4765), .Q (new_AGEMA_signal_4766) ) ;
    buf_clk new_AGEMA_reg_buffer_1337 ( .C (clk), .D (new_AGEMA_signal_4767), .Q (new_AGEMA_signal_4768) ) ;
    buf_clk new_AGEMA_reg_buffer_1339 ( .C (clk), .D (new_AGEMA_signal_4769), .Q (new_AGEMA_signal_4770) ) ;
    buf_clk new_AGEMA_reg_buffer_1341 ( .C (clk), .D (new_AGEMA_signal_4771), .Q (new_AGEMA_signal_4772) ) ;
    buf_clk new_AGEMA_reg_buffer_1343 ( .C (clk), .D (new_AGEMA_signal_4773), .Q (new_AGEMA_signal_4774) ) ;
    buf_clk new_AGEMA_reg_buffer_1345 ( .C (clk), .D (new_AGEMA_signal_4775), .Q (new_AGEMA_signal_4776) ) ;
    buf_clk new_AGEMA_reg_buffer_1347 ( .C (clk), .D (new_AGEMA_signal_4777), .Q (new_AGEMA_signal_4778) ) ;
    buf_clk new_AGEMA_reg_buffer_1349 ( .C (clk), .D (new_AGEMA_signal_4779), .Q (new_AGEMA_signal_4780) ) ;
    buf_clk new_AGEMA_reg_buffer_1351 ( .C (clk), .D (new_AGEMA_signal_4781), .Q (new_AGEMA_signal_4782) ) ;
    buf_clk new_AGEMA_reg_buffer_1353 ( .C (clk), .D (new_AGEMA_signal_4783), .Q (new_AGEMA_signal_4784) ) ;
    buf_clk new_AGEMA_reg_buffer_1355 ( .C (clk), .D (new_AGEMA_signal_4785), .Q (new_AGEMA_signal_4786) ) ;
    buf_clk new_AGEMA_reg_buffer_1357 ( .C (clk), .D (new_AGEMA_signal_4787), .Q (new_AGEMA_signal_4788) ) ;
    buf_clk new_AGEMA_reg_buffer_1359 ( .C (clk), .D (new_AGEMA_signal_4789), .Q (new_AGEMA_signal_4790) ) ;
    buf_clk new_AGEMA_reg_buffer_1361 ( .C (clk), .D (new_AGEMA_signal_4791), .Q (new_AGEMA_signal_4792) ) ;
    buf_clk new_AGEMA_reg_buffer_1363 ( .C (clk), .D (new_AGEMA_signal_4793), .Q (new_AGEMA_signal_4794) ) ;
    buf_clk new_AGEMA_reg_buffer_1365 ( .C (clk), .D (new_AGEMA_signal_4795), .Q (new_AGEMA_signal_4796) ) ;
    buf_clk new_AGEMA_reg_buffer_1367 ( .C (clk), .D (new_AGEMA_signal_4797), .Q (new_AGEMA_signal_4798) ) ;
    buf_clk new_AGEMA_reg_buffer_1369 ( .C (clk), .D (new_AGEMA_signal_4799), .Q (new_AGEMA_signal_4800) ) ;
    buf_clk new_AGEMA_reg_buffer_1371 ( .C (clk), .D (new_AGEMA_signal_4801), .Q (new_AGEMA_signal_4802) ) ;
    buf_clk new_AGEMA_reg_buffer_1373 ( .C (clk), .D (new_AGEMA_signal_4803), .Q (new_AGEMA_signal_4804) ) ;
    buf_clk new_AGEMA_reg_buffer_1375 ( .C (clk), .D (new_AGEMA_signal_4805), .Q (new_AGEMA_signal_4806) ) ;
    buf_clk new_AGEMA_reg_buffer_1377 ( .C (clk), .D (new_AGEMA_signal_4807), .Q (new_AGEMA_signal_4808) ) ;
    buf_clk new_AGEMA_reg_buffer_1379 ( .C (clk), .D (new_AGEMA_signal_4809), .Q (new_AGEMA_signal_4810) ) ;
    buf_clk new_AGEMA_reg_buffer_1381 ( .C (clk), .D (new_AGEMA_signal_4811), .Q (new_AGEMA_signal_4812) ) ;
    buf_clk new_AGEMA_reg_buffer_1383 ( .C (clk), .D (new_AGEMA_signal_4813), .Q (new_AGEMA_signal_4814) ) ;
    buf_clk new_AGEMA_reg_buffer_1385 ( .C (clk), .D (new_AGEMA_signal_4815), .Q (new_AGEMA_signal_4816) ) ;
    buf_clk new_AGEMA_reg_buffer_1387 ( .C (clk), .D (new_AGEMA_signal_4817), .Q (new_AGEMA_signal_4818) ) ;
    buf_clk new_AGEMA_reg_buffer_1389 ( .C (clk), .D (new_AGEMA_signal_4819), .Q (new_AGEMA_signal_4820) ) ;
    buf_clk new_AGEMA_reg_buffer_1391 ( .C (clk), .D (new_AGEMA_signal_4821), .Q (new_AGEMA_signal_4822) ) ;
    buf_clk new_AGEMA_reg_buffer_1393 ( .C (clk), .D (new_AGEMA_signal_4823), .Q (new_AGEMA_signal_4824) ) ;
    buf_clk new_AGEMA_reg_buffer_1395 ( .C (clk), .D (new_AGEMA_signal_4825), .Q (new_AGEMA_signal_4826) ) ;
    buf_clk new_AGEMA_reg_buffer_1397 ( .C (clk), .D (new_AGEMA_signal_4827), .Q (new_AGEMA_signal_4828) ) ;
    buf_clk new_AGEMA_reg_buffer_1399 ( .C (clk), .D (new_AGEMA_signal_4829), .Q (new_AGEMA_signal_4830) ) ;
    buf_clk new_AGEMA_reg_buffer_1401 ( .C (clk), .D (new_AGEMA_signal_4831), .Q (new_AGEMA_signal_4832) ) ;
    buf_clk new_AGEMA_reg_buffer_1403 ( .C (clk), .D (new_AGEMA_signal_4833), .Q (new_AGEMA_signal_4834) ) ;
    buf_clk new_AGEMA_reg_buffer_1405 ( .C (clk), .D (new_AGEMA_signal_4835), .Q (new_AGEMA_signal_4836) ) ;
    buf_clk new_AGEMA_reg_buffer_1407 ( .C (clk), .D (new_AGEMA_signal_4837), .Q (new_AGEMA_signal_4838) ) ;
    buf_clk new_AGEMA_reg_buffer_1409 ( .C (clk), .D (new_AGEMA_signal_4839), .Q (new_AGEMA_signal_4840) ) ;
    buf_clk new_AGEMA_reg_buffer_1411 ( .C (clk), .D (new_AGEMA_signal_4841), .Q (new_AGEMA_signal_4842) ) ;
    buf_clk new_AGEMA_reg_buffer_1413 ( .C (clk), .D (new_AGEMA_signal_4843), .Q (new_AGEMA_signal_4844) ) ;
    buf_clk new_AGEMA_reg_buffer_1415 ( .C (clk), .D (new_AGEMA_signal_4845), .Q (new_AGEMA_signal_4846) ) ;
    buf_clk new_AGEMA_reg_buffer_1417 ( .C (clk), .D (new_AGEMA_signal_4847), .Q (new_AGEMA_signal_4848) ) ;
    buf_clk new_AGEMA_reg_buffer_1419 ( .C (clk), .D (new_AGEMA_signal_4849), .Q (new_AGEMA_signal_4850) ) ;
    buf_clk new_AGEMA_reg_buffer_1421 ( .C (clk), .D (new_AGEMA_signal_4851), .Q (new_AGEMA_signal_4852) ) ;
    buf_clk new_AGEMA_reg_buffer_1423 ( .C (clk), .D (new_AGEMA_signal_4853), .Q (new_AGEMA_signal_4854) ) ;
    buf_clk new_AGEMA_reg_buffer_1425 ( .C (clk), .D (new_AGEMA_signal_4855), .Q (new_AGEMA_signal_4856) ) ;
    buf_clk new_AGEMA_reg_buffer_1427 ( .C (clk), .D (new_AGEMA_signal_4857), .Q (new_AGEMA_signal_4858) ) ;
    buf_clk new_AGEMA_reg_buffer_1429 ( .C (clk), .D (new_AGEMA_signal_4859), .Q (new_AGEMA_signal_4860) ) ;
    buf_clk new_AGEMA_reg_buffer_1431 ( .C (clk), .D (new_AGEMA_signal_4861), .Q (new_AGEMA_signal_4862) ) ;
    buf_clk new_AGEMA_reg_buffer_1433 ( .C (clk), .D (new_AGEMA_signal_4863), .Q (new_AGEMA_signal_4864) ) ;
    buf_clk new_AGEMA_reg_buffer_1435 ( .C (clk), .D (new_AGEMA_signal_4865), .Q (new_AGEMA_signal_4866) ) ;
    buf_clk new_AGEMA_reg_buffer_1437 ( .C (clk), .D (new_AGEMA_signal_4867), .Q (new_AGEMA_signal_4868) ) ;
    buf_clk new_AGEMA_reg_buffer_1439 ( .C (clk), .D (new_AGEMA_signal_4869), .Q (new_AGEMA_signal_4870) ) ;
    buf_clk new_AGEMA_reg_buffer_1441 ( .C (clk), .D (new_AGEMA_signal_4871), .Q (new_AGEMA_signal_4872) ) ;
    buf_clk new_AGEMA_reg_buffer_1443 ( .C (clk), .D (new_AGEMA_signal_4873), .Q (new_AGEMA_signal_4874) ) ;
    buf_clk new_AGEMA_reg_buffer_1445 ( .C (clk), .D (new_AGEMA_signal_4875), .Q (new_AGEMA_signal_4876) ) ;
    buf_clk new_AGEMA_reg_buffer_1447 ( .C (clk), .D (new_AGEMA_signal_4877), .Q (new_AGEMA_signal_4878) ) ;
    buf_clk new_AGEMA_reg_buffer_1449 ( .C (clk), .D (new_AGEMA_signal_4879), .Q (new_AGEMA_signal_4880) ) ;
    buf_clk new_AGEMA_reg_buffer_1451 ( .C (clk), .D (new_AGEMA_signal_4881), .Q (new_AGEMA_signal_4882) ) ;
    buf_clk new_AGEMA_reg_buffer_1453 ( .C (clk), .D (new_AGEMA_signal_4883), .Q (new_AGEMA_signal_4884) ) ;
    buf_clk new_AGEMA_reg_buffer_1455 ( .C (clk), .D (new_AGEMA_signal_4885), .Q (new_AGEMA_signal_4886) ) ;
    buf_clk new_AGEMA_reg_buffer_1457 ( .C (clk), .D (new_AGEMA_signal_4887), .Q (new_AGEMA_signal_4888) ) ;
    buf_clk new_AGEMA_reg_buffer_1459 ( .C (clk), .D (new_AGEMA_signal_4889), .Q (new_AGEMA_signal_4890) ) ;
    buf_clk new_AGEMA_reg_buffer_1461 ( .C (clk), .D (new_AGEMA_signal_4891), .Q (new_AGEMA_signal_4892) ) ;
    buf_clk new_AGEMA_reg_buffer_1463 ( .C (clk), .D (new_AGEMA_signal_4893), .Q (new_AGEMA_signal_4894) ) ;
    buf_clk new_AGEMA_reg_buffer_1465 ( .C (clk), .D (new_AGEMA_signal_4895), .Q (new_AGEMA_signal_4896) ) ;
    buf_clk new_AGEMA_reg_buffer_1467 ( .C (clk), .D (new_AGEMA_signal_4897), .Q (new_AGEMA_signal_4898) ) ;
    buf_clk new_AGEMA_reg_buffer_1469 ( .C (clk), .D (new_AGEMA_signal_4899), .Q (new_AGEMA_signal_4900) ) ;
    buf_clk new_AGEMA_reg_buffer_1471 ( .C (clk), .D (new_AGEMA_signal_4901), .Q (new_AGEMA_signal_4902) ) ;
    buf_clk new_AGEMA_reg_buffer_1473 ( .C (clk), .D (new_AGEMA_signal_4903), .Q (new_AGEMA_signal_4904) ) ;
    buf_clk new_AGEMA_reg_buffer_1475 ( .C (clk), .D (new_AGEMA_signal_4905), .Q (new_AGEMA_signal_4906) ) ;
    buf_clk new_AGEMA_reg_buffer_1477 ( .C (clk), .D (new_AGEMA_signal_4907), .Q (new_AGEMA_signal_4908) ) ;
    buf_clk new_AGEMA_reg_buffer_1479 ( .C (clk), .D (new_AGEMA_signal_4909), .Q (new_AGEMA_signal_4910) ) ;
    buf_clk new_AGEMA_reg_buffer_1481 ( .C (clk), .D (new_AGEMA_signal_4911), .Q (new_AGEMA_signal_4912) ) ;
    buf_clk new_AGEMA_reg_buffer_1483 ( .C (clk), .D (new_AGEMA_signal_4913), .Q (new_AGEMA_signal_4914) ) ;
    buf_clk new_AGEMA_reg_buffer_1485 ( .C (clk), .D (new_AGEMA_signal_4915), .Q (new_AGEMA_signal_4916) ) ;
    buf_clk new_AGEMA_reg_buffer_1487 ( .C (clk), .D (new_AGEMA_signal_4917), .Q (new_AGEMA_signal_4918) ) ;
    buf_clk new_AGEMA_reg_buffer_1489 ( .C (clk), .D (new_AGEMA_signal_4919), .Q (new_AGEMA_signal_4920) ) ;
    buf_clk new_AGEMA_reg_buffer_1491 ( .C (clk), .D (new_AGEMA_signal_4921), .Q (new_AGEMA_signal_4922) ) ;
    buf_clk new_AGEMA_reg_buffer_1493 ( .C (clk), .D (new_AGEMA_signal_4923), .Q (new_AGEMA_signal_4924) ) ;
    buf_clk new_AGEMA_reg_buffer_1495 ( .C (clk), .D (new_AGEMA_signal_4925), .Q (new_AGEMA_signal_4926) ) ;
    buf_clk new_AGEMA_reg_buffer_1497 ( .C (clk), .D (new_AGEMA_signal_4927), .Q (new_AGEMA_signal_4928) ) ;
    buf_clk new_AGEMA_reg_buffer_1499 ( .C (clk), .D (new_AGEMA_signal_4929), .Q (new_AGEMA_signal_4930) ) ;
    buf_clk new_AGEMA_reg_buffer_1501 ( .C (clk), .D (new_AGEMA_signal_4931), .Q (new_AGEMA_signal_4932) ) ;
    buf_clk new_AGEMA_reg_buffer_1503 ( .C (clk), .D (new_AGEMA_signal_4933), .Q (new_AGEMA_signal_4934) ) ;
    buf_clk new_AGEMA_reg_buffer_1505 ( .C (clk), .D (new_AGEMA_signal_4935), .Q (new_AGEMA_signal_4936) ) ;
    buf_clk new_AGEMA_reg_buffer_1507 ( .C (clk), .D (new_AGEMA_signal_4937), .Q (new_AGEMA_signal_4938) ) ;
    buf_clk new_AGEMA_reg_buffer_1509 ( .C (clk), .D (new_AGEMA_signal_4939), .Q (new_AGEMA_signal_4940) ) ;
    buf_clk new_AGEMA_reg_buffer_1511 ( .C (clk), .D (new_AGEMA_signal_4941), .Q (new_AGEMA_signal_4942) ) ;
    buf_clk new_AGEMA_reg_buffer_1513 ( .C (clk), .D (new_AGEMA_signal_4943), .Q (new_AGEMA_signal_4944) ) ;
    buf_clk new_AGEMA_reg_buffer_1515 ( .C (clk), .D (new_AGEMA_signal_4945), .Q (new_AGEMA_signal_4946) ) ;
    buf_clk new_AGEMA_reg_buffer_1517 ( .C (clk), .D (new_AGEMA_signal_4947), .Q (new_AGEMA_signal_4948) ) ;
    buf_clk new_AGEMA_reg_buffer_1519 ( .C (clk), .D (new_AGEMA_signal_4949), .Q (new_AGEMA_signal_4950) ) ;
    buf_clk new_AGEMA_reg_buffer_1521 ( .C (clk), .D (new_AGEMA_signal_4951), .Q (new_AGEMA_signal_4952) ) ;
    buf_clk new_AGEMA_reg_buffer_1523 ( .C (clk), .D (new_AGEMA_signal_4953), .Q (new_AGEMA_signal_4954) ) ;
    buf_clk new_AGEMA_reg_buffer_1525 ( .C (clk), .D (new_AGEMA_signal_4955), .Q (new_AGEMA_signal_4956) ) ;
    buf_clk new_AGEMA_reg_buffer_1527 ( .C (clk), .D (new_AGEMA_signal_4957), .Q (new_AGEMA_signal_4958) ) ;
    buf_clk new_AGEMA_reg_buffer_1529 ( .C (clk), .D (new_AGEMA_signal_4959), .Q (new_AGEMA_signal_4960) ) ;
    buf_clk new_AGEMA_reg_buffer_1531 ( .C (clk), .D (new_AGEMA_signal_4961), .Q (new_AGEMA_signal_4962) ) ;
    buf_clk new_AGEMA_reg_buffer_1533 ( .C (clk), .D (new_AGEMA_signal_4963), .Q (new_AGEMA_signal_4964) ) ;
    buf_clk new_AGEMA_reg_buffer_1535 ( .C (clk), .D (new_AGEMA_signal_4965), .Q (new_AGEMA_signal_4966) ) ;
    buf_clk new_AGEMA_reg_buffer_1537 ( .C (clk), .D (new_AGEMA_signal_4967), .Q (new_AGEMA_signal_4968) ) ;
    buf_clk new_AGEMA_reg_buffer_1539 ( .C (clk), .D (new_AGEMA_signal_4969), .Q (new_AGEMA_signal_4970) ) ;
    buf_clk new_AGEMA_reg_buffer_1541 ( .C (clk), .D (new_AGEMA_signal_4971), .Q (new_AGEMA_signal_4972) ) ;
    buf_clk new_AGEMA_reg_buffer_1543 ( .C (clk), .D (new_AGEMA_signal_4973), .Q (new_AGEMA_signal_4974) ) ;
    buf_clk new_AGEMA_reg_buffer_1545 ( .C (clk), .D (new_AGEMA_signal_4975), .Q (new_AGEMA_signal_4976) ) ;
    buf_clk new_AGEMA_reg_buffer_1547 ( .C (clk), .D (new_AGEMA_signal_4977), .Q (new_AGEMA_signal_4978) ) ;
    buf_clk new_AGEMA_reg_buffer_1549 ( .C (clk), .D (new_AGEMA_signal_4979), .Q (new_AGEMA_signal_4980) ) ;
    buf_clk new_AGEMA_reg_buffer_1551 ( .C (clk), .D (new_AGEMA_signal_4981), .Q (new_AGEMA_signal_4982) ) ;
    buf_clk new_AGEMA_reg_buffer_1553 ( .C (clk), .D (new_AGEMA_signal_4983), .Q (new_AGEMA_signal_4984) ) ;
    buf_clk new_AGEMA_reg_buffer_1555 ( .C (clk), .D (new_AGEMA_signal_4985), .Q (new_AGEMA_signal_4986) ) ;
    buf_clk new_AGEMA_reg_buffer_1557 ( .C (clk), .D (new_AGEMA_signal_4987), .Q (new_AGEMA_signal_4988) ) ;
    buf_clk new_AGEMA_reg_buffer_1559 ( .C (clk), .D (new_AGEMA_signal_4989), .Q (new_AGEMA_signal_4990) ) ;
    buf_clk new_AGEMA_reg_buffer_1561 ( .C (clk), .D (new_AGEMA_signal_4991), .Q (new_AGEMA_signal_4992) ) ;
    buf_clk new_AGEMA_reg_buffer_1563 ( .C (clk), .D (new_AGEMA_signal_4993), .Q (new_AGEMA_signal_4994) ) ;
    buf_clk new_AGEMA_reg_buffer_1565 ( .C (clk), .D (new_AGEMA_signal_4995), .Q (new_AGEMA_signal_4996) ) ;
    buf_clk new_AGEMA_reg_buffer_1567 ( .C (clk), .D (new_AGEMA_signal_4997), .Q (new_AGEMA_signal_4998) ) ;
    buf_clk new_AGEMA_reg_buffer_1569 ( .C (clk), .D (new_AGEMA_signal_4999), .Q (new_AGEMA_signal_5000) ) ;
    buf_clk new_AGEMA_reg_buffer_1571 ( .C (clk), .D (new_AGEMA_signal_5001), .Q (new_AGEMA_signal_5002) ) ;
    buf_clk new_AGEMA_reg_buffer_1573 ( .C (clk), .D (new_AGEMA_signal_5003), .Q (new_AGEMA_signal_5004) ) ;
    buf_clk new_AGEMA_reg_buffer_1575 ( .C (clk), .D (new_AGEMA_signal_5005), .Q (new_AGEMA_signal_5006) ) ;
    buf_clk new_AGEMA_reg_buffer_1577 ( .C (clk), .D (new_AGEMA_signal_5007), .Q (new_AGEMA_signal_5008) ) ;
    buf_clk new_AGEMA_reg_buffer_1579 ( .C (clk), .D (new_AGEMA_signal_5009), .Q (new_AGEMA_signal_5010) ) ;
    buf_clk new_AGEMA_reg_buffer_1581 ( .C (clk), .D (new_AGEMA_signal_5011), .Q (new_AGEMA_signal_5012) ) ;
    buf_clk new_AGEMA_reg_buffer_1583 ( .C (clk), .D (new_AGEMA_signal_5013), .Q (new_AGEMA_signal_5014) ) ;
    buf_clk new_AGEMA_reg_buffer_1585 ( .C (clk), .D (new_AGEMA_signal_5015), .Q (new_AGEMA_signal_5016) ) ;
    buf_clk new_AGEMA_reg_buffer_1587 ( .C (clk), .D (new_AGEMA_signal_5017), .Q (new_AGEMA_signal_5018) ) ;
    buf_clk new_AGEMA_reg_buffer_1589 ( .C (clk), .D (new_AGEMA_signal_5019), .Q (new_AGEMA_signal_5020) ) ;
    buf_clk new_AGEMA_reg_buffer_1591 ( .C (clk), .D (new_AGEMA_signal_5021), .Q (new_AGEMA_signal_5022) ) ;
    buf_clk new_AGEMA_reg_buffer_1593 ( .C (clk), .D (new_AGEMA_signal_5023), .Q (new_AGEMA_signal_5024) ) ;
    buf_clk new_AGEMA_reg_buffer_1595 ( .C (clk), .D (new_AGEMA_signal_5025), .Q (new_AGEMA_signal_5026) ) ;
    buf_clk new_AGEMA_reg_buffer_1597 ( .C (clk), .D (new_AGEMA_signal_5027), .Q (new_AGEMA_signal_5028) ) ;
    buf_clk new_AGEMA_reg_buffer_1599 ( .C (clk), .D (new_AGEMA_signal_5029), .Q (new_AGEMA_signal_5030) ) ;
    buf_clk new_AGEMA_reg_buffer_1601 ( .C (clk), .D (new_AGEMA_signal_5031), .Q (new_AGEMA_signal_5032) ) ;
    buf_clk new_AGEMA_reg_buffer_1603 ( .C (clk), .D (new_AGEMA_signal_5033), .Q (new_AGEMA_signal_5034) ) ;
    buf_clk new_AGEMA_reg_buffer_1605 ( .C (clk), .D (new_AGEMA_signal_5035), .Q (new_AGEMA_signal_5036) ) ;
    buf_clk new_AGEMA_reg_buffer_1607 ( .C (clk), .D (new_AGEMA_signal_5037), .Q (new_AGEMA_signal_5038) ) ;
    buf_clk new_AGEMA_reg_buffer_1609 ( .C (clk), .D (new_AGEMA_signal_5039), .Q (new_AGEMA_signal_5040) ) ;
    buf_clk new_AGEMA_reg_buffer_1611 ( .C (clk), .D (new_AGEMA_signal_5041), .Q (new_AGEMA_signal_5042) ) ;
    buf_clk new_AGEMA_reg_buffer_1613 ( .C (clk), .D (new_AGEMA_signal_5043), .Q (new_AGEMA_signal_5044) ) ;
    buf_clk new_AGEMA_reg_buffer_1615 ( .C (clk), .D (new_AGEMA_signal_5045), .Q (new_AGEMA_signal_5046) ) ;
    buf_clk new_AGEMA_reg_buffer_1617 ( .C (clk), .D (new_AGEMA_signal_5047), .Q (new_AGEMA_signal_5048) ) ;
    buf_clk new_AGEMA_reg_buffer_1619 ( .C (clk), .D (new_AGEMA_signal_5049), .Q (new_AGEMA_signal_5050) ) ;
    buf_clk new_AGEMA_reg_buffer_1621 ( .C (clk), .D (new_AGEMA_signal_5051), .Q (new_AGEMA_signal_5052) ) ;
    buf_clk new_AGEMA_reg_buffer_1623 ( .C (clk), .D (new_AGEMA_signal_5053), .Q (new_AGEMA_signal_5054) ) ;
    buf_clk new_AGEMA_reg_buffer_1625 ( .C (clk), .D (new_AGEMA_signal_5055), .Q (new_AGEMA_signal_5056) ) ;
    buf_clk new_AGEMA_reg_buffer_1627 ( .C (clk), .D (new_AGEMA_signal_5057), .Q (new_AGEMA_signal_5058) ) ;
    buf_clk new_AGEMA_reg_buffer_1629 ( .C (clk), .D (new_AGEMA_signal_5059), .Q (new_AGEMA_signal_5060) ) ;
    buf_clk new_AGEMA_reg_buffer_1631 ( .C (clk), .D (new_AGEMA_signal_5061), .Q (new_AGEMA_signal_5062) ) ;
    buf_clk new_AGEMA_reg_buffer_1633 ( .C (clk), .D (new_AGEMA_signal_5063), .Q (new_AGEMA_signal_5064) ) ;
    buf_clk new_AGEMA_reg_buffer_1635 ( .C (clk), .D (new_AGEMA_signal_5065), .Q (new_AGEMA_signal_5066) ) ;
    buf_clk new_AGEMA_reg_buffer_1637 ( .C (clk), .D (new_AGEMA_signal_5067), .Q (new_AGEMA_signal_5068) ) ;
    buf_clk new_AGEMA_reg_buffer_1639 ( .C (clk), .D (new_AGEMA_signal_5069), .Q (new_AGEMA_signal_5070) ) ;
    buf_clk new_AGEMA_reg_buffer_1641 ( .C (clk), .D (new_AGEMA_signal_5071), .Q (new_AGEMA_signal_5072) ) ;
    buf_clk new_AGEMA_reg_buffer_1643 ( .C (clk), .D (new_AGEMA_signal_5073), .Q (new_AGEMA_signal_5074) ) ;
    buf_clk new_AGEMA_reg_buffer_1645 ( .C (clk), .D (new_AGEMA_signal_5075), .Q (new_AGEMA_signal_5076) ) ;
    buf_clk new_AGEMA_reg_buffer_1647 ( .C (clk), .D (new_AGEMA_signal_5077), .Q (new_AGEMA_signal_5078) ) ;
    buf_clk new_AGEMA_reg_buffer_1649 ( .C (clk), .D (new_AGEMA_signal_5079), .Q (new_AGEMA_signal_5080) ) ;
    buf_clk new_AGEMA_reg_buffer_1651 ( .C (clk), .D (new_AGEMA_signal_5081), .Q (new_AGEMA_signal_5082) ) ;
    buf_clk new_AGEMA_reg_buffer_1653 ( .C (clk), .D (new_AGEMA_signal_5083), .Q (new_AGEMA_signal_5084) ) ;
    buf_clk new_AGEMA_reg_buffer_1655 ( .C (clk), .D (new_AGEMA_signal_5085), .Q (new_AGEMA_signal_5086) ) ;
    buf_clk new_AGEMA_reg_buffer_1657 ( .C (clk), .D (new_AGEMA_signal_5087), .Q (new_AGEMA_signal_5088) ) ;
    buf_clk new_AGEMA_reg_buffer_1659 ( .C (clk), .D (new_AGEMA_signal_5089), .Q (new_AGEMA_signal_5090) ) ;
    buf_clk new_AGEMA_reg_buffer_1661 ( .C (clk), .D (new_AGEMA_signal_5091), .Q (new_AGEMA_signal_5092) ) ;
    buf_clk new_AGEMA_reg_buffer_1663 ( .C (clk), .D (new_AGEMA_signal_5093), .Q (new_AGEMA_signal_5094) ) ;
    buf_clk new_AGEMA_reg_buffer_1665 ( .C (clk), .D (new_AGEMA_signal_5095), .Q (new_AGEMA_signal_5096) ) ;
    buf_clk new_AGEMA_reg_buffer_1667 ( .C (clk), .D (new_AGEMA_signal_5097), .Q (new_AGEMA_signal_5098) ) ;
    buf_clk new_AGEMA_reg_buffer_1669 ( .C (clk), .D (new_AGEMA_signal_5099), .Q (new_AGEMA_signal_5100) ) ;
    buf_clk new_AGEMA_reg_buffer_1671 ( .C (clk), .D (new_AGEMA_signal_5101), .Q (new_AGEMA_signal_5102) ) ;
    buf_clk new_AGEMA_reg_buffer_1673 ( .C (clk), .D (new_AGEMA_signal_5103), .Q (new_AGEMA_signal_5104) ) ;
    buf_clk new_AGEMA_reg_buffer_1675 ( .C (clk), .D (new_AGEMA_signal_5105), .Q (new_AGEMA_signal_5106) ) ;
    buf_clk new_AGEMA_reg_buffer_1677 ( .C (clk), .D (new_AGEMA_signal_5107), .Q (new_AGEMA_signal_5108) ) ;
    buf_clk new_AGEMA_reg_buffer_1679 ( .C (clk), .D (new_AGEMA_signal_5109), .Q (new_AGEMA_signal_5110) ) ;
    buf_clk new_AGEMA_reg_buffer_1681 ( .C (clk), .D (new_AGEMA_signal_5111), .Q (new_AGEMA_signal_5112) ) ;
    buf_clk new_AGEMA_reg_buffer_1683 ( .C (clk), .D (new_AGEMA_signal_5113), .Q (new_AGEMA_signal_5114) ) ;
    buf_clk new_AGEMA_reg_buffer_1685 ( .C (clk), .D (new_AGEMA_signal_5115), .Q (new_AGEMA_signal_5116) ) ;
    buf_clk new_AGEMA_reg_buffer_1687 ( .C (clk), .D (new_AGEMA_signal_5117), .Q (new_AGEMA_signal_5118) ) ;
    buf_clk new_AGEMA_reg_buffer_1689 ( .C (clk), .D (new_AGEMA_signal_5119), .Q (new_AGEMA_signal_5120) ) ;
    buf_clk new_AGEMA_reg_buffer_1691 ( .C (clk), .D (new_AGEMA_signal_5121), .Q (new_AGEMA_signal_5122) ) ;
    buf_clk new_AGEMA_reg_buffer_1693 ( .C (clk), .D (new_AGEMA_signal_5123), .Q (new_AGEMA_signal_5124) ) ;
    buf_clk new_AGEMA_reg_buffer_1695 ( .C (clk), .D (new_AGEMA_signal_5125), .Q (new_AGEMA_signal_5126) ) ;
    buf_clk new_AGEMA_reg_buffer_1697 ( .C (clk), .D (new_AGEMA_signal_5127), .Q (new_AGEMA_signal_5128) ) ;
    buf_clk new_AGEMA_reg_buffer_1699 ( .C (clk), .D (new_AGEMA_signal_5129), .Q (new_AGEMA_signal_5130) ) ;
    buf_clk new_AGEMA_reg_buffer_1701 ( .C (clk), .D (new_AGEMA_signal_5131), .Q (new_AGEMA_signal_5132) ) ;
    buf_clk new_AGEMA_reg_buffer_1703 ( .C (clk), .D (new_AGEMA_signal_5133), .Q (new_AGEMA_signal_5134) ) ;
    buf_clk new_AGEMA_reg_buffer_1705 ( .C (clk), .D (new_AGEMA_signal_5135), .Q (new_AGEMA_signal_5136) ) ;
    buf_clk new_AGEMA_reg_buffer_1707 ( .C (clk), .D (new_AGEMA_signal_5137), .Q (new_AGEMA_signal_5138) ) ;
    buf_clk new_AGEMA_reg_buffer_1709 ( .C (clk), .D (new_AGEMA_signal_5139), .Q (new_AGEMA_signal_5140) ) ;
    buf_clk new_AGEMA_reg_buffer_1711 ( .C (clk), .D (new_AGEMA_signal_5141), .Q (new_AGEMA_signal_5142) ) ;
    buf_clk new_AGEMA_reg_buffer_1713 ( .C (clk), .D (new_AGEMA_signal_5143), .Q (new_AGEMA_signal_5144) ) ;
    buf_clk new_AGEMA_reg_buffer_1715 ( .C (clk), .D (new_AGEMA_signal_5145), .Q (new_AGEMA_signal_5146) ) ;
    buf_clk new_AGEMA_reg_buffer_1717 ( .C (clk), .D (new_AGEMA_signal_5147), .Q (new_AGEMA_signal_5148) ) ;
    buf_clk new_AGEMA_reg_buffer_1719 ( .C (clk), .D (new_AGEMA_signal_5149), .Q (new_AGEMA_signal_5150) ) ;
    buf_clk new_AGEMA_reg_buffer_1721 ( .C (clk), .D (new_AGEMA_signal_5151), .Q (new_AGEMA_signal_5152) ) ;
    buf_clk new_AGEMA_reg_buffer_1723 ( .C (clk), .D (new_AGEMA_signal_5153), .Q (new_AGEMA_signal_5154) ) ;
    buf_clk new_AGEMA_reg_buffer_1725 ( .C (clk), .D (new_AGEMA_signal_5155), .Q (new_AGEMA_signal_5156) ) ;
    buf_clk new_AGEMA_reg_buffer_1727 ( .C (clk), .D (new_AGEMA_signal_5157), .Q (new_AGEMA_signal_5158) ) ;
    buf_clk new_AGEMA_reg_buffer_1729 ( .C (clk), .D (new_AGEMA_signal_5159), .Q (new_AGEMA_signal_5160) ) ;
    buf_clk new_AGEMA_reg_buffer_1731 ( .C (clk), .D (new_AGEMA_signal_5161), .Q (new_AGEMA_signal_5162) ) ;
    buf_clk new_AGEMA_reg_buffer_1733 ( .C (clk), .D (new_AGEMA_signal_5163), .Q (new_AGEMA_signal_5164) ) ;
    buf_clk new_AGEMA_reg_buffer_1735 ( .C (clk), .D (new_AGEMA_signal_5165), .Q (new_AGEMA_signal_5166) ) ;
    buf_clk new_AGEMA_reg_buffer_1737 ( .C (clk), .D (new_AGEMA_signal_5167), .Q (new_AGEMA_signal_5168) ) ;
    buf_clk new_AGEMA_reg_buffer_1739 ( .C (clk), .D (new_AGEMA_signal_5169), .Q (new_AGEMA_signal_5170) ) ;
    buf_clk new_AGEMA_reg_buffer_1741 ( .C (clk), .D (new_AGEMA_signal_5171), .Q (new_AGEMA_signal_5172) ) ;
    buf_clk new_AGEMA_reg_buffer_1743 ( .C (clk), .D (new_AGEMA_signal_5173), .Q (new_AGEMA_signal_5174) ) ;
    buf_clk new_AGEMA_reg_buffer_1745 ( .C (clk), .D (new_AGEMA_signal_5175), .Q (new_AGEMA_signal_5176) ) ;
    buf_clk new_AGEMA_reg_buffer_1747 ( .C (clk), .D (new_AGEMA_signal_5177), .Q (new_AGEMA_signal_5178) ) ;
    buf_clk new_AGEMA_reg_buffer_1749 ( .C (clk), .D (new_AGEMA_signal_5179), .Q (new_AGEMA_signal_5180) ) ;
    buf_clk new_AGEMA_reg_buffer_1751 ( .C (clk), .D (new_AGEMA_signal_5181), .Q (new_AGEMA_signal_5182) ) ;
    buf_clk new_AGEMA_reg_buffer_1753 ( .C (clk), .D (new_AGEMA_signal_5183), .Q (new_AGEMA_signal_5184) ) ;
    buf_clk new_AGEMA_reg_buffer_1755 ( .C (clk), .D (new_AGEMA_signal_5185), .Q (new_AGEMA_signal_5186) ) ;
    buf_clk new_AGEMA_reg_buffer_1757 ( .C (clk), .D (new_AGEMA_signal_5187), .Q (new_AGEMA_signal_5188) ) ;
    buf_clk new_AGEMA_reg_buffer_1759 ( .C (clk), .D (new_AGEMA_signal_5189), .Q (new_AGEMA_signal_5190) ) ;
    buf_clk new_AGEMA_reg_buffer_1761 ( .C (clk), .D (new_AGEMA_signal_5191), .Q (new_AGEMA_signal_5192) ) ;
    buf_clk new_AGEMA_reg_buffer_1763 ( .C (clk), .D (new_AGEMA_signal_5193), .Q (new_AGEMA_signal_5194) ) ;
    buf_clk new_AGEMA_reg_buffer_1765 ( .C (clk), .D (new_AGEMA_signal_5195), .Q (new_AGEMA_signal_5196) ) ;
    buf_clk new_AGEMA_reg_buffer_1767 ( .C (clk), .D (new_AGEMA_signal_5197), .Q (new_AGEMA_signal_5198) ) ;
    buf_clk new_AGEMA_reg_buffer_1769 ( .C (clk), .D (new_AGEMA_signal_5199), .Q (new_AGEMA_signal_5200) ) ;
    buf_clk new_AGEMA_reg_buffer_1771 ( .C (clk), .D (new_AGEMA_signal_5201), .Q (new_AGEMA_signal_5202) ) ;
    buf_clk new_AGEMA_reg_buffer_1773 ( .C (clk), .D (new_AGEMA_signal_5203), .Q (new_AGEMA_signal_5204) ) ;
    buf_clk new_AGEMA_reg_buffer_1775 ( .C (clk), .D (new_AGEMA_signal_5205), .Q (new_AGEMA_signal_5206) ) ;
    buf_clk new_AGEMA_reg_buffer_1777 ( .C (clk), .D (new_AGEMA_signal_5207), .Q (new_AGEMA_signal_5208) ) ;
    buf_clk new_AGEMA_reg_buffer_1779 ( .C (clk), .D (new_AGEMA_signal_5209), .Q (new_AGEMA_signal_5210) ) ;
    buf_clk new_AGEMA_reg_buffer_1781 ( .C (clk), .D (new_AGEMA_signal_5211), .Q (new_AGEMA_signal_5212) ) ;
    buf_clk new_AGEMA_reg_buffer_1783 ( .C (clk), .D (new_AGEMA_signal_5213), .Q (new_AGEMA_signal_5214) ) ;
    buf_clk new_AGEMA_reg_buffer_1785 ( .C (clk), .D (new_AGEMA_signal_5215), .Q (new_AGEMA_signal_5216) ) ;
    buf_clk new_AGEMA_reg_buffer_1787 ( .C (clk), .D (new_AGEMA_signal_5217), .Q (new_AGEMA_signal_5218) ) ;
    buf_clk new_AGEMA_reg_buffer_1789 ( .C (clk), .D (new_AGEMA_signal_5219), .Q (new_AGEMA_signal_5220) ) ;
    buf_clk new_AGEMA_reg_buffer_1791 ( .C (clk), .D (new_AGEMA_signal_5221), .Q (new_AGEMA_signal_5222) ) ;
    buf_clk new_AGEMA_reg_buffer_1793 ( .C (clk), .D (new_AGEMA_signal_5223), .Q (new_AGEMA_signal_5224) ) ;
    buf_clk new_AGEMA_reg_buffer_1795 ( .C (clk), .D (new_AGEMA_signal_5225), .Q (new_AGEMA_signal_5226) ) ;
    buf_clk new_AGEMA_reg_buffer_1797 ( .C (clk), .D (new_AGEMA_signal_5227), .Q (new_AGEMA_signal_5228) ) ;
    buf_clk new_AGEMA_reg_buffer_1799 ( .C (clk), .D (new_AGEMA_signal_5229), .Q (new_AGEMA_signal_5230) ) ;
    buf_clk new_AGEMA_reg_buffer_1801 ( .C (clk), .D (new_AGEMA_signal_5231), .Q (new_AGEMA_signal_5232) ) ;
    buf_clk new_AGEMA_reg_buffer_1803 ( .C (clk), .D (new_AGEMA_signal_5233), .Q (new_AGEMA_signal_5234) ) ;
    buf_clk new_AGEMA_reg_buffer_1805 ( .C (clk), .D (new_AGEMA_signal_5235), .Q (new_AGEMA_signal_5236) ) ;
    buf_clk new_AGEMA_reg_buffer_1807 ( .C (clk), .D (new_AGEMA_signal_5237), .Q (new_AGEMA_signal_5238) ) ;
    buf_clk new_AGEMA_reg_buffer_1809 ( .C (clk), .D (new_AGEMA_signal_5239), .Q (new_AGEMA_signal_5240) ) ;
    buf_clk new_AGEMA_reg_buffer_1811 ( .C (clk), .D (new_AGEMA_signal_5241), .Q (new_AGEMA_signal_5242) ) ;
    buf_clk new_AGEMA_reg_buffer_1813 ( .C (clk), .D (new_AGEMA_signal_5243), .Q (new_AGEMA_signal_5244) ) ;
    buf_clk new_AGEMA_reg_buffer_1815 ( .C (clk), .D (new_AGEMA_signal_5245), .Q (new_AGEMA_signal_5246) ) ;
    buf_clk new_AGEMA_reg_buffer_1817 ( .C (clk), .D (new_AGEMA_signal_5247), .Q (new_AGEMA_signal_5248) ) ;
    buf_clk new_AGEMA_reg_buffer_1819 ( .C (clk), .D (new_AGEMA_signal_5249), .Q (new_AGEMA_signal_5250) ) ;
    buf_clk new_AGEMA_reg_buffer_1821 ( .C (clk), .D (new_AGEMA_signal_5251), .Q (new_AGEMA_signal_5252) ) ;
    buf_clk new_AGEMA_reg_buffer_1823 ( .C (clk), .D (new_AGEMA_signal_5253), .Q (new_AGEMA_signal_5254) ) ;
    buf_clk new_AGEMA_reg_buffer_1825 ( .C (clk), .D (new_AGEMA_signal_5255), .Q (new_AGEMA_signal_5256) ) ;
    buf_clk new_AGEMA_reg_buffer_1827 ( .C (clk), .D (new_AGEMA_signal_5257), .Q (new_AGEMA_signal_5258) ) ;
    buf_clk new_AGEMA_reg_buffer_1829 ( .C (clk), .D (new_AGEMA_signal_5259), .Q (new_AGEMA_signal_5260) ) ;
    buf_clk new_AGEMA_reg_buffer_1831 ( .C (clk), .D (new_AGEMA_signal_5261), .Q (new_AGEMA_signal_5262) ) ;
    buf_clk new_AGEMA_reg_buffer_1833 ( .C (clk), .D (new_AGEMA_signal_5263), .Q (new_AGEMA_signal_5264) ) ;
    buf_clk new_AGEMA_reg_buffer_1835 ( .C (clk), .D (new_AGEMA_signal_5265), .Q (new_AGEMA_signal_5266) ) ;
    buf_clk new_AGEMA_reg_buffer_1837 ( .C (clk), .D (new_AGEMA_signal_5267), .Q (new_AGEMA_signal_5268) ) ;
    buf_clk new_AGEMA_reg_buffer_1839 ( .C (clk), .D (new_AGEMA_signal_5269), .Q (new_AGEMA_signal_5270) ) ;
    buf_clk new_AGEMA_reg_buffer_1841 ( .C (clk), .D (new_AGEMA_signal_5271), .Q (new_AGEMA_signal_5272) ) ;
    buf_clk new_AGEMA_reg_buffer_1843 ( .C (clk), .D (new_AGEMA_signal_5273), .Q (new_AGEMA_signal_5274) ) ;
    buf_clk new_AGEMA_reg_buffer_1845 ( .C (clk), .D (new_AGEMA_signal_5275), .Q (new_AGEMA_signal_5276) ) ;
    buf_clk new_AGEMA_reg_buffer_1847 ( .C (clk), .D (new_AGEMA_signal_5277), .Q (new_AGEMA_signal_5278) ) ;
    buf_clk new_AGEMA_reg_buffer_1849 ( .C (clk), .D (new_AGEMA_signal_5279), .Q (new_AGEMA_signal_5280) ) ;
    buf_clk new_AGEMA_reg_buffer_1851 ( .C (clk), .D (new_AGEMA_signal_5281), .Q (new_AGEMA_signal_5282) ) ;
    buf_clk new_AGEMA_reg_buffer_1853 ( .C (clk), .D (new_AGEMA_signal_5283), .Q (new_AGEMA_signal_5284) ) ;
    buf_clk new_AGEMA_reg_buffer_1855 ( .C (clk), .D (new_AGEMA_signal_5285), .Q (new_AGEMA_signal_5286) ) ;
    buf_clk new_AGEMA_reg_buffer_1857 ( .C (clk), .D (new_AGEMA_signal_5287), .Q (new_AGEMA_signal_5288) ) ;
    buf_clk new_AGEMA_reg_buffer_1859 ( .C (clk), .D (new_AGEMA_signal_5289), .Q (new_AGEMA_signal_5290) ) ;
    buf_clk new_AGEMA_reg_buffer_1861 ( .C (clk), .D (new_AGEMA_signal_5291), .Q (new_AGEMA_signal_5292) ) ;
    buf_clk new_AGEMA_reg_buffer_1863 ( .C (clk), .D (new_AGEMA_signal_5293), .Q (new_AGEMA_signal_5294) ) ;
    buf_clk new_AGEMA_reg_buffer_1865 ( .C (clk), .D (new_AGEMA_signal_5295), .Q (new_AGEMA_signal_5296) ) ;
    buf_clk new_AGEMA_reg_buffer_1867 ( .C (clk), .D (new_AGEMA_signal_5297), .Q (new_AGEMA_signal_5298) ) ;
    buf_clk new_AGEMA_reg_buffer_1869 ( .C (clk), .D (new_AGEMA_signal_5299), .Q (new_AGEMA_signal_5300) ) ;
    buf_clk new_AGEMA_reg_buffer_1871 ( .C (clk), .D (new_AGEMA_signal_5301), .Q (new_AGEMA_signal_5302) ) ;
    buf_clk new_AGEMA_reg_buffer_1873 ( .C (clk), .D (new_AGEMA_signal_5303), .Q (new_AGEMA_signal_5304) ) ;
    buf_clk new_AGEMA_reg_buffer_1875 ( .C (clk), .D (new_AGEMA_signal_5305), .Q (new_AGEMA_signal_5306) ) ;
    buf_clk new_AGEMA_reg_buffer_1877 ( .C (clk), .D (new_AGEMA_signal_5307), .Q (new_AGEMA_signal_5308) ) ;
    buf_clk new_AGEMA_reg_buffer_1879 ( .C (clk), .D (new_AGEMA_signal_5309), .Q (new_AGEMA_signal_5310) ) ;
    buf_clk new_AGEMA_reg_buffer_1881 ( .C (clk), .D (new_AGEMA_signal_5311), .Q (new_AGEMA_signal_5312) ) ;
    buf_clk new_AGEMA_reg_buffer_1883 ( .C (clk), .D (new_AGEMA_signal_5313), .Q (new_AGEMA_signal_5314) ) ;
    buf_clk new_AGEMA_reg_buffer_1885 ( .C (clk), .D (new_AGEMA_signal_5315), .Q (new_AGEMA_signal_5316) ) ;
    buf_clk new_AGEMA_reg_buffer_1887 ( .C (clk), .D (new_AGEMA_signal_5317), .Q (new_AGEMA_signal_5318) ) ;
    buf_clk new_AGEMA_reg_buffer_1889 ( .C (clk), .D (new_AGEMA_signal_5319), .Q (new_AGEMA_signal_5320) ) ;
    buf_clk new_AGEMA_reg_buffer_1891 ( .C (clk), .D (new_AGEMA_signal_5321), .Q (new_AGEMA_signal_5322) ) ;
    buf_clk new_AGEMA_reg_buffer_1893 ( .C (clk), .D (new_AGEMA_signal_5323), .Q (new_AGEMA_signal_5324) ) ;
    buf_clk new_AGEMA_reg_buffer_1895 ( .C (clk), .D (new_AGEMA_signal_5325), .Q (new_AGEMA_signal_5326) ) ;
    buf_clk new_AGEMA_reg_buffer_1897 ( .C (clk), .D (new_AGEMA_signal_5327), .Q (new_AGEMA_signal_5328) ) ;
    buf_clk new_AGEMA_reg_buffer_1899 ( .C (clk), .D (new_AGEMA_signal_5329), .Q (new_AGEMA_signal_5330) ) ;
    buf_clk new_AGEMA_reg_buffer_1901 ( .C (clk), .D (new_AGEMA_signal_5331), .Q (new_AGEMA_signal_5332) ) ;
    buf_clk new_AGEMA_reg_buffer_1905 ( .C (clk), .D (new_AGEMA_signal_5335), .Q (new_AGEMA_signal_5336) ) ;
    buf_clk new_AGEMA_reg_buffer_1909 ( .C (clk), .D (new_AGEMA_signal_5339), .Q (new_AGEMA_signal_5340) ) ;
    buf_clk new_AGEMA_reg_buffer_1913 ( .C (clk), .D (new_AGEMA_signal_5343), .Q (new_AGEMA_signal_5344) ) ;
    buf_clk new_AGEMA_reg_buffer_1917 ( .C (clk), .D (new_AGEMA_signal_5347), .Q (new_AGEMA_signal_5348) ) ;
    buf_clk new_AGEMA_reg_buffer_1921 ( .C (clk), .D (new_AGEMA_signal_5351), .Q (new_AGEMA_signal_5352) ) ;
    buf_clk new_AGEMA_reg_buffer_1925 ( .C (clk), .D (new_AGEMA_signal_5355), .Q (new_AGEMA_signal_5356) ) ;
    buf_clk new_AGEMA_reg_buffer_1929 ( .C (clk), .D (new_AGEMA_signal_5359), .Q (new_AGEMA_signal_5360) ) ;
    buf_clk new_AGEMA_reg_buffer_1933 ( .C (clk), .D (new_AGEMA_signal_5363), .Q (new_AGEMA_signal_5364) ) ;
    buf_clk new_AGEMA_reg_buffer_1937 ( .C (clk), .D (new_AGEMA_signal_5367), .Q (new_AGEMA_signal_5368) ) ;
    buf_clk new_AGEMA_reg_buffer_1941 ( .C (clk), .D (new_AGEMA_signal_5371), .Q (new_AGEMA_signal_5372) ) ;
    buf_clk new_AGEMA_reg_buffer_1945 ( .C (clk), .D (new_AGEMA_signal_5375), .Q (new_AGEMA_signal_5376) ) ;
    buf_clk new_AGEMA_reg_buffer_1949 ( .C (clk), .D (new_AGEMA_signal_5379), .Q (new_AGEMA_signal_5380) ) ;
    buf_clk new_AGEMA_reg_buffer_1953 ( .C (clk), .D (new_AGEMA_signal_5383), .Q (new_AGEMA_signal_5384) ) ;
    buf_clk new_AGEMA_reg_buffer_1957 ( .C (clk), .D (new_AGEMA_signal_5387), .Q (new_AGEMA_signal_5388) ) ;
    buf_clk new_AGEMA_reg_buffer_1961 ( .C (clk), .D (new_AGEMA_signal_5391), .Q (new_AGEMA_signal_5392) ) ;
    buf_clk new_AGEMA_reg_buffer_1965 ( .C (clk), .D (new_AGEMA_signal_5395), .Q (new_AGEMA_signal_5396) ) ;
    buf_clk new_AGEMA_reg_buffer_1969 ( .C (clk), .D (new_AGEMA_signal_5399), .Q (new_AGEMA_signal_5400) ) ;
    buf_clk new_AGEMA_reg_buffer_1973 ( .C (clk), .D (new_AGEMA_signal_5403), .Q (new_AGEMA_signal_5404) ) ;
    buf_clk new_AGEMA_reg_buffer_1977 ( .C (clk), .D (new_AGEMA_signal_5407), .Q (new_AGEMA_signal_5408) ) ;
    buf_clk new_AGEMA_reg_buffer_1981 ( .C (clk), .D (new_AGEMA_signal_5411), .Q (new_AGEMA_signal_5412) ) ;
    buf_clk new_AGEMA_reg_buffer_1985 ( .C (clk), .D (new_AGEMA_signal_5415), .Q (new_AGEMA_signal_5416) ) ;
    buf_clk new_AGEMA_reg_buffer_1989 ( .C (clk), .D (new_AGEMA_signal_5419), .Q (new_AGEMA_signal_5420) ) ;
    buf_clk new_AGEMA_reg_buffer_1993 ( .C (clk), .D (new_AGEMA_signal_5423), .Q (new_AGEMA_signal_5424) ) ;
    buf_clk new_AGEMA_reg_buffer_1997 ( .C (clk), .D (new_AGEMA_signal_5427), .Q (new_AGEMA_signal_5428) ) ;
    buf_clk new_AGEMA_reg_buffer_2001 ( .C (clk), .D (new_AGEMA_signal_5431), .Q (new_AGEMA_signal_5432) ) ;
    buf_clk new_AGEMA_reg_buffer_2005 ( .C (clk), .D (new_AGEMA_signal_5435), .Q (new_AGEMA_signal_5436) ) ;
    buf_clk new_AGEMA_reg_buffer_2009 ( .C (clk), .D (new_AGEMA_signal_5439), .Q (new_AGEMA_signal_5440) ) ;
    buf_clk new_AGEMA_reg_buffer_2013 ( .C (clk), .D (new_AGEMA_signal_5443), .Q (new_AGEMA_signal_5444) ) ;
    buf_clk new_AGEMA_reg_buffer_2017 ( .C (clk), .D (new_AGEMA_signal_5447), .Q (new_AGEMA_signal_5448) ) ;
    buf_clk new_AGEMA_reg_buffer_2021 ( .C (clk), .D (new_AGEMA_signal_5451), .Q (new_AGEMA_signal_5452) ) ;
    buf_clk new_AGEMA_reg_buffer_2025 ( .C (clk), .D (new_AGEMA_signal_5455), .Q (new_AGEMA_signal_5456) ) ;
    buf_clk new_AGEMA_reg_buffer_2029 ( .C (clk), .D (new_AGEMA_signal_5459), .Q (new_AGEMA_signal_5460) ) ;
    buf_clk new_AGEMA_reg_buffer_2033 ( .C (clk), .D (new_AGEMA_signal_5463), .Q (new_AGEMA_signal_5464) ) ;
    buf_clk new_AGEMA_reg_buffer_2037 ( .C (clk), .D (new_AGEMA_signal_5467), .Q (new_AGEMA_signal_5468) ) ;
    buf_clk new_AGEMA_reg_buffer_2041 ( .C (clk), .D (new_AGEMA_signal_5471), .Q (new_AGEMA_signal_5472) ) ;
    buf_clk new_AGEMA_reg_buffer_2045 ( .C (clk), .D (new_AGEMA_signal_5475), .Q (new_AGEMA_signal_5476) ) ;
    buf_clk new_AGEMA_reg_buffer_2049 ( .C (clk), .D (new_AGEMA_signal_5479), .Q (new_AGEMA_signal_5480) ) ;
    buf_clk new_AGEMA_reg_buffer_2053 ( .C (clk), .D (new_AGEMA_signal_5483), .Q (new_AGEMA_signal_5484) ) ;
    buf_clk new_AGEMA_reg_buffer_2057 ( .C (clk), .D (new_AGEMA_signal_5487), .Q (new_AGEMA_signal_5488) ) ;
    buf_clk new_AGEMA_reg_buffer_2061 ( .C (clk), .D (new_AGEMA_signal_5491), .Q (new_AGEMA_signal_5492) ) ;
    buf_clk new_AGEMA_reg_buffer_2065 ( .C (clk), .D (new_AGEMA_signal_5495), .Q (new_AGEMA_signal_5496) ) ;
    buf_clk new_AGEMA_reg_buffer_2069 ( .C (clk), .D (new_AGEMA_signal_5499), .Q (new_AGEMA_signal_5500) ) ;
    buf_clk new_AGEMA_reg_buffer_2073 ( .C (clk), .D (new_AGEMA_signal_5503), .Q (new_AGEMA_signal_5504) ) ;
    buf_clk new_AGEMA_reg_buffer_2077 ( .C (clk), .D (new_AGEMA_signal_5507), .Q (new_AGEMA_signal_5508) ) ;
    buf_clk new_AGEMA_reg_buffer_2081 ( .C (clk), .D (new_AGEMA_signal_5511), .Q (new_AGEMA_signal_5512) ) ;
    buf_clk new_AGEMA_reg_buffer_2085 ( .C (clk), .D (new_AGEMA_signal_5515), .Q (new_AGEMA_signal_5516) ) ;
    buf_clk new_AGEMA_reg_buffer_2089 ( .C (clk), .D (new_AGEMA_signal_5519), .Q (new_AGEMA_signal_5520) ) ;
    buf_clk new_AGEMA_reg_buffer_2093 ( .C (clk), .D (new_AGEMA_signal_5523), .Q (new_AGEMA_signal_5524) ) ;
    buf_clk new_AGEMA_reg_buffer_2097 ( .C (clk), .D (new_AGEMA_signal_5527), .Q (new_AGEMA_signal_5528) ) ;
    buf_clk new_AGEMA_reg_buffer_2101 ( .C (clk), .D (new_AGEMA_signal_5531), .Q (new_AGEMA_signal_5532) ) ;
    buf_clk new_AGEMA_reg_buffer_2105 ( .C (clk), .D (new_AGEMA_signal_5535), .Q (new_AGEMA_signal_5536) ) ;
    buf_clk new_AGEMA_reg_buffer_2109 ( .C (clk), .D (new_AGEMA_signal_5539), .Q (new_AGEMA_signal_5540) ) ;
    buf_clk new_AGEMA_reg_buffer_2113 ( .C (clk), .D (new_AGEMA_signal_5543), .Q (new_AGEMA_signal_5544) ) ;
    buf_clk new_AGEMA_reg_buffer_2117 ( .C (clk), .D (new_AGEMA_signal_5547), .Q (new_AGEMA_signal_5548) ) ;
    buf_clk new_AGEMA_reg_buffer_2121 ( .C (clk), .D (new_AGEMA_signal_5551), .Q (new_AGEMA_signal_5552) ) ;
    buf_clk new_AGEMA_reg_buffer_2125 ( .C (clk), .D (new_AGEMA_signal_5555), .Q (new_AGEMA_signal_5556) ) ;
    buf_clk new_AGEMA_reg_buffer_2129 ( .C (clk), .D (new_AGEMA_signal_5559), .Q (new_AGEMA_signal_5560) ) ;
    buf_clk new_AGEMA_reg_buffer_2133 ( .C (clk), .D (new_AGEMA_signal_5563), .Q (new_AGEMA_signal_5564) ) ;
    buf_clk new_AGEMA_reg_buffer_2137 ( .C (clk), .D (new_AGEMA_signal_5567), .Q (new_AGEMA_signal_5568) ) ;
    buf_clk new_AGEMA_reg_buffer_2141 ( .C (clk), .D (new_AGEMA_signal_5571), .Q (new_AGEMA_signal_5572) ) ;
    buf_clk new_AGEMA_reg_buffer_2145 ( .C (clk), .D (new_AGEMA_signal_5575), .Q (new_AGEMA_signal_5576) ) ;
    buf_clk new_AGEMA_reg_buffer_2149 ( .C (clk), .D (new_AGEMA_signal_5579), .Q (new_AGEMA_signal_5580) ) ;
    buf_clk new_AGEMA_reg_buffer_2153 ( .C (clk), .D (new_AGEMA_signal_5583), .Q (new_AGEMA_signal_5584) ) ;
    buf_clk new_AGEMA_reg_buffer_2157 ( .C (clk), .D (new_AGEMA_signal_5587), .Q (new_AGEMA_signal_5588) ) ;
    buf_clk new_AGEMA_reg_buffer_2161 ( .C (clk), .D (new_AGEMA_signal_5591), .Q (new_AGEMA_signal_5592) ) ;
    buf_clk new_AGEMA_reg_buffer_2165 ( .C (clk), .D (new_AGEMA_signal_5595), .Q (new_AGEMA_signal_5596) ) ;
    buf_clk new_AGEMA_reg_buffer_2169 ( .C (clk), .D (new_AGEMA_signal_5599), .Q (new_AGEMA_signal_5600) ) ;
    buf_clk new_AGEMA_reg_buffer_2173 ( .C (clk), .D (new_AGEMA_signal_5603), .Q (new_AGEMA_signal_5604) ) ;
    buf_clk new_AGEMA_reg_buffer_2177 ( .C (clk), .D (new_AGEMA_signal_5607), .Q (new_AGEMA_signal_5608) ) ;
    buf_clk new_AGEMA_reg_buffer_2181 ( .C (clk), .D (new_AGEMA_signal_5611), .Q (new_AGEMA_signal_5612) ) ;
    buf_clk new_AGEMA_reg_buffer_2185 ( .C (clk), .D (new_AGEMA_signal_5615), .Q (new_AGEMA_signal_5616) ) ;
    buf_clk new_AGEMA_reg_buffer_2189 ( .C (clk), .D (new_AGEMA_signal_5619), .Q (new_AGEMA_signal_5620) ) ;
    buf_clk new_AGEMA_reg_buffer_2193 ( .C (clk), .D (new_AGEMA_signal_5623), .Q (new_AGEMA_signal_5624) ) ;
    buf_clk new_AGEMA_reg_buffer_2197 ( .C (clk), .D (new_AGEMA_signal_5627), .Q (new_AGEMA_signal_5628) ) ;
    buf_clk new_AGEMA_reg_buffer_2201 ( .C (clk), .D (new_AGEMA_signal_5631), .Q (new_AGEMA_signal_5632) ) ;
    buf_clk new_AGEMA_reg_buffer_2205 ( .C (clk), .D (new_AGEMA_signal_5635), .Q (new_AGEMA_signal_5636) ) ;
    buf_clk new_AGEMA_reg_buffer_2209 ( .C (clk), .D (new_AGEMA_signal_5639), .Q (new_AGEMA_signal_5640) ) ;
    buf_clk new_AGEMA_reg_buffer_2213 ( .C (clk), .D (new_AGEMA_signal_5643), .Q (new_AGEMA_signal_5644) ) ;
    buf_clk new_AGEMA_reg_buffer_2217 ( .C (clk), .D (new_AGEMA_signal_5647), .Q (new_AGEMA_signal_5648) ) ;
    buf_clk new_AGEMA_reg_buffer_2221 ( .C (clk), .D (new_AGEMA_signal_5651), .Q (new_AGEMA_signal_5652) ) ;
    buf_clk new_AGEMA_reg_buffer_2225 ( .C (clk), .D (new_AGEMA_signal_5655), .Q (new_AGEMA_signal_5656) ) ;
    buf_clk new_AGEMA_reg_buffer_2229 ( .C (clk), .D (new_AGEMA_signal_5659), .Q (new_AGEMA_signal_5660) ) ;
    buf_clk new_AGEMA_reg_buffer_2233 ( .C (clk), .D (new_AGEMA_signal_5663), .Q (new_AGEMA_signal_5664) ) ;
    buf_clk new_AGEMA_reg_buffer_2237 ( .C (clk), .D (new_AGEMA_signal_5667), .Q (new_AGEMA_signal_5668) ) ;
    buf_clk new_AGEMA_reg_buffer_2241 ( .C (clk), .D (new_AGEMA_signal_5671), .Q (new_AGEMA_signal_5672) ) ;
    buf_clk new_AGEMA_reg_buffer_2245 ( .C (clk), .D (new_AGEMA_signal_5675), .Q (new_AGEMA_signal_5676) ) ;
    buf_clk new_AGEMA_reg_buffer_2249 ( .C (clk), .D (new_AGEMA_signal_5679), .Q (new_AGEMA_signal_5680) ) ;
    buf_clk new_AGEMA_reg_buffer_2253 ( .C (clk), .D (new_AGEMA_signal_5683), .Q (new_AGEMA_signal_5684) ) ;
    buf_clk new_AGEMA_reg_buffer_2257 ( .C (clk), .D (new_AGEMA_signal_5687), .Q (new_AGEMA_signal_5688) ) ;
    buf_clk new_AGEMA_reg_buffer_2261 ( .C (clk), .D (new_AGEMA_signal_5691), .Q (new_AGEMA_signal_5692) ) ;
    buf_clk new_AGEMA_reg_buffer_2265 ( .C (clk), .D (new_AGEMA_signal_5695), .Q (new_AGEMA_signal_5696) ) ;
    buf_clk new_AGEMA_reg_buffer_2269 ( .C (clk), .D (new_AGEMA_signal_5699), .Q (new_AGEMA_signal_5700) ) ;
    buf_clk new_AGEMA_reg_buffer_2273 ( .C (clk), .D (new_AGEMA_signal_5703), .Q (new_AGEMA_signal_5704) ) ;
    buf_clk new_AGEMA_reg_buffer_2277 ( .C (clk), .D (new_AGEMA_signal_5707), .Q (new_AGEMA_signal_5708) ) ;
    buf_clk new_AGEMA_reg_buffer_2281 ( .C (clk), .D (new_AGEMA_signal_5711), .Q (new_AGEMA_signal_5712) ) ;
    buf_clk new_AGEMA_reg_buffer_2285 ( .C (clk), .D (new_AGEMA_signal_5715), .Q (new_AGEMA_signal_5716) ) ;
    buf_clk new_AGEMA_reg_buffer_2289 ( .C (clk), .D (new_AGEMA_signal_5719), .Q (new_AGEMA_signal_5720) ) ;
    buf_clk new_AGEMA_reg_buffer_2293 ( .C (clk), .D (new_AGEMA_signal_5723), .Q (new_AGEMA_signal_5724) ) ;
    buf_clk new_AGEMA_reg_buffer_2297 ( .C (clk), .D (new_AGEMA_signal_5727), .Q (new_AGEMA_signal_5728) ) ;
    buf_clk new_AGEMA_reg_buffer_2301 ( .C (clk), .D (new_AGEMA_signal_5731), .Q (new_AGEMA_signal_5732) ) ;
    buf_clk new_AGEMA_reg_buffer_2305 ( .C (clk), .D (new_AGEMA_signal_5735), .Q (new_AGEMA_signal_5736) ) ;
    buf_clk new_AGEMA_reg_buffer_2309 ( .C (clk), .D (new_AGEMA_signal_5739), .Q (new_AGEMA_signal_5740) ) ;
    buf_clk new_AGEMA_reg_buffer_2313 ( .C (clk), .D (new_AGEMA_signal_5743), .Q (new_AGEMA_signal_5744) ) ;
    buf_clk new_AGEMA_reg_buffer_2317 ( .C (clk), .D (new_AGEMA_signal_5747), .Q (new_AGEMA_signal_5748) ) ;
    buf_clk new_AGEMA_reg_buffer_2321 ( .C (clk), .D (new_AGEMA_signal_5751), .Q (new_AGEMA_signal_5752) ) ;
    buf_clk new_AGEMA_reg_buffer_2325 ( .C (clk), .D (new_AGEMA_signal_5755), .Q (new_AGEMA_signal_5756) ) ;
    buf_clk new_AGEMA_reg_buffer_2329 ( .C (clk), .D (new_AGEMA_signal_5759), .Q (new_AGEMA_signal_5760) ) ;
    buf_clk new_AGEMA_reg_buffer_2333 ( .C (clk), .D (new_AGEMA_signal_5763), .Q (new_AGEMA_signal_5764) ) ;
    buf_clk new_AGEMA_reg_buffer_2337 ( .C (clk), .D (new_AGEMA_signal_5767), .Q (new_AGEMA_signal_5768) ) ;
    buf_clk new_AGEMA_reg_buffer_2341 ( .C (clk), .D (new_AGEMA_signal_5771), .Q (new_AGEMA_signal_5772) ) ;
    buf_clk new_AGEMA_reg_buffer_2345 ( .C (clk), .D (new_AGEMA_signal_5775), .Q (new_AGEMA_signal_5776) ) ;
    buf_clk new_AGEMA_reg_buffer_2349 ( .C (clk), .D (new_AGEMA_signal_5779), .Q (new_AGEMA_signal_5780) ) ;
    buf_clk new_AGEMA_reg_buffer_2353 ( .C (clk), .D (new_AGEMA_signal_5783), .Q (new_AGEMA_signal_5784) ) ;
    buf_clk new_AGEMA_reg_buffer_2357 ( .C (clk), .D (new_AGEMA_signal_5787), .Q (new_AGEMA_signal_5788) ) ;
    buf_clk new_AGEMA_reg_buffer_2361 ( .C (clk), .D (new_AGEMA_signal_5791), .Q (new_AGEMA_signal_5792) ) ;
    buf_clk new_AGEMA_reg_buffer_2365 ( .C (clk), .D (new_AGEMA_signal_5795), .Q (new_AGEMA_signal_5796) ) ;
    buf_clk new_AGEMA_reg_buffer_2369 ( .C (clk), .D (new_AGEMA_signal_5799), .Q (new_AGEMA_signal_5800) ) ;
    buf_clk new_AGEMA_reg_buffer_2373 ( .C (clk), .D (new_AGEMA_signal_5803), .Q (new_AGEMA_signal_5804) ) ;
    buf_clk new_AGEMA_reg_buffer_2377 ( .C (clk), .D (new_AGEMA_signal_5807), .Q (new_AGEMA_signal_5808) ) ;
    buf_clk new_AGEMA_reg_buffer_2381 ( .C (clk), .D (new_AGEMA_signal_5811), .Q (new_AGEMA_signal_5812) ) ;
    buf_clk new_AGEMA_reg_buffer_2385 ( .C (clk), .D (new_AGEMA_signal_5815), .Q (new_AGEMA_signal_5816) ) ;
    buf_clk new_AGEMA_reg_buffer_2389 ( .C (clk), .D (new_AGEMA_signal_5819), .Q (new_AGEMA_signal_5820) ) ;
    buf_clk new_AGEMA_reg_buffer_2393 ( .C (clk), .D (new_AGEMA_signal_5823), .Q (new_AGEMA_signal_5824) ) ;
    buf_clk new_AGEMA_reg_buffer_2397 ( .C (clk), .D (new_AGEMA_signal_5827), .Q (new_AGEMA_signal_5828) ) ;
    buf_clk new_AGEMA_reg_buffer_2401 ( .C (clk), .D (new_AGEMA_signal_5831), .Q (new_AGEMA_signal_5832) ) ;
    buf_clk new_AGEMA_reg_buffer_2405 ( .C (clk), .D (new_AGEMA_signal_5835), .Q (new_AGEMA_signal_5836) ) ;
    buf_clk new_AGEMA_reg_buffer_2409 ( .C (clk), .D (new_AGEMA_signal_5839), .Q (new_AGEMA_signal_5840) ) ;
    buf_clk new_AGEMA_reg_buffer_2413 ( .C (clk), .D (new_AGEMA_signal_5843), .Q (new_AGEMA_signal_5844) ) ;
    buf_clk new_AGEMA_reg_buffer_2417 ( .C (clk), .D (new_AGEMA_signal_5847), .Q (new_AGEMA_signal_5848) ) ;
    buf_clk new_AGEMA_reg_buffer_2419 ( .C (clk), .D (new_AGEMA_signal_5849), .Q (new_AGEMA_signal_5850) ) ;
    buf_clk new_AGEMA_reg_buffer_2421 ( .C (clk), .D (new_AGEMA_signal_5851), .Q (new_AGEMA_signal_5852) ) ;
    buf_clk new_AGEMA_reg_buffer_2423 ( .C (clk), .D (new_AGEMA_signal_5853), .Q (new_AGEMA_signal_5854) ) ;
    buf_clk new_AGEMA_reg_buffer_2433 ( .C (clk), .D (new_AGEMA_signal_5863), .Q (new_AGEMA_signal_5864) ) ;
    buf_clk new_AGEMA_reg_buffer_2435 ( .C (clk), .D (new_AGEMA_signal_5865), .Q (new_AGEMA_signal_5866) ) ;
    buf_clk new_AGEMA_reg_buffer_2437 ( .C (clk), .D (new_AGEMA_signal_5867), .Q (new_AGEMA_signal_5868) ) ;
    buf_clk new_AGEMA_reg_buffer_2439 ( .C (clk), .D (new_AGEMA_signal_5869), .Q (new_AGEMA_signal_5870) ) ;
    buf_clk new_AGEMA_reg_buffer_2441 ( .C (clk), .D (new_AGEMA_signal_5871), .Q (new_AGEMA_signal_5872) ) ;
    buf_clk new_AGEMA_reg_buffer_2445 ( .C (clk), .D (new_AGEMA_signal_5875), .Q (new_AGEMA_signal_5876) ) ;
    buf_clk new_AGEMA_reg_buffer_2449 ( .C (clk), .D (new_AGEMA_signal_5879), .Q (new_AGEMA_signal_5880) ) ;
    buf_clk new_AGEMA_reg_buffer_2453 ( .C (clk), .D (new_AGEMA_signal_5883), .Q (new_AGEMA_signal_5884) ) ;
    buf_clk new_AGEMA_reg_buffer_2465 ( .C (clk), .D (new_AGEMA_signal_5895), .Q (new_AGEMA_signal_5896) ) ;
    buf_clk new_AGEMA_reg_buffer_2467 ( .C (clk), .D (new_AGEMA_signal_5897), .Q (new_AGEMA_signal_5898) ) ;
    buf_clk new_AGEMA_reg_buffer_2469 ( .C (clk), .D (new_AGEMA_signal_5899), .Q (new_AGEMA_signal_5900) ) ;
    buf_clk new_AGEMA_reg_buffer_2471 ( .C (clk), .D (new_AGEMA_signal_5901), .Q (new_AGEMA_signal_5902) ) ;
    buf_clk new_AGEMA_reg_buffer_2481 ( .C (clk), .D (new_AGEMA_signal_5911), .Q (new_AGEMA_signal_5912) ) ;
    buf_clk new_AGEMA_reg_buffer_2483 ( .C (clk), .D (new_AGEMA_signal_5913), .Q (new_AGEMA_signal_5914) ) ;
    buf_clk new_AGEMA_reg_buffer_2485 ( .C (clk), .D (new_AGEMA_signal_5915), .Q (new_AGEMA_signal_5916) ) ;
    buf_clk new_AGEMA_reg_buffer_2487 ( .C (clk), .D (new_AGEMA_signal_5917), .Q (new_AGEMA_signal_5918) ) ;
    buf_clk new_AGEMA_reg_buffer_2489 ( .C (clk), .D (new_AGEMA_signal_5919), .Q (new_AGEMA_signal_5920) ) ;
    buf_clk new_AGEMA_reg_buffer_2493 ( .C (clk), .D (new_AGEMA_signal_5923), .Q (new_AGEMA_signal_5924) ) ;
    buf_clk new_AGEMA_reg_buffer_2497 ( .C (clk), .D (new_AGEMA_signal_5927), .Q (new_AGEMA_signal_5928) ) ;
    buf_clk new_AGEMA_reg_buffer_2501 ( .C (clk), .D (new_AGEMA_signal_5931), .Q (new_AGEMA_signal_5932) ) ;
    buf_clk new_AGEMA_reg_buffer_2513 ( .C (clk), .D (new_AGEMA_signal_5943), .Q (new_AGEMA_signal_5944) ) ;
    buf_clk new_AGEMA_reg_buffer_2515 ( .C (clk), .D (new_AGEMA_signal_5945), .Q (new_AGEMA_signal_5946) ) ;
    buf_clk new_AGEMA_reg_buffer_2517 ( .C (clk), .D (new_AGEMA_signal_5947), .Q (new_AGEMA_signal_5948) ) ;
    buf_clk new_AGEMA_reg_buffer_2519 ( .C (clk), .D (new_AGEMA_signal_5949), .Q (new_AGEMA_signal_5950) ) ;
    buf_clk new_AGEMA_reg_buffer_2529 ( .C (clk), .D (new_AGEMA_signal_5959), .Q (new_AGEMA_signal_5960) ) ;
    buf_clk new_AGEMA_reg_buffer_2531 ( .C (clk), .D (new_AGEMA_signal_5961), .Q (new_AGEMA_signal_5962) ) ;
    buf_clk new_AGEMA_reg_buffer_2533 ( .C (clk), .D (new_AGEMA_signal_5963), .Q (new_AGEMA_signal_5964) ) ;
    buf_clk new_AGEMA_reg_buffer_2535 ( .C (clk), .D (new_AGEMA_signal_5965), .Q (new_AGEMA_signal_5966) ) ;
    buf_clk new_AGEMA_reg_buffer_2537 ( .C (clk), .D (new_AGEMA_signal_5967), .Q (new_AGEMA_signal_5968) ) ;
    buf_clk new_AGEMA_reg_buffer_2541 ( .C (clk), .D (new_AGEMA_signal_5971), .Q (new_AGEMA_signal_5972) ) ;
    buf_clk new_AGEMA_reg_buffer_2545 ( .C (clk), .D (new_AGEMA_signal_5975), .Q (new_AGEMA_signal_5976) ) ;
    buf_clk new_AGEMA_reg_buffer_2549 ( .C (clk), .D (new_AGEMA_signal_5979), .Q (new_AGEMA_signal_5980) ) ;
    buf_clk new_AGEMA_reg_buffer_2561 ( .C (clk), .D (new_AGEMA_signal_5991), .Q (new_AGEMA_signal_5992) ) ;
    buf_clk new_AGEMA_reg_buffer_2563 ( .C (clk), .D (new_AGEMA_signal_5993), .Q (new_AGEMA_signal_5994) ) ;
    buf_clk new_AGEMA_reg_buffer_2565 ( .C (clk), .D (new_AGEMA_signal_5995), .Q (new_AGEMA_signal_5996) ) ;
    buf_clk new_AGEMA_reg_buffer_2567 ( .C (clk), .D (new_AGEMA_signal_5997), .Q (new_AGEMA_signal_5998) ) ;
    buf_clk new_AGEMA_reg_buffer_2577 ( .C (clk), .D (new_AGEMA_signal_6007), .Q (new_AGEMA_signal_6008) ) ;
    buf_clk new_AGEMA_reg_buffer_2579 ( .C (clk), .D (new_AGEMA_signal_6009), .Q (new_AGEMA_signal_6010) ) ;
    buf_clk new_AGEMA_reg_buffer_2581 ( .C (clk), .D (new_AGEMA_signal_6011), .Q (new_AGEMA_signal_6012) ) ;
    buf_clk new_AGEMA_reg_buffer_2583 ( .C (clk), .D (new_AGEMA_signal_6013), .Q (new_AGEMA_signal_6014) ) ;
    buf_clk new_AGEMA_reg_buffer_2585 ( .C (clk), .D (new_AGEMA_signal_6015), .Q (new_AGEMA_signal_6016) ) ;
    buf_clk new_AGEMA_reg_buffer_2589 ( .C (clk), .D (new_AGEMA_signal_6019), .Q (new_AGEMA_signal_6020) ) ;
    buf_clk new_AGEMA_reg_buffer_2593 ( .C (clk), .D (new_AGEMA_signal_6023), .Q (new_AGEMA_signal_6024) ) ;
    buf_clk new_AGEMA_reg_buffer_2597 ( .C (clk), .D (new_AGEMA_signal_6027), .Q (new_AGEMA_signal_6028) ) ;
    buf_clk new_AGEMA_reg_buffer_2609 ( .C (clk), .D (new_AGEMA_signal_6039), .Q (new_AGEMA_signal_6040) ) ;
    buf_clk new_AGEMA_reg_buffer_2611 ( .C (clk), .D (new_AGEMA_signal_6041), .Q (new_AGEMA_signal_6042) ) ;
    buf_clk new_AGEMA_reg_buffer_2613 ( .C (clk), .D (new_AGEMA_signal_6043), .Q (new_AGEMA_signal_6044) ) ;
    buf_clk new_AGEMA_reg_buffer_2615 ( .C (clk), .D (new_AGEMA_signal_6045), .Q (new_AGEMA_signal_6046) ) ;
    buf_clk new_AGEMA_reg_buffer_2625 ( .C (clk), .D (new_AGEMA_signal_6055), .Q (new_AGEMA_signal_6056) ) ;
    buf_clk new_AGEMA_reg_buffer_2627 ( .C (clk), .D (new_AGEMA_signal_6057), .Q (new_AGEMA_signal_6058) ) ;
    buf_clk new_AGEMA_reg_buffer_2629 ( .C (clk), .D (new_AGEMA_signal_6059), .Q (new_AGEMA_signal_6060) ) ;
    buf_clk new_AGEMA_reg_buffer_2631 ( .C (clk), .D (new_AGEMA_signal_6061), .Q (new_AGEMA_signal_6062) ) ;
    buf_clk new_AGEMA_reg_buffer_2633 ( .C (clk), .D (new_AGEMA_signal_6063), .Q (new_AGEMA_signal_6064) ) ;
    buf_clk new_AGEMA_reg_buffer_2637 ( .C (clk), .D (new_AGEMA_signal_6067), .Q (new_AGEMA_signal_6068) ) ;
    buf_clk new_AGEMA_reg_buffer_2641 ( .C (clk), .D (new_AGEMA_signal_6071), .Q (new_AGEMA_signal_6072) ) ;
    buf_clk new_AGEMA_reg_buffer_2645 ( .C (clk), .D (new_AGEMA_signal_6075), .Q (new_AGEMA_signal_6076) ) ;
    buf_clk new_AGEMA_reg_buffer_2657 ( .C (clk), .D (new_AGEMA_signal_6087), .Q (new_AGEMA_signal_6088) ) ;
    buf_clk new_AGEMA_reg_buffer_2659 ( .C (clk), .D (new_AGEMA_signal_6089), .Q (new_AGEMA_signal_6090) ) ;
    buf_clk new_AGEMA_reg_buffer_2661 ( .C (clk), .D (new_AGEMA_signal_6091), .Q (new_AGEMA_signal_6092) ) ;
    buf_clk new_AGEMA_reg_buffer_2663 ( .C (clk), .D (new_AGEMA_signal_6093), .Q (new_AGEMA_signal_6094) ) ;
    buf_clk new_AGEMA_reg_buffer_2673 ( .C (clk), .D (new_AGEMA_signal_6103), .Q (new_AGEMA_signal_6104) ) ;
    buf_clk new_AGEMA_reg_buffer_2675 ( .C (clk), .D (new_AGEMA_signal_6105), .Q (new_AGEMA_signal_6106) ) ;
    buf_clk new_AGEMA_reg_buffer_2677 ( .C (clk), .D (new_AGEMA_signal_6107), .Q (new_AGEMA_signal_6108) ) ;
    buf_clk new_AGEMA_reg_buffer_2679 ( .C (clk), .D (new_AGEMA_signal_6109), .Q (new_AGEMA_signal_6110) ) ;
    buf_clk new_AGEMA_reg_buffer_2681 ( .C (clk), .D (new_AGEMA_signal_6111), .Q (new_AGEMA_signal_6112) ) ;
    buf_clk new_AGEMA_reg_buffer_2685 ( .C (clk), .D (new_AGEMA_signal_6115), .Q (new_AGEMA_signal_6116) ) ;
    buf_clk new_AGEMA_reg_buffer_2689 ( .C (clk), .D (new_AGEMA_signal_6119), .Q (new_AGEMA_signal_6120) ) ;
    buf_clk new_AGEMA_reg_buffer_2693 ( .C (clk), .D (new_AGEMA_signal_6123), .Q (new_AGEMA_signal_6124) ) ;
    buf_clk new_AGEMA_reg_buffer_2705 ( .C (clk), .D (new_AGEMA_signal_6135), .Q (new_AGEMA_signal_6136) ) ;
    buf_clk new_AGEMA_reg_buffer_2707 ( .C (clk), .D (new_AGEMA_signal_6137), .Q (new_AGEMA_signal_6138) ) ;
    buf_clk new_AGEMA_reg_buffer_2709 ( .C (clk), .D (new_AGEMA_signal_6139), .Q (new_AGEMA_signal_6140) ) ;
    buf_clk new_AGEMA_reg_buffer_2711 ( .C (clk), .D (new_AGEMA_signal_6141), .Q (new_AGEMA_signal_6142) ) ;
    buf_clk new_AGEMA_reg_buffer_2721 ( .C (clk), .D (new_AGEMA_signal_6151), .Q (new_AGEMA_signal_6152) ) ;
    buf_clk new_AGEMA_reg_buffer_2723 ( .C (clk), .D (new_AGEMA_signal_6153), .Q (new_AGEMA_signal_6154) ) ;
    buf_clk new_AGEMA_reg_buffer_2725 ( .C (clk), .D (new_AGEMA_signal_6155), .Q (new_AGEMA_signal_6156) ) ;
    buf_clk new_AGEMA_reg_buffer_2727 ( .C (clk), .D (new_AGEMA_signal_6157), .Q (new_AGEMA_signal_6158) ) ;
    buf_clk new_AGEMA_reg_buffer_2729 ( .C (clk), .D (new_AGEMA_signal_6159), .Q (new_AGEMA_signal_6160) ) ;
    buf_clk new_AGEMA_reg_buffer_2733 ( .C (clk), .D (new_AGEMA_signal_6163), .Q (new_AGEMA_signal_6164) ) ;
    buf_clk new_AGEMA_reg_buffer_2737 ( .C (clk), .D (new_AGEMA_signal_6167), .Q (new_AGEMA_signal_6168) ) ;
    buf_clk new_AGEMA_reg_buffer_2741 ( .C (clk), .D (new_AGEMA_signal_6171), .Q (new_AGEMA_signal_6172) ) ;
    buf_clk new_AGEMA_reg_buffer_2753 ( .C (clk), .D (new_AGEMA_signal_6183), .Q (new_AGEMA_signal_6184) ) ;
    buf_clk new_AGEMA_reg_buffer_2755 ( .C (clk), .D (new_AGEMA_signal_6185), .Q (new_AGEMA_signal_6186) ) ;
    buf_clk new_AGEMA_reg_buffer_2757 ( .C (clk), .D (new_AGEMA_signal_6187), .Q (new_AGEMA_signal_6188) ) ;
    buf_clk new_AGEMA_reg_buffer_2759 ( .C (clk), .D (new_AGEMA_signal_6189), .Q (new_AGEMA_signal_6190) ) ;
    buf_clk new_AGEMA_reg_buffer_2769 ( .C (clk), .D (new_AGEMA_signal_6199), .Q (new_AGEMA_signal_6200) ) ;
    buf_clk new_AGEMA_reg_buffer_2771 ( .C (clk), .D (new_AGEMA_signal_6201), .Q (new_AGEMA_signal_6202) ) ;
    buf_clk new_AGEMA_reg_buffer_2773 ( .C (clk), .D (new_AGEMA_signal_6203), .Q (new_AGEMA_signal_6204) ) ;
    buf_clk new_AGEMA_reg_buffer_2775 ( .C (clk), .D (new_AGEMA_signal_6205), .Q (new_AGEMA_signal_6206) ) ;
    buf_clk new_AGEMA_reg_buffer_2777 ( .C (clk), .D (new_AGEMA_signal_6207), .Q (new_AGEMA_signal_6208) ) ;
    buf_clk new_AGEMA_reg_buffer_2781 ( .C (clk), .D (new_AGEMA_signal_6211), .Q (new_AGEMA_signal_6212) ) ;
    buf_clk new_AGEMA_reg_buffer_2785 ( .C (clk), .D (new_AGEMA_signal_6215), .Q (new_AGEMA_signal_6216) ) ;
    buf_clk new_AGEMA_reg_buffer_2789 ( .C (clk), .D (new_AGEMA_signal_6219), .Q (new_AGEMA_signal_6220) ) ;
    buf_clk new_AGEMA_reg_buffer_2801 ( .C (clk), .D (new_AGEMA_signal_6231), .Q (new_AGEMA_signal_6232) ) ;
    buf_clk new_AGEMA_reg_buffer_2803 ( .C (clk), .D (new_AGEMA_signal_6233), .Q (new_AGEMA_signal_6234) ) ;
    buf_clk new_AGEMA_reg_buffer_2805 ( .C (clk), .D (new_AGEMA_signal_6235), .Q (new_AGEMA_signal_6236) ) ;
    buf_clk new_AGEMA_reg_buffer_2807 ( .C (clk), .D (new_AGEMA_signal_6237), .Q (new_AGEMA_signal_6238) ) ;
    buf_clk new_AGEMA_reg_buffer_2817 ( .C (clk), .D (new_AGEMA_signal_6247), .Q (new_AGEMA_signal_6248) ) ;
    buf_clk new_AGEMA_reg_buffer_2819 ( .C (clk), .D (new_AGEMA_signal_6249), .Q (new_AGEMA_signal_6250) ) ;
    buf_clk new_AGEMA_reg_buffer_2821 ( .C (clk), .D (new_AGEMA_signal_6251), .Q (new_AGEMA_signal_6252) ) ;
    buf_clk new_AGEMA_reg_buffer_2823 ( .C (clk), .D (new_AGEMA_signal_6253), .Q (new_AGEMA_signal_6254) ) ;
    buf_clk new_AGEMA_reg_buffer_2825 ( .C (clk), .D (new_AGEMA_signal_6255), .Q (new_AGEMA_signal_6256) ) ;
    buf_clk new_AGEMA_reg_buffer_2829 ( .C (clk), .D (new_AGEMA_signal_6259), .Q (new_AGEMA_signal_6260) ) ;
    buf_clk new_AGEMA_reg_buffer_2833 ( .C (clk), .D (new_AGEMA_signal_6263), .Q (new_AGEMA_signal_6264) ) ;
    buf_clk new_AGEMA_reg_buffer_2837 ( .C (clk), .D (new_AGEMA_signal_6267), .Q (new_AGEMA_signal_6268) ) ;
    buf_clk new_AGEMA_reg_buffer_2849 ( .C (clk), .D (new_AGEMA_signal_6279), .Q (new_AGEMA_signal_6280) ) ;
    buf_clk new_AGEMA_reg_buffer_2851 ( .C (clk), .D (new_AGEMA_signal_6281), .Q (new_AGEMA_signal_6282) ) ;
    buf_clk new_AGEMA_reg_buffer_2853 ( .C (clk), .D (new_AGEMA_signal_6283), .Q (new_AGEMA_signal_6284) ) ;
    buf_clk new_AGEMA_reg_buffer_2855 ( .C (clk), .D (new_AGEMA_signal_6285), .Q (new_AGEMA_signal_6286) ) ;
    buf_clk new_AGEMA_reg_buffer_2865 ( .C (clk), .D (new_AGEMA_signal_6295), .Q (new_AGEMA_signal_6296) ) ;
    buf_clk new_AGEMA_reg_buffer_2867 ( .C (clk), .D (new_AGEMA_signal_6297), .Q (new_AGEMA_signal_6298) ) ;
    buf_clk new_AGEMA_reg_buffer_2869 ( .C (clk), .D (new_AGEMA_signal_6299), .Q (new_AGEMA_signal_6300) ) ;
    buf_clk new_AGEMA_reg_buffer_2871 ( .C (clk), .D (new_AGEMA_signal_6301), .Q (new_AGEMA_signal_6302) ) ;
    buf_clk new_AGEMA_reg_buffer_2873 ( .C (clk), .D (new_AGEMA_signal_6303), .Q (new_AGEMA_signal_6304) ) ;
    buf_clk new_AGEMA_reg_buffer_2877 ( .C (clk), .D (new_AGEMA_signal_6307), .Q (new_AGEMA_signal_6308) ) ;
    buf_clk new_AGEMA_reg_buffer_2881 ( .C (clk), .D (new_AGEMA_signal_6311), .Q (new_AGEMA_signal_6312) ) ;
    buf_clk new_AGEMA_reg_buffer_2885 ( .C (clk), .D (new_AGEMA_signal_6315), .Q (new_AGEMA_signal_6316) ) ;
    buf_clk new_AGEMA_reg_buffer_2897 ( .C (clk), .D (new_AGEMA_signal_6327), .Q (new_AGEMA_signal_6328) ) ;
    buf_clk new_AGEMA_reg_buffer_2899 ( .C (clk), .D (new_AGEMA_signal_6329), .Q (new_AGEMA_signal_6330) ) ;
    buf_clk new_AGEMA_reg_buffer_2901 ( .C (clk), .D (new_AGEMA_signal_6331), .Q (new_AGEMA_signal_6332) ) ;
    buf_clk new_AGEMA_reg_buffer_2903 ( .C (clk), .D (new_AGEMA_signal_6333), .Q (new_AGEMA_signal_6334) ) ;
    buf_clk new_AGEMA_reg_buffer_2913 ( .C (clk), .D (new_AGEMA_signal_6343), .Q (new_AGEMA_signal_6344) ) ;
    buf_clk new_AGEMA_reg_buffer_2915 ( .C (clk), .D (new_AGEMA_signal_6345), .Q (new_AGEMA_signal_6346) ) ;
    buf_clk new_AGEMA_reg_buffer_2917 ( .C (clk), .D (new_AGEMA_signal_6347), .Q (new_AGEMA_signal_6348) ) ;
    buf_clk new_AGEMA_reg_buffer_2919 ( .C (clk), .D (new_AGEMA_signal_6349), .Q (new_AGEMA_signal_6350) ) ;
    buf_clk new_AGEMA_reg_buffer_2921 ( .C (clk), .D (new_AGEMA_signal_6351), .Q (new_AGEMA_signal_6352) ) ;
    buf_clk new_AGEMA_reg_buffer_2925 ( .C (clk), .D (new_AGEMA_signal_6355), .Q (new_AGEMA_signal_6356) ) ;
    buf_clk new_AGEMA_reg_buffer_2929 ( .C (clk), .D (new_AGEMA_signal_6359), .Q (new_AGEMA_signal_6360) ) ;
    buf_clk new_AGEMA_reg_buffer_2933 ( .C (clk), .D (new_AGEMA_signal_6363), .Q (new_AGEMA_signal_6364) ) ;
    buf_clk new_AGEMA_reg_buffer_2945 ( .C (clk), .D (new_AGEMA_signal_6375), .Q (new_AGEMA_signal_6376) ) ;
    buf_clk new_AGEMA_reg_buffer_2947 ( .C (clk), .D (new_AGEMA_signal_6377), .Q (new_AGEMA_signal_6378) ) ;
    buf_clk new_AGEMA_reg_buffer_2949 ( .C (clk), .D (new_AGEMA_signal_6379), .Q (new_AGEMA_signal_6380) ) ;
    buf_clk new_AGEMA_reg_buffer_2951 ( .C (clk), .D (new_AGEMA_signal_6381), .Q (new_AGEMA_signal_6382) ) ;
    buf_clk new_AGEMA_reg_buffer_2961 ( .C (clk), .D (new_AGEMA_signal_6391), .Q (new_AGEMA_signal_6392) ) ;
    buf_clk new_AGEMA_reg_buffer_2963 ( .C (clk), .D (new_AGEMA_signal_6393), .Q (new_AGEMA_signal_6394) ) ;
    buf_clk new_AGEMA_reg_buffer_2965 ( .C (clk), .D (new_AGEMA_signal_6395), .Q (new_AGEMA_signal_6396) ) ;
    buf_clk new_AGEMA_reg_buffer_2967 ( .C (clk), .D (new_AGEMA_signal_6397), .Q (new_AGEMA_signal_6398) ) ;
    buf_clk new_AGEMA_reg_buffer_2969 ( .C (clk), .D (new_AGEMA_signal_6399), .Q (new_AGEMA_signal_6400) ) ;
    buf_clk new_AGEMA_reg_buffer_2973 ( .C (clk), .D (new_AGEMA_signal_6403), .Q (new_AGEMA_signal_6404) ) ;
    buf_clk new_AGEMA_reg_buffer_2977 ( .C (clk), .D (new_AGEMA_signal_6407), .Q (new_AGEMA_signal_6408) ) ;
    buf_clk new_AGEMA_reg_buffer_2981 ( .C (clk), .D (new_AGEMA_signal_6411), .Q (new_AGEMA_signal_6412) ) ;
    buf_clk new_AGEMA_reg_buffer_2993 ( .C (clk), .D (new_AGEMA_signal_6423), .Q (new_AGEMA_signal_6424) ) ;
    buf_clk new_AGEMA_reg_buffer_2995 ( .C (clk), .D (new_AGEMA_signal_6425), .Q (new_AGEMA_signal_6426) ) ;
    buf_clk new_AGEMA_reg_buffer_2997 ( .C (clk), .D (new_AGEMA_signal_6427), .Q (new_AGEMA_signal_6428) ) ;
    buf_clk new_AGEMA_reg_buffer_2999 ( .C (clk), .D (new_AGEMA_signal_6429), .Q (new_AGEMA_signal_6430) ) ;
    buf_clk new_AGEMA_reg_buffer_3009 ( .C (clk), .D (new_AGEMA_signal_6439), .Q (new_AGEMA_signal_6440) ) ;
    buf_clk new_AGEMA_reg_buffer_3011 ( .C (clk), .D (new_AGEMA_signal_6441), .Q (new_AGEMA_signal_6442) ) ;
    buf_clk new_AGEMA_reg_buffer_3013 ( .C (clk), .D (new_AGEMA_signal_6443), .Q (new_AGEMA_signal_6444) ) ;
    buf_clk new_AGEMA_reg_buffer_3015 ( .C (clk), .D (new_AGEMA_signal_6445), .Q (new_AGEMA_signal_6446) ) ;
    buf_clk new_AGEMA_reg_buffer_3017 ( .C (clk), .D (new_AGEMA_signal_6447), .Q (new_AGEMA_signal_6448) ) ;
    buf_clk new_AGEMA_reg_buffer_3021 ( .C (clk), .D (new_AGEMA_signal_6451), .Q (new_AGEMA_signal_6452) ) ;
    buf_clk new_AGEMA_reg_buffer_3025 ( .C (clk), .D (new_AGEMA_signal_6455), .Q (new_AGEMA_signal_6456) ) ;
    buf_clk new_AGEMA_reg_buffer_3029 ( .C (clk), .D (new_AGEMA_signal_6459), .Q (new_AGEMA_signal_6460) ) ;
    buf_clk new_AGEMA_reg_buffer_3041 ( .C (clk), .D (new_AGEMA_signal_6471), .Q (new_AGEMA_signal_6472) ) ;
    buf_clk new_AGEMA_reg_buffer_3043 ( .C (clk), .D (new_AGEMA_signal_6473), .Q (new_AGEMA_signal_6474) ) ;
    buf_clk new_AGEMA_reg_buffer_3045 ( .C (clk), .D (new_AGEMA_signal_6475), .Q (new_AGEMA_signal_6476) ) ;
    buf_clk new_AGEMA_reg_buffer_3047 ( .C (clk), .D (new_AGEMA_signal_6477), .Q (new_AGEMA_signal_6478) ) ;
    buf_clk new_AGEMA_reg_buffer_3057 ( .C (clk), .D (new_AGEMA_signal_6487), .Q (new_AGEMA_signal_6488) ) ;
    buf_clk new_AGEMA_reg_buffer_3059 ( .C (clk), .D (new_AGEMA_signal_6489), .Q (new_AGEMA_signal_6490) ) ;
    buf_clk new_AGEMA_reg_buffer_3061 ( .C (clk), .D (new_AGEMA_signal_6491), .Q (new_AGEMA_signal_6492) ) ;
    buf_clk new_AGEMA_reg_buffer_3063 ( .C (clk), .D (new_AGEMA_signal_6493), .Q (new_AGEMA_signal_6494) ) ;
    buf_clk new_AGEMA_reg_buffer_3065 ( .C (clk), .D (new_AGEMA_signal_6495), .Q (new_AGEMA_signal_6496) ) ;
    buf_clk new_AGEMA_reg_buffer_3069 ( .C (clk), .D (new_AGEMA_signal_6499), .Q (new_AGEMA_signal_6500) ) ;
    buf_clk new_AGEMA_reg_buffer_3073 ( .C (clk), .D (new_AGEMA_signal_6503), .Q (new_AGEMA_signal_6504) ) ;
    buf_clk new_AGEMA_reg_buffer_3077 ( .C (clk), .D (new_AGEMA_signal_6507), .Q (new_AGEMA_signal_6508) ) ;
    buf_clk new_AGEMA_reg_buffer_3089 ( .C (clk), .D (new_AGEMA_signal_6519), .Q (new_AGEMA_signal_6520) ) ;
    buf_clk new_AGEMA_reg_buffer_3091 ( .C (clk), .D (new_AGEMA_signal_6521), .Q (new_AGEMA_signal_6522) ) ;
    buf_clk new_AGEMA_reg_buffer_3093 ( .C (clk), .D (new_AGEMA_signal_6523), .Q (new_AGEMA_signal_6524) ) ;
    buf_clk new_AGEMA_reg_buffer_3095 ( .C (clk), .D (new_AGEMA_signal_6525), .Q (new_AGEMA_signal_6526) ) ;
    buf_clk new_AGEMA_reg_buffer_3105 ( .C (clk), .D (new_AGEMA_signal_6535), .Q (new_AGEMA_signal_6536) ) ;
    buf_clk new_AGEMA_reg_buffer_3107 ( .C (clk), .D (new_AGEMA_signal_6537), .Q (new_AGEMA_signal_6538) ) ;
    buf_clk new_AGEMA_reg_buffer_3109 ( .C (clk), .D (new_AGEMA_signal_6539), .Q (new_AGEMA_signal_6540) ) ;
    buf_clk new_AGEMA_reg_buffer_3111 ( .C (clk), .D (new_AGEMA_signal_6541), .Q (new_AGEMA_signal_6542) ) ;
    buf_clk new_AGEMA_reg_buffer_3113 ( .C (clk), .D (new_AGEMA_signal_6543), .Q (new_AGEMA_signal_6544) ) ;
    buf_clk new_AGEMA_reg_buffer_3117 ( .C (clk), .D (new_AGEMA_signal_6547), .Q (new_AGEMA_signal_6548) ) ;
    buf_clk new_AGEMA_reg_buffer_3121 ( .C (clk), .D (new_AGEMA_signal_6551), .Q (new_AGEMA_signal_6552) ) ;
    buf_clk new_AGEMA_reg_buffer_3125 ( .C (clk), .D (new_AGEMA_signal_6555), .Q (new_AGEMA_signal_6556) ) ;
    buf_clk new_AGEMA_reg_buffer_3137 ( .C (clk), .D (new_AGEMA_signal_6567), .Q (new_AGEMA_signal_6568) ) ;
    buf_clk new_AGEMA_reg_buffer_3139 ( .C (clk), .D (new_AGEMA_signal_6569), .Q (new_AGEMA_signal_6570) ) ;
    buf_clk new_AGEMA_reg_buffer_3141 ( .C (clk), .D (new_AGEMA_signal_6571), .Q (new_AGEMA_signal_6572) ) ;
    buf_clk new_AGEMA_reg_buffer_3143 ( .C (clk), .D (new_AGEMA_signal_6573), .Q (new_AGEMA_signal_6574) ) ;
    buf_clk new_AGEMA_reg_buffer_3153 ( .C (clk), .D (new_AGEMA_signal_6583), .Q (new_AGEMA_signal_6584) ) ;
    buf_clk new_AGEMA_reg_buffer_3155 ( .C (clk), .D (new_AGEMA_signal_6585), .Q (new_AGEMA_signal_6586) ) ;
    buf_clk new_AGEMA_reg_buffer_3157 ( .C (clk), .D (new_AGEMA_signal_6587), .Q (new_AGEMA_signal_6588) ) ;
    buf_clk new_AGEMA_reg_buffer_3159 ( .C (clk), .D (new_AGEMA_signal_6589), .Q (new_AGEMA_signal_6590) ) ;
    buf_clk new_AGEMA_reg_buffer_3161 ( .C (clk), .D (new_AGEMA_signal_6591), .Q (new_AGEMA_signal_6592) ) ;
    buf_clk new_AGEMA_reg_buffer_3165 ( .C (clk), .D (new_AGEMA_signal_6595), .Q (new_AGEMA_signal_6596) ) ;
    buf_clk new_AGEMA_reg_buffer_3169 ( .C (clk), .D (new_AGEMA_signal_6599), .Q (new_AGEMA_signal_6600) ) ;
    buf_clk new_AGEMA_reg_buffer_3173 ( .C (clk), .D (new_AGEMA_signal_6603), .Q (new_AGEMA_signal_6604) ) ;
    buf_clk new_AGEMA_reg_buffer_3185 ( .C (clk), .D (new_AGEMA_signal_6615), .Q (new_AGEMA_signal_6616) ) ;
    buf_clk new_AGEMA_reg_buffer_3189 ( .C (clk), .D (new_AGEMA_signal_6619), .Q (new_AGEMA_signal_6620) ) ;
    buf_clk new_AGEMA_reg_buffer_3193 ( .C (clk), .D (new_AGEMA_signal_6623), .Q (new_AGEMA_signal_6624) ) ;
    buf_clk new_AGEMA_reg_buffer_3197 ( .C (clk), .D (new_AGEMA_signal_6627), .Q (new_AGEMA_signal_6628) ) ;
    buf_clk new_AGEMA_reg_buffer_3201 ( .C (clk), .D (new_AGEMA_signal_6631), .Q (new_AGEMA_signal_6632) ) ;
    buf_clk new_AGEMA_reg_buffer_3205 ( .C (clk), .D (new_AGEMA_signal_6635), .Q (new_AGEMA_signal_6636) ) ;
    buf_clk new_AGEMA_reg_buffer_3209 ( .C (clk), .D (new_AGEMA_signal_6639), .Q (new_AGEMA_signal_6640) ) ;
    buf_clk new_AGEMA_reg_buffer_3213 ( .C (clk), .D (new_AGEMA_signal_6643), .Q (new_AGEMA_signal_6644) ) ;
    buf_clk new_AGEMA_reg_buffer_3217 ( .C (clk), .D (new_AGEMA_signal_6647), .Q (new_AGEMA_signal_6648) ) ;
    buf_clk new_AGEMA_reg_buffer_3221 ( .C (clk), .D (new_AGEMA_signal_6651), .Q (new_AGEMA_signal_6652) ) ;
    buf_clk new_AGEMA_reg_buffer_3225 ( .C (clk), .D (new_AGEMA_signal_6655), .Q (new_AGEMA_signal_6656) ) ;
    buf_clk new_AGEMA_reg_buffer_3229 ( .C (clk), .D (new_AGEMA_signal_6659), .Q (new_AGEMA_signal_6660) ) ;
    buf_clk new_AGEMA_reg_buffer_3233 ( .C (clk), .D (new_AGEMA_signal_6663), .Q (new_AGEMA_signal_6664) ) ;
    buf_clk new_AGEMA_reg_buffer_3237 ( .C (clk), .D (new_AGEMA_signal_6667), .Q (new_AGEMA_signal_6668) ) ;
    buf_clk new_AGEMA_reg_buffer_3241 ( .C (clk), .D (new_AGEMA_signal_6671), .Q (new_AGEMA_signal_6672) ) ;
    buf_clk new_AGEMA_reg_buffer_3245 ( .C (clk), .D (new_AGEMA_signal_6675), .Q (new_AGEMA_signal_6676) ) ;
    buf_clk new_AGEMA_reg_buffer_3249 ( .C (clk), .D (new_AGEMA_signal_6679), .Q (new_AGEMA_signal_6680) ) ;
    buf_clk new_AGEMA_reg_buffer_3253 ( .C (clk), .D (new_AGEMA_signal_6683), .Q (new_AGEMA_signal_6684) ) ;
    buf_clk new_AGEMA_reg_buffer_3257 ( .C (clk), .D (new_AGEMA_signal_6687), .Q (new_AGEMA_signal_6688) ) ;
    buf_clk new_AGEMA_reg_buffer_3261 ( .C (clk), .D (new_AGEMA_signal_6691), .Q (new_AGEMA_signal_6692) ) ;
    buf_clk new_AGEMA_reg_buffer_3265 ( .C (clk), .D (new_AGEMA_signal_6695), .Q (new_AGEMA_signal_6696) ) ;
    buf_clk new_AGEMA_reg_buffer_3269 ( .C (clk), .D (new_AGEMA_signal_6699), .Q (new_AGEMA_signal_6700) ) ;
    buf_clk new_AGEMA_reg_buffer_3273 ( .C (clk), .D (new_AGEMA_signal_6703), .Q (new_AGEMA_signal_6704) ) ;
    buf_clk new_AGEMA_reg_buffer_3277 ( .C (clk), .D (new_AGEMA_signal_6707), .Q (new_AGEMA_signal_6708) ) ;
    buf_clk new_AGEMA_reg_buffer_3281 ( .C (clk), .D (new_AGEMA_signal_6711), .Q (new_AGEMA_signal_6712) ) ;
    buf_clk new_AGEMA_reg_buffer_3285 ( .C (clk), .D (new_AGEMA_signal_6715), .Q (new_AGEMA_signal_6716) ) ;
    buf_clk new_AGEMA_reg_buffer_3289 ( .C (clk), .D (new_AGEMA_signal_6719), .Q (new_AGEMA_signal_6720) ) ;
    buf_clk new_AGEMA_reg_buffer_3293 ( .C (clk), .D (new_AGEMA_signal_6723), .Q (new_AGEMA_signal_6724) ) ;
    buf_clk new_AGEMA_reg_buffer_3297 ( .C (clk), .D (new_AGEMA_signal_6727), .Q (new_AGEMA_signal_6728) ) ;
    buf_clk new_AGEMA_reg_buffer_3301 ( .C (clk), .D (new_AGEMA_signal_6731), .Q (new_AGEMA_signal_6732) ) ;
    buf_clk new_AGEMA_reg_buffer_3305 ( .C (clk), .D (new_AGEMA_signal_6735), .Q (new_AGEMA_signal_6736) ) ;
    buf_clk new_AGEMA_reg_buffer_3309 ( .C (clk), .D (new_AGEMA_signal_6739), .Q (new_AGEMA_signal_6740) ) ;
    buf_clk new_AGEMA_reg_buffer_3313 ( .C (clk), .D (new_AGEMA_signal_6743), .Q (new_AGEMA_signal_6744) ) ;
    buf_clk new_AGEMA_reg_buffer_3317 ( .C (clk), .D (new_AGEMA_signal_6747), .Q (new_AGEMA_signal_6748) ) ;
    buf_clk new_AGEMA_reg_buffer_3321 ( .C (clk), .D (new_AGEMA_signal_6751), .Q (new_AGEMA_signal_6752) ) ;
    buf_clk new_AGEMA_reg_buffer_3325 ( .C (clk), .D (new_AGEMA_signal_6755), .Q (new_AGEMA_signal_6756) ) ;
    buf_clk new_AGEMA_reg_buffer_3329 ( .C (clk), .D (new_AGEMA_signal_6759), .Q (new_AGEMA_signal_6760) ) ;
    buf_clk new_AGEMA_reg_buffer_3333 ( .C (clk), .D (new_AGEMA_signal_6763), .Q (new_AGEMA_signal_6764) ) ;
    buf_clk new_AGEMA_reg_buffer_3337 ( .C (clk), .D (new_AGEMA_signal_6767), .Q (new_AGEMA_signal_6768) ) ;
    buf_clk new_AGEMA_reg_buffer_3341 ( .C (clk), .D (new_AGEMA_signal_6771), .Q (new_AGEMA_signal_6772) ) ;
    buf_clk new_AGEMA_reg_buffer_3345 ( .C (clk), .D (new_AGEMA_signal_6775), .Q (new_AGEMA_signal_6776) ) ;
    buf_clk new_AGEMA_reg_buffer_3349 ( .C (clk), .D (new_AGEMA_signal_6779), .Q (new_AGEMA_signal_6780) ) ;
    buf_clk new_AGEMA_reg_buffer_3353 ( .C (clk), .D (new_AGEMA_signal_6783), .Q (new_AGEMA_signal_6784) ) ;
    buf_clk new_AGEMA_reg_buffer_3357 ( .C (clk), .D (new_AGEMA_signal_6787), .Q (new_AGEMA_signal_6788) ) ;
    buf_clk new_AGEMA_reg_buffer_3361 ( .C (clk), .D (new_AGEMA_signal_6791), .Q (new_AGEMA_signal_6792) ) ;
    buf_clk new_AGEMA_reg_buffer_3365 ( .C (clk), .D (new_AGEMA_signal_6795), .Q (new_AGEMA_signal_6796) ) ;
    buf_clk new_AGEMA_reg_buffer_3369 ( .C (clk), .D (new_AGEMA_signal_6799), .Q (new_AGEMA_signal_6800) ) ;
    buf_clk new_AGEMA_reg_buffer_3373 ( .C (clk), .D (new_AGEMA_signal_6803), .Q (new_AGEMA_signal_6804) ) ;
    buf_clk new_AGEMA_reg_buffer_3377 ( .C (clk), .D (new_AGEMA_signal_6807), .Q (new_AGEMA_signal_6808) ) ;
    buf_clk new_AGEMA_reg_buffer_3381 ( .C (clk), .D (new_AGEMA_signal_6811), .Q (new_AGEMA_signal_6812) ) ;
    buf_clk new_AGEMA_reg_buffer_3385 ( .C (clk), .D (new_AGEMA_signal_6815), .Q (new_AGEMA_signal_6816) ) ;
    buf_clk new_AGEMA_reg_buffer_3389 ( .C (clk), .D (new_AGEMA_signal_6819), .Q (new_AGEMA_signal_6820) ) ;
    buf_clk new_AGEMA_reg_buffer_3393 ( .C (clk), .D (new_AGEMA_signal_6823), .Q (new_AGEMA_signal_6824) ) ;
    buf_clk new_AGEMA_reg_buffer_3397 ( .C (clk), .D (new_AGEMA_signal_6827), .Q (new_AGEMA_signal_6828) ) ;
    buf_clk new_AGEMA_reg_buffer_3401 ( .C (clk), .D (new_AGEMA_signal_6831), .Q (new_AGEMA_signal_6832) ) ;
    buf_clk new_AGEMA_reg_buffer_3405 ( .C (clk), .D (new_AGEMA_signal_6835), .Q (new_AGEMA_signal_6836) ) ;
    buf_clk new_AGEMA_reg_buffer_3409 ( .C (clk), .D (new_AGEMA_signal_6839), .Q (new_AGEMA_signal_6840) ) ;
    buf_clk new_AGEMA_reg_buffer_3413 ( .C (clk), .D (new_AGEMA_signal_6843), .Q (new_AGEMA_signal_6844) ) ;
    buf_clk new_AGEMA_reg_buffer_3417 ( .C (clk), .D (new_AGEMA_signal_6847), .Q (new_AGEMA_signal_6848) ) ;
    buf_clk new_AGEMA_reg_buffer_3421 ( .C (clk), .D (new_AGEMA_signal_6851), .Q (new_AGEMA_signal_6852) ) ;
    buf_clk new_AGEMA_reg_buffer_3425 ( .C (clk), .D (new_AGEMA_signal_6855), .Q (new_AGEMA_signal_6856) ) ;
    buf_clk new_AGEMA_reg_buffer_3429 ( .C (clk), .D (new_AGEMA_signal_6859), .Q (new_AGEMA_signal_6860) ) ;
    buf_clk new_AGEMA_reg_buffer_3433 ( .C (clk), .D (new_AGEMA_signal_6863), .Q (new_AGEMA_signal_6864) ) ;
    buf_clk new_AGEMA_reg_buffer_3437 ( .C (clk), .D (new_AGEMA_signal_6867), .Q (new_AGEMA_signal_6868) ) ;
    buf_clk new_AGEMA_reg_buffer_3441 ( .C (clk), .D (new_AGEMA_signal_6871), .Q (new_AGEMA_signal_6872) ) ;
    buf_clk new_AGEMA_reg_buffer_3445 ( .C (clk), .D (new_AGEMA_signal_6875), .Q (new_AGEMA_signal_6876) ) ;
    buf_clk new_AGEMA_reg_buffer_3449 ( .C (clk), .D (new_AGEMA_signal_6879), .Q (new_AGEMA_signal_6880) ) ;
    buf_clk new_AGEMA_reg_buffer_3453 ( .C (clk), .D (new_AGEMA_signal_6883), .Q (new_AGEMA_signal_6884) ) ;
    buf_clk new_AGEMA_reg_buffer_3713 ( .C (clk), .D (new_AGEMA_signal_7143), .Q (new_AGEMA_signal_7144) ) ;
    buf_clk new_AGEMA_reg_buffer_3717 ( .C (clk), .D (new_AGEMA_signal_7147), .Q (new_AGEMA_signal_7148) ) ;
    buf_clk new_AGEMA_reg_buffer_3721 ( .C (clk), .D (new_AGEMA_signal_7151), .Q (new_AGEMA_signal_7152) ) ;
    buf_clk new_AGEMA_reg_buffer_3725 ( .C (clk), .D (new_AGEMA_signal_7155), .Q (new_AGEMA_signal_7156) ) ;
    buf_clk new_AGEMA_reg_buffer_3729 ( .C (clk), .D (new_AGEMA_signal_7159), .Q (new_AGEMA_signal_7160) ) ;
    buf_clk new_AGEMA_reg_buffer_3733 ( .C (clk), .D (new_AGEMA_signal_7163), .Q (new_AGEMA_signal_7164) ) ;
    buf_clk new_AGEMA_reg_buffer_3737 ( .C (clk), .D (new_AGEMA_signal_7167), .Q (new_AGEMA_signal_7168) ) ;
    buf_clk new_AGEMA_reg_buffer_3741 ( .C (clk), .D (new_AGEMA_signal_7171), .Q (new_AGEMA_signal_7172) ) ;
    buf_clk new_AGEMA_reg_buffer_3745 ( .C (clk), .D (new_AGEMA_signal_7175), .Q (new_AGEMA_signal_7176) ) ;
    buf_clk new_AGEMA_reg_buffer_3749 ( .C (clk), .D (new_AGEMA_signal_7179), .Q (new_AGEMA_signal_7180) ) ;
    buf_clk new_AGEMA_reg_buffer_3753 ( .C (clk), .D (new_AGEMA_signal_7183), .Q (new_AGEMA_signal_7184) ) ;
    buf_clk new_AGEMA_reg_buffer_3757 ( .C (clk), .D (new_AGEMA_signal_7187), .Q (new_AGEMA_signal_7188) ) ;
    buf_clk new_AGEMA_reg_buffer_3761 ( .C (clk), .D (new_AGEMA_signal_7191), .Q (new_AGEMA_signal_7192) ) ;
    buf_clk new_AGEMA_reg_buffer_3765 ( .C (clk), .D (new_AGEMA_signal_7195), .Q (new_AGEMA_signal_7196) ) ;
    buf_clk new_AGEMA_reg_buffer_3769 ( .C (clk), .D (new_AGEMA_signal_7199), .Q (new_AGEMA_signal_7200) ) ;
    buf_clk new_AGEMA_reg_buffer_3773 ( .C (clk), .D (new_AGEMA_signal_7203), .Q (new_AGEMA_signal_7204) ) ;
    buf_clk new_AGEMA_reg_buffer_3777 ( .C (clk), .D (new_AGEMA_signal_7207), .Q (new_AGEMA_signal_7208) ) ;
    buf_clk new_AGEMA_reg_buffer_3781 ( .C (clk), .D (new_AGEMA_signal_7211), .Q (new_AGEMA_signal_7212) ) ;
    buf_clk new_AGEMA_reg_buffer_3785 ( .C (clk), .D (new_AGEMA_signal_7215), .Q (new_AGEMA_signal_7216) ) ;
    buf_clk new_AGEMA_reg_buffer_3789 ( .C (clk), .D (new_AGEMA_signal_7219), .Q (new_AGEMA_signal_7220) ) ;
    buf_clk new_AGEMA_reg_buffer_3793 ( .C (clk), .D (new_AGEMA_signal_7223), .Q (new_AGEMA_signal_7224) ) ;
    buf_clk new_AGEMA_reg_buffer_3797 ( .C (clk), .D (new_AGEMA_signal_7227), .Q (new_AGEMA_signal_7228) ) ;
    buf_clk new_AGEMA_reg_buffer_3801 ( .C (clk), .D (new_AGEMA_signal_7231), .Q (new_AGEMA_signal_7232) ) ;
    buf_clk new_AGEMA_reg_buffer_3805 ( .C (clk), .D (new_AGEMA_signal_7235), .Q (new_AGEMA_signal_7236) ) ;
    buf_clk new_AGEMA_reg_buffer_3809 ( .C (clk), .D (new_AGEMA_signal_7239), .Q (new_AGEMA_signal_7240) ) ;
    buf_clk new_AGEMA_reg_buffer_3813 ( .C (clk), .D (new_AGEMA_signal_7243), .Q (new_AGEMA_signal_7244) ) ;
    buf_clk new_AGEMA_reg_buffer_3817 ( .C (clk), .D (new_AGEMA_signal_7247), .Q (new_AGEMA_signal_7248) ) ;
    buf_clk new_AGEMA_reg_buffer_3821 ( .C (clk), .D (new_AGEMA_signal_7251), .Q (new_AGEMA_signal_7252) ) ;
    buf_clk new_AGEMA_reg_buffer_3825 ( .C (clk), .D (new_AGEMA_signal_7255), .Q (new_AGEMA_signal_7256) ) ;
    buf_clk new_AGEMA_reg_buffer_3829 ( .C (clk), .D (new_AGEMA_signal_7259), .Q (new_AGEMA_signal_7260) ) ;
    buf_clk new_AGEMA_reg_buffer_3833 ( .C (clk), .D (new_AGEMA_signal_7263), .Q (new_AGEMA_signal_7264) ) ;
    buf_clk new_AGEMA_reg_buffer_3837 ( .C (clk), .D (new_AGEMA_signal_7267), .Q (new_AGEMA_signal_7268) ) ;
    buf_clk new_AGEMA_reg_buffer_3841 ( .C (clk), .D (new_AGEMA_signal_7271), .Q (new_AGEMA_signal_7272) ) ;
    buf_clk new_AGEMA_reg_buffer_3845 ( .C (clk), .D (new_AGEMA_signal_7275), .Q (new_AGEMA_signal_7276) ) ;
    buf_clk new_AGEMA_reg_buffer_3849 ( .C (clk), .D (new_AGEMA_signal_7279), .Q (new_AGEMA_signal_7280) ) ;
    buf_clk new_AGEMA_reg_buffer_3853 ( .C (clk), .D (new_AGEMA_signal_7283), .Q (new_AGEMA_signal_7284) ) ;
    buf_clk new_AGEMA_reg_buffer_3857 ( .C (clk), .D (new_AGEMA_signal_7287), .Q (new_AGEMA_signal_7288) ) ;
    buf_clk new_AGEMA_reg_buffer_3861 ( .C (clk), .D (new_AGEMA_signal_7291), .Q (new_AGEMA_signal_7292) ) ;
    buf_clk new_AGEMA_reg_buffer_3865 ( .C (clk), .D (new_AGEMA_signal_7295), .Q (new_AGEMA_signal_7296) ) ;
    buf_clk new_AGEMA_reg_buffer_3869 ( .C (clk), .D (new_AGEMA_signal_7299), .Q (new_AGEMA_signal_7300) ) ;
    buf_clk new_AGEMA_reg_buffer_3873 ( .C (clk), .D (new_AGEMA_signal_7303), .Q (new_AGEMA_signal_7304) ) ;
    buf_clk new_AGEMA_reg_buffer_3877 ( .C (clk), .D (new_AGEMA_signal_7307), .Q (new_AGEMA_signal_7308) ) ;
    buf_clk new_AGEMA_reg_buffer_3881 ( .C (clk), .D (new_AGEMA_signal_7311), .Q (new_AGEMA_signal_7312) ) ;
    buf_clk new_AGEMA_reg_buffer_3885 ( .C (clk), .D (new_AGEMA_signal_7315), .Q (new_AGEMA_signal_7316) ) ;
    buf_clk new_AGEMA_reg_buffer_3889 ( .C (clk), .D (new_AGEMA_signal_7319), .Q (new_AGEMA_signal_7320) ) ;
    buf_clk new_AGEMA_reg_buffer_3893 ( .C (clk), .D (new_AGEMA_signal_7323), .Q (new_AGEMA_signal_7324) ) ;
    buf_clk new_AGEMA_reg_buffer_3897 ( .C (clk), .D (new_AGEMA_signal_7327), .Q (new_AGEMA_signal_7328) ) ;
    buf_clk new_AGEMA_reg_buffer_3901 ( .C (clk), .D (new_AGEMA_signal_7331), .Q (new_AGEMA_signal_7332) ) ;
    buf_clk new_AGEMA_reg_buffer_3905 ( .C (clk), .D (new_AGEMA_signal_7335), .Q (new_AGEMA_signal_7336) ) ;
    buf_clk new_AGEMA_reg_buffer_3909 ( .C (clk), .D (new_AGEMA_signal_7339), .Q (new_AGEMA_signal_7340) ) ;
    buf_clk new_AGEMA_reg_buffer_3913 ( .C (clk), .D (new_AGEMA_signal_7343), .Q (new_AGEMA_signal_7344) ) ;
    buf_clk new_AGEMA_reg_buffer_3917 ( .C (clk), .D (new_AGEMA_signal_7347), .Q (new_AGEMA_signal_7348) ) ;
    buf_clk new_AGEMA_reg_buffer_3921 ( .C (clk), .D (new_AGEMA_signal_7351), .Q (new_AGEMA_signal_7352) ) ;
    buf_clk new_AGEMA_reg_buffer_3925 ( .C (clk), .D (new_AGEMA_signal_7355), .Q (new_AGEMA_signal_7356) ) ;
    buf_clk new_AGEMA_reg_buffer_3929 ( .C (clk), .D (new_AGEMA_signal_7359), .Q (new_AGEMA_signal_7360) ) ;
    buf_clk new_AGEMA_reg_buffer_3933 ( .C (clk), .D (new_AGEMA_signal_7363), .Q (new_AGEMA_signal_7364) ) ;
    buf_clk new_AGEMA_reg_buffer_3937 ( .C (clk), .D (new_AGEMA_signal_7367), .Q (new_AGEMA_signal_7368) ) ;
    buf_clk new_AGEMA_reg_buffer_3941 ( .C (clk), .D (new_AGEMA_signal_7371), .Q (new_AGEMA_signal_7372) ) ;
    buf_clk new_AGEMA_reg_buffer_3945 ( .C (clk), .D (new_AGEMA_signal_7375), .Q (new_AGEMA_signal_7376) ) ;
    buf_clk new_AGEMA_reg_buffer_3949 ( .C (clk), .D (new_AGEMA_signal_7379), .Q (new_AGEMA_signal_7380) ) ;
    buf_clk new_AGEMA_reg_buffer_3953 ( .C (clk), .D (new_AGEMA_signal_7383), .Q (new_AGEMA_signal_7384) ) ;
    buf_clk new_AGEMA_reg_buffer_3957 ( .C (clk), .D (new_AGEMA_signal_7387), .Q (new_AGEMA_signal_7388) ) ;
    buf_clk new_AGEMA_reg_buffer_3961 ( .C (clk), .D (new_AGEMA_signal_7391), .Q (new_AGEMA_signal_7392) ) ;
    buf_clk new_AGEMA_reg_buffer_3965 ( .C (clk), .D (new_AGEMA_signal_7395), .Q (new_AGEMA_signal_7396) ) ;
    buf_clk new_AGEMA_reg_buffer_3969 ( .C (clk), .D (new_AGEMA_signal_7399), .Q (new_AGEMA_signal_7400) ) ;
    buf_clk new_AGEMA_reg_buffer_3973 ( .C (clk), .D (new_AGEMA_signal_7403), .Q (new_AGEMA_signal_7404) ) ;
    buf_clk new_AGEMA_reg_buffer_3977 ( .C (clk), .D (new_AGEMA_signal_7407), .Q (new_AGEMA_signal_7408) ) ;
    buf_clk new_AGEMA_reg_buffer_3981 ( .C (clk), .D (new_AGEMA_signal_7411), .Q (new_AGEMA_signal_7412) ) ;
    buf_clk new_AGEMA_reg_buffer_3985 ( .C (clk), .D (new_AGEMA_signal_7415), .Q (new_AGEMA_signal_7416) ) ;
    buf_clk new_AGEMA_reg_buffer_3989 ( .C (clk), .D (new_AGEMA_signal_7419), .Q (new_AGEMA_signal_7420) ) ;
    buf_clk new_AGEMA_reg_buffer_3993 ( .C (clk), .D (new_AGEMA_signal_7423), .Q (new_AGEMA_signal_7424) ) ;
    buf_clk new_AGEMA_reg_buffer_3997 ( .C (clk), .D (new_AGEMA_signal_7427), .Q (new_AGEMA_signal_7428) ) ;
    buf_clk new_AGEMA_reg_buffer_4001 ( .C (clk), .D (new_AGEMA_signal_7431), .Q (new_AGEMA_signal_7432) ) ;
    buf_clk new_AGEMA_reg_buffer_4005 ( .C (clk), .D (new_AGEMA_signal_7435), .Q (new_AGEMA_signal_7436) ) ;
    buf_clk new_AGEMA_reg_buffer_4009 ( .C (clk), .D (new_AGEMA_signal_7439), .Q (new_AGEMA_signal_7440) ) ;
    buf_clk new_AGEMA_reg_buffer_4013 ( .C (clk), .D (new_AGEMA_signal_7443), .Q (new_AGEMA_signal_7444) ) ;
    buf_clk new_AGEMA_reg_buffer_4017 ( .C (clk), .D (new_AGEMA_signal_7447), .Q (new_AGEMA_signal_7448) ) ;
    buf_clk new_AGEMA_reg_buffer_4021 ( .C (clk), .D (new_AGEMA_signal_7451), .Q (new_AGEMA_signal_7452) ) ;
    buf_clk new_AGEMA_reg_buffer_4025 ( .C (clk), .D (new_AGEMA_signal_7455), .Q (new_AGEMA_signal_7456) ) ;
    buf_clk new_AGEMA_reg_buffer_4029 ( .C (clk), .D (new_AGEMA_signal_7459), .Q (new_AGEMA_signal_7460) ) ;
    buf_clk new_AGEMA_reg_buffer_4033 ( .C (clk), .D (new_AGEMA_signal_7463), .Q (new_AGEMA_signal_7464) ) ;
    buf_clk new_AGEMA_reg_buffer_4037 ( .C (clk), .D (new_AGEMA_signal_7467), .Q (new_AGEMA_signal_7468) ) ;
    buf_clk new_AGEMA_reg_buffer_4041 ( .C (clk), .D (new_AGEMA_signal_7471), .Q (new_AGEMA_signal_7472) ) ;
    buf_clk new_AGEMA_reg_buffer_4045 ( .C (clk), .D (new_AGEMA_signal_7475), .Q (new_AGEMA_signal_7476) ) ;
    buf_clk new_AGEMA_reg_buffer_4049 ( .C (clk), .D (new_AGEMA_signal_7479), .Q (new_AGEMA_signal_7480) ) ;
    buf_clk new_AGEMA_reg_buffer_4053 ( .C (clk), .D (new_AGEMA_signal_7483), .Q (new_AGEMA_signal_7484) ) ;
    buf_clk new_AGEMA_reg_buffer_4057 ( .C (clk), .D (new_AGEMA_signal_7487), .Q (new_AGEMA_signal_7488) ) ;
    buf_clk new_AGEMA_reg_buffer_4061 ( .C (clk), .D (new_AGEMA_signal_7491), .Q (new_AGEMA_signal_7492) ) ;
    buf_clk new_AGEMA_reg_buffer_4065 ( .C (clk), .D (new_AGEMA_signal_7495), .Q (new_AGEMA_signal_7496) ) ;
    buf_clk new_AGEMA_reg_buffer_4069 ( .C (clk), .D (new_AGEMA_signal_7499), .Q (new_AGEMA_signal_7500) ) ;
    buf_clk new_AGEMA_reg_buffer_4073 ( .C (clk), .D (new_AGEMA_signal_7503), .Q (new_AGEMA_signal_7504) ) ;
    buf_clk new_AGEMA_reg_buffer_4077 ( .C (clk), .D (new_AGEMA_signal_7507), .Q (new_AGEMA_signal_7508) ) ;
    buf_clk new_AGEMA_reg_buffer_4081 ( .C (clk), .D (new_AGEMA_signal_7511), .Q (new_AGEMA_signal_7512) ) ;
    buf_clk new_AGEMA_reg_buffer_4085 ( .C (clk), .D (new_AGEMA_signal_7515), .Q (new_AGEMA_signal_7516) ) ;
    buf_clk new_AGEMA_reg_buffer_4089 ( .C (clk), .D (new_AGEMA_signal_7519), .Q (new_AGEMA_signal_7520) ) ;
    buf_clk new_AGEMA_reg_buffer_4093 ( .C (clk), .D (new_AGEMA_signal_7523), .Q (new_AGEMA_signal_7524) ) ;
    buf_clk new_AGEMA_reg_buffer_4097 ( .C (clk), .D (new_AGEMA_signal_7527), .Q (new_AGEMA_signal_7528) ) ;
    buf_clk new_AGEMA_reg_buffer_4101 ( .C (clk), .D (new_AGEMA_signal_7531), .Q (new_AGEMA_signal_7532) ) ;
    buf_clk new_AGEMA_reg_buffer_4105 ( .C (clk), .D (new_AGEMA_signal_7535), .Q (new_AGEMA_signal_7536) ) ;
    buf_clk new_AGEMA_reg_buffer_4109 ( .C (clk), .D (new_AGEMA_signal_7539), .Q (new_AGEMA_signal_7540) ) ;
    buf_clk new_AGEMA_reg_buffer_4113 ( .C (clk), .D (new_AGEMA_signal_7543), .Q (new_AGEMA_signal_7544) ) ;
    buf_clk new_AGEMA_reg_buffer_4117 ( .C (clk), .D (new_AGEMA_signal_7547), .Q (new_AGEMA_signal_7548) ) ;
    buf_clk new_AGEMA_reg_buffer_4121 ( .C (clk), .D (new_AGEMA_signal_7551), .Q (new_AGEMA_signal_7552) ) ;
    buf_clk new_AGEMA_reg_buffer_4125 ( .C (clk), .D (new_AGEMA_signal_7555), .Q (new_AGEMA_signal_7556) ) ;
    buf_clk new_AGEMA_reg_buffer_4129 ( .C (clk), .D (new_AGEMA_signal_7559), .Q (new_AGEMA_signal_7560) ) ;
    buf_clk new_AGEMA_reg_buffer_4133 ( .C (clk), .D (new_AGEMA_signal_7563), .Q (new_AGEMA_signal_7564) ) ;
    buf_clk new_AGEMA_reg_buffer_4137 ( .C (clk), .D (new_AGEMA_signal_7567), .Q (new_AGEMA_signal_7568) ) ;
    buf_clk new_AGEMA_reg_buffer_4141 ( .C (clk), .D (new_AGEMA_signal_7571), .Q (new_AGEMA_signal_7572) ) ;
    buf_clk new_AGEMA_reg_buffer_4145 ( .C (clk), .D (new_AGEMA_signal_7575), .Q (new_AGEMA_signal_7576) ) ;
    buf_clk new_AGEMA_reg_buffer_4149 ( .C (clk), .D (new_AGEMA_signal_7579), .Q (new_AGEMA_signal_7580) ) ;
    buf_clk new_AGEMA_reg_buffer_4153 ( .C (clk), .D (new_AGEMA_signal_7583), .Q (new_AGEMA_signal_7584) ) ;
    buf_clk new_AGEMA_reg_buffer_4157 ( .C (clk), .D (new_AGEMA_signal_7587), .Q (new_AGEMA_signal_7588) ) ;
    buf_clk new_AGEMA_reg_buffer_4161 ( .C (clk), .D (new_AGEMA_signal_7591), .Q (new_AGEMA_signal_7592) ) ;
    buf_clk new_AGEMA_reg_buffer_4165 ( .C (clk), .D (new_AGEMA_signal_7595), .Q (new_AGEMA_signal_7596) ) ;
    buf_clk new_AGEMA_reg_buffer_4169 ( .C (clk), .D (new_AGEMA_signal_7599), .Q (new_AGEMA_signal_7600) ) ;
    buf_clk new_AGEMA_reg_buffer_4173 ( .C (clk), .D (new_AGEMA_signal_7603), .Q (new_AGEMA_signal_7604) ) ;
    buf_clk new_AGEMA_reg_buffer_4177 ( .C (clk), .D (new_AGEMA_signal_7607), .Q (new_AGEMA_signal_7608) ) ;
    buf_clk new_AGEMA_reg_buffer_4181 ( .C (clk), .D (new_AGEMA_signal_7611), .Q (new_AGEMA_signal_7612) ) ;
    buf_clk new_AGEMA_reg_buffer_4185 ( .C (clk), .D (new_AGEMA_signal_7615), .Q (new_AGEMA_signal_7616) ) ;
    buf_clk new_AGEMA_reg_buffer_4189 ( .C (clk), .D (new_AGEMA_signal_7619), .Q (new_AGEMA_signal_7620) ) ;
    buf_clk new_AGEMA_reg_buffer_4193 ( .C (clk), .D (new_AGEMA_signal_7623), .Q (new_AGEMA_signal_7624) ) ;
    buf_clk new_AGEMA_reg_buffer_4197 ( .C (clk), .D (new_AGEMA_signal_7627), .Q (new_AGEMA_signal_7628) ) ;
    buf_clk new_AGEMA_reg_buffer_4201 ( .C (clk), .D (new_AGEMA_signal_7631), .Q (new_AGEMA_signal_7632) ) ;
    buf_clk new_AGEMA_reg_buffer_4205 ( .C (clk), .D (new_AGEMA_signal_7635), .Q (new_AGEMA_signal_7636) ) ;
    buf_clk new_AGEMA_reg_buffer_4209 ( .C (clk), .D (new_AGEMA_signal_7639), .Q (new_AGEMA_signal_7640) ) ;
    buf_clk new_AGEMA_reg_buffer_4213 ( .C (clk), .D (new_AGEMA_signal_7643), .Q (new_AGEMA_signal_7644) ) ;
    buf_clk new_AGEMA_reg_buffer_4217 ( .C (clk), .D (new_AGEMA_signal_7647), .Q (new_AGEMA_signal_7648) ) ;
    buf_clk new_AGEMA_reg_buffer_4221 ( .C (clk), .D (new_AGEMA_signal_7651), .Q (new_AGEMA_signal_7652) ) ;
    buf_clk new_AGEMA_reg_buffer_4225 ( .C (clk), .D (new_AGEMA_signal_7655), .Q (new_AGEMA_signal_7656) ) ;
    buf_clk new_AGEMA_reg_buffer_4229 ( .C (clk), .D (new_AGEMA_signal_7659), .Q (new_AGEMA_signal_7660) ) ;
    buf_clk new_AGEMA_reg_buffer_4233 ( .C (clk), .D (new_AGEMA_signal_7663), .Q (new_AGEMA_signal_7664) ) ;
    buf_clk new_AGEMA_reg_buffer_4237 ( .C (clk), .D (new_AGEMA_signal_7667), .Q (new_AGEMA_signal_7668) ) ;
    buf_clk new_AGEMA_reg_buffer_4241 ( .C (clk), .D (new_AGEMA_signal_7671), .Q (new_AGEMA_signal_7672) ) ;
    buf_clk new_AGEMA_reg_buffer_4245 ( .C (clk), .D (new_AGEMA_signal_7675), .Q (new_AGEMA_signal_7676) ) ;
    buf_clk new_AGEMA_reg_buffer_4249 ( .C (clk), .D (new_AGEMA_signal_7679), .Q (new_AGEMA_signal_7680) ) ;
    buf_clk new_AGEMA_reg_buffer_4253 ( .C (clk), .D (new_AGEMA_signal_7683), .Q (new_AGEMA_signal_7684) ) ;
    buf_clk new_AGEMA_reg_buffer_4257 ( .C (clk), .D (new_AGEMA_signal_7687), .Q (new_AGEMA_signal_7688) ) ;
    buf_clk new_AGEMA_reg_buffer_4261 ( .C (clk), .D (new_AGEMA_signal_7691), .Q (new_AGEMA_signal_7692) ) ;
    buf_clk new_AGEMA_reg_buffer_4265 ( .C (clk), .D (new_AGEMA_signal_7695), .Q (new_AGEMA_signal_7696) ) ;
    buf_clk new_AGEMA_reg_buffer_4269 ( .C (clk), .D (new_AGEMA_signal_7699), .Q (new_AGEMA_signal_7700) ) ;
    buf_clk new_AGEMA_reg_buffer_4273 ( .C (clk), .D (new_AGEMA_signal_7703), .Q (new_AGEMA_signal_7704) ) ;
    buf_clk new_AGEMA_reg_buffer_4277 ( .C (clk), .D (new_AGEMA_signal_7707), .Q (new_AGEMA_signal_7708) ) ;
    buf_clk new_AGEMA_reg_buffer_4281 ( .C (clk), .D (new_AGEMA_signal_7711), .Q (new_AGEMA_signal_7712) ) ;
    buf_clk new_AGEMA_reg_buffer_4285 ( .C (clk), .D (new_AGEMA_signal_7715), .Q (new_AGEMA_signal_7716) ) ;
    buf_clk new_AGEMA_reg_buffer_4289 ( .C (clk), .D (new_AGEMA_signal_7719), .Q (new_AGEMA_signal_7720) ) ;
    buf_clk new_AGEMA_reg_buffer_4293 ( .C (clk), .D (new_AGEMA_signal_7723), .Q (new_AGEMA_signal_7724) ) ;
    buf_clk new_AGEMA_reg_buffer_4297 ( .C (clk), .D (new_AGEMA_signal_7727), .Q (new_AGEMA_signal_7728) ) ;
    buf_clk new_AGEMA_reg_buffer_4301 ( .C (clk), .D (new_AGEMA_signal_7731), .Q (new_AGEMA_signal_7732) ) ;
    buf_clk new_AGEMA_reg_buffer_4305 ( .C (clk), .D (new_AGEMA_signal_7735), .Q (new_AGEMA_signal_7736) ) ;
    buf_clk new_AGEMA_reg_buffer_4309 ( .C (clk), .D (new_AGEMA_signal_7739), .Q (new_AGEMA_signal_7740) ) ;
    buf_clk new_AGEMA_reg_buffer_4313 ( .C (clk), .D (new_AGEMA_signal_7743), .Q (new_AGEMA_signal_7744) ) ;
    buf_clk new_AGEMA_reg_buffer_4317 ( .C (clk), .D (new_AGEMA_signal_7747), .Q (new_AGEMA_signal_7748) ) ;
    buf_clk new_AGEMA_reg_buffer_4321 ( .C (clk), .D (new_AGEMA_signal_7751), .Q (new_AGEMA_signal_7752) ) ;
    buf_clk new_AGEMA_reg_buffer_4325 ( .C (clk), .D (new_AGEMA_signal_7755), .Q (new_AGEMA_signal_7756) ) ;
    buf_clk new_AGEMA_reg_buffer_4329 ( .C (clk), .D (new_AGEMA_signal_7759), .Q (new_AGEMA_signal_7760) ) ;
    buf_clk new_AGEMA_reg_buffer_4333 ( .C (clk), .D (new_AGEMA_signal_7763), .Q (new_AGEMA_signal_7764) ) ;
    buf_clk new_AGEMA_reg_buffer_4337 ( .C (clk), .D (new_AGEMA_signal_7767), .Q (new_AGEMA_signal_7768) ) ;
    buf_clk new_AGEMA_reg_buffer_4341 ( .C (clk), .D (new_AGEMA_signal_7771), .Q (new_AGEMA_signal_7772) ) ;
    buf_clk new_AGEMA_reg_buffer_4345 ( .C (clk), .D (new_AGEMA_signal_7775), .Q (new_AGEMA_signal_7776) ) ;
    buf_clk new_AGEMA_reg_buffer_4349 ( .C (clk), .D (new_AGEMA_signal_7779), .Q (new_AGEMA_signal_7780) ) ;
    buf_clk new_AGEMA_reg_buffer_4353 ( .C (clk), .D (new_AGEMA_signal_7783), .Q (new_AGEMA_signal_7784) ) ;
    buf_clk new_AGEMA_reg_buffer_4357 ( .C (clk), .D (new_AGEMA_signal_7787), .Q (new_AGEMA_signal_7788) ) ;
    buf_clk new_AGEMA_reg_buffer_4361 ( .C (clk), .D (new_AGEMA_signal_7791), .Q (new_AGEMA_signal_7792) ) ;
    buf_clk new_AGEMA_reg_buffer_4365 ( .C (clk), .D (new_AGEMA_signal_7795), .Q (new_AGEMA_signal_7796) ) ;
    buf_clk new_AGEMA_reg_buffer_4369 ( .C (clk), .D (new_AGEMA_signal_7799), .Q (new_AGEMA_signal_7800) ) ;
    buf_clk new_AGEMA_reg_buffer_4373 ( .C (clk), .D (new_AGEMA_signal_7803), .Q (new_AGEMA_signal_7804) ) ;
    buf_clk new_AGEMA_reg_buffer_4377 ( .C (clk), .D (new_AGEMA_signal_7807), .Q (new_AGEMA_signal_7808) ) ;
    buf_clk new_AGEMA_reg_buffer_4381 ( .C (clk), .D (new_AGEMA_signal_7811), .Q (new_AGEMA_signal_7812) ) ;
    buf_clk new_AGEMA_reg_buffer_4385 ( .C (clk), .D (new_AGEMA_signal_7815), .Q (new_AGEMA_signal_7816) ) ;
    buf_clk new_AGEMA_reg_buffer_4389 ( .C (clk), .D (new_AGEMA_signal_7819), .Q (new_AGEMA_signal_7820) ) ;
    buf_clk new_AGEMA_reg_buffer_4393 ( .C (clk), .D (new_AGEMA_signal_7823), .Q (new_AGEMA_signal_7824) ) ;
    buf_clk new_AGEMA_reg_buffer_4397 ( .C (clk), .D (new_AGEMA_signal_7827), .Q (new_AGEMA_signal_7828) ) ;
    buf_clk new_AGEMA_reg_buffer_4401 ( .C (clk), .D (new_AGEMA_signal_7831), .Q (new_AGEMA_signal_7832) ) ;
    buf_clk new_AGEMA_reg_buffer_4405 ( .C (clk), .D (new_AGEMA_signal_7835), .Q (new_AGEMA_signal_7836) ) ;
    buf_clk new_AGEMA_reg_buffer_4409 ( .C (clk), .D (new_AGEMA_signal_7839), .Q (new_AGEMA_signal_7840) ) ;
    buf_clk new_AGEMA_reg_buffer_4413 ( .C (clk), .D (new_AGEMA_signal_7843), .Q (new_AGEMA_signal_7844) ) ;
    buf_clk new_AGEMA_reg_buffer_4417 ( .C (clk), .D (new_AGEMA_signal_7847), .Q (new_AGEMA_signal_7848) ) ;
    buf_clk new_AGEMA_reg_buffer_4421 ( .C (clk), .D (new_AGEMA_signal_7851), .Q (new_AGEMA_signal_7852) ) ;
    buf_clk new_AGEMA_reg_buffer_4425 ( .C (clk), .D (new_AGEMA_signal_7855), .Q (new_AGEMA_signal_7856) ) ;
    buf_clk new_AGEMA_reg_buffer_4429 ( .C (clk), .D (new_AGEMA_signal_7859), .Q (new_AGEMA_signal_7860) ) ;
    buf_clk new_AGEMA_reg_buffer_4433 ( .C (clk), .D (new_AGEMA_signal_7863), .Q (new_AGEMA_signal_7864) ) ;
    buf_clk new_AGEMA_reg_buffer_4437 ( .C (clk), .D (new_AGEMA_signal_7867), .Q (new_AGEMA_signal_7868) ) ;
    buf_clk new_AGEMA_reg_buffer_4441 ( .C (clk), .D (new_AGEMA_signal_7871), .Q (new_AGEMA_signal_7872) ) ;
    buf_clk new_AGEMA_reg_buffer_4445 ( .C (clk), .D (new_AGEMA_signal_7875), .Q (new_AGEMA_signal_7876) ) ;
    buf_clk new_AGEMA_reg_buffer_4449 ( .C (clk), .D (new_AGEMA_signal_7879), .Q (new_AGEMA_signal_7880) ) ;
    buf_clk new_AGEMA_reg_buffer_4453 ( .C (clk), .D (new_AGEMA_signal_7883), .Q (new_AGEMA_signal_7884) ) ;
    buf_clk new_AGEMA_reg_buffer_4457 ( .C (clk), .D (new_AGEMA_signal_7887), .Q (new_AGEMA_signal_7888) ) ;
    buf_clk new_AGEMA_reg_buffer_4461 ( .C (clk), .D (new_AGEMA_signal_7891), .Q (new_AGEMA_signal_7892) ) ;
    buf_clk new_AGEMA_reg_buffer_4465 ( .C (clk), .D (new_AGEMA_signal_7895), .Q (new_AGEMA_signal_7896) ) ;
    buf_clk new_AGEMA_reg_buffer_4469 ( .C (clk), .D (new_AGEMA_signal_7899), .Q (new_AGEMA_signal_7900) ) ;
    buf_clk new_AGEMA_reg_buffer_4473 ( .C (clk), .D (new_AGEMA_signal_7903), .Q (new_AGEMA_signal_7904) ) ;
    buf_clk new_AGEMA_reg_buffer_4477 ( .C (clk), .D (new_AGEMA_signal_7907), .Q (new_AGEMA_signal_7908) ) ;
    buf_clk new_AGEMA_reg_buffer_4481 ( .C (clk), .D (new_AGEMA_signal_7911), .Q (new_AGEMA_signal_7912) ) ;
    buf_clk new_AGEMA_reg_buffer_4485 ( .C (clk), .D (new_AGEMA_signal_7915), .Q (new_AGEMA_signal_7916) ) ;
    buf_clk new_AGEMA_reg_buffer_4489 ( .C (clk), .D (new_AGEMA_signal_7919), .Q (new_AGEMA_signal_7920) ) ;
    buf_clk new_AGEMA_reg_buffer_4493 ( .C (clk), .D (new_AGEMA_signal_7923), .Q (new_AGEMA_signal_7924) ) ;
    buf_clk new_AGEMA_reg_buffer_4497 ( .C (clk), .D (new_AGEMA_signal_7927), .Q (new_AGEMA_signal_7928) ) ;
    buf_clk new_AGEMA_reg_buffer_4501 ( .C (clk), .D (new_AGEMA_signal_7931), .Q (new_AGEMA_signal_7932) ) ;
    buf_clk new_AGEMA_reg_buffer_4505 ( .C (clk), .D (new_AGEMA_signal_7935), .Q (new_AGEMA_signal_7936) ) ;
    buf_clk new_AGEMA_reg_buffer_4509 ( .C (clk), .D (new_AGEMA_signal_7939), .Q (new_AGEMA_signal_7940) ) ;
    buf_clk new_AGEMA_reg_buffer_4513 ( .C (clk), .D (new_AGEMA_signal_7943), .Q (new_AGEMA_signal_7944) ) ;
    buf_clk new_AGEMA_reg_buffer_4517 ( .C (clk), .D (new_AGEMA_signal_7947), .Q (new_AGEMA_signal_7948) ) ;
    buf_clk new_AGEMA_reg_buffer_4521 ( .C (clk), .D (new_AGEMA_signal_7951), .Q (new_AGEMA_signal_7952) ) ;
    buf_clk new_AGEMA_reg_buffer_4525 ( .C (clk), .D (new_AGEMA_signal_7955), .Q (new_AGEMA_signal_7956) ) ;
    buf_clk new_AGEMA_reg_buffer_4529 ( .C (clk), .D (new_AGEMA_signal_7959), .Q (new_AGEMA_signal_7960) ) ;
    buf_clk new_AGEMA_reg_buffer_4533 ( .C (clk), .D (new_AGEMA_signal_7963), .Q (new_AGEMA_signal_7964) ) ;
    buf_clk new_AGEMA_reg_buffer_4537 ( .C (clk), .D (new_AGEMA_signal_7967), .Q (new_AGEMA_signal_7968) ) ;
    buf_clk new_AGEMA_reg_buffer_4541 ( .C (clk), .D (new_AGEMA_signal_7971), .Q (new_AGEMA_signal_7972) ) ;
    buf_clk new_AGEMA_reg_buffer_4545 ( .C (clk), .D (new_AGEMA_signal_7975), .Q (new_AGEMA_signal_7976) ) ;
    buf_clk new_AGEMA_reg_buffer_4549 ( .C (clk), .D (new_AGEMA_signal_7979), .Q (new_AGEMA_signal_7980) ) ;
    buf_clk new_AGEMA_reg_buffer_4553 ( .C (clk), .D (new_AGEMA_signal_7983), .Q (new_AGEMA_signal_7984) ) ;
    buf_clk new_AGEMA_reg_buffer_4557 ( .C (clk), .D (new_AGEMA_signal_7987), .Q (new_AGEMA_signal_7988) ) ;
    buf_clk new_AGEMA_reg_buffer_4561 ( .C (clk), .D (new_AGEMA_signal_7991), .Q (new_AGEMA_signal_7992) ) ;
    buf_clk new_AGEMA_reg_buffer_4565 ( .C (clk), .D (new_AGEMA_signal_7995), .Q (new_AGEMA_signal_7996) ) ;
    buf_clk new_AGEMA_reg_buffer_4569 ( .C (clk), .D (new_AGEMA_signal_7999), .Q (new_AGEMA_signal_8000) ) ;
    buf_clk new_AGEMA_reg_buffer_4573 ( .C (clk), .D (new_AGEMA_signal_8003), .Q (new_AGEMA_signal_8004) ) ;
    buf_clk new_AGEMA_reg_buffer_4577 ( .C (clk), .D (new_AGEMA_signal_8007), .Q (new_AGEMA_signal_8008) ) ;
    buf_clk new_AGEMA_reg_buffer_4581 ( .C (clk), .D (new_AGEMA_signal_8011), .Q (new_AGEMA_signal_8012) ) ;
    buf_clk new_AGEMA_reg_buffer_4585 ( .C (clk), .D (new_AGEMA_signal_8015), .Q (new_AGEMA_signal_8016) ) ;
    buf_clk new_AGEMA_reg_buffer_4589 ( .C (clk), .D (new_AGEMA_signal_8019), .Q (new_AGEMA_signal_8020) ) ;
    buf_clk new_AGEMA_reg_buffer_4593 ( .C (clk), .D (new_AGEMA_signal_8023), .Q (new_AGEMA_signal_8024) ) ;
    buf_clk new_AGEMA_reg_buffer_4597 ( .C (clk), .D (new_AGEMA_signal_8027), .Q (new_AGEMA_signal_8028) ) ;
    buf_clk new_AGEMA_reg_buffer_4601 ( .C (clk), .D (new_AGEMA_signal_8031), .Q (new_AGEMA_signal_8032) ) ;
    buf_clk new_AGEMA_reg_buffer_4605 ( .C (clk), .D (new_AGEMA_signal_8035), .Q (new_AGEMA_signal_8036) ) ;
    buf_clk new_AGEMA_reg_buffer_4609 ( .C (clk), .D (new_AGEMA_signal_8039), .Q (new_AGEMA_signal_8040) ) ;
    buf_clk new_AGEMA_reg_buffer_4613 ( .C (clk), .D (new_AGEMA_signal_8043), .Q (new_AGEMA_signal_8044) ) ;
    buf_clk new_AGEMA_reg_buffer_4617 ( .C (clk), .D (new_AGEMA_signal_8047), .Q (new_AGEMA_signal_8048) ) ;
    buf_clk new_AGEMA_reg_buffer_4621 ( .C (clk), .D (new_AGEMA_signal_8051), .Q (new_AGEMA_signal_8052) ) ;
    buf_clk new_AGEMA_reg_buffer_4625 ( .C (clk), .D (new_AGEMA_signal_8055), .Q (new_AGEMA_signal_8056) ) ;
    buf_clk new_AGEMA_reg_buffer_4629 ( .C (clk), .D (new_AGEMA_signal_8059), .Q (new_AGEMA_signal_8060) ) ;
    buf_clk new_AGEMA_reg_buffer_4633 ( .C (clk), .D (new_AGEMA_signal_8063), .Q (new_AGEMA_signal_8064) ) ;
    buf_clk new_AGEMA_reg_buffer_4637 ( .C (clk), .D (new_AGEMA_signal_8067), .Q (new_AGEMA_signal_8068) ) ;
    buf_clk new_AGEMA_reg_buffer_4641 ( .C (clk), .D (new_AGEMA_signal_8071), .Q (new_AGEMA_signal_8072) ) ;
    buf_clk new_AGEMA_reg_buffer_4645 ( .C (clk), .D (new_AGEMA_signal_8075), .Q (new_AGEMA_signal_8076) ) ;
    buf_clk new_AGEMA_reg_buffer_4649 ( .C (clk), .D (new_AGEMA_signal_8079), .Q (new_AGEMA_signal_8080) ) ;
    buf_clk new_AGEMA_reg_buffer_4653 ( .C (clk), .D (new_AGEMA_signal_8083), .Q (new_AGEMA_signal_8084) ) ;
    buf_clk new_AGEMA_reg_buffer_4657 ( .C (clk), .D (new_AGEMA_signal_8087), .Q (new_AGEMA_signal_8088) ) ;
    buf_clk new_AGEMA_reg_buffer_4661 ( .C (clk), .D (new_AGEMA_signal_8091), .Q (new_AGEMA_signal_8092) ) ;
    buf_clk new_AGEMA_reg_buffer_4665 ( .C (clk), .D (new_AGEMA_signal_8095), .Q (new_AGEMA_signal_8096) ) ;
    buf_clk new_AGEMA_reg_buffer_4669 ( .C (clk), .D (new_AGEMA_signal_8099), .Q (new_AGEMA_signal_8100) ) ;
    buf_clk new_AGEMA_reg_buffer_4673 ( .C (clk), .D (new_AGEMA_signal_8103), .Q (new_AGEMA_signal_8104) ) ;
    buf_clk new_AGEMA_reg_buffer_4677 ( .C (clk), .D (new_AGEMA_signal_8107), .Q (new_AGEMA_signal_8108) ) ;
    buf_clk new_AGEMA_reg_buffer_4681 ( .C (clk), .D (new_AGEMA_signal_8111), .Q (new_AGEMA_signal_8112) ) ;
    buf_clk new_AGEMA_reg_buffer_4685 ( .C (clk), .D (new_AGEMA_signal_8115), .Q (new_AGEMA_signal_8116) ) ;
    buf_clk new_AGEMA_reg_buffer_4689 ( .C (clk), .D (new_AGEMA_signal_8119), .Q (new_AGEMA_signal_8120) ) ;
    buf_clk new_AGEMA_reg_buffer_4693 ( .C (clk), .D (new_AGEMA_signal_8123), .Q (new_AGEMA_signal_8124) ) ;
    buf_clk new_AGEMA_reg_buffer_4697 ( .C (clk), .D (new_AGEMA_signal_8127), .Q (new_AGEMA_signal_8128) ) ;
    buf_clk new_AGEMA_reg_buffer_4701 ( .C (clk), .D (new_AGEMA_signal_8131), .Q (new_AGEMA_signal_8132) ) ;
    buf_clk new_AGEMA_reg_buffer_4705 ( .C (clk), .D (new_AGEMA_signal_8135), .Q (new_AGEMA_signal_8136) ) ;
    buf_clk new_AGEMA_reg_buffer_4709 ( .C (clk), .D (new_AGEMA_signal_8139), .Q (new_AGEMA_signal_8140) ) ;
    buf_clk new_AGEMA_reg_buffer_4713 ( .C (clk), .D (new_AGEMA_signal_8143), .Q (new_AGEMA_signal_8144) ) ;
    buf_clk new_AGEMA_reg_buffer_4717 ( .C (clk), .D (new_AGEMA_signal_8147), .Q (new_AGEMA_signal_8148) ) ;
    buf_clk new_AGEMA_reg_buffer_4721 ( .C (clk), .D (new_AGEMA_signal_8151), .Q (new_AGEMA_signal_8152) ) ;
    buf_clk new_AGEMA_reg_buffer_4725 ( .C (clk), .D (new_AGEMA_signal_8155), .Q (new_AGEMA_signal_8156) ) ;
    buf_clk new_AGEMA_reg_buffer_4729 ( .C (clk), .D (new_AGEMA_signal_8159), .Q (new_AGEMA_signal_8160) ) ;
    buf_clk new_AGEMA_reg_buffer_4733 ( .C (clk), .D (new_AGEMA_signal_8163), .Q (new_AGEMA_signal_8164) ) ;
    buf_clk new_AGEMA_reg_buffer_4737 ( .C (clk), .D (new_AGEMA_signal_8167), .Q (new_AGEMA_signal_8168) ) ;
    buf_clk new_AGEMA_reg_buffer_4741 ( .C (clk), .D (new_AGEMA_signal_8171), .Q (new_AGEMA_signal_8172) ) ;
    buf_clk new_AGEMA_reg_buffer_4745 ( .C (clk), .D (new_AGEMA_signal_8175), .Q (new_AGEMA_signal_8176) ) ;
    buf_clk new_AGEMA_reg_buffer_4749 ( .C (clk), .D (new_AGEMA_signal_8179), .Q (new_AGEMA_signal_8180) ) ;
    buf_clk new_AGEMA_reg_buffer_4753 ( .C (clk), .D (new_AGEMA_signal_8183), .Q (new_AGEMA_signal_8184) ) ;
    buf_clk new_AGEMA_reg_buffer_4757 ( .C (clk), .D (new_AGEMA_signal_8187), .Q (new_AGEMA_signal_8188) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_1902 ( .C (clk), .D (new_AGEMA_signal_4432), .Q (new_AGEMA_signal_5333) ) ;
    buf_clk new_AGEMA_reg_buffer_1906 ( .C (clk), .D (new_AGEMA_signal_5336), .Q (new_AGEMA_signal_5337) ) ;
    buf_clk new_AGEMA_reg_buffer_1910 ( .C (clk), .D (new_AGEMA_signal_5340), .Q (new_AGEMA_signal_5341) ) ;
    buf_clk new_AGEMA_reg_buffer_1914 ( .C (clk), .D (new_AGEMA_signal_5344), .Q (new_AGEMA_signal_5345) ) ;
    buf_clk new_AGEMA_reg_buffer_1918 ( .C (clk), .D (new_AGEMA_signal_5348), .Q (new_AGEMA_signal_5349) ) ;
    buf_clk new_AGEMA_reg_buffer_1922 ( .C (clk), .D (new_AGEMA_signal_5352), .Q (new_AGEMA_signal_5353) ) ;
    buf_clk new_AGEMA_reg_buffer_1926 ( .C (clk), .D (new_AGEMA_signal_5356), .Q (new_AGEMA_signal_5357) ) ;
    buf_clk new_AGEMA_reg_buffer_1930 ( .C (clk), .D (new_AGEMA_signal_5360), .Q (new_AGEMA_signal_5361) ) ;
    buf_clk new_AGEMA_reg_buffer_1934 ( .C (clk), .D (new_AGEMA_signal_5364), .Q (new_AGEMA_signal_5365) ) ;
    buf_clk new_AGEMA_reg_buffer_1938 ( .C (clk), .D (new_AGEMA_signal_5368), .Q (new_AGEMA_signal_5369) ) ;
    buf_clk new_AGEMA_reg_buffer_1942 ( .C (clk), .D (new_AGEMA_signal_5372), .Q (new_AGEMA_signal_5373) ) ;
    buf_clk new_AGEMA_reg_buffer_1946 ( .C (clk), .D (new_AGEMA_signal_5376), .Q (new_AGEMA_signal_5377) ) ;
    buf_clk new_AGEMA_reg_buffer_1950 ( .C (clk), .D (new_AGEMA_signal_5380), .Q (new_AGEMA_signal_5381) ) ;
    buf_clk new_AGEMA_reg_buffer_1954 ( .C (clk), .D (new_AGEMA_signal_5384), .Q (new_AGEMA_signal_5385) ) ;
    buf_clk new_AGEMA_reg_buffer_1958 ( .C (clk), .D (new_AGEMA_signal_5388), .Q (new_AGEMA_signal_5389) ) ;
    buf_clk new_AGEMA_reg_buffer_1962 ( .C (clk), .D (new_AGEMA_signal_5392), .Q (new_AGEMA_signal_5393) ) ;
    buf_clk new_AGEMA_reg_buffer_1966 ( .C (clk), .D (new_AGEMA_signal_5396), .Q (new_AGEMA_signal_5397) ) ;
    buf_clk new_AGEMA_reg_buffer_1970 ( .C (clk), .D (new_AGEMA_signal_5400), .Q (new_AGEMA_signal_5401) ) ;
    buf_clk new_AGEMA_reg_buffer_1974 ( .C (clk), .D (new_AGEMA_signal_5404), .Q (new_AGEMA_signal_5405) ) ;
    buf_clk new_AGEMA_reg_buffer_1978 ( .C (clk), .D (new_AGEMA_signal_5408), .Q (new_AGEMA_signal_5409) ) ;
    buf_clk new_AGEMA_reg_buffer_1982 ( .C (clk), .D (new_AGEMA_signal_5412), .Q (new_AGEMA_signal_5413) ) ;
    buf_clk new_AGEMA_reg_buffer_1986 ( .C (clk), .D (new_AGEMA_signal_5416), .Q (new_AGEMA_signal_5417) ) ;
    buf_clk new_AGEMA_reg_buffer_1990 ( .C (clk), .D (new_AGEMA_signal_5420), .Q (new_AGEMA_signal_5421) ) ;
    buf_clk new_AGEMA_reg_buffer_1994 ( .C (clk), .D (new_AGEMA_signal_5424), .Q (new_AGEMA_signal_5425) ) ;
    buf_clk new_AGEMA_reg_buffer_1998 ( .C (clk), .D (new_AGEMA_signal_5428), .Q (new_AGEMA_signal_5429) ) ;
    buf_clk new_AGEMA_reg_buffer_2002 ( .C (clk), .D (new_AGEMA_signal_5432), .Q (new_AGEMA_signal_5433) ) ;
    buf_clk new_AGEMA_reg_buffer_2006 ( .C (clk), .D (new_AGEMA_signal_5436), .Q (new_AGEMA_signal_5437) ) ;
    buf_clk new_AGEMA_reg_buffer_2010 ( .C (clk), .D (new_AGEMA_signal_5440), .Q (new_AGEMA_signal_5441) ) ;
    buf_clk new_AGEMA_reg_buffer_2014 ( .C (clk), .D (new_AGEMA_signal_5444), .Q (new_AGEMA_signal_5445) ) ;
    buf_clk new_AGEMA_reg_buffer_2018 ( .C (clk), .D (new_AGEMA_signal_5448), .Q (new_AGEMA_signal_5449) ) ;
    buf_clk new_AGEMA_reg_buffer_2022 ( .C (clk), .D (new_AGEMA_signal_5452), .Q (new_AGEMA_signal_5453) ) ;
    buf_clk new_AGEMA_reg_buffer_2026 ( .C (clk), .D (new_AGEMA_signal_5456), .Q (new_AGEMA_signal_5457) ) ;
    buf_clk new_AGEMA_reg_buffer_2030 ( .C (clk), .D (new_AGEMA_signal_5460), .Q (new_AGEMA_signal_5461) ) ;
    buf_clk new_AGEMA_reg_buffer_2034 ( .C (clk), .D (new_AGEMA_signal_5464), .Q (new_AGEMA_signal_5465) ) ;
    buf_clk new_AGEMA_reg_buffer_2038 ( .C (clk), .D (new_AGEMA_signal_5468), .Q (new_AGEMA_signal_5469) ) ;
    buf_clk new_AGEMA_reg_buffer_2042 ( .C (clk), .D (new_AGEMA_signal_5472), .Q (new_AGEMA_signal_5473) ) ;
    buf_clk new_AGEMA_reg_buffer_2046 ( .C (clk), .D (new_AGEMA_signal_5476), .Q (new_AGEMA_signal_5477) ) ;
    buf_clk new_AGEMA_reg_buffer_2050 ( .C (clk), .D (new_AGEMA_signal_5480), .Q (new_AGEMA_signal_5481) ) ;
    buf_clk new_AGEMA_reg_buffer_2054 ( .C (clk), .D (new_AGEMA_signal_5484), .Q (new_AGEMA_signal_5485) ) ;
    buf_clk new_AGEMA_reg_buffer_2058 ( .C (clk), .D (new_AGEMA_signal_5488), .Q (new_AGEMA_signal_5489) ) ;
    buf_clk new_AGEMA_reg_buffer_2062 ( .C (clk), .D (new_AGEMA_signal_5492), .Q (new_AGEMA_signal_5493) ) ;
    buf_clk new_AGEMA_reg_buffer_2066 ( .C (clk), .D (new_AGEMA_signal_5496), .Q (new_AGEMA_signal_5497) ) ;
    buf_clk new_AGEMA_reg_buffer_2070 ( .C (clk), .D (new_AGEMA_signal_5500), .Q (new_AGEMA_signal_5501) ) ;
    buf_clk new_AGEMA_reg_buffer_2074 ( .C (clk), .D (new_AGEMA_signal_5504), .Q (new_AGEMA_signal_5505) ) ;
    buf_clk new_AGEMA_reg_buffer_2078 ( .C (clk), .D (new_AGEMA_signal_5508), .Q (new_AGEMA_signal_5509) ) ;
    buf_clk new_AGEMA_reg_buffer_2082 ( .C (clk), .D (new_AGEMA_signal_5512), .Q (new_AGEMA_signal_5513) ) ;
    buf_clk new_AGEMA_reg_buffer_2086 ( .C (clk), .D (new_AGEMA_signal_5516), .Q (new_AGEMA_signal_5517) ) ;
    buf_clk new_AGEMA_reg_buffer_2090 ( .C (clk), .D (new_AGEMA_signal_5520), .Q (new_AGEMA_signal_5521) ) ;
    buf_clk new_AGEMA_reg_buffer_2094 ( .C (clk), .D (new_AGEMA_signal_5524), .Q (new_AGEMA_signal_5525) ) ;
    buf_clk new_AGEMA_reg_buffer_2098 ( .C (clk), .D (new_AGEMA_signal_5528), .Q (new_AGEMA_signal_5529) ) ;
    buf_clk new_AGEMA_reg_buffer_2102 ( .C (clk), .D (new_AGEMA_signal_5532), .Q (new_AGEMA_signal_5533) ) ;
    buf_clk new_AGEMA_reg_buffer_2106 ( .C (clk), .D (new_AGEMA_signal_5536), .Q (new_AGEMA_signal_5537) ) ;
    buf_clk new_AGEMA_reg_buffer_2110 ( .C (clk), .D (new_AGEMA_signal_5540), .Q (new_AGEMA_signal_5541) ) ;
    buf_clk new_AGEMA_reg_buffer_2114 ( .C (clk), .D (new_AGEMA_signal_5544), .Q (new_AGEMA_signal_5545) ) ;
    buf_clk new_AGEMA_reg_buffer_2118 ( .C (clk), .D (new_AGEMA_signal_5548), .Q (new_AGEMA_signal_5549) ) ;
    buf_clk new_AGEMA_reg_buffer_2122 ( .C (clk), .D (new_AGEMA_signal_5552), .Q (new_AGEMA_signal_5553) ) ;
    buf_clk new_AGEMA_reg_buffer_2126 ( .C (clk), .D (new_AGEMA_signal_5556), .Q (new_AGEMA_signal_5557) ) ;
    buf_clk new_AGEMA_reg_buffer_2130 ( .C (clk), .D (new_AGEMA_signal_5560), .Q (new_AGEMA_signal_5561) ) ;
    buf_clk new_AGEMA_reg_buffer_2134 ( .C (clk), .D (new_AGEMA_signal_5564), .Q (new_AGEMA_signal_5565) ) ;
    buf_clk new_AGEMA_reg_buffer_2138 ( .C (clk), .D (new_AGEMA_signal_5568), .Q (new_AGEMA_signal_5569) ) ;
    buf_clk new_AGEMA_reg_buffer_2142 ( .C (clk), .D (new_AGEMA_signal_5572), .Q (new_AGEMA_signal_5573) ) ;
    buf_clk new_AGEMA_reg_buffer_2146 ( .C (clk), .D (new_AGEMA_signal_5576), .Q (new_AGEMA_signal_5577) ) ;
    buf_clk new_AGEMA_reg_buffer_2150 ( .C (clk), .D (new_AGEMA_signal_5580), .Q (new_AGEMA_signal_5581) ) ;
    buf_clk new_AGEMA_reg_buffer_2154 ( .C (clk), .D (new_AGEMA_signal_5584), .Q (new_AGEMA_signal_5585) ) ;
    buf_clk new_AGEMA_reg_buffer_2158 ( .C (clk), .D (new_AGEMA_signal_5588), .Q (new_AGEMA_signal_5589) ) ;
    buf_clk new_AGEMA_reg_buffer_2162 ( .C (clk), .D (new_AGEMA_signal_5592), .Q (new_AGEMA_signal_5593) ) ;
    buf_clk new_AGEMA_reg_buffer_2166 ( .C (clk), .D (new_AGEMA_signal_5596), .Q (new_AGEMA_signal_5597) ) ;
    buf_clk new_AGEMA_reg_buffer_2170 ( .C (clk), .D (new_AGEMA_signal_5600), .Q (new_AGEMA_signal_5601) ) ;
    buf_clk new_AGEMA_reg_buffer_2174 ( .C (clk), .D (new_AGEMA_signal_5604), .Q (new_AGEMA_signal_5605) ) ;
    buf_clk new_AGEMA_reg_buffer_2178 ( .C (clk), .D (new_AGEMA_signal_5608), .Q (new_AGEMA_signal_5609) ) ;
    buf_clk new_AGEMA_reg_buffer_2182 ( .C (clk), .D (new_AGEMA_signal_5612), .Q (new_AGEMA_signal_5613) ) ;
    buf_clk new_AGEMA_reg_buffer_2186 ( .C (clk), .D (new_AGEMA_signal_5616), .Q (new_AGEMA_signal_5617) ) ;
    buf_clk new_AGEMA_reg_buffer_2190 ( .C (clk), .D (new_AGEMA_signal_5620), .Q (new_AGEMA_signal_5621) ) ;
    buf_clk new_AGEMA_reg_buffer_2194 ( .C (clk), .D (new_AGEMA_signal_5624), .Q (new_AGEMA_signal_5625) ) ;
    buf_clk new_AGEMA_reg_buffer_2198 ( .C (clk), .D (new_AGEMA_signal_5628), .Q (new_AGEMA_signal_5629) ) ;
    buf_clk new_AGEMA_reg_buffer_2202 ( .C (clk), .D (new_AGEMA_signal_5632), .Q (new_AGEMA_signal_5633) ) ;
    buf_clk new_AGEMA_reg_buffer_2206 ( .C (clk), .D (new_AGEMA_signal_5636), .Q (new_AGEMA_signal_5637) ) ;
    buf_clk new_AGEMA_reg_buffer_2210 ( .C (clk), .D (new_AGEMA_signal_5640), .Q (new_AGEMA_signal_5641) ) ;
    buf_clk new_AGEMA_reg_buffer_2214 ( .C (clk), .D (new_AGEMA_signal_5644), .Q (new_AGEMA_signal_5645) ) ;
    buf_clk new_AGEMA_reg_buffer_2218 ( .C (clk), .D (new_AGEMA_signal_5648), .Q (new_AGEMA_signal_5649) ) ;
    buf_clk new_AGEMA_reg_buffer_2222 ( .C (clk), .D (new_AGEMA_signal_5652), .Q (new_AGEMA_signal_5653) ) ;
    buf_clk new_AGEMA_reg_buffer_2226 ( .C (clk), .D (new_AGEMA_signal_5656), .Q (new_AGEMA_signal_5657) ) ;
    buf_clk new_AGEMA_reg_buffer_2230 ( .C (clk), .D (new_AGEMA_signal_5660), .Q (new_AGEMA_signal_5661) ) ;
    buf_clk new_AGEMA_reg_buffer_2234 ( .C (clk), .D (new_AGEMA_signal_5664), .Q (new_AGEMA_signal_5665) ) ;
    buf_clk new_AGEMA_reg_buffer_2238 ( .C (clk), .D (new_AGEMA_signal_5668), .Q (new_AGEMA_signal_5669) ) ;
    buf_clk new_AGEMA_reg_buffer_2242 ( .C (clk), .D (new_AGEMA_signal_5672), .Q (new_AGEMA_signal_5673) ) ;
    buf_clk new_AGEMA_reg_buffer_2246 ( .C (clk), .D (new_AGEMA_signal_5676), .Q (new_AGEMA_signal_5677) ) ;
    buf_clk new_AGEMA_reg_buffer_2250 ( .C (clk), .D (new_AGEMA_signal_5680), .Q (new_AGEMA_signal_5681) ) ;
    buf_clk new_AGEMA_reg_buffer_2254 ( .C (clk), .D (new_AGEMA_signal_5684), .Q (new_AGEMA_signal_5685) ) ;
    buf_clk new_AGEMA_reg_buffer_2258 ( .C (clk), .D (new_AGEMA_signal_5688), .Q (new_AGEMA_signal_5689) ) ;
    buf_clk new_AGEMA_reg_buffer_2262 ( .C (clk), .D (new_AGEMA_signal_5692), .Q (new_AGEMA_signal_5693) ) ;
    buf_clk new_AGEMA_reg_buffer_2266 ( .C (clk), .D (new_AGEMA_signal_5696), .Q (new_AGEMA_signal_5697) ) ;
    buf_clk new_AGEMA_reg_buffer_2270 ( .C (clk), .D (new_AGEMA_signal_5700), .Q (new_AGEMA_signal_5701) ) ;
    buf_clk new_AGEMA_reg_buffer_2274 ( .C (clk), .D (new_AGEMA_signal_5704), .Q (new_AGEMA_signal_5705) ) ;
    buf_clk new_AGEMA_reg_buffer_2278 ( .C (clk), .D (new_AGEMA_signal_5708), .Q (new_AGEMA_signal_5709) ) ;
    buf_clk new_AGEMA_reg_buffer_2282 ( .C (clk), .D (new_AGEMA_signal_5712), .Q (new_AGEMA_signal_5713) ) ;
    buf_clk new_AGEMA_reg_buffer_2286 ( .C (clk), .D (new_AGEMA_signal_5716), .Q (new_AGEMA_signal_5717) ) ;
    buf_clk new_AGEMA_reg_buffer_2290 ( .C (clk), .D (new_AGEMA_signal_5720), .Q (new_AGEMA_signal_5721) ) ;
    buf_clk new_AGEMA_reg_buffer_2294 ( .C (clk), .D (new_AGEMA_signal_5724), .Q (new_AGEMA_signal_5725) ) ;
    buf_clk new_AGEMA_reg_buffer_2298 ( .C (clk), .D (new_AGEMA_signal_5728), .Q (new_AGEMA_signal_5729) ) ;
    buf_clk new_AGEMA_reg_buffer_2302 ( .C (clk), .D (new_AGEMA_signal_5732), .Q (new_AGEMA_signal_5733) ) ;
    buf_clk new_AGEMA_reg_buffer_2306 ( .C (clk), .D (new_AGEMA_signal_5736), .Q (new_AGEMA_signal_5737) ) ;
    buf_clk new_AGEMA_reg_buffer_2310 ( .C (clk), .D (new_AGEMA_signal_5740), .Q (new_AGEMA_signal_5741) ) ;
    buf_clk new_AGEMA_reg_buffer_2314 ( .C (clk), .D (new_AGEMA_signal_5744), .Q (new_AGEMA_signal_5745) ) ;
    buf_clk new_AGEMA_reg_buffer_2318 ( .C (clk), .D (new_AGEMA_signal_5748), .Q (new_AGEMA_signal_5749) ) ;
    buf_clk new_AGEMA_reg_buffer_2322 ( .C (clk), .D (new_AGEMA_signal_5752), .Q (new_AGEMA_signal_5753) ) ;
    buf_clk new_AGEMA_reg_buffer_2326 ( .C (clk), .D (new_AGEMA_signal_5756), .Q (new_AGEMA_signal_5757) ) ;
    buf_clk new_AGEMA_reg_buffer_2330 ( .C (clk), .D (new_AGEMA_signal_5760), .Q (new_AGEMA_signal_5761) ) ;
    buf_clk new_AGEMA_reg_buffer_2334 ( .C (clk), .D (new_AGEMA_signal_5764), .Q (new_AGEMA_signal_5765) ) ;
    buf_clk new_AGEMA_reg_buffer_2338 ( .C (clk), .D (new_AGEMA_signal_5768), .Q (new_AGEMA_signal_5769) ) ;
    buf_clk new_AGEMA_reg_buffer_2342 ( .C (clk), .D (new_AGEMA_signal_5772), .Q (new_AGEMA_signal_5773) ) ;
    buf_clk new_AGEMA_reg_buffer_2346 ( .C (clk), .D (new_AGEMA_signal_5776), .Q (new_AGEMA_signal_5777) ) ;
    buf_clk new_AGEMA_reg_buffer_2350 ( .C (clk), .D (new_AGEMA_signal_5780), .Q (new_AGEMA_signal_5781) ) ;
    buf_clk new_AGEMA_reg_buffer_2354 ( .C (clk), .D (new_AGEMA_signal_5784), .Q (new_AGEMA_signal_5785) ) ;
    buf_clk new_AGEMA_reg_buffer_2358 ( .C (clk), .D (new_AGEMA_signal_5788), .Q (new_AGEMA_signal_5789) ) ;
    buf_clk new_AGEMA_reg_buffer_2362 ( .C (clk), .D (new_AGEMA_signal_5792), .Q (new_AGEMA_signal_5793) ) ;
    buf_clk new_AGEMA_reg_buffer_2366 ( .C (clk), .D (new_AGEMA_signal_5796), .Q (new_AGEMA_signal_5797) ) ;
    buf_clk new_AGEMA_reg_buffer_2370 ( .C (clk), .D (new_AGEMA_signal_5800), .Q (new_AGEMA_signal_5801) ) ;
    buf_clk new_AGEMA_reg_buffer_2374 ( .C (clk), .D (new_AGEMA_signal_5804), .Q (new_AGEMA_signal_5805) ) ;
    buf_clk new_AGEMA_reg_buffer_2378 ( .C (clk), .D (new_AGEMA_signal_5808), .Q (new_AGEMA_signal_5809) ) ;
    buf_clk new_AGEMA_reg_buffer_2382 ( .C (clk), .D (new_AGEMA_signal_5812), .Q (new_AGEMA_signal_5813) ) ;
    buf_clk new_AGEMA_reg_buffer_2386 ( .C (clk), .D (new_AGEMA_signal_5816), .Q (new_AGEMA_signal_5817) ) ;
    buf_clk new_AGEMA_reg_buffer_2390 ( .C (clk), .D (new_AGEMA_signal_5820), .Q (new_AGEMA_signal_5821) ) ;
    buf_clk new_AGEMA_reg_buffer_2394 ( .C (clk), .D (new_AGEMA_signal_5824), .Q (new_AGEMA_signal_5825) ) ;
    buf_clk new_AGEMA_reg_buffer_2398 ( .C (clk), .D (new_AGEMA_signal_5828), .Q (new_AGEMA_signal_5829) ) ;
    buf_clk new_AGEMA_reg_buffer_2402 ( .C (clk), .D (new_AGEMA_signal_5832), .Q (new_AGEMA_signal_5833) ) ;
    buf_clk new_AGEMA_reg_buffer_2406 ( .C (clk), .D (new_AGEMA_signal_5836), .Q (new_AGEMA_signal_5837) ) ;
    buf_clk new_AGEMA_reg_buffer_2410 ( .C (clk), .D (new_AGEMA_signal_5840), .Q (new_AGEMA_signal_5841) ) ;
    buf_clk new_AGEMA_reg_buffer_2414 ( .C (clk), .D (new_AGEMA_signal_5844), .Q (new_AGEMA_signal_5845) ) ;
    buf_clk new_AGEMA_reg_buffer_2424 ( .C (clk), .D (SubCellInst_SboxInst_0_T2), .Q (new_AGEMA_signal_5855) ) ;
    buf_clk new_AGEMA_reg_buffer_2426 ( .C (clk), .D (new_AGEMA_signal_2319), .Q (new_AGEMA_signal_5857) ) ;
    buf_clk new_AGEMA_reg_buffer_2428 ( .C (clk), .D (new_AGEMA_signal_2320), .Q (new_AGEMA_signal_5859) ) ;
    buf_clk new_AGEMA_reg_buffer_2430 ( .C (clk), .D (new_AGEMA_signal_2321), .Q (new_AGEMA_signal_5861) ) ;
    buf_clk new_AGEMA_reg_buffer_2442 ( .C (clk), .D (new_AGEMA_signal_5872), .Q (new_AGEMA_signal_5873) ) ;
    buf_clk new_AGEMA_reg_buffer_2446 ( .C (clk), .D (new_AGEMA_signal_5876), .Q (new_AGEMA_signal_5877) ) ;
    buf_clk new_AGEMA_reg_buffer_2450 ( .C (clk), .D (new_AGEMA_signal_5880), .Q (new_AGEMA_signal_5881) ) ;
    buf_clk new_AGEMA_reg_buffer_2454 ( .C (clk), .D (new_AGEMA_signal_5884), .Q (new_AGEMA_signal_5885) ) ;
    buf_clk new_AGEMA_reg_buffer_2456 ( .C (clk), .D (SubCellInst_SboxInst_0_YY_1_), .Q (new_AGEMA_signal_5887) ) ;
    buf_clk new_AGEMA_reg_buffer_2458 ( .C (clk), .D (new_AGEMA_signal_2661), .Q (new_AGEMA_signal_5889) ) ;
    buf_clk new_AGEMA_reg_buffer_2460 ( .C (clk), .D (new_AGEMA_signal_2662), .Q (new_AGEMA_signal_5891) ) ;
    buf_clk new_AGEMA_reg_buffer_2462 ( .C (clk), .D (new_AGEMA_signal_2663), .Q (new_AGEMA_signal_5893) ) ;
    buf_clk new_AGEMA_reg_buffer_2472 ( .C (clk), .D (SubCellInst_SboxInst_1_T2), .Q (new_AGEMA_signal_5903) ) ;
    buf_clk new_AGEMA_reg_buffer_2474 ( .C (clk), .D (new_AGEMA_signal_2328), .Q (new_AGEMA_signal_5905) ) ;
    buf_clk new_AGEMA_reg_buffer_2476 ( .C (clk), .D (new_AGEMA_signal_2329), .Q (new_AGEMA_signal_5907) ) ;
    buf_clk new_AGEMA_reg_buffer_2478 ( .C (clk), .D (new_AGEMA_signal_2330), .Q (new_AGEMA_signal_5909) ) ;
    buf_clk new_AGEMA_reg_buffer_2490 ( .C (clk), .D (new_AGEMA_signal_5920), .Q (new_AGEMA_signal_5921) ) ;
    buf_clk new_AGEMA_reg_buffer_2494 ( .C (clk), .D (new_AGEMA_signal_5924), .Q (new_AGEMA_signal_5925) ) ;
    buf_clk new_AGEMA_reg_buffer_2498 ( .C (clk), .D (new_AGEMA_signal_5928), .Q (new_AGEMA_signal_5929) ) ;
    buf_clk new_AGEMA_reg_buffer_2502 ( .C (clk), .D (new_AGEMA_signal_5932), .Q (new_AGEMA_signal_5933) ) ;
    buf_clk new_AGEMA_reg_buffer_2504 ( .C (clk), .D (SubCellInst_SboxInst_1_YY_1_), .Q (new_AGEMA_signal_5935) ) ;
    buf_clk new_AGEMA_reg_buffer_2506 ( .C (clk), .D (new_AGEMA_signal_2673), .Q (new_AGEMA_signal_5937) ) ;
    buf_clk new_AGEMA_reg_buffer_2508 ( .C (clk), .D (new_AGEMA_signal_2674), .Q (new_AGEMA_signal_5939) ) ;
    buf_clk new_AGEMA_reg_buffer_2510 ( .C (clk), .D (new_AGEMA_signal_2675), .Q (new_AGEMA_signal_5941) ) ;
    buf_clk new_AGEMA_reg_buffer_2520 ( .C (clk), .D (SubCellInst_SboxInst_2_T2), .Q (new_AGEMA_signal_5951) ) ;
    buf_clk new_AGEMA_reg_buffer_2522 ( .C (clk), .D (new_AGEMA_signal_2337), .Q (new_AGEMA_signal_5953) ) ;
    buf_clk new_AGEMA_reg_buffer_2524 ( .C (clk), .D (new_AGEMA_signal_2338), .Q (new_AGEMA_signal_5955) ) ;
    buf_clk new_AGEMA_reg_buffer_2526 ( .C (clk), .D (new_AGEMA_signal_2339), .Q (new_AGEMA_signal_5957) ) ;
    buf_clk new_AGEMA_reg_buffer_2538 ( .C (clk), .D (new_AGEMA_signal_5968), .Q (new_AGEMA_signal_5969) ) ;
    buf_clk new_AGEMA_reg_buffer_2542 ( .C (clk), .D (new_AGEMA_signal_5972), .Q (new_AGEMA_signal_5973) ) ;
    buf_clk new_AGEMA_reg_buffer_2546 ( .C (clk), .D (new_AGEMA_signal_5976), .Q (new_AGEMA_signal_5977) ) ;
    buf_clk new_AGEMA_reg_buffer_2550 ( .C (clk), .D (new_AGEMA_signal_5980), .Q (new_AGEMA_signal_5981) ) ;
    buf_clk new_AGEMA_reg_buffer_2552 ( .C (clk), .D (SubCellInst_SboxInst_2_YY_1_), .Q (new_AGEMA_signal_5983) ) ;
    buf_clk new_AGEMA_reg_buffer_2554 ( .C (clk), .D (new_AGEMA_signal_2685), .Q (new_AGEMA_signal_5985) ) ;
    buf_clk new_AGEMA_reg_buffer_2556 ( .C (clk), .D (new_AGEMA_signal_2686), .Q (new_AGEMA_signal_5987) ) ;
    buf_clk new_AGEMA_reg_buffer_2558 ( .C (clk), .D (new_AGEMA_signal_2687), .Q (new_AGEMA_signal_5989) ) ;
    buf_clk new_AGEMA_reg_buffer_2568 ( .C (clk), .D (SubCellInst_SboxInst_3_T2), .Q (new_AGEMA_signal_5999) ) ;
    buf_clk new_AGEMA_reg_buffer_2570 ( .C (clk), .D (new_AGEMA_signal_2346), .Q (new_AGEMA_signal_6001) ) ;
    buf_clk new_AGEMA_reg_buffer_2572 ( .C (clk), .D (new_AGEMA_signal_2347), .Q (new_AGEMA_signal_6003) ) ;
    buf_clk new_AGEMA_reg_buffer_2574 ( .C (clk), .D (new_AGEMA_signal_2348), .Q (new_AGEMA_signal_6005) ) ;
    buf_clk new_AGEMA_reg_buffer_2586 ( .C (clk), .D (new_AGEMA_signal_6016), .Q (new_AGEMA_signal_6017) ) ;
    buf_clk new_AGEMA_reg_buffer_2590 ( .C (clk), .D (new_AGEMA_signal_6020), .Q (new_AGEMA_signal_6021) ) ;
    buf_clk new_AGEMA_reg_buffer_2594 ( .C (clk), .D (new_AGEMA_signal_6024), .Q (new_AGEMA_signal_6025) ) ;
    buf_clk new_AGEMA_reg_buffer_2598 ( .C (clk), .D (new_AGEMA_signal_6028), .Q (new_AGEMA_signal_6029) ) ;
    buf_clk new_AGEMA_reg_buffer_2600 ( .C (clk), .D (SubCellInst_SboxInst_3_YY_1_), .Q (new_AGEMA_signal_6031) ) ;
    buf_clk new_AGEMA_reg_buffer_2602 ( .C (clk), .D (new_AGEMA_signal_2697), .Q (new_AGEMA_signal_6033) ) ;
    buf_clk new_AGEMA_reg_buffer_2604 ( .C (clk), .D (new_AGEMA_signal_2698), .Q (new_AGEMA_signal_6035) ) ;
    buf_clk new_AGEMA_reg_buffer_2606 ( .C (clk), .D (new_AGEMA_signal_2699), .Q (new_AGEMA_signal_6037) ) ;
    buf_clk new_AGEMA_reg_buffer_2616 ( .C (clk), .D (SubCellInst_SboxInst_4_T2), .Q (new_AGEMA_signal_6047) ) ;
    buf_clk new_AGEMA_reg_buffer_2618 ( .C (clk), .D (new_AGEMA_signal_2355), .Q (new_AGEMA_signal_6049) ) ;
    buf_clk new_AGEMA_reg_buffer_2620 ( .C (clk), .D (new_AGEMA_signal_2356), .Q (new_AGEMA_signal_6051) ) ;
    buf_clk new_AGEMA_reg_buffer_2622 ( .C (clk), .D (new_AGEMA_signal_2357), .Q (new_AGEMA_signal_6053) ) ;
    buf_clk new_AGEMA_reg_buffer_2634 ( .C (clk), .D (new_AGEMA_signal_6064), .Q (new_AGEMA_signal_6065) ) ;
    buf_clk new_AGEMA_reg_buffer_2638 ( .C (clk), .D (new_AGEMA_signal_6068), .Q (new_AGEMA_signal_6069) ) ;
    buf_clk new_AGEMA_reg_buffer_2642 ( .C (clk), .D (new_AGEMA_signal_6072), .Q (new_AGEMA_signal_6073) ) ;
    buf_clk new_AGEMA_reg_buffer_2646 ( .C (clk), .D (new_AGEMA_signal_6076), .Q (new_AGEMA_signal_6077) ) ;
    buf_clk new_AGEMA_reg_buffer_2648 ( .C (clk), .D (SubCellInst_SboxInst_4_YY_1_), .Q (new_AGEMA_signal_6079) ) ;
    buf_clk new_AGEMA_reg_buffer_2650 ( .C (clk), .D (new_AGEMA_signal_2709), .Q (new_AGEMA_signal_6081) ) ;
    buf_clk new_AGEMA_reg_buffer_2652 ( .C (clk), .D (new_AGEMA_signal_2710), .Q (new_AGEMA_signal_6083) ) ;
    buf_clk new_AGEMA_reg_buffer_2654 ( .C (clk), .D (new_AGEMA_signal_2711), .Q (new_AGEMA_signal_6085) ) ;
    buf_clk new_AGEMA_reg_buffer_2664 ( .C (clk), .D (SubCellInst_SboxInst_5_T2), .Q (new_AGEMA_signal_6095) ) ;
    buf_clk new_AGEMA_reg_buffer_2666 ( .C (clk), .D (new_AGEMA_signal_2364), .Q (new_AGEMA_signal_6097) ) ;
    buf_clk new_AGEMA_reg_buffer_2668 ( .C (clk), .D (new_AGEMA_signal_2365), .Q (new_AGEMA_signal_6099) ) ;
    buf_clk new_AGEMA_reg_buffer_2670 ( .C (clk), .D (new_AGEMA_signal_2366), .Q (new_AGEMA_signal_6101) ) ;
    buf_clk new_AGEMA_reg_buffer_2682 ( .C (clk), .D (new_AGEMA_signal_6112), .Q (new_AGEMA_signal_6113) ) ;
    buf_clk new_AGEMA_reg_buffer_2686 ( .C (clk), .D (new_AGEMA_signal_6116), .Q (new_AGEMA_signal_6117) ) ;
    buf_clk new_AGEMA_reg_buffer_2690 ( .C (clk), .D (new_AGEMA_signal_6120), .Q (new_AGEMA_signal_6121) ) ;
    buf_clk new_AGEMA_reg_buffer_2694 ( .C (clk), .D (new_AGEMA_signal_6124), .Q (new_AGEMA_signal_6125) ) ;
    buf_clk new_AGEMA_reg_buffer_2696 ( .C (clk), .D (SubCellInst_SboxInst_5_YY_1_), .Q (new_AGEMA_signal_6127) ) ;
    buf_clk new_AGEMA_reg_buffer_2698 ( .C (clk), .D (new_AGEMA_signal_2721), .Q (new_AGEMA_signal_6129) ) ;
    buf_clk new_AGEMA_reg_buffer_2700 ( .C (clk), .D (new_AGEMA_signal_2722), .Q (new_AGEMA_signal_6131) ) ;
    buf_clk new_AGEMA_reg_buffer_2702 ( .C (clk), .D (new_AGEMA_signal_2723), .Q (new_AGEMA_signal_6133) ) ;
    buf_clk new_AGEMA_reg_buffer_2712 ( .C (clk), .D (SubCellInst_SboxInst_6_T2), .Q (new_AGEMA_signal_6143) ) ;
    buf_clk new_AGEMA_reg_buffer_2714 ( .C (clk), .D (new_AGEMA_signal_2373), .Q (new_AGEMA_signal_6145) ) ;
    buf_clk new_AGEMA_reg_buffer_2716 ( .C (clk), .D (new_AGEMA_signal_2374), .Q (new_AGEMA_signal_6147) ) ;
    buf_clk new_AGEMA_reg_buffer_2718 ( .C (clk), .D (new_AGEMA_signal_2375), .Q (new_AGEMA_signal_6149) ) ;
    buf_clk new_AGEMA_reg_buffer_2730 ( .C (clk), .D (new_AGEMA_signal_6160), .Q (new_AGEMA_signal_6161) ) ;
    buf_clk new_AGEMA_reg_buffer_2734 ( .C (clk), .D (new_AGEMA_signal_6164), .Q (new_AGEMA_signal_6165) ) ;
    buf_clk new_AGEMA_reg_buffer_2738 ( .C (clk), .D (new_AGEMA_signal_6168), .Q (new_AGEMA_signal_6169) ) ;
    buf_clk new_AGEMA_reg_buffer_2742 ( .C (clk), .D (new_AGEMA_signal_6172), .Q (new_AGEMA_signal_6173) ) ;
    buf_clk new_AGEMA_reg_buffer_2744 ( .C (clk), .D (SubCellInst_SboxInst_6_YY_1_), .Q (new_AGEMA_signal_6175) ) ;
    buf_clk new_AGEMA_reg_buffer_2746 ( .C (clk), .D (new_AGEMA_signal_2733), .Q (new_AGEMA_signal_6177) ) ;
    buf_clk new_AGEMA_reg_buffer_2748 ( .C (clk), .D (new_AGEMA_signal_2734), .Q (new_AGEMA_signal_6179) ) ;
    buf_clk new_AGEMA_reg_buffer_2750 ( .C (clk), .D (new_AGEMA_signal_2735), .Q (new_AGEMA_signal_6181) ) ;
    buf_clk new_AGEMA_reg_buffer_2760 ( .C (clk), .D (SubCellInst_SboxInst_7_T2), .Q (new_AGEMA_signal_6191) ) ;
    buf_clk new_AGEMA_reg_buffer_2762 ( .C (clk), .D (new_AGEMA_signal_2382), .Q (new_AGEMA_signal_6193) ) ;
    buf_clk new_AGEMA_reg_buffer_2764 ( .C (clk), .D (new_AGEMA_signal_2383), .Q (new_AGEMA_signal_6195) ) ;
    buf_clk new_AGEMA_reg_buffer_2766 ( .C (clk), .D (new_AGEMA_signal_2384), .Q (new_AGEMA_signal_6197) ) ;
    buf_clk new_AGEMA_reg_buffer_2778 ( .C (clk), .D (new_AGEMA_signal_6208), .Q (new_AGEMA_signal_6209) ) ;
    buf_clk new_AGEMA_reg_buffer_2782 ( .C (clk), .D (new_AGEMA_signal_6212), .Q (new_AGEMA_signal_6213) ) ;
    buf_clk new_AGEMA_reg_buffer_2786 ( .C (clk), .D (new_AGEMA_signal_6216), .Q (new_AGEMA_signal_6217) ) ;
    buf_clk new_AGEMA_reg_buffer_2790 ( .C (clk), .D (new_AGEMA_signal_6220), .Q (new_AGEMA_signal_6221) ) ;
    buf_clk new_AGEMA_reg_buffer_2792 ( .C (clk), .D (SubCellInst_SboxInst_7_YY_1_), .Q (new_AGEMA_signal_6223) ) ;
    buf_clk new_AGEMA_reg_buffer_2794 ( .C (clk), .D (new_AGEMA_signal_2745), .Q (new_AGEMA_signal_6225) ) ;
    buf_clk new_AGEMA_reg_buffer_2796 ( .C (clk), .D (new_AGEMA_signal_2746), .Q (new_AGEMA_signal_6227) ) ;
    buf_clk new_AGEMA_reg_buffer_2798 ( .C (clk), .D (new_AGEMA_signal_2747), .Q (new_AGEMA_signal_6229) ) ;
    buf_clk new_AGEMA_reg_buffer_2808 ( .C (clk), .D (SubCellInst_SboxInst_8_T2), .Q (new_AGEMA_signal_6239) ) ;
    buf_clk new_AGEMA_reg_buffer_2810 ( .C (clk), .D (new_AGEMA_signal_2391), .Q (new_AGEMA_signal_6241) ) ;
    buf_clk new_AGEMA_reg_buffer_2812 ( .C (clk), .D (new_AGEMA_signal_2392), .Q (new_AGEMA_signal_6243) ) ;
    buf_clk new_AGEMA_reg_buffer_2814 ( .C (clk), .D (new_AGEMA_signal_2393), .Q (new_AGEMA_signal_6245) ) ;
    buf_clk new_AGEMA_reg_buffer_2826 ( .C (clk), .D (new_AGEMA_signal_6256), .Q (new_AGEMA_signal_6257) ) ;
    buf_clk new_AGEMA_reg_buffer_2830 ( .C (clk), .D (new_AGEMA_signal_6260), .Q (new_AGEMA_signal_6261) ) ;
    buf_clk new_AGEMA_reg_buffer_2834 ( .C (clk), .D (new_AGEMA_signal_6264), .Q (new_AGEMA_signal_6265) ) ;
    buf_clk new_AGEMA_reg_buffer_2838 ( .C (clk), .D (new_AGEMA_signal_6268), .Q (new_AGEMA_signal_6269) ) ;
    buf_clk new_AGEMA_reg_buffer_2840 ( .C (clk), .D (SubCellInst_SboxInst_8_YY_1_), .Q (new_AGEMA_signal_6271) ) ;
    buf_clk new_AGEMA_reg_buffer_2842 ( .C (clk), .D (new_AGEMA_signal_2757), .Q (new_AGEMA_signal_6273) ) ;
    buf_clk new_AGEMA_reg_buffer_2844 ( .C (clk), .D (new_AGEMA_signal_2758), .Q (new_AGEMA_signal_6275) ) ;
    buf_clk new_AGEMA_reg_buffer_2846 ( .C (clk), .D (new_AGEMA_signal_2759), .Q (new_AGEMA_signal_6277) ) ;
    buf_clk new_AGEMA_reg_buffer_2856 ( .C (clk), .D (SubCellInst_SboxInst_9_T2), .Q (new_AGEMA_signal_6287) ) ;
    buf_clk new_AGEMA_reg_buffer_2858 ( .C (clk), .D (new_AGEMA_signal_2400), .Q (new_AGEMA_signal_6289) ) ;
    buf_clk new_AGEMA_reg_buffer_2860 ( .C (clk), .D (new_AGEMA_signal_2401), .Q (new_AGEMA_signal_6291) ) ;
    buf_clk new_AGEMA_reg_buffer_2862 ( .C (clk), .D (new_AGEMA_signal_2402), .Q (new_AGEMA_signal_6293) ) ;
    buf_clk new_AGEMA_reg_buffer_2874 ( .C (clk), .D (new_AGEMA_signal_6304), .Q (new_AGEMA_signal_6305) ) ;
    buf_clk new_AGEMA_reg_buffer_2878 ( .C (clk), .D (new_AGEMA_signal_6308), .Q (new_AGEMA_signal_6309) ) ;
    buf_clk new_AGEMA_reg_buffer_2882 ( .C (clk), .D (new_AGEMA_signal_6312), .Q (new_AGEMA_signal_6313) ) ;
    buf_clk new_AGEMA_reg_buffer_2886 ( .C (clk), .D (new_AGEMA_signal_6316), .Q (new_AGEMA_signal_6317) ) ;
    buf_clk new_AGEMA_reg_buffer_2888 ( .C (clk), .D (SubCellInst_SboxInst_9_YY_1_), .Q (new_AGEMA_signal_6319) ) ;
    buf_clk new_AGEMA_reg_buffer_2890 ( .C (clk), .D (new_AGEMA_signal_2769), .Q (new_AGEMA_signal_6321) ) ;
    buf_clk new_AGEMA_reg_buffer_2892 ( .C (clk), .D (new_AGEMA_signal_2770), .Q (new_AGEMA_signal_6323) ) ;
    buf_clk new_AGEMA_reg_buffer_2894 ( .C (clk), .D (new_AGEMA_signal_2771), .Q (new_AGEMA_signal_6325) ) ;
    buf_clk new_AGEMA_reg_buffer_2904 ( .C (clk), .D (SubCellInst_SboxInst_10_T2), .Q (new_AGEMA_signal_6335) ) ;
    buf_clk new_AGEMA_reg_buffer_2906 ( .C (clk), .D (new_AGEMA_signal_2409), .Q (new_AGEMA_signal_6337) ) ;
    buf_clk new_AGEMA_reg_buffer_2908 ( .C (clk), .D (new_AGEMA_signal_2410), .Q (new_AGEMA_signal_6339) ) ;
    buf_clk new_AGEMA_reg_buffer_2910 ( .C (clk), .D (new_AGEMA_signal_2411), .Q (new_AGEMA_signal_6341) ) ;
    buf_clk new_AGEMA_reg_buffer_2922 ( .C (clk), .D (new_AGEMA_signal_6352), .Q (new_AGEMA_signal_6353) ) ;
    buf_clk new_AGEMA_reg_buffer_2926 ( .C (clk), .D (new_AGEMA_signal_6356), .Q (new_AGEMA_signal_6357) ) ;
    buf_clk new_AGEMA_reg_buffer_2930 ( .C (clk), .D (new_AGEMA_signal_6360), .Q (new_AGEMA_signal_6361) ) ;
    buf_clk new_AGEMA_reg_buffer_2934 ( .C (clk), .D (new_AGEMA_signal_6364), .Q (new_AGEMA_signal_6365) ) ;
    buf_clk new_AGEMA_reg_buffer_2936 ( .C (clk), .D (SubCellInst_SboxInst_10_YY_1_), .Q (new_AGEMA_signal_6367) ) ;
    buf_clk new_AGEMA_reg_buffer_2938 ( .C (clk), .D (new_AGEMA_signal_2781), .Q (new_AGEMA_signal_6369) ) ;
    buf_clk new_AGEMA_reg_buffer_2940 ( .C (clk), .D (new_AGEMA_signal_2782), .Q (new_AGEMA_signal_6371) ) ;
    buf_clk new_AGEMA_reg_buffer_2942 ( .C (clk), .D (new_AGEMA_signal_2783), .Q (new_AGEMA_signal_6373) ) ;
    buf_clk new_AGEMA_reg_buffer_2952 ( .C (clk), .D (SubCellInst_SboxInst_11_T2), .Q (new_AGEMA_signal_6383) ) ;
    buf_clk new_AGEMA_reg_buffer_2954 ( .C (clk), .D (new_AGEMA_signal_2418), .Q (new_AGEMA_signal_6385) ) ;
    buf_clk new_AGEMA_reg_buffer_2956 ( .C (clk), .D (new_AGEMA_signal_2419), .Q (new_AGEMA_signal_6387) ) ;
    buf_clk new_AGEMA_reg_buffer_2958 ( .C (clk), .D (new_AGEMA_signal_2420), .Q (new_AGEMA_signal_6389) ) ;
    buf_clk new_AGEMA_reg_buffer_2970 ( .C (clk), .D (new_AGEMA_signal_6400), .Q (new_AGEMA_signal_6401) ) ;
    buf_clk new_AGEMA_reg_buffer_2974 ( .C (clk), .D (new_AGEMA_signal_6404), .Q (new_AGEMA_signal_6405) ) ;
    buf_clk new_AGEMA_reg_buffer_2978 ( .C (clk), .D (new_AGEMA_signal_6408), .Q (new_AGEMA_signal_6409) ) ;
    buf_clk new_AGEMA_reg_buffer_2982 ( .C (clk), .D (new_AGEMA_signal_6412), .Q (new_AGEMA_signal_6413) ) ;
    buf_clk new_AGEMA_reg_buffer_2984 ( .C (clk), .D (SubCellInst_SboxInst_11_YY_1_), .Q (new_AGEMA_signal_6415) ) ;
    buf_clk new_AGEMA_reg_buffer_2986 ( .C (clk), .D (new_AGEMA_signal_2793), .Q (new_AGEMA_signal_6417) ) ;
    buf_clk new_AGEMA_reg_buffer_2988 ( .C (clk), .D (new_AGEMA_signal_2794), .Q (new_AGEMA_signal_6419) ) ;
    buf_clk new_AGEMA_reg_buffer_2990 ( .C (clk), .D (new_AGEMA_signal_2795), .Q (new_AGEMA_signal_6421) ) ;
    buf_clk new_AGEMA_reg_buffer_3000 ( .C (clk), .D (SubCellInst_SboxInst_12_T2), .Q (new_AGEMA_signal_6431) ) ;
    buf_clk new_AGEMA_reg_buffer_3002 ( .C (clk), .D (new_AGEMA_signal_2427), .Q (new_AGEMA_signal_6433) ) ;
    buf_clk new_AGEMA_reg_buffer_3004 ( .C (clk), .D (new_AGEMA_signal_2428), .Q (new_AGEMA_signal_6435) ) ;
    buf_clk new_AGEMA_reg_buffer_3006 ( .C (clk), .D (new_AGEMA_signal_2429), .Q (new_AGEMA_signal_6437) ) ;
    buf_clk new_AGEMA_reg_buffer_3018 ( .C (clk), .D (new_AGEMA_signal_6448), .Q (new_AGEMA_signal_6449) ) ;
    buf_clk new_AGEMA_reg_buffer_3022 ( .C (clk), .D (new_AGEMA_signal_6452), .Q (new_AGEMA_signal_6453) ) ;
    buf_clk new_AGEMA_reg_buffer_3026 ( .C (clk), .D (new_AGEMA_signal_6456), .Q (new_AGEMA_signal_6457) ) ;
    buf_clk new_AGEMA_reg_buffer_3030 ( .C (clk), .D (new_AGEMA_signal_6460), .Q (new_AGEMA_signal_6461) ) ;
    buf_clk new_AGEMA_reg_buffer_3032 ( .C (clk), .D (SubCellInst_SboxInst_12_YY_1_), .Q (new_AGEMA_signal_6463) ) ;
    buf_clk new_AGEMA_reg_buffer_3034 ( .C (clk), .D (new_AGEMA_signal_2805), .Q (new_AGEMA_signal_6465) ) ;
    buf_clk new_AGEMA_reg_buffer_3036 ( .C (clk), .D (new_AGEMA_signal_2806), .Q (new_AGEMA_signal_6467) ) ;
    buf_clk new_AGEMA_reg_buffer_3038 ( .C (clk), .D (new_AGEMA_signal_2807), .Q (new_AGEMA_signal_6469) ) ;
    buf_clk new_AGEMA_reg_buffer_3048 ( .C (clk), .D (SubCellInst_SboxInst_13_T2), .Q (new_AGEMA_signal_6479) ) ;
    buf_clk new_AGEMA_reg_buffer_3050 ( .C (clk), .D (new_AGEMA_signal_2436), .Q (new_AGEMA_signal_6481) ) ;
    buf_clk new_AGEMA_reg_buffer_3052 ( .C (clk), .D (new_AGEMA_signal_2437), .Q (new_AGEMA_signal_6483) ) ;
    buf_clk new_AGEMA_reg_buffer_3054 ( .C (clk), .D (new_AGEMA_signal_2438), .Q (new_AGEMA_signal_6485) ) ;
    buf_clk new_AGEMA_reg_buffer_3066 ( .C (clk), .D (new_AGEMA_signal_6496), .Q (new_AGEMA_signal_6497) ) ;
    buf_clk new_AGEMA_reg_buffer_3070 ( .C (clk), .D (new_AGEMA_signal_6500), .Q (new_AGEMA_signal_6501) ) ;
    buf_clk new_AGEMA_reg_buffer_3074 ( .C (clk), .D (new_AGEMA_signal_6504), .Q (new_AGEMA_signal_6505) ) ;
    buf_clk new_AGEMA_reg_buffer_3078 ( .C (clk), .D (new_AGEMA_signal_6508), .Q (new_AGEMA_signal_6509) ) ;
    buf_clk new_AGEMA_reg_buffer_3080 ( .C (clk), .D (SubCellInst_SboxInst_13_YY_1_), .Q (new_AGEMA_signal_6511) ) ;
    buf_clk new_AGEMA_reg_buffer_3082 ( .C (clk), .D (new_AGEMA_signal_2817), .Q (new_AGEMA_signal_6513) ) ;
    buf_clk new_AGEMA_reg_buffer_3084 ( .C (clk), .D (new_AGEMA_signal_2818), .Q (new_AGEMA_signal_6515) ) ;
    buf_clk new_AGEMA_reg_buffer_3086 ( .C (clk), .D (new_AGEMA_signal_2819), .Q (new_AGEMA_signal_6517) ) ;
    buf_clk new_AGEMA_reg_buffer_3096 ( .C (clk), .D (SubCellInst_SboxInst_14_T2), .Q (new_AGEMA_signal_6527) ) ;
    buf_clk new_AGEMA_reg_buffer_3098 ( .C (clk), .D (new_AGEMA_signal_2445), .Q (new_AGEMA_signal_6529) ) ;
    buf_clk new_AGEMA_reg_buffer_3100 ( .C (clk), .D (new_AGEMA_signal_2446), .Q (new_AGEMA_signal_6531) ) ;
    buf_clk new_AGEMA_reg_buffer_3102 ( .C (clk), .D (new_AGEMA_signal_2447), .Q (new_AGEMA_signal_6533) ) ;
    buf_clk new_AGEMA_reg_buffer_3114 ( .C (clk), .D (new_AGEMA_signal_6544), .Q (new_AGEMA_signal_6545) ) ;
    buf_clk new_AGEMA_reg_buffer_3118 ( .C (clk), .D (new_AGEMA_signal_6548), .Q (new_AGEMA_signal_6549) ) ;
    buf_clk new_AGEMA_reg_buffer_3122 ( .C (clk), .D (new_AGEMA_signal_6552), .Q (new_AGEMA_signal_6553) ) ;
    buf_clk new_AGEMA_reg_buffer_3126 ( .C (clk), .D (new_AGEMA_signal_6556), .Q (new_AGEMA_signal_6557) ) ;
    buf_clk new_AGEMA_reg_buffer_3128 ( .C (clk), .D (SubCellInst_SboxInst_14_YY_1_), .Q (new_AGEMA_signal_6559) ) ;
    buf_clk new_AGEMA_reg_buffer_3130 ( .C (clk), .D (new_AGEMA_signal_2829), .Q (new_AGEMA_signal_6561) ) ;
    buf_clk new_AGEMA_reg_buffer_3132 ( .C (clk), .D (new_AGEMA_signal_2830), .Q (new_AGEMA_signal_6563) ) ;
    buf_clk new_AGEMA_reg_buffer_3134 ( .C (clk), .D (new_AGEMA_signal_2831), .Q (new_AGEMA_signal_6565) ) ;
    buf_clk new_AGEMA_reg_buffer_3144 ( .C (clk), .D (SubCellInst_SboxInst_15_T2), .Q (new_AGEMA_signal_6575) ) ;
    buf_clk new_AGEMA_reg_buffer_3146 ( .C (clk), .D (new_AGEMA_signal_2454), .Q (new_AGEMA_signal_6577) ) ;
    buf_clk new_AGEMA_reg_buffer_3148 ( .C (clk), .D (new_AGEMA_signal_2455), .Q (new_AGEMA_signal_6579) ) ;
    buf_clk new_AGEMA_reg_buffer_3150 ( .C (clk), .D (new_AGEMA_signal_2456), .Q (new_AGEMA_signal_6581) ) ;
    buf_clk new_AGEMA_reg_buffer_3162 ( .C (clk), .D (new_AGEMA_signal_6592), .Q (new_AGEMA_signal_6593) ) ;
    buf_clk new_AGEMA_reg_buffer_3166 ( .C (clk), .D (new_AGEMA_signal_6596), .Q (new_AGEMA_signal_6597) ) ;
    buf_clk new_AGEMA_reg_buffer_3170 ( .C (clk), .D (new_AGEMA_signal_6600), .Q (new_AGEMA_signal_6601) ) ;
    buf_clk new_AGEMA_reg_buffer_3174 ( .C (clk), .D (new_AGEMA_signal_6604), .Q (new_AGEMA_signal_6605) ) ;
    buf_clk new_AGEMA_reg_buffer_3176 ( .C (clk), .D (SubCellInst_SboxInst_15_YY_1_), .Q (new_AGEMA_signal_6607) ) ;
    buf_clk new_AGEMA_reg_buffer_3178 ( .C (clk), .D (new_AGEMA_signal_2841), .Q (new_AGEMA_signal_6609) ) ;
    buf_clk new_AGEMA_reg_buffer_3180 ( .C (clk), .D (new_AGEMA_signal_2842), .Q (new_AGEMA_signal_6611) ) ;
    buf_clk new_AGEMA_reg_buffer_3182 ( .C (clk), .D (new_AGEMA_signal_2843), .Q (new_AGEMA_signal_6613) ) ;
    buf_clk new_AGEMA_reg_buffer_3186 ( .C (clk), .D (new_AGEMA_signal_6616), .Q (new_AGEMA_signal_6617) ) ;
    buf_clk new_AGEMA_reg_buffer_3190 ( .C (clk), .D (new_AGEMA_signal_6620), .Q (new_AGEMA_signal_6621) ) ;
    buf_clk new_AGEMA_reg_buffer_3194 ( .C (clk), .D (new_AGEMA_signal_6624), .Q (new_AGEMA_signal_6625) ) ;
    buf_clk new_AGEMA_reg_buffer_3198 ( .C (clk), .D (new_AGEMA_signal_6628), .Q (new_AGEMA_signal_6629) ) ;
    buf_clk new_AGEMA_reg_buffer_3202 ( .C (clk), .D (new_AGEMA_signal_6632), .Q (new_AGEMA_signal_6633) ) ;
    buf_clk new_AGEMA_reg_buffer_3206 ( .C (clk), .D (new_AGEMA_signal_6636), .Q (new_AGEMA_signal_6637) ) ;
    buf_clk new_AGEMA_reg_buffer_3210 ( .C (clk), .D (new_AGEMA_signal_6640), .Q (new_AGEMA_signal_6641) ) ;
    buf_clk new_AGEMA_reg_buffer_3214 ( .C (clk), .D (new_AGEMA_signal_6644), .Q (new_AGEMA_signal_6645) ) ;
    buf_clk new_AGEMA_reg_buffer_3218 ( .C (clk), .D (new_AGEMA_signal_6648), .Q (new_AGEMA_signal_6649) ) ;
    buf_clk new_AGEMA_reg_buffer_3222 ( .C (clk), .D (new_AGEMA_signal_6652), .Q (new_AGEMA_signal_6653) ) ;
    buf_clk new_AGEMA_reg_buffer_3226 ( .C (clk), .D (new_AGEMA_signal_6656), .Q (new_AGEMA_signal_6657) ) ;
    buf_clk new_AGEMA_reg_buffer_3230 ( .C (clk), .D (new_AGEMA_signal_6660), .Q (new_AGEMA_signal_6661) ) ;
    buf_clk new_AGEMA_reg_buffer_3234 ( .C (clk), .D (new_AGEMA_signal_6664), .Q (new_AGEMA_signal_6665) ) ;
    buf_clk new_AGEMA_reg_buffer_3238 ( .C (clk), .D (new_AGEMA_signal_6668), .Q (new_AGEMA_signal_6669) ) ;
    buf_clk new_AGEMA_reg_buffer_3242 ( .C (clk), .D (new_AGEMA_signal_6672), .Q (new_AGEMA_signal_6673) ) ;
    buf_clk new_AGEMA_reg_buffer_3246 ( .C (clk), .D (new_AGEMA_signal_6676), .Q (new_AGEMA_signal_6677) ) ;
    buf_clk new_AGEMA_reg_buffer_3250 ( .C (clk), .D (new_AGEMA_signal_6680), .Q (new_AGEMA_signal_6681) ) ;
    buf_clk new_AGEMA_reg_buffer_3254 ( .C (clk), .D (new_AGEMA_signal_6684), .Q (new_AGEMA_signal_6685) ) ;
    buf_clk new_AGEMA_reg_buffer_3258 ( .C (clk), .D (new_AGEMA_signal_6688), .Q (new_AGEMA_signal_6689) ) ;
    buf_clk new_AGEMA_reg_buffer_3262 ( .C (clk), .D (new_AGEMA_signal_6692), .Q (new_AGEMA_signal_6693) ) ;
    buf_clk new_AGEMA_reg_buffer_3266 ( .C (clk), .D (new_AGEMA_signal_6696), .Q (new_AGEMA_signal_6697) ) ;
    buf_clk new_AGEMA_reg_buffer_3270 ( .C (clk), .D (new_AGEMA_signal_6700), .Q (new_AGEMA_signal_6701) ) ;
    buf_clk new_AGEMA_reg_buffer_3274 ( .C (clk), .D (new_AGEMA_signal_6704), .Q (new_AGEMA_signal_6705) ) ;
    buf_clk new_AGEMA_reg_buffer_3278 ( .C (clk), .D (new_AGEMA_signal_6708), .Q (new_AGEMA_signal_6709) ) ;
    buf_clk new_AGEMA_reg_buffer_3282 ( .C (clk), .D (new_AGEMA_signal_6712), .Q (new_AGEMA_signal_6713) ) ;
    buf_clk new_AGEMA_reg_buffer_3286 ( .C (clk), .D (new_AGEMA_signal_6716), .Q (new_AGEMA_signal_6717) ) ;
    buf_clk new_AGEMA_reg_buffer_3290 ( .C (clk), .D (new_AGEMA_signal_6720), .Q (new_AGEMA_signal_6721) ) ;
    buf_clk new_AGEMA_reg_buffer_3294 ( .C (clk), .D (new_AGEMA_signal_6724), .Q (new_AGEMA_signal_6725) ) ;
    buf_clk new_AGEMA_reg_buffer_3298 ( .C (clk), .D (new_AGEMA_signal_6728), .Q (new_AGEMA_signal_6729) ) ;
    buf_clk new_AGEMA_reg_buffer_3302 ( .C (clk), .D (new_AGEMA_signal_6732), .Q (new_AGEMA_signal_6733) ) ;
    buf_clk new_AGEMA_reg_buffer_3306 ( .C (clk), .D (new_AGEMA_signal_6736), .Q (new_AGEMA_signal_6737) ) ;
    buf_clk new_AGEMA_reg_buffer_3310 ( .C (clk), .D (new_AGEMA_signal_6740), .Q (new_AGEMA_signal_6741) ) ;
    buf_clk new_AGEMA_reg_buffer_3314 ( .C (clk), .D (new_AGEMA_signal_6744), .Q (new_AGEMA_signal_6745) ) ;
    buf_clk new_AGEMA_reg_buffer_3318 ( .C (clk), .D (new_AGEMA_signal_6748), .Q (new_AGEMA_signal_6749) ) ;
    buf_clk new_AGEMA_reg_buffer_3322 ( .C (clk), .D (new_AGEMA_signal_6752), .Q (new_AGEMA_signal_6753) ) ;
    buf_clk new_AGEMA_reg_buffer_3326 ( .C (clk), .D (new_AGEMA_signal_6756), .Q (new_AGEMA_signal_6757) ) ;
    buf_clk new_AGEMA_reg_buffer_3330 ( .C (clk), .D (new_AGEMA_signal_6760), .Q (new_AGEMA_signal_6761) ) ;
    buf_clk new_AGEMA_reg_buffer_3334 ( .C (clk), .D (new_AGEMA_signal_6764), .Q (new_AGEMA_signal_6765) ) ;
    buf_clk new_AGEMA_reg_buffer_3338 ( .C (clk), .D (new_AGEMA_signal_6768), .Q (new_AGEMA_signal_6769) ) ;
    buf_clk new_AGEMA_reg_buffer_3342 ( .C (clk), .D (new_AGEMA_signal_6772), .Q (new_AGEMA_signal_6773) ) ;
    buf_clk new_AGEMA_reg_buffer_3346 ( .C (clk), .D (new_AGEMA_signal_6776), .Q (new_AGEMA_signal_6777) ) ;
    buf_clk new_AGEMA_reg_buffer_3350 ( .C (clk), .D (new_AGEMA_signal_6780), .Q (new_AGEMA_signal_6781) ) ;
    buf_clk new_AGEMA_reg_buffer_3354 ( .C (clk), .D (new_AGEMA_signal_6784), .Q (new_AGEMA_signal_6785) ) ;
    buf_clk new_AGEMA_reg_buffer_3358 ( .C (clk), .D (new_AGEMA_signal_6788), .Q (new_AGEMA_signal_6789) ) ;
    buf_clk new_AGEMA_reg_buffer_3362 ( .C (clk), .D (new_AGEMA_signal_6792), .Q (new_AGEMA_signal_6793) ) ;
    buf_clk new_AGEMA_reg_buffer_3366 ( .C (clk), .D (new_AGEMA_signal_6796), .Q (new_AGEMA_signal_6797) ) ;
    buf_clk new_AGEMA_reg_buffer_3370 ( .C (clk), .D (new_AGEMA_signal_6800), .Q (new_AGEMA_signal_6801) ) ;
    buf_clk new_AGEMA_reg_buffer_3374 ( .C (clk), .D (new_AGEMA_signal_6804), .Q (new_AGEMA_signal_6805) ) ;
    buf_clk new_AGEMA_reg_buffer_3378 ( .C (clk), .D (new_AGEMA_signal_6808), .Q (new_AGEMA_signal_6809) ) ;
    buf_clk new_AGEMA_reg_buffer_3382 ( .C (clk), .D (new_AGEMA_signal_6812), .Q (new_AGEMA_signal_6813) ) ;
    buf_clk new_AGEMA_reg_buffer_3386 ( .C (clk), .D (new_AGEMA_signal_6816), .Q (new_AGEMA_signal_6817) ) ;
    buf_clk new_AGEMA_reg_buffer_3390 ( .C (clk), .D (new_AGEMA_signal_6820), .Q (new_AGEMA_signal_6821) ) ;
    buf_clk new_AGEMA_reg_buffer_3394 ( .C (clk), .D (new_AGEMA_signal_6824), .Q (new_AGEMA_signal_6825) ) ;
    buf_clk new_AGEMA_reg_buffer_3398 ( .C (clk), .D (new_AGEMA_signal_6828), .Q (new_AGEMA_signal_6829) ) ;
    buf_clk new_AGEMA_reg_buffer_3402 ( .C (clk), .D (new_AGEMA_signal_6832), .Q (new_AGEMA_signal_6833) ) ;
    buf_clk new_AGEMA_reg_buffer_3406 ( .C (clk), .D (new_AGEMA_signal_6836), .Q (new_AGEMA_signal_6837) ) ;
    buf_clk new_AGEMA_reg_buffer_3410 ( .C (clk), .D (new_AGEMA_signal_6840), .Q (new_AGEMA_signal_6841) ) ;
    buf_clk new_AGEMA_reg_buffer_3414 ( .C (clk), .D (new_AGEMA_signal_6844), .Q (new_AGEMA_signal_6845) ) ;
    buf_clk new_AGEMA_reg_buffer_3418 ( .C (clk), .D (new_AGEMA_signal_6848), .Q (new_AGEMA_signal_6849) ) ;
    buf_clk new_AGEMA_reg_buffer_3422 ( .C (clk), .D (new_AGEMA_signal_6852), .Q (new_AGEMA_signal_6853) ) ;
    buf_clk new_AGEMA_reg_buffer_3426 ( .C (clk), .D (new_AGEMA_signal_6856), .Q (new_AGEMA_signal_6857) ) ;
    buf_clk new_AGEMA_reg_buffer_3430 ( .C (clk), .D (new_AGEMA_signal_6860), .Q (new_AGEMA_signal_6861) ) ;
    buf_clk new_AGEMA_reg_buffer_3434 ( .C (clk), .D (new_AGEMA_signal_6864), .Q (new_AGEMA_signal_6865) ) ;
    buf_clk new_AGEMA_reg_buffer_3438 ( .C (clk), .D (new_AGEMA_signal_6868), .Q (new_AGEMA_signal_6869) ) ;
    buf_clk new_AGEMA_reg_buffer_3442 ( .C (clk), .D (new_AGEMA_signal_6872), .Q (new_AGEMA_signal_6873) ) ;
    buf_clk new_AGEMA_reg_buffer_3446 ( .C (clk), .D (new_AGEMA_signal_6876), .Q (new_AGEMA_signal_6877) ) ;
    buf_clk new_AGEMA_reg_buffer_3450 ( .C (clk), .D (new_AGEMA_signal_6880), .Q (new_AGEMA_signal_6881) ) ;
    buf_clk new_AGEMA_reg_buffer_3454 ( .C (clk), .D (new_AGEMA_signal_6884), .Q (new_AGEMA_signal_6885) ) ;
    buf_clk new_AGEMA_reg_buffer_3456 ( .C (clk), .D (StateRegInput[63]), .Q (new_AGEMA_signal_6887) ) ;
    buf_clk new_AGEMA_reg_buffer_3458 ( .C (clk), .D (new_AGEMA_signal_3981), .Q (new_AGEMA_signal_6889) ) ;
    buf_clk new_AGEMA_reg_buffer_3460 ( .C (clk), .D (new_AGEMA_signal_3982), .Q (new_AGEMA_signal_6891) ) ;
    buf_clk new_AGEMA_reg_buffer_3462 ( .C (clk), .D (new_AGEMA_signal_3983), .Q (new_AGEMA_signal_6893) ) ;
    buf_clk new_AGEMA_reg_buffer_3464 ( .C (clk), .D (StateRegInput[62]), .Q (new_AGEMA_signal_6895) ) ;
    buf_clk new_AGEMA_reg_buffer_3466 ( .C (clk), .D (new_AGEMA_signal_3852), .Q (new_AGEMA_signal_6897) ) ;
    buf_clk new_AGEMA_reg_buffer_3468 ( .C (clk), .D (new_AGEMA_signal_3853), .Q (new_AGEMA_signal_6899) ) ;
    buf_clk new_AGEMA_reg_buffer_3470 ( .C (clk), .D (new_AGEMA_signal_3854), .Q (new_AGEMA_signal_6901) ) ;
    buf_clk new_AGEMA_reg_buffer_3472 ( .C (clk), .D (StateRegInput[59]), .Q (new_AGEMA_signal_6903) ) ;
    buf_clk new_AGEMA_reg_buffer_3474 ( .C (clk), .D (new_AGEMA_signal_3690), .Q (new_AGEMA_signal_6905) ) ;
    buf_clk new_AGEMA_reg_buffer_3476 ( .C (clk), .D (new_AGEMA_signal_3691), .Q (new_AGEMA_signal_6907) ) ;
    buf_clk new_AGEMA_reg_buffer_3478 ( .C (clk), .D (new_AGEMA_signal_3692), .Q (new_AGEMA_signal_6909) ) ;
    buf_clk new_AGEMA_reg_buffer_3480 ( .C (clk), .D (StateRegInput[58]), .Q (new_AGEMA_signal_6911) ) ;
    buf_clk new_AGEMA_reg_buffer_3482 ( .C (clk), .D (new_AGEMA_signal_3510), .Q (new_AGEMA_signal_6913) ) ;
    buf_clk new_AGEMA_reg_buffer_3484 ( .C (clk), .D (new_AGEMA_signal_3511), .Q (new_AGEMA_signal_6915) ) ;
    buf_clk new_AGEMA_reg_buffer_3486 ( .C (clk), .D (new_AGEMA_signal_3512), .Q (new_AGEMA_signal_6917) ) ;
    buf_clk new_AGEMA_reg_buffer_3488 ( .C (clk), .D (StateRegInput[55]), .Q (new_AGEMA_signal_6919) ) ;
    buf_clk new_AGEMA_reg_buffer_3490 ( .C (clk), .D (new_AGEMA_signal_3684), .Q (new_AGEMA_signal_6921) ) ;
    buf_clk new_AGEMA_reg_buffer_3492 ( .C (clk), .D (new_AGEMA_signal_3685), .Q (new_AGEMA_signal_6923) ) ;
    buf_clk new_AGEMA_reg_buffer_3494 ( .C (clk), .D (new_AGEMA_signal_3686), .Q (new_AGEMA_signal_6925) ) ;
    buf_clk new_AGEMA_reg_buffer_3496 ( .C (clk), .D (StateRegInput[54]), .Q (new_AGEMA_signal_6927) ) ;
    buf_clk new_AGEMA_reg_buffer_3498 ( .C (clk), .D (new_AGEMA_signal_3504), .Q (new_AGEMA_signal_6929) ) ;
    buf_clk new_AGEMA_reg_buffer_3500 ( .C (clk), .D (new_AGEMA_signal_3505), .Q (new_AGEMA_signal_6931) ) ;
    buf_clk new_AGEMA_reg_buffer_3502 ( .C (clk), .D (new_AGEMA_signal_3506), .Q (new_AGEMA_signal_6933) ) ;
    buf_clk new_AGEMA_reg_buffer_3504 ( .C (clk), .D (StateRegInput[51]), .Q (new_AGEMA_signal_6935) ) ;
    buf_clk new_AGEMA_reg_buffer_3506 ( .C (clk), .D (new_AGEMA_signal_3678), .Q (new_AGEMA_signal_6937) ) ;
    buf_clk new_AGEMA_reg_buffer_3508 ( .C (clk), .D (new_AGEMA_signal_3679), .Q (new_AGEMA_signal_6939) ) ;
    buf_clk new_AGEMA_reg_buffer_3510 ( .C (clk), .D (new_AGEMA_signal_3680), .Q (new_AGEMA_signal_6941) ) ;
    buf_clk new_AGEMA_reg_buffer_3512 ( .C (clk), .D (StateRegInput[50]), .Q (new_AGEMA_signal_6943) ) ;
    buf_clk new_AGEMA_reg_buffer_3514 ( .C (clk), .D (new_AGEMA_signal_3498), .Q (new_AGEMA_signal_6945) ) ;
    buf_clk new_AGEMA_reg_buffer_3516 ( .C (clk), .D (new_AGEMA_signal_3499), .Q (new_AGEMA_signal_6947) ) ;
    buf_clk new_AGEMA_reg_buffer_3518 ( .C (clk), .D (new_AGEMA_signal_3500), .Q (new_AGEMA_signal_6949) ) ;
    buf_clk new_AGEMA_reg_buffer_3520 ( .C (clk), .D (StateRegInput[47]), .Q (new_AGEMA_signal_6951) ) ;
    buf_clk new_AGEMA_reg_buffer_3522 ( .C (clk), .D (new_AGEMA_signal_3672), .Q (new_AGEMA_signal_6953) ) ;
    buf_clk new_AGEMA_reg_buffer_3524 ( .C (clk), .D (new_AGEMA_signal_3673), .Q (new_AGEMA_signal_6955) ) ;
    buf_clk new_AGEMA_reg_buffer_3526 ( .C (clk), .D (new_AGEMA_signal_3674), .Q (new_AGEMA_signal_6957) ) ;
    buf_clk new_AGEMA_reg_buffer_3528 ( .C (clk), .D (StateRegInput[46]), .Q (new_AGEMA_signal_6959) ) ;
    buf_clk new_AGEMA_reg_buffer_3530 ( .C (clk), .D (new_AGEMA_signal_3492), .Q (new_AGEMA_signal_6961) ) ;
    buf_clk new_AGEMA_reg_buffer_3532 ( .C (clk), .D (new_AGEMA_signal_3493), .Q (new_AGEMA_signal_6963) ) ;
    buf_clk new_AGEMA_reg_buffer_3534 ( .C (clk), .D (new_AGEMA_signal_3494), .Q (new_AGEMA_signal_6965) ) ;
    buf_clk new_AGEMA_reg_buffer_3536 ( .C (clk), .D (StateRegInput[43]), .Q (new_AGEMA_signal_6967) ) ;
    buf_clk new_AGEMA_reg_buffer_3538 ( .C (clk), .D (new_AGEMA_signal_3306), .Q (new_AGEMA_signal_6969) ) ;
    buf_clk new_AGEMA_reg_buffer_3540 ( .C (clk), .D (new_AGEMA_signal_3307), .Q (new_AGEMA_signal_6971) ) ;
    buf_clk new_AGEMA_reg_buffer_3542 ( .C (clk), .D (new_AGEMA_signal_3308), .Q (new_AGEMA_signal_6973) ) ;
    buf_clk new_AGEMA_reg_buffer_3544 ( .C (clk), .D (StateRegInput[42]), .Q (new_AGEMA_signal_6975) ) ;
    buf_clk new_AGEMA_reg_buffer_3546 ( .C (clk), .D (new_AGEMA_signal_3147), .Q (new_AGEMA_signal_6977) ) ;
    buf_clk new_AGEMA_reg_buffer_3548 ( .C (clk), .D (new_AGEMA_signal_3148), .Q (new_AGEMA_signal_6979) ) ;
    buf_clk new_AGEMA_reg_buffer_3550 ( .C (clk), .D (new_AGEMA_signal_3149), .Q (new_AGEMA_signal_6981) ) ;
    buf_clk new_AGEMA_reg_buffer_3552 ( .C (clk), .D (StateRegInput[39]), .Q (new_AGEMA_signal_6983) ) ;
    buf_clk new_AGEMA_reg_buffer_3554 ( .C (clk), .D (new_AGEMA_signal_3300), .Q (new_AGEMA_signal_6985) ) ;
    buf_clk new_AGEMA_reg_buffer_3556 ( .C (clk), .D (new_AGEMA_signal_3301), .Q (new_AGEMA_signal_6987) ) ;
    buf_clk new_AGEMA_reg_buffer_3558 ( .C (clk), .D (new_AGEMA_signal_3302), .Q (new_AGEMA_signal_6989) ) ;
    buf_clk new_AGEMA_reg_buffer_3560 ( .C (clk), .D (StateRegInput[38]), .Q (new_AGEMA_signal_6991) ) ;
    buf_clk new_AGEMA_reg_buffer_3562 ( .C (clk), .D (new_AGEMA_signal_3141), .Q (new_AGEMA_signal_6993) ) ;
    buf_clk new_AGEMA_reg_buffer_3564 ( .C (clk), .D (new_AGEMA_signal_3142), .Q (new_AGEMA_signal_6995) ) ;
    buf_clk new_AGEMA_reg_buffer_3566 ( .C (clk), .D (new_AGEMA_signal_3143), .Q (new_AGEMA_signal_6997) ) ;
    buf_clk new_AGEMA_reg_buffer_3568 ( .C (clk), .D (StateRegInput[35]), .Q (new_AGEMA_signal_6999) ) ;
    buf_clk new_AGEMA_reg_buffer_3570 ( .C (clk), .D (new_AGEMA_signal_3294), .Q (new_AGEMA_signal_7001) ) ;
    buf_clk new_AGEMA_reg_buffer_3572 ( .C (clk), .D (new_AGEMA_signal_3295), .Q (new_AGEMA_signal_7003) ) ;
    buf_clk new_AGEMA_reg_buffer_3574 ( .C (clk), .D (new_AGEMA_signal_3296), .Q (new_AGEMA_signal_7005) ) ;
    buf_clk new_AGEMA_reg_buffer_3576 ( .C (clk), .D (StateRegInput[34]), .Q (new_AGEMA_signal_7007) ) ;
    buf_clk new_AGEMA_reg_buffer_3578 ( .C (clk), .D (new_AGEMA_signal_3135), .Q (new_AGEMA_signal_7009) ) ;
    buf_clk new_AGEMA_reg_buffer_3580 ( .C (clk), .D (new_AGEMA_signal_3136), .Q (new_AGEMA_signal_7011) ) ;
    buf_clk new_AGEMA_reg_buffer_3582 ( .C (clk), .D (new_AGEMA_signal_3137), .Q (new_AGEMA_signal_7013) ) ;
    buf_clk new_AGEMA_reg_buffer_3584 ( .C (clk), .D (StateRegInput[31]), .Q (new_AGEMA_signal_7015) ) ;
    buf_clk new_AGEMA_reg_buffer_3586 ( .C (clk), .D (new_AGEMA_signal_3648), .Q (new_AGEMA_signal_7017) ) ;
    buf_clk new_AGEMA_reg_buffer_3588 ( .C (clk), .D (new_AGEMA_signal_3649), .Q (new_AGEMA_signal_7019) ) ;
    buf_clk new_AGEMA_reg_buffer_3590 ( .C (clk), .D (new_AGEMA_signal_3650), .Q (new_AGEMA_signal_7021) ) ;
    buf_clk new_AGEMA_reg_buffer_3592 ( .C (clk), .D (StateRegInput[30]), .Q (new_AGEMA_signal_7023) ) ;
    buf_clk new_AGEMA_reg_buffer_3594 ( .C (clk), .D (new_AGEMA_signal_3468), .Q (new_AGEMA_signal_7025) ) ;
    buf_clk new_AGEMA_reg_buffer_3596 ( .C (clk), .D (new_AGEMA_signal_3469), .Q (new_AGEMA_signal_7027) ) ;
    buf_clk new_AGEMA_reg_buffer_3598 ( .C (clk), .D (new_AGEMA_signal_3470), .Q (new_AGEMA_signal_7029) ) ;
    buf_clk new_AGEMA_reg_buffer_3600 ( .C (clk), .D (StateRegInput[27]), .Q (new_AGEMA_signal_7031) ) ;
    buf_clk new_AGEMA_reg_buffer_3602 ( .C (clk), .D (new_AGEMA_signal_3945), .Q (new_AGEMA_signal_7033) ) ;
    buf_clk new_AGEMA_reg_buffer_3604 ( .C (clk), .D (new_AGEMA_signal_3946), .Q (new_AGEMA_signal_7035) ) ;
    buf_clk new_AGEMA_reg_buffer_3606 ( .C (clk), .D (new_AGEMA_signal_3947), .Q (new_AGEMA_signal_7037) ) ;
    buf_clk new_AGEMA_reg_buffer_3608 ( .C (clk), .D (StateRegInput[26]), .Q (new_AGEMA_signal_7039) ) ;
    buf_clk new_AGEMA_reg_buffer_3610 ( .C (clk), .D (new_AGEMA_signal_3816), .Q (new_AGEMA_signal_7041) ) ;
    buf_clk new_AGEMA_reg_buffer_3612 ( .C (clk), .D (new_AGEMA_signal_3817), .Q (new_AGEMA_signal_7043) ) ;
    buf_clk new_AGEMA_reg_buffer_3614 ( .C (clk), .D (new_AGEMA_signal_3818), .Q (new_AGEMA_signal_7045) ) ;
    buf_clk new_AGEMA_reg_buffer_3616 ( .C (clk), .D (StateRegInput[23]), .Q (new_AGEMA_signal_7047) ) ;
    buf_clk new_AGEMA_reg_buffer_3618 ( .C (clk), .D (new_AGEMA_signal_3642), .Q (new_AGEMA_signal_7049) ) ;
    buf_clk new_AGEMA_reg_buffer_3620 ( .C (clk), .D (new_AGEMA_signal_3643), .Q (new_AGEMA_signal_7051) ) ;
    buf_clk new_AGEMA_reg_buffer_3622 ( .C (clk), .D (new_AGEMA_signal_3644), .Q (new_AGEMA_signal_7053) ) ;
    buf_clk new_AGEMA_reg_buffer_3624 ( .C (clk), .D (StateRegInput[22]), .Q (new_AGEMA_signal_7055) ) ;
    buf_clk new_AGEMA_reg_buffer_3626 ( .C (clk), .D (new_AGEMA_signal_3462), .Q (new_AGEMA_signal_7057) ) ;
    buf_clk new_AGEMA_reg_buffer_3628 ( .C (clk), .D (new_AGEMA_signal_3463), .Q (new_AGEMA_signal_7059) ) ;
    buf_clk new_AGEMA_reg_buffer_3630 ( .C (clk), .D (new_AGEMA_signal_3464), .Q (new_AGEMA_signal_7061) ) ;
    buf_clk new_AGEMA_reg_buffer_3632 ( .C (clk), .D (StateRegInput[19]), .Q (new_AGEMA_signal_7063) ) ;
    buf_clk new_AGEMA_reg_buffer_3634 ( .C (clk), .D (new_AGEMA_signal_3636), .Q (new_AGEMA_signal_7065) ) ;
    buf_clk new_AGEMA_reg_buffer_3636 ( .C (clk), .D (new_AGEMA_signal_3637), .Q (new_AGEMA_signal_7067) ) ;
    buf_clk new_AGEMA_reg_buffer_3638 ( .C (clk), .D (new_AGEMA_signal_3638), .Q (new_AGEMA_signal_7069) ) ;
    buf_clk new_AGEMA_reg_buffer_3640 ( .C (clk), .D (StateRegInput[18]), .Q (new_AGEMA_signal_7071) ) ;
    buf_clk new_AGEMA_reg_buffer_3642 ( .C (clk), .D (new_AGEMA_signal_3456), .Q (new_AGEMA_signal_7073) ) ;
    buf_clk new_AGEMA_reg_buffer_3644 ( .C (clk), .D (new_AGEMA_signal_3457), .Q (new_AGEMA_signal_7075) ) ;
    buf_clk new_AGEMA_reg_buffer_3646 ( .C (clk), .D (new_AGEMA_signal_3458), .Q (new_AGEMA_signal_7077) ) ;
    buf_clk new_AGEMA_reg_buffer_3648 ( .C (clk), .D (StateRegInput[15]), .Q (new_AGEMA_signal_7079) ) ;
    buf_clk new_AGEMA_reg_buffer_3650 ( .C (clk), .D (new_AGEMA_signal_3927), .Q (new_AGEMA_signal_7081) ) ;
    buf_clk new_AGEMA_reg_buffer_3652 ( .C (clk), .D (new_AGEMA_signal_3928), .Q (new_AGEMA_signal_7083) ) ;
    buf_clk new_AGEMA_reg_buffer_3654 ( .C (clk), .D (new_AGEMA_signal_3929), .Q (new_AGEMA_signal_7085) ) ;
    buf_clk new_AGEMA_reg_buffer_3656 ( .C (clk), .D (StateRegInput[14]), .Q (new_AGEMA_signal_7087) ) ;
    buf_clk new_AGEMA_reg_buffer_3658 ( .C (clk), .D (new_AGEMA_signal_3798), .Q (new_AGEMA_signal_7089) ) ;
    buf_clk new_AGEMA_reg_buffer_3660 ( .C (clk), .D (new_AGEMA_signal_3799), .Q (new_AGEMA_signal_7091) ) ;
    buf_clk new_AGEMA_reg_buffer_3662 ( .C (clk), .D (new_AGEMA_signal_3800), .Q (new_AGEMA_signal_7093) ) ;
    buf_clk new_AGEMA_reg_buffer_3664 ( .C (clk), .D (StateRegInput[11]), .Q (new_AGEMA_signal_7095) ) ;
    buf_clk new_AGEMA_reg_buffer_3666 ( .C (clk), .D (new_AGEMA_signal_3630), .Q (new_AGEMA_signal_7097) ) ;
    buf_clk new_AGEMA_reg_buffer_3668 ( .C (clk), .D (new_AGEMA_signal_3631), .Q (new_AGEMA_signal_7099) ) ;
    buf_clk new_AGEMA_reg_buffer_3670 ( .C (clk), .D (new_AGEMA_signal_3632), .Q (new_AGEMA_signal_7101) ) ;
    buf_clk new_AGEMA_reg_buffer_3672 ( .C (clk), .D (StateRegInput[10]), .Q (new_AGEMA_signal_7103) ) ;
    buf_clk new_AGEMA_reg_buffer_3674 ( .C (clk), .D (new_AGEMA_signal_3450), .Q (new_AGEMA_signal_7105) ) ;
    buf_clk new_AGEMA_reg_buffer_3676 ( .C (clk), .D (new_AGEMA_signal_3451), .Q (new_AGEMA_signal_7107) ) ;
    buf_clk new_AGEMA_reg_buffer_3678 ( .C (clk), .D (new_AGEMA_signal_3452), .Q (new_AGEMA_signal_7109) ) ;
    buf_clk new_AGEMA_reg_buffer_3680 ( .C (clk), .D (StateRegInput[7]), .Q (new_AGEMA_signal_7111) ) ;
    buf_clk new_AGEMA_reg_buffer_3682 ( .C (clk), .D (new_AGEMA_signal_3624), .Q (new_AGEMA_signal_7113) ) ;
    buf_clk new_AGEMA_reg_buffer_3684 ( .C (clk), .D (new_AGEMA_signal_3625), .Q (new_AGEMA_signal_7115) ) ;
    buf_clk new_AGEMA_reg_buffer_3686 ( .C (clk), .D (new_AGEMA_signal_3626), .Q (new_AGEMA_signal_7117) ) ;
    buf_clk new_AGEMA_reg_buffer_3688 ( .C (clk), .D (StateRegInput[6]), .Q (new_AGEMA_signal_7119) ) ;
    buf_clk new_AGEMA_reg_buffer_3690 ( .C (clk), .D (new_AGEMA_signal_3444), .Q (new_AGEMA_signal_7121) ) ;
    buf_clk new_AGEMA_reg_buffer_3692 ( .C (clk), .D (new_AGEMA_signal_3445), .Q (new_AGEMA_signal_7123) ) ;
    buf_clk new_AGEMA_reg_buffer_3694 ( .C (clk), .D (new_AGEMA_signal_3446), .Q (new_AGEMA_signal_7125) ) ;
    buf_clk new_AGEMA_reg_buffer_3696 ( .C (clk), .D (StateRegInput[3]), .Q (new_AGEMA_signal_7127) ) ;
    buf_clk new_AGEMA_reg_buffer_3698 ( .C (clk), .D (new_AGEMA_signal_3618), .Q (new_AGEMA_signal_7129) ) ;
    buf_clk new_AGEMA_reg_buffer_3700 ( .C (clk), .D (new_AGEMA_signal_3619), .Q (new_AGEMA_signal_7131) ) ;
    buf_clk new_AGEMA_reg_buffer_3702 ( .C (clk), .D (new_AGEMA_signal_3620), .Q (new_AGEMA_signal_7133) ) ;
    buf_clk new_AGEMA_reg_buffer_3704 ( .C (clk), .D (StateRegInput[2]), .Q (new_AGEMA_signal_7135) ) ;
    buf_clk new_AGEMA_reg_buffer_3706 ( .C (clk), .D (new_AGEMA_signal_3438), .Q (new_AGEMA_signal_7137) ) ;
    buf_clk new_AGEMA_reg_buffer_3708 ( .C (clk), .D (new_AGEMA_signal_3439), .Q (new_AGEMA_signal_7139) ) ;
    buf_clk new_AGEMA_reg_buffer_3710 ( .C (clk), .D (new_AGEMA_signal_3440), .Q (new_AGEMA_signal_7141) ) ;
    buf_clk new_AGEMA_reg_buffer_3714 ( .C (clk), .D (new_AGEMA_signal_7144), .Q (new_AGEMA_signal_7145) ) ;
    buf_clk new_AGEMA_reg_buffer_3718 ( .C (clk), .D (new_AGEMA_signal_7148), .Q (new_AGEMA_signal_7149) ) ;
    buf_clk new_AGEMA_reg_buffer_3722 ( .C (clk), .D (new_AGEMA_signal_7152), .Q (new_AGEMA_signal_7153) ) ;
    buf_clk new_AGEMA_reg_buffer_3726 ( .C (clk), .D (new_AGEMA_signal_7156), .Q (new_AGEMA_signal_7157) ) ;
    buf_clk new_AGEMA_reg_buffer_3730 ( .C (clk), .D (new_AGEMA_signal_7160), .Q (new_AGEMA_signal_7161) ) ;
    buf_clk new_AGEMA_reg_buffer_3734 ( .C (clk), .D (new_AGEMA_signal_7164), .Q (new_AGEMA_signal_7165) ) ;
    buf_clk new_AGEMA_reg_buffer_3738 ( .C (clk), .D (new_AGEMA_signal_7168), .Q (new_AGEMA_signal_7169) ) ;
    buf_clk new_AGEMA_reg_buffer_3742 ( .C (clk), .D (new_AGEMA_signal_7172), .Q (new_AGEMA_signal_7173) ) ;
    buf_clk new_AGEMA_reg_buffer_3746 ( .C (clk), .D (new_AGEMA_signal_7176), .Q (new_AGEMA_signal_7177) ) ;
    buf_clk new_AGEMA_reg_buffer_3750 ( .C (clk), .D (new_AGEMA_signal_7180), .Q (new_AGEMA_signal_7181) ) ;
    buf_clk new_AGEMA_reg_buffer_3754 ( .C (clk), .D (new_AGEMA_signal_7184), .Q (new_AGEMA_signal_7185) ) ;
    buf_clk new_AGEMA_reg_buffer_3758 ( .C (clk), .D (new_AGEMA_signal_7188), .Q (new_AGEMA_signal_7189) ) ;
    buf_clk new_AGEMA_reg_buffer_3762 ( .C (clk), .D (new_AGEMA_signal_7192), .Q (new_AGEMA_signal_7193) ) ;
    buf_clk new_AGEMA_reg_buffer_3766 ( .C (clk), .D (new_AGEMA_signal_7196), .Q (new_AGEMA_signal_7197) ) ;
    buf_clk new_AGEMA_reg_buffer_3770 ( .C (clk), .D (new_AGEMA_signal_7200), .Q (new_AGEMA_signal_7201) ) ;
    buf_clk new_AGEMA_reg_buffer_3774 ( .C (clk), .D (new_AGEMA_signal_7204), .Q (new_AGEMA_signal_7205) ) ;
    buf_clk new_AGEMA_reg_buffer_3778 ( .C (clk), .D (new_AGEMA_signal_7208), .Q (new_AGEMA_signal_7209) ) ;
    buf_clk new_AGEMA_reg_buffer_3782 ( .C (clk), .D (new_AGEMA_signal_7212), .Q (new_AGEMA_signal_7213) ) ;
    buf_clk new_AGEMA_reg_buffer_3786 ( .C (clk), .D (new_AGEMA_signal_7216), .Q (new_AGEMA_signal_7217) ) ;
    buf_clk new_AGEMA_reg_buffer_3790 ( .C (clk), .D (new_AGEMA_signal_7220), .Q (new_AGEMA_signal_7221) ) ;
    buf_clk new_AGEMA_reg_buffer_3794 ( .C (clk), .D (new_AGEMA_signal_7224), .Q (new_AGEMA_signal_7225) ) ;
    buf_clk new_AGEMA_reg_buffer_3798 ( .C (clk), .D (new_AGEMA_signal_7228), .Q (new_AGEMA_signal_7229) ) ;
    buf_clk new_AGEMA_reg_buffer_3802 ( .C (clk), .D (new_AGEMA_signal_7232), .Q (new_AGEMA_signal_7233) ) ;
    buf_clk new_AGEMA_reg_buffer_3806 ( .C (clk), .D (new_AGEMA_signal_7236), .Q (new_AGEMA_signal_7237) ) ;
    buf_clk new_AGEMA_reg_buffer_3810 ( .C (clk), .D (new_AGEMA_signal_7240), .Q (new_AGEMA_signal_7241) ) ;
    buf_clk new_AGEMA_reg_buffer_3814 ( .C (clk), .D (new_AGEMA_signal_7244), .Q (new_AGEMA_signal_7245) ) ;
    buf_clk new_AGEMA_reg_buffer_3818 ( .C (clk), .D (new_AGEMA_signal_7248), .Q (new_AGEMA_signal_7249) ) ;
    buf_clk new_AGEMA_reg_buffer_3822 ( .C (clk), .D (new_AGEMA_signal_7252), .Q (new_AGEMA_signal_7253) ) ;
    buf_clk new_AGEMA_reg_buffer_3826 ( .C (clk), .D (new_AGEMA_signal_7256), .Q (new_AGEMA_signal_7257) ) ;
    buf_clk new_AGEMA_reg_buffer_3830 ( .C (clk), .D (new_AGEMA_signal_7260), .Q (new_AGEMA_signal_7261) ) ;
    buf_clk new_AGEMA_reg_buffer_3834 ( .C (clk), .D (new_AGEMA_signal_7264), .Q (new_AGEMA_signal_7265) ) ;
    buf_clk new_AGEMA_reg_buffer_3838 ( .C (clk), .D (new_AGEMA_signal_7268), .Q (new_AGEMA_signal_7269) ) ;
    buf_clk new_AGEMA_reg_buffer_3842 ( .C (clk), .D (new_AGEMA_signal_7272), .Q (new_AGEMA_signal_7273) ) ;
    buf_clk new_AGEMA_reg_buffer_3846 ( .C (clk), .D (new_AGEMA_signal_7276), .Q (new_AGEMA_signal_7277) ) ;
    buf_clk new_AGEMA_reg_buffer_3850 ( .C (clk), .D (new_AGEMA_signal_7280), .Q (new_AGEMA_signal_7281) ) ;
    buf_clk new_AGEMA_reg_buffer_3854 ( .C (clk), .D (new_AGEMA_signal_7284), .Q (new_AGEMA_signal_7285) ) ;
    buf_clk new_AGEMA_reg_buffer_3858 ( .C (clk), .D (new_AGEMA_signal_7288), .Q (new_AGEMA_signal_7289) ) ;
    buf_clk new_AGEMA_reg_buffer_3862 ( .C (clk), .D (new_AGEMA_signal_7292), .Q (new_AGEMA_signal_7293) ) ;
    buf_clk new_AGEMA_reg_buffer_3866 ( .C (clk), .D (new_AGEMA_signal_7296), .Q (new_AGEMA_signal_7297) ) ;
    buf_clk new_AGEMA_reg_buffer_3870 ( .C (clk), .D (new_AGEMA_signal_7300), .Q (new_AGEMA_signal_7301) ) ;
    buf_clk new_AGEMA_reg_buffer_3874 ( .C (clk), .D (new_AGEMA_signal_7304), .Q (new_AGEMA_signal_7305) ) ;
    buf_clk new_AGEMA_reg_buffer_3878 ( .C (clk), .D (new_AGEMA_signal_7308), .Q (new_AGEMA_signal_7309) ) ;
    buf_clk new_AGEMA_reg_buffer_3882 ( .C (clk), .D (new_AGEMA_signal_7312), .Q (new_AGEMA_signal_7313) ) ;
    buf_clk new_AGEMA_reg_buffer_3886 ( .C (clk), .D (new_AGEMA_signal_7316), .Q (new_AGEMA_signal_7317) ) ;
    buf_clk new_AGEMA_reg_buffer_3890 ( .C (clk), .D (new_AGEMA_signal_7320), .Q (new_AGEMA_signal_7321) ) ;
    buf_clk new_AGEMA_reg_buffer_3894 ( .C (clk), .D (new_AGEMA_signal_7324), .Q (new_AGEMA_signal_7325) ) ;
    buf_clk new_AGEMA_reg_buffer_3898 ( .C (clk), .D (new_AGEMA_signal_7328), .Q (new_AGEMA_signal_7329) ) ;
    buf_clk new_AGEMA_reg_buffer_3902 ( .C (clk), .D (new_AGEMA_signal_7332), .Q (new_AGEMA_signal_7333) ) ;
    buf_clk new_AGEMA_reg_buffer_3906 ( .C (clk), .D (new_AGEMA_signal_7336), .Q (new_AGEMA_signal_7337) ) ;
    buf_clk new_AGEMA_reg_buffer_3910 ( .C (clk), .D (new_AGEMA_signal_7340), .Q (new_AGEMA_signal_7341) ) ;
    buf_clk new_AGEMA_reg_buffer_3914 ( .C (clk), .D (new_AGEMA_signal_7344), .Q (new_AGEMA_signal_7345) ) ;
    buf_clk new_AGEMA_reg_buffer_3918 ( .C (clk), .D (new_AGEMA_signal_7348), .Q (new_AGEMA_signal_7349) ) ;
    buf_clk new_AGEMA_reg_buffer_3922 ( .C (clk), .D (new_AGEMA_signal_7352), .Q (new_AGEMA_signal_7353) ) ;
    buf_clk new_AGEMA_reg_buffer_3926 ( .C (clk), .D (new_AGEMA_signal_7356), .Q (new_AGEMA_signal_7357) ) ;
    buf_clk new_AGEMA_reg_buffer_3930 ( .C (clk), .D (new_AGEMA_signal_7360), .Q (new_AGEMA_signal_7361) ) ;
    buf_clk new_AGEMA_reg_buffer_3934 ( .C (clk), .D (new_AGEMA_signal_7364), .Q (new_AGEMA_signal_7365) ) ;
    buf_clk new_AGEMA_reg_buffer_3938 ( .C (clk), .D (new_AGEMA_signal_7368), .Q (new_AGEMA_signal_7369) ) ;
    buf_clk new_AGEMA_reg_buffer_3942 ( .C (clk), .D (new_AGEMA_signal_7372), .Q (new_AGEMA_signal_7373) ) ;
    buf_clk new_AGEMA_reg_buffer_3946 ( .C (clk), .D (new_AGEMA_signal_7376), .Q (new_AGEMA_signal_7377) ) ;
    buf_clk new_AGEMA_reg_buffer_3950 ( .C (clk), .D (new_AGEMA_signal_7380), .Q (new_AGEMA_signal_7381) ) ;
    buf_clk new_AGEMA_reg_buffer_3954 ( .C (clk), .D (new_AGEMA_signal_7384), .Q (new_AGEMA_signal_7385) ) ;
    buf_clk new_AGEMA_reg_buffer_3958 ( .C (clk), .D (new_AGEMA_signal_7388), .Q (new_AGEMA_signal_7389) ) ;
    buf_clk new_AGEMA_reg_buffer_3962 ( .C (clk), .D (new_AGEMA_signal_7392), .Q (new_AGEMA_signal_7393) ) ;
    buf_clk new_AGEMA_reg_buffer_3966 ( .C (clk), .D (new_AGEMA_signal_7396), .Q (new_AGEMA_signal_7397) ) ;
    buf_clk new_AGEMA_reg_buffer_3970 ( .C (clk), .D (new_AGEMA_signal_7400), .Q (new_AGEMA_signal_7401) ) ;
    buf_clk new_AGEMA_reg_buffer_3974 ( .C (clk), .D (new_AGEMA_signal_7404), .Q (new_AGEMA_signal_7405) ) ;
    buf_clk new_AGEMA_reg_buffer_3978 ( .C (clk), .D (new_AGEMA_signal_7408), .Q (new_AGEMA_signal_7409) ) ;
    buf_clk new_AGEMA_reg_buffer_3982 ( .C (clk), .D (new_AGEMA_signal_7412), .Q (new_AGEMA_signal_7413) ) ;
    buf_clk new_AGEMA_reg_buffer_3986 ( .C (clk), .D (new_AGEMA_signal_7416), .Q (new_AGEMA_signal_7417) ) ;
    buf_clk new_AGEMA_reg_buffer_3990 ( .C (clk), .D (new_AGEMA_signal_7420), .Q (new_AGEMA_signal_7421) ) ;
    buf_clk new_AGEMA_reg_buffer_3994 ( .C (clk), .D (new_AGEMA_signal_7424), .Q (new_AGEMA_signal_7425) ) ;
    buf_clk new_AGEMA_reg_buffer_3998 ( .C (clk), .D (new_AGEMA_signal_7428), .Q (new_AGEMA_signal_7429) ) ;
    buf_clk new_AGEMA_reg_buffer_4002 ( .C (clk), .D (new_AGEMA_signal_7432), .Q (new_AGEMA_signal_7433) ) ;
    buf_clk new_AGEMA_reg_buffer_4006 ( .C (clk), .D (new_AGEMA_signal_7436), .Q (new_AGEMA_signal_7437) ) ;
    buf_clk new_AGEMA_reg_buffer_4010 ( .C (clk), .D (new_AGEMA_signal_7440), .Q (new_AGEMA_signal_7441) ) ;
    buf_clk new_AGEMA_reg_buffer_4014 ( .C (clk), .D (new_AGEMA_signal_7444), .Q (new_AGEMA_signal_7445) ) ;
    buf_clk new_AGEMA_reg_buffer_4018 ( .C (clk), .D (new_AGEMA_signal_7448), .Q (new_AGEMA_signal_7449) ) ;
    buf_clk new_AGEMA_reg_buffer_4022 ( .C (clk), .D (new_AGEMA_signal_7452), .Q (new_AGEMA_signal_7453) ) ;
    buf_clk new_AGEMA_reg_buffer_4026 ( .C (clk), .D (new_AGEMA_signal_7456), .Q (new_AGEMA_signal_7457) ) ;
    buf_clk new_AGEMA_reg_buffer_4030 ( .C (clk), .D (new_AGEMA_signal_7460), .Q (new_AGEMA_signal_7461) ) ;
    buf_clk new_AGEMA_reg_buffer_4034 ( .C (clk), .D (new_AGEMA_signal_7464), .Q (new_AGEMA_signal_7465) ) ;
    buf_clk new_AGEMA_reg_buffer_4038 ( .C (clk), .D (new_AGEMA_signal_7468), .Q (new_AGEMA_signal_7469) ) ;
    buf_clk new_AGEMA_reg_buffer_4042 ( .C (clk), .D (new_AGEMA_signal_7472), .Q (new_AGEMA_signal_7473) ) ;
    buf_clk new_AGEMA_reg_buffer_4046 ( .C (clk), .D (new_AGEMA_signal_7476), .Q (new_AGEMA_signal_7477) ) ;
    buf_clk new_AGEMA_reg_buffer_4050 ( .C (clk), .D (new_AGEMA_signal_7480), .Q (new_AGEMA_signal_7481) ) ;
    buf_clk new_AGEMA_reg_buffer_4054 ( .C (clk), .D (new_AGEMA_signal_7484), .Q (new_AGEMA_signal_7485) ) ;
    buf_clk new_AGEMA_reg_buffer_4058 ( .C (clk), .D (new_AGEMA_signal_7488), .Q (new_AGEMA_signal_7489) ) ;
    buf_clk new_AGEMA_reg_buffer_4062 ( .C (clk), .D (new_AGEMA_signal_7492), .Q (new_AGEMA_signal_7493) ) ;
    buf_clk new_AGEMA_reg_buffer_4066 ( .C (clk), .D (new_AGEMA_signal_7496), .Q (new_AGEMA_signal_7497) ) ;
    buf_clk new_AGEMA_reg_buffer_4070 ( .C (clk), .D (new_AGEMA_signal_7500), .Q (new_AGEMA_signal_7501) ) ;
    buf_clk new_AGEMA_reg_buffer_4074 ( .C (clk), .D (new_AGEMA_signal_7504), .Q (new_AGEMA_signal_7505) ) ;
    buf_clk new_AGEMA_reg_buffer_4078 ( .C (clk), .D (new_AGEMA_signal_7508), .Q (new_AGEMA_signal_7509) ) ;
    buf_clk new_AGEMA_reg_buffer_4082 ( .C (clk), .D (new_AGEMA_signal_7512), .Q (new_AGEMA_signal_7513) ) ;
    buf_clk new_AGEMA_reg_buffer_4086 ( .C (clk), .D (new_AGEMA_signal_7516), .Q (new_AGEMA_signal_7517) ) ;
    buf_clk new_AGEMA_reg_buffer_4090 ( .C (clk), .D (new_AGEMA_signal_7520), .Q (new_AGEMA_signal_7521) ) ;
    buf_clk new_AGEMA_reg_buffer_4094 ( .C (clk), .D (new_AGEMA_signal_7524), .Q (new_AGEMA_signal_7525) ) ;
    buf_clk new_AGEMA_reg_buffer_4098 ( .C (clk), .D (new_AGEMA_signal_7528), .Q (new_AGEMA_signal_7529) ) ;
    buf_clk new_AGEMA_reg_buffer_4102 ( .C (clk), .D (new_AGEMA_signal_7532), .Q (new_AGEMA_signal_7533) ) ;
    buf_clk new_AGEMA_reg_buffer_4106 ( .C (clk), .D (new_AGEMA_signal_7536), .Q (new_AGEMA_signal_7537) ) ;
    buf_clk new_AGEMA_reg_buffer_4110 ( .C (clk), .D (new_AGEMA_signal_7540), .Q (new_AGEMA_signal_7541) ) ;
    buf_clk new_AGEMA_reg_buffer_4114 ( .C (clk), .D (new_AGEMA_signal_7544), .Q (new_AGEMA_signal_7545) ) ;
    buf_clk new_AGEMA_reg_buffer_4118 ( .C (clk), .D (new_AGEMA_signal_7548), .Q (new_AGEMA_signal_7549) ) ;
    buf_clk new_AGEMA_reg_buffer_4122 ( .C (clk), .D (new_AGEMA_signal_7552), .Q (new_AGEMA_signal_7553) ) ;
    buf_clk new_AGEMA_reg_buffer_4126 ( .C (clk), .D (new_AGEMA_signal_7556), .Q (new_AGEMA_signal_7557) ) ;
    buf_clk new_AGEMA_reg_buffer_4130 ( .C (clk), .D (new_AGEMA_signal_7560), .Q (new_AGEMA_signal_7561) ) ;
    buf_clk new_AGEMA_reg_buffer_4134 ( .C (clk), .D (new_AGEMA_signal_7564), .Q (new_AGEMA_signal_7565) ) ;
    buf_clk new_AGEMA_reg_buffer_4138 ( .C (clk), .D (new_AGEMA_signal_7568), .Q (new_AGEMA_signal_7569) ) ;
    buf_clk new_AGEMA_reg_buffer_4142 ( .C (clk), .D (new_AGEMA_signal_7572), .Q (new_AGEMA_signal_7573) ) ;
    buf_clk new_AGEMA_reg_buffer_4146 ( .C (clk), .D (new_AGEMA_signal_7576), .Q (new_AGEMA_signal_7577) ) ;
    buf_clk new_AGEMA_reg_buffer_4150 ( .C (clk), .D (new_AGEMA_signal_7580), .Q (new_AGEMA_signal_7581) ) ;
    buf_clk new_AGEMA_reg_buffer_4154 ( .C (clk), .D (new_AGEMA_signal_7584), .Q (new_AGEMA_signal_7585) ) ;
    buf_clk new_AGEMA_reg_buffer_4158 ( .C (clk), .D (new_AGEMA_signal_7588), .Q (new_AGEMA_signal_7589) ) ;
    buf_clk new_AGEMA_reg_buffer_4162 ( .C (clk), .D (new_AGEMA_signal_7592), .Q (new_AGEMA_signal_7593) ) ;
    buf_clk new_AGEMA_reg_buffer_4166 ( .C (clk), .D (new_AGEMA_signal_7596), .Q (new_AGEMA_signal_7597) ) ;
    buf_clk new_AGEMA_reg_buffer_4170 ( .C (clk), .D (new_AGEMA_signal_7600), .Q (new_AGEMA_signal_7601) ) ;
    buf_clk new_AGEMA_reg_buffer_4174 ( .C (clk), .D (new_AGEMA_signal_7604), .Q (new_AGEMA_signal_7605) ) ;
    buf_clk new_AGEMA_reg_buffer_4178 ( .C (clk), .D (new_AGEMA_signal_7608), .Q (new_AGEMA_signal_7609) ) ;
    buf_clk new_AGEMA_reg_buffer_4182 ( .C (clk), .D (new_AGEMA_signal_7612), .Q (new_AGEMA_signal_7613) ) ;
    buf_clk new_AGEMA_reg_buffer_4186 ( .C (clk), .D (new_AGEMA_signal_7616), .Q (new_AGEMA_signal_7617) ) ;
    buf_clk new_AGEMA_reg_buffer_4190 ( .C (clk), .D (new_AGEMA_signal_7620), .Q (new_AGEMA_signal_7621) ) ;
    buf_clk new_AGEMA_reg_buffer_4194 ( .C (clk), .D (new_AGEMA_signal_7624), .Q (new_AGEMA_signal_7625) ) ;
    buf_clk new_AGEMA_reg_buffer_4198 ( .C (clk), .D (new_AGEMA_signal_7628), .Q (new_AGEMA_signal_7629) ) ;
    buf_clk new_AGEMA_reg_buffer_4202 ( .C (clk), .D (new_AGEMA_signal_7632), .Q (new_AGEMA_signal_7633) ) ;
    buf_clk new_AGEMA_reg_buffer_4206 ( .C (clk), .D (new_AGEMA_signal_7636), .Q (new_AGEMA_signal_7637) ) ;
    buf_clk new_AGEMA_reg_buffer_4210 ( .C (clk), .D (new_AGEMA_signal_7640), .Q (new_AGEMA_signal_7641) ) ;
    buf_clk new_AGEMA_reg_buffer_4214 ( .C (clk), .D (new_AGEMA_signal_7644), .Q (new_AGEMA_signal_7645) ) ;
    buf_clk new_AGEMA_reg_buffer_4218 ( .C (clk), .D (new_AGEMA_signal_7648), .Q (new_AGEMA_signal_7649) ) ;
    buf_clk new_AGEMA_reg_buffer_4222 ( .C (clk), .D (new_AGEMA_signal_7652), .Q (new_AGEMA_signal_7653) ) ;
    buf_clk new_AGEMA_reg_buffer_4226 ( .C (clk), .D (new_AGEMA_signal_7656), .Q (new_AGEMA_signal_7657) ) ;
    buf_clk new_AGEMA_reg_buffer_4230 ( .C (clk), .D (new_AGEMA_signal_7660), .Q (new_AGEMA_signal_7661) ) ;
    buf_clk new_AGEMA_reg_buffer_4234 ( .C (clk), .D (new_AGEMA_signal_7664), .Q (new_AGEMA_signal_7665) ) ;
    buf_clk new_AGEMA_reg_buffer_4238 ( .C (clk), .D (new_AGEMA_signal_7668), .Q (new_AGEMA_signal_7669) ) ;
    buf_clk new_AGEMA_reg_buffer_4242 ( .C (clk), .D (new_AGEMA_signal_7672), .Q (new_AGEMA_signal_7673) ) ;
    buf_clk new_AGEMA_reg_buffer_4246 ( .C (clk), .D (new_AGEMA_signal_7676), .Q (new_AGEMA_signal_7677) ) ;
    buf_clk new_AGEMA_reg_buffer_4250 ( .C (clk), .D (new_AGEMA_signal_7680), .Q (new_AGEMA_signal_7681) ) ;
    buf_clk new_AGEMA_reg_buffer_4254 ( .C (clk), .D (new_AGEMA_signal_7684), .Q (new_AGEMA_signal_7685) ) ;
    buf_clk new_AGEMA_reg_buffer_4258 ( .C (clk), .D (new_AGEMA_signal_7688), .Q (new_AGEMA_signal_7689) ) ;
    buf_clk new_AGEMA_reg_buffer_4262 ( .C (clk), .D (new_AGEMA_signal_7692), .Q (new_AGEMA_signal_7693) ) ;
    buf_clk new_AGEMA_reg_buffer_4266 ( .C (clk), .D (new_AGEMA_signal_7696), .Q (new_AGEMA_signal_7697) ) ;
    buf_clk new_AGEMA_reg_buffer_4270 ( .C (clk), .D (new_AGEMA_signal_7700), .Q (new_AGEMA_signal_7701) ) ;
    buf_clk new_AGEMA_reg_buffer_4274 ( .C (clk), .D (new_AGEMA_signal_7704), .Q (new_AGEMA_signal_7705) ) ;
    buf_clk new_AGEMA_reg_buffer_4278 ( .C (clk), .D (new_AGEMA_signal_7708), .Q (new_AGEMA_signal_7709) ) ;
    buf_clk new_AGEMA_reg_buffer_4282 ( .C (clk), .D (new_AGEMA_signal_7712), .Q (new_AGEMA_signal_7713) ) ;
    buf_clk new_AGEMA_reg_buffer_4286 ( .C (clk), .D (new_AGEMA_signal_7716), .Q (new_AGEMA_signal_7717) ) ;
    buf_clk new_AGEMA_reg_buffer_4290 ( .C (clk), .D (new_AGEMA_signal_7720), .Q (new_AGEMA_signal_7721) ) ;
    buf_clk new_AGEMA_reg_buffer_4294 ( .C (clk), .D (new_AGEMA_signal_7724), .Q (new_AGEMA_signal_7725) ) ;
    buf_clk new_AGEMA_reg_buffer_4298 ( .C (clk), .D (new_AGEMA_signal_7728), .Q (new_AGEMA_signal_7729) ) ;
    buf_clk new_AGEMA_reg_buffer_4302 ( .C (clk), .D (new_AGEMA_signal_7732), .Q (new_AGEMA_signal_7733) ) ;
    buf_clk new_AGEMA_reg_buffer_4306 ( .C (clk), .D (new_AGEMA_signal_7736), .Q (new_AGEMA_signal_7737) ) ;
    buf_clk new_AGEMA_reg_buffer_4310 ( .C (clk), .D (new_AGEMA_signal_7740), .Q (new_AGEMA_signal_7741) ) ;
    buf_clk new_AGEMA_reg_buffer_4314 ( .C (clk), .D (new_AGEMA_signal_7744), .Q (new_AGEMA_signal_7745) ) ;
    buf_clk new_AGEMA_reg_buffer_4318 ( .C (clk), .D (new_AGEMA_signal_7748), .Q (new_AGEMA_signal_7749) ) ;
    buf_clk new_AGEMA_reg_buffer_4322 ( .C (clk), .D (new_AGEMA_signal_7752), .Q (new_AGEMA_signal_7753) ) ;
    buf_clk new_AGEMA_reg_buffer_4326 ( .C (clk), .D (new_AGEMA_signal_7756), .Q (new_AGEMA_signal_7757) ) ;
    buf_clk new_AGEMA_reg_buffer_4330 ( .C (clk), .D (new_AGEMA_signal_7760), .Q (new_AGEMA_signal_7761) ) ;
    buf_clk new_AGEMA_reg_buffer_4334 ( .C (clk), .D (new_AGEMA_signal_7764), .Q (new_AGEMA_signal_7765) ) ;
    buf_clk new_AGEMA_reg_buffer_4338 ( .C (clk), .D (new_AGEMA_signal_7768), .Q (new_AGEMA_signal_7769) ) ;
    buf_clk new_AGEMA_reg_buffer_4342 ( .C (clk), .D (new_AGEMA_signal_7772), .Q (new_AGEMA_signal_7773) ) ;
    buf_clk new_AGEMA_reg_buffer_4346 ( .C (clk), .D (new_AGEMA_signal_7776), .Q (new_AGEMA_signal_7777) ) ;
    buf_clk new_AGEMA_reg_buffer_4350 ( .C (clk), .D (new_AGEMA_signal_7780), .Q (new_AGEMA_signal_7781) ) ;
    buf_clk new_AGEMA_reg_buffer_4354 ( .C (clk), .D (new_AGEMA_signal_7784), .Q (new_AGEMA_signal_7785) ) ;
    buf_clk new_AGEMA_reg_buffer_4358 ( .C (clk), .D (new_AGEMA_signal_7788), .Q (new_AGEMA_signal_7789) ) ;
    buf_clk new_AGEMA_reg_buffer_4362 ( .C (clk), .D (new_AGEMA_signal_7792), .Q (new_AGEMA_signal_7793) ) ;
    buf_clk new_AGEMA_reg_buffer_4366 ( .C (clk), .D (new_AGEMA_signal_7796), .Q (new_AGEMA_signal_7797) ) ;
    buf_clk new_AGEMA_reg_buffer_4370 ( .C (clk), .D (new_AGEMA_signal_7800), .Q (new_AGEMA_signal_7801) ) ;
    buf_clk new_AGEMA_reg_buffer_4374 ( .C (clk), .D (new_AGEMA_signal_7804), .Q (new_AGEMA_signal_7805) ) ;
    buf_clk new_AGEMA_reg_buffer_4378 ( .C (clk), .D (new_AGEMA_signal_7808), .Q (new_AGEMA_signal_7809) ) ;
    buf_clk new_AGEMA_reg_buffer_4382 ( .C (clk), .D (new_AGEMA_signal_7812), .Q (new_AGEMA_signal_7813) ) ;
    buf_clk new_AGEMA_reg_buffer_4386 ( .C (clk), .D (new_AGEMA_signal_7816), .Q (new_AGEMA_signal_7817) ) ;
    buf_clk new_AGEMA_reg_buffer_4390 ( .C (clk), .D (new_AGEMA_signal_7820), .Q (new_AGEMA_signal_7821) ) ;
    buf_clk new_AGEMA_reg_buffer_4394 ( .C (clk), .D (new_AGEMA_signal_7824), .Q (new_AGEMA_signal_7825) ) ;
    buf_clk new_AGEMA_reg_buffer_4398 ( .C (clk), .D (new_AGEMA_signal_7828), .Q (new_AGEMA_signal_7829) ) ;
    buf_clk new_AGEMA_reg_buffer_4402 ( .C (clk), .D (new_AGEMA_signal_7832), .Q (new_AGEMA_signal_7833) ) ;
    buf_clk new_AGEMA_reg_buffer_4406 ( .C (clk), .D (new_AGEMA_signal_7836), .Q (new_AGEMA_signal_7837) ) ;
    buf_clk new_AGEMA_reg_buffer_4410 ( .C (clk), .D (new_AGEMA_signal_7840), .Q (new_AGEMA_signal_7841) ) ;
    buf_clk new_AGEMA_reg_buffer_4414 ( .C (clk), .D (new_AGEMA_signal_7844), .Q (new_AGEMA_signal_7845) ) ;
    buf_clk new_AGEMA_reg_buffer_4418 ( .C (clk), .D (new_AGEMA_signal_7848), .Q (new_AGEMA_signal_7849) ) ;
    buf_clk new_AGEMA_reg_buffer_4422 ( .C (clk), .D (new_AGEMA_signal_7852), .Q (new_AGEMA_signal_7853) ) ;
    buf_clk new_AGEMA_reg_buffer_4426 ( .C (clk), .D (new_AGEMA_signal_7856), .Q (new_AGEMA_signal_7857) ) ;
    buf_clk new_AGEMA_reg_buffer_4430 ( .C (clk), .D (new_AGEMA_signal_7860), .Q (new_AGEMA_signal_7861) ) ;
    buf_clk new_AGEMA_reg_buffer_4434 ( .C (clk), .D (new_AGEMA_signal_7864), .Q (new_AGEMA_signal_7865) ) ;
    buf_clk new_AGEMA_reg_buffer_4438 ( .C (clk), .D (new_AGEMA_signal_7868), .Q (new_AGEMA_signal_7869) ) ;
    buf_clk new_AGEMA_reg_buffer_4442 ( .C (clk), .D (new_AGEMA_signal_7872), .Q (new_AGEMA_signal_7873) ) ;
    buf_clk new_AGEMA_reg_buffer_4446 ( .C (clk), .D (new_AGEMA_signal_7876), .Q (new_AGEMA_signal_7877) ) ;
    buf_clk new_AGEMA_reg_buffer_4450 ( .C (clk), .D (new_AGEMA_signal_7880), .Q (new_AGEMA_signal_7881) ) ;
    buf_clk new_AGEMA_reg_buffer_4454 ( .C (clk), .D (new_AGEMA_signal_7884), .Q (new_AGEMA_signal_7885) ) ;
    buf_clk new_AGEMA_reg_buffer_4458 ( .C (clk), .D (new_AGEMA_signal_7888), .Q (new_AGEMA_signal_7889) ) ;
    buf_clk new_AGEMA_reg_buffer_4462 ( .C (clk), .D (new_AGEMA_signal_7892), .Q (new_AGEMA_signal_7893) ) ;
    buf_clk new_AGEMA_reg_buffer_4466 ( .C (clk), .D (new_AGEMA_signal_7896), .Q (new_AGEMA_signal_7897) ) ;
    buf_clk new_AGEMA_reg_buffer_4470 ( .C (clk), .D (new_AGEMA_signal_7900), .Q (new_AGEMA_signal_7901) ) ;
    buf_clk new_AGEMA_reg_buffer_4474 ( .C (clk), .D (new_AGEMA_signal_7904), .Q (new_AGEMA_signal_7905) ) ;
    buf_clk new_AGEMA_reg_buffer_4478 ( .C (clk), .D (new_AGEMA_signal_7908), .Q (new_AGEMA_signal_7909) ) ;
    buf_clk new_AGEMA_reg_buffer_4482 ( .C (clk), .D (new_AGEMA_signal_7912), .Q (new_AGEMA_signal_7913) ) ;
    buf_clk new_AGEMA_reg_buffer_4486 ( .C (clk), .D (new_AGEMA_signal_7916), .Q (new_AGEMA_signal_7917) ) ;
    buf_clk new_AGEMA_reg_buffer_4490 ( .C (clk), .D (new_AGEMA_signal_7920), .Q (new_AGEMA_signal_7921) ) ;
    buf_clk new_AGEMA_reg_buffer_4494 ( .C (clk), .D (new_AGEMA_signal_7924), .Q (new_AGEMA_signal_7925) ) ;
    buf_clk new_AGEMA_reg_buffer_4498 ( .C (clk), .D (new_AGEMA_signal_7928), .Q (new_AGEMA_signal_7929) ) ;
    buf_clk new_AGEMA_reg_buffer_4502 ( .C (clk), .D (new_AGEMA_signal_7932), .Q (new_AGEMA_signal_7933) ) ;
    buf_clk new_AGEMA_reg_buffer_4506 ( .C (clk), .D (new_AGEMA_signal_7936), .Q (new_AGEMA_signal_7937) ) ;
    buf_clk new_AGEMA_reg_buffer_4510 ( .C (clk), .D (new_AGEMA_signal_7940), .Q (new_AGEMA_signal_7941) ) ;
    buf_clk new_AGEMA_reg_buffer_4514 ( .C (clk), .D (new_AGEMA_signal_7944), .Q (new_AGEMA_signal_7945) ) ;
    buf_clk new_AGEMA_reg_buffer_4518 ( .C (clk), .D (new_AGEMA_signal_7948), .Q (new_AGEMA_signal_7949) ) ;
    buf_clk new_AGEMA_reg_buffer_4522 ( .C (clk), .D (new_AGEMA_signal_7952), .Q (new_AGEMA_signal_7953) ) ;
    buf_clk new_AGEMA_reg_buffer_4526 ( .C (clk), .D (new_AGEMA_signal_7956), .Q (new_AGEMA_signal_7957) ) ;
    buf_clk new_AGEMA_reg_buffer_4530 ( .C (clk), .D (new_AGEMA_signal_7960), .Q (new_AGEMA_signal_7961) ) ;
    buf_clk new_AGEMA_reg_buffer_4534 ( .C (clk), .D (new_AGEMA_signal_7964), .Q (new_AGEMA_signal_7965) ) ;
    buf_clk new_AGEMA_reg_buffer_4538 ( .C (clk), .D (new_AGEMA_signal_7968), .Q (new_AGEMA_signal_7969) ) ;
    buf_clk new_AGEMA_reg_buffer_4542 ( .C (clk), .D (new_AGEMA_signal_7972), .Q (new_AGEMA_signal_7973) ) ;
    buf_clk new_AGEMA_reg_buffer_4546 ( .C (clk), .D (new_AGEMA_signal_7976), .Q (new_AGEMA_signal_7977) ) ;
    buf_clk new_AGEMA_reg_buffer_4550 ( .C (clk), .D (new_AGEMA_signal_7980), .Q (new_AGEMA_signal_7981) ) ;
    buf_clk new_AGEMA_reg_buffer_4554 ( .C (clk), .D (new_AGEMA_signal_7984), .Q (new_AGEMA_signal_7985) ) ;
    buf_clk new_AGEMA_reg_buffer_4558 ( .C (clk), .D (new_AGEMA_signal_7988), .Q (new_AGEMA_signal_7989) ) ;
    buf_clk new_AGEMA_reg_buffer_4562 ( .C (clk), .D (new_AGEMA_signal_7992), .Q (new_AGEMA_signal_7993) ) ;
    buf_clk new_AGEMA_reg_buffer_4566 ( .C (clk), .D (new_AGEMA_signal_7996), .Q (new_AGEMA_signal_7997) ) ;
    buf_clk new_AGEMA_reg_buffer_4570 ( .C (clk), .D (new_AGEMA_signal_8000), .Q (new_AGEMA_signal_8001) ) ;
    buf_clk new_AGEMA_reg_buffer_4574 ( .C (clk), .D (new_AGEMA_signal_8004), .Q (new_AGEMA_signal_8005) ) ;
    buf_clk new_AGEMA_reg_buffer_4578 ( .C (clk), .D (new_AGEMA_signal_8008), .Q (new_AGEMA_signal_8009) ) ;
    buf_clk new_AGEMA_reg_buffer_4582 ( .C (clk), .D (new_AGEMA_signal_8012), .Q (new_AGEMA_signal_8013) ) ;
    buf_clk new_AGEMA_reg_buffer_4586 ( .C (clk), .D (new_AGEMA_signal_8016), .Q (new_AGEMA_signal_8017) ) ;
    buf_clk new_AGEMA_reg_buffer_4590 ( .C (clk), .D (new_AGEMA_signal_8020), .Q (new_AGEMA_signal_8021) ) ;
    buf_clk new_AGEMA_reg_buffer_4594 ( .C (clk), .D (new_AGEMA_signal_8024), .Q (new_AGEMA_signal_8025) ) ;
    buf_clk new_AGEMA_reg_buffer_4598 ( .C (clk), .D (new_AGEMA_signal_8028), .Q (new_AGEMA_signal_8029) ) ;
    buf_clk new_AGEMA_reg_buffer_4602 ( .C (clk), .D (new_AGEMA_signal_8032), .Q (new_AGEMA_signal_8033) ) ;
    buf_clk new_AGEMA_reg_buffer_4606 ( .C (clk), .D (new_AGEMA_signal_8036), .Q (new_AGEMA_signal_8037) ) ;
    buf_clk new_AGEMA_reg_buffer_4610 ( .C (clk), .D (new_AGEMA_signal_8040), .Q (new_AGEMA_signal_8041) ) ;
    buf_clk new_AGEMA_reg_buffer_4614 ( .C (clk), .D (new_AGEMA_signal_8044), .Q (new_AGEMA_signal_8045) ) ;
    buf_clk new_AGEMA_reg_buffer_4618 ( .C (clk), .D (new_AGEMA_signal_8048), .Q (new_AGEMA_signal_8049) ) ;
    buf_clk new_AGEMA_reg_buffer_4622 ( .C (clk), .D (new_AGEMA_signal_8052), .Q (new_AGEMA_signal_8053) ) ;
    buf_clk new_AGEMA_reg_buffer_4626 ( .C (clk), .D (new_AGEMA_signal_8056), .Q (new_AGEMA_signal_8057) ) ;
    buf_clk new_AGEMA_reg_buffer_4630 ( .C (clk), .D (new_AGEMA_signal_8060), .Q (new_AGEMA_signal_8061) ) ;
    buf_clk new_AGEMA_reg_buffer_4634 ( .C (clk), .D (new_AGEMA_signal_8064), .Q (new_AGEMA_signal_8065) ) ;
    buf_clk new_AGEMA_reg_buffer_4638 ( .C (clk), .D (new_AGEMA_signal_8068), .Q (new_AGEMA_signal_8069) ) ;
    buf_clk new_AGEMA_reg_buffer_4642 ( .C (clk), .D (new_AGEMA_signal_8072), .Q (new_AGEMA_signal_8073) ) ;
    buf_clk new_AGEMA_reg_buffer_4646 ( .C (clk), .D (new_AGEMA_signal_8076), .Q (new_AGEMA_signal_8077) ) ;
    buf_clk new_AGEMA_reg_buffer_4650 ( .C (clk), .D (new_AGEMA_signal_8080), .Q (new_AGEMA_signal_8081) ) ;
    buf_clk new_AGEMA_reg_buffer_4654 ( .C (clk), .D (new_AGEMA_signal_8084), .Q (new_AGEMA_signal_8085) ) ;
    buf_clk new_AGEMA_reg_buffer_4658 ( .C (clk), .D (new_AGEMA_signal_8088), .Q (new_AGEMA_signal_8089) ) ;
    buf_clk new_AGEMA_reg_buffer_4662 ( .C (clk), .D (new_AGEMA_signal_8092), .Q (new_AGEMA_signal_8093) ) ;
    buf_clk new_AGEMA_reg_buffer_4666 ( .C (clk), .D (new_AGEMA_signal_8096), .Q (new_AGEMA_signal_8097) ) ;
    buf_clk new_AGEMA_reg_buffer_4670 ( .C (clk), .D (new_AGEMA_signal_8100), .Q (new_AGEMA_signal_8101) ) ;
    buf_clk new_AGEMA_reg_buffer_4674 ( .C (clk), .D (new_AGEMA_signal_8104), .Q (new_AGEMA_signal_8105) ) ;
    buf_clk new_AGEMA_reg_buffer_4678 ( .C (clk), .D (new_AGEMA_signal_8108), .Q (new_AGEMA_signal_8109) ) ;
    buf_clk new_AGEMA_reg_buffer_4682 ( .C (clk), .D (new_AGEMA_signal_8112), .Q (new_AGEMA_signal_8113) ) ;
    buf_clk new_AGEMA_reg_buffer_4686 ( .C (clk), .D (new_AGEMA_signal_8116), .Q (new_AGEMA_signal_8117) ) ;
    buf_clk new_AGEMA_reg_buffer_4690 ( .C (clk), .D (new_AGEMA_signal_8120), .Q (new_AGEMA_signal_8121) ) ;
    buf_clk new_AGEMA_reg_buffer_4694 ( .C (clk), .D (new_AGEMA_signal_8124), .Q (new_AGEMA_signal_8125) ) ;
    buf_clk new_AGEMA_reg_buffer_4698 ( .C (clk), .D (new_AGEMA_signal_8128), .Q (new_AGEMA_signal_8129) ) ;
    buf_clk new_AGEMA_reg_buffer_4702 ( .C (clk), .D (new_AGEMA_signal_8132), .Q (new_AGEMA_signal_8133) ) ;
    buf_clk new_AGEMA_reg_buffer_4706 ( .C (clk), .D (new_AGEMA_signal_8136), .Q (new_AGEMA_signal_8137) ) ;
    buf_clk new_AGEMA_reg_buffer_4710 ( .C (clk), .D (new_AGEMA_signal_8140), .Q (new_AGEMA_signal_8141) ) ;
    buf_clk new_AGEMA_reg_buffer_4714 ( .C (clk), .D (new_AGEMA_signal_8144), .Q (new_AGEMA_signal_8145) ) ;
    buf_clk new_AGEMA_reg_buffer_4718 ( .C (clk), .D (new_AGEMA_signal_8148), .Q (new_AGEMA_signal_8149) ) ;
    buf_clk new_AGEMA_reg_buffer_4722 ( .C (clk), .D (new_AGEMA_signal_8152), .Q (new_AGEMA_signal_8153) ) ;
    buf_clk new_AGEMA_reg_buffer_4726 ( .C (clk), .D (new_AGEMA_signal_8156), .Q (new_AGEMA_signal_8157) ) ;
    buf_clk new_AGEMA_reg_buffer_4730 ( .C (clk), .D (new_AGEMA_signal_8160), .Q (new_AGEMA_signal_8161) ) ;
    buf_clk new_AGEMA_reg_buffer_4734 ( .C (clk), .D (new_AGEMA_signal_8164), .Q (new_AGEMA_signal_8165) ) ;
    buf_clk new_AGEMA_reg_buffer_4738 ( .C (clk), .D (new_AGEMA_signal_8168), .Q (new_AGEMA_signal_8169) ) ;
    buf_clk new_AGEMA_reg_buffer_4742 ( .C (clk), .D (new_AGEMA_signal_8172), .Q (new_AGEMA_signal_8173) ) ;
    buf_clk new_AGEMA_reg_buffer_4746 ( .C (clk), .D (new_AGEMA_signal_8176), .Q (new_AGEMA_signal_8177) ) ;
    buf_clk new_AGEMA_reg_buffer_4750 ( .C (clk), .D (new_AGEMA_signal_8180), .Q (new_AGEMA_signal_8181) ) ;
    buf_clk new_AGEMA_reg_buffer_4754 ( .C (clk), .D (new_AGEMA_signal_8184), .Q (new_AGEMA_signal_8185) ) ;
    buf_clk new_AGEMA_reg_buffer_4758 ( .C (clk), .D (new_AGEMA_signal_8188), .Q (new_AGEMA_signal_8189) ) ;

    /* cells in depth 4 */
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_0_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, new_AGEMA_signal_3753, MCOutput[0]}), .a ({new_AGEMA_signal_5350, new_AGEMA_signal_5346, new_AGEMA_signal_5342, new_AGEMA_signal_5338}), .c ({new_AGEMA_signal_3782, new_AGEMA_signal_3781, new_AGEMA_signal_3780, StateRegInput[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_1_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, new_AGEMA_signal_3891, MCOutput[1]}), .a ({new_AGEMA_signal_5366, new_AGEMA_signal_5362, new_AGEMA_signal_5358, new_AGEMA_signal_5354}), .c ({new_AGEMA_signal_3911, new_AGEMA_signal_3910, new_AGEMA_signal_3909, StateRegInput[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_4_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, new_AGEMA_signal_3759, MCOutput[4]}), .a ({new_AGEMA_signal_5382, new_AGEMA_signal_5378, new_AGEMA_signal_5374, new_AGEMA_signal_5370}), .c ({new_AGEMA_signal_3788, new_AGEMA_signal_3787, new_AGEMA_signal_3786, StateRegInput[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_5_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3896, new_AGEMA_signal_3895, new_AGEMA_signal_3894, MCOutput[5]}), .a ({new_AGEMA_signal_5398, new_AGEMA_signal_5394, new_AGEMA_signal_5390, new_AGEMA_signal_5386}), .c ({new_AGEMA_signal_3917, new_AGEMA_signal_3916, new_AGEMA_signal_3915, StateRegInput[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_8_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, new_AGEMA_signal_3765, MCOutput[8]}), .a ({new_AGEMA_signal_5414, new_AGEMA_signal_5410, new_AGEMA_signal_5406, new_AGEMA_signal_5402}), .c ({new_AGEMA_signal_3794, new_AGEMA_signal_3793, new_AGEMA_signal_3792, StateRegInput[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_9_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3899, new_AGEMA_signal_3898, new_AGEMA_signal_3897, MCOutput[9]}), .a ({new_AGEMA_signal_5430, new_AGEMA_signal_5426, new_AGEMA_signal_5422, new_AGEMA_signal_5418}), .c ({new_AGEMA_signal_3923, new_AGEMA_signal_3922, new_AGEMA_signal_3921, StateRegInput[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_12_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3998, new_AGEMA_signal_3997, new_AGEMA_signal_3996, MCOutput[12]}), .a ({new_AGEMA_signal_5446, new_AGEMA_signal_5442, new_AGEMA_signal_5438, new_AGEMA_signal_5434}), .c ({new_AGEMA_signal_4007, new_AGEMA_signal_4006, new_AGEMA_signal_4005, StateRegInput[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_13_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_4028, new_AGEMA_signal_4027, new_AGEMA_signal_4026, MCOutput[13]}), .a ({new_AGEMA_signal_5462, new_AGEMA_signal_5458, new_AGEMA_signal_5454, new_AGEMA_signal_5450}), .c ({new_AGEMA_signal_4034, new_AGEMA_signal_4033, new_AGEMA_signal_4032, StateRegInput[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_16_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3731, new_AGEMA_signal_3730, new_AGEMA_signal_3729, MCOutput[16]}), .a ({new_AGEMA_signal_5478, new_AGEMA_signal_5474, new_AGEMA_signal_5470, new_AGEMA_signal_5466}), .c ({new_AGEMA_signal_3806, new_AGEMA_signal_3805, new_AGEMA_signal_3804, StateRegInput[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_17_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3878, new_AGEMA_signal_3877, new_AGEMA_signal_3876, MCOutput[17]}), .a ({new_AGEMA_signal_5494, new_AGEMA_signal_5490, new_AGEMA_signal_5486, new_AGEMA_signal_5482}), .c ({new_AGEMA_signal_3935, new_AGEMA_signal_3934, new_AGEMA_signal_3933, StateRegInput[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_20_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3737, new_AGEMA_signal_3736, new_AGEMA_signal_3735, MCOutput[20]}), .a ({new_AGEMA_signal_5510, new_AGEMA_signal_5506, new_AGEMA_signal_5502, new_AGEMA_signal_5498}), .c ({new_AGEMA_signal_3812, new_AGEMA_signal_3811, new_AGEMA_signal_3810, StateRegInput[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_21_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, new_AGEMA_signal_3879, MCOutput[21]}), .a ({new_AGEMA_signal_5526, new_AGEMA_signal_5522, new_AGEMA_signal_5518, new_AGEMA_signal_5514}), .c ({new_AGEMA_signal_3941, new_AGEMA_signal_3940, new_AGEMA_signal_3939, StateRegInput[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_24_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3992, new_AGEMA_signal_3991, new_AGEMA_signal_3990, MCOutput[24]}), .a ({new_AGEMA_signal_5542, new_AGEMA_signal_5538, new_AGEMA_signal_5534, new_AGEMA_signal_5530}), .c ({new_AGEMA_signal_4013, new_AGEMA_signal_4012, new_AGEMA_signal_4011, StateRegInput[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_25_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_4025, new_AGEMA_signal_4024, new_AGEMA_signal_4023, MCOutput[25]}), .a ({new_AGEMA_signal_5558, new_AGEMA_signal_5554, new_AGEMA_signal_5550, new_AGEMA_signal_5546}), .c ({new_AGEMA_signal_4040, new_AGEMA_signal_4039, new_AGEMA_signal_4038, StateRegInput[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_28_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, new_AGEMA_signal_3747, MCOutput[28]}), .a ({new_AGEMA_signal_5574, new_AGEMA_signal_5570, new_AGEMA_signal_5566, new_AGEMA_signal_5562}), .c ({new_AGEMA_signal_3824, new_AGEMA_signal_3823, new_AGEMA_signal_3822, StateRegInput[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_29_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3890, new_AGEMA_signal_3889, new_AGEMA_signal_3888, MCOutput[29]}), .a ({new_AGEMA_signal_5590, new_AGEMA_signal_5586, new_AGEMA_signal_5582, new_AGEMA_signal_5578}), .c ({new_AGEMA_signal_3953, new_AGEMA_signal_3952, new_AGEMA_signal_3951, StateRegInput[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_32_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3350, new_AGEMA_signal_3349, new_AGEMA_signal_3348, MCOutput[32]}), .a ({new_AGEMA_signal_5606, new_AGEMA_signal_5602, new_AGEMA_signal_5598, new_AGEMA_signal_5594}), .c ({new_AGEMA_signal_3476, new_AGEMA_signal_3475, new_AGEMA_signal_3474, StateRegInput[32]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_33_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3536, new_AGEMA_signal_3535, new_AGEMA_signal_3534, MCOutput[33]}), .a ({new_AGEMA_signal_5622, new_AGEMA_signal_5618, new_AGEMA_signal_5614, new_AGEMA_signal_5610}), .c ({new_AGEMA_signal_3656, new_AGEMA_signal_3655, new_AGEMA_signal_3654, StateRegInput[33]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_36_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3356, new_AGEMA_signal_3355, new_AGEMA_signal_3354, MCOutput[36]}), .a ({new_AGEMA_signal_5638, new_AGEMA_signal_5634, new_AGEMA_signal_5630, new_AGEMA_signal_5626}), .c ({new_AGEMA_signal_3482, new_AGEMA_signal_3481, new_AGEMA_signal_3480, StateRegInput[36]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_37_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, new_AGEMA_signal_3537, MCOutput[37]}), .a ({new_AGEMA_signal_5654, new_AGEMA_signal_5650, new_AGEMA_signal_5646, new_AGEMA_signal_5642}), .c ({new_AGEMA_signal_3662, new_AGEMA_signal_3661, new_AGEMA_signal_3660, StateRegInput[37]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_40_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3362, new_AGEMA_signal_3361, new_AGEMA_signal_3360, MCOutput[40]}), .a ({new_AGEMA_signal_5670, new_AGEMA_signal_5666, new_AGEMA_signal_5662, new_AGEMA_signal_5658}), .c ({new_AGEMA_signal_3488, new_AGEMA_signal_3487, new_AGEMA_signal_3486, StateRegInput[40]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_41_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3542, new_AGEMA_signal_3541, new_AGEMA_signal_3540, MCOutput[41]}), .a ({new_AGEMA_signal_5686, new_AGEMA_signal_5682, new_AGEMA_signal_5678, new_AGEMA_signal_5674}), .c ({new_AGEMA_signal_3668, new_AGEMA_signal_3667, new_AGEMA_signal_3666, StateRegInput[41]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_44_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, new_AGEMA_signal_3699, MCOutput[44]}), .a ({new_AGEMA_signal_5702, new_AGEMA_signal_5698, new_AGEMA_signal_5694, new_AGEMA_signal_5690}), .c ({new_AGEMA_signal_3830, new_AGEMA_signal_3829, new_AGEMA_signal_3828, StateRegInput[44]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_45_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3860, new_AGEMA_signal_3859, new_AGEMA_signal_3858, MCOutput[45]}), .a ({new_AGEMA_signal_5718, new_AGEMA_signal_5714, new_AGEMA_signal_5710, new_AGEMA_signal_5706}), .c ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, new_AGEMA_signal_3957, StateRegInput[45]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_48_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, new_AGEMA_signal_3705, MCOutput[48]}), .a ({new_AGEMA_signal_5734, new_AGEMA_signal_5730, new_AGEMA_signal_5726, new_AGEMA_signal_5722}), .c ({new_AGEMA_signal_3836, new_AGEMA_signal_3835, new_AGEMA_signal_3834, StateRegInput[48]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_49_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3863, new_AGEMA_signal_3862, new_AGEMA_signal_3861, MCOutput[49]}), .a ({new_AGEMA_signal_5750, new_AGEMA_signal_5746, new_AGEMA_signal_5742, new_AGEMA_signal_5738}), .c ({new_AGEMA_signal_3965, new_AGEMA_signal_3964, new_AGEMA_signal_3963, StateRegInput[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_52_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, new_AGEMA_signal_3711, MCOutput[52]}), .a ({new_AGEMA_signal_5766, new_AGEMA_signal_5762, new_AGEMA_signal_5758, new_AGEMA_signal_5754}), .c ({new_AGEMA_signal_3842, new_AGEMA_signal_3841, new_AGEMA_signal_3840, StateRegInput[52]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_53_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3866, new_AGEMA_signal_3865, new_AGEMA_signal_3864, MCOutput[53]}), .a ({new_AGEMA_signal_5782, new_AGEMA_signal_5778, new_AGEMA_signal_5774, new_AGEMA_signal_5770}), .c ({new_AGEMA_signal_3971, new_AGEMA_signal_3970, new_AGEMA_signal_3969, StateRegInput[53]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_56_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, new_AGEMA_signal_3717, MCOutput[56]}), .a ({new_AGEMA_signal_5798, new_AGEMA_signal_5794, new_AGEMA_signal_5790, new_AGEMA_signal_5786}), .c ({new_AGEMA_signal_3848, new_AGEMA_signal_3847, new_AGEMA_signal_3846, StateRegInput[56]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_57_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, new_AGEMA_signal_3867, MCOutput[57]}), .a ({new_AGEMA_signal_5814, new_AGEMA_signal_5810, new_AGEMA_signal_5806, new_AGEMA_signal_5802}), .c ({new_AGEMA_signal_3977, new_AGEMA_signal_3976, new_AGEMA_signal_3975, StateRegInput[57]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_60_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_3986, new_AGEMA_signal_3985, new_AGEMA_signal_3984, MCOutput[60]}), .a ({new_AGEMA_signal_5830, new_AGEMA_signal_5826, new_AGEMA_signal_5822, new_AGEMA_signal_5818}), .c ({new_AGEMA_signal_4019, new_AGEMA_signal_4018, new_AGEMA_signal_4017, StateRegInput[60]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) PlaintextMUX_MUXInst_61_U1 ( .s (new_AGEMA_signal_5334), .b ({new_AGEMA_signal_4022, new_AGEMA_signal_4021, new_AGEMA_signal_4020, MCOutput[61]}), .a ({new_AGEMA_signal_5846, new_AGEMA_signal_5842, new_AGEMA_signal_5838, new_AGEMA_signal_5834}), .c ({new_AGEMA_signal_4046, new_AGEMA_signal_4045, new_AGEMA_signal_4044, StateRegInput[61]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_AND2_U1 ( .a ({new_AGEMA_signal_5854, new_AGEMA_signal_5852, new_AGEMA_signal_5850, new_AGEMA_signal_5848}), .b ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, new_AGEMA_signal_2460, SubCellInst_SboxInst_0_Q2}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, new_AGEMA_signal_2655, SubCellInst_SboxInst_0_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_XOR4_U1 ( .a ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, new_AGEMA_signal_2655, SubCellInst_SboxInst_0_T1}), .b ({new_AGEMA_signal_5862, new_AGEMA_signal_5860, new_AGEMA_signal_5858, new_AGEMA_signal_5856}), .c ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, new_AGEMA_signal_2847, SubCellInst_SboxInst_0_L0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_AND4_U1 ( .a ({new_AGEMA_signal_5870, new_AGEMA_signal_5868, new_AGEMA_signal_5866, new_AGEMA_signal_5864}), .b ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, new_AGEMA_signal_2463, SubCellInst_SboxInst_0_Q7}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_2660, new_AGEMA_signal_2659, new_AGEMA_signal_2658, SubCellInst_SboxInst_0_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_XOR9_U1 ( .a ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, new_AGEMA_signal_2847, SubCellInst_SboxInst_0_L0}), .b ({new_AGEMA_signal_5886, new_AGEMA_signal_5882, new_AGEMA_signal_5878, new_AGEMA_signal_5874}), .c ({new_AGEMA_signal_2978, new_AGEMA_signal_2977, new_AGEMA_signal_2976, SubCellInst_SboxInst_0_YY_3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_XOR10_U1 ( .a ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, new_AGEMA_signal_2847, SubCellInst_SboxInst_0_L0}), .b ({new_AGEMA_signal_2660, new_AGEMA_signal_2659, new_AGEMA_signal_2658, SubCellInst_SboxInst_0_T3}), .c ({new_AGEMA_signal_2981, new_AGEMA_signal_2980, new_AGEMA_signal_2979, ShiftRowsOutput[4]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_0_XOR_o1_U1 ( .a ({new_AGEMA_signal_5894, new_AGEMA_signal_5892, new_AGEMA_signal_5890, new_AGEMA_signal_5888}), .b ({new_AGEMA_signal_2978, new_AGEMA_signal_2977, new_AGEMA_signal_2976, SubCellInst_SboxInst_0_YY_3}), .c ({new_AGEMA_signal_3152, new_AGEMA_signal_3151, new_AGEMA_signal_3150, ShiftRowsOutput[5]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_AND2_U1 ( .a ({new_AGEMA_signal_5902, new_AGEMA_signal_5900, new_AGEMA_signal_5898, new_AGEMA_signal_5896}), .b ({new_AGEMA_signal_2474, new_AGEMA_signal_2473, new_AGEMA_signal_2472, SubCellInst_SboxInst_1_Q2}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, new_AGEMA_signal_2667, SubCellInst_SboxInst_1_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_XOR4_U1 ( .a ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, new_AGEMA_signal_2667, SubCellInst_SboxInst_1_T1}), .b ({new_AGEMA_signal_5910, new_AGEMA_signal_5908, new_AGEMA_signal_5906, new_AGEMA_signal_5904}), .c ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, new_AGEMA_signal_2853, SubCellInst_SboxInst_1_L0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_AND4_U1 ( .a ({new_AGEMA_signal_5918, new_AGEMA_signal_5916, new_AGEMA_signal_5914, new_AGEMA_signal_5912}), .b ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, new_AGEMA_signal_2475, SubCellInst_SboxInst_1_Q7}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_2672, new_AGEMA_signal_2671, new_AGEMA_signal_2670, SubCellInst_SboxInst_1_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_XOR9_U1 ( .a ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, new_AGEMA_signal_2853, SubCellInst_SboxInst_1_L0}), .b ({new_AGEMA_signal_5934, new_AGEMA_signal_5930, new_AGEMA_signal_5926, new_AGEMA_signal_5922}), .c ({new_AGEMA_signal_2984, new_AGEMA_signal_2983, new_AGEMA_signal_2982, SubCellInst_SboxInst_1_YY_3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_XOR10_U1 ( .a ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, new_AGEMA_signal_2853, SubCellInst_SboxInst_1_L0}), .b ({new_AGEMA_signal_2672, new_AGEMA_signal_2671, new_AGEMA_signal_2670, SubCellInst_SboxInst_1_T3}), .c ({new_AGEMA_signal_2987, new_AGEMA_signal_2986, new_AGEMA_signal_2985, ShiftRowsOutput[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_1_XOR_o1_U1 ( .a ({new_AGEMA_signal_5942, new_AGEMA_signal_5940, new_AGEMA_signal_5938, new_AGEMA_signal_5936}), .b ({new_AGEMA_signal_2984, new_AGEMA_signal_2983, new_AGEMA_signal_2982, SubCellInst_SboxInst_1_YY_3}), .c ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, new_AGEMA_signal_3153, ShiftRowsOutput[9]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_AND2_U1 ( .a ({new_AGEMA_signal_5950, new_AGEMA_signal_5948, new_AGEMA_signal_5946, new_AGEMA_signal_5944}), .b ({new_AGEMA_signal_2486, new_AGEMA_signal_2485, new_AGEMA_signal_2484, SubCellInst_SboxInst_2_Q2}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, new_AGEMA_signal_2679, SubCellInst_SboxInst_2_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_XOR4_U1 ( .a ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, new_AGEMA_signal_2679, SubCellInst_SboxInst_2_T1}), .b ({new_AGEMA_signal_5958, new_AGEMA_signal_5956, new_AGEMA_signal_5954, new_AGEMA_signal_5952}), .c ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, new_AGEMA_signal_2859, SubCellInst_SboxInst_2_L0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_AND4_U1 ( .a ({new_AGEMA_signal_5966, new_AGEMA_signal_5964, new_AGEMA_signal_5962, new_AGEMA_signal_5960}), .b ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, new_AGEMA_signal_2487, SubCellInst_SboxInst_2_Q7}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_2684, new_AGEMA_signal_2683, new_AGEMA_signal_2682, SubCellInst_SboxInst_2_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_XOR9_U1 ( .a ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, new_AGEMA_signal_2859, SubCellInst_SboxInst_2_L0}), .b ({new_AGEMA_signal_5982, new_AGEMA_signal_5978, new_AGEMA_signal_5974, new_AGEMA_signal_5970}), .c ({new_AGEMA_signal_2990, new_AGEMA_signal_2989, new_AGEMA_signal_2988, SubCellInst_SboxInst_2_YY_3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_XOR10_U1 ( .a ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, new_AGEMA_signal_2859, SubCellInst_SboxInst_2_L0}), .b ({new_AGEMA_signal_2684, new_AGEMA_signal_2683, new_AGEMA_signal_2682, SubCellInst_SboxInst_2_T3}), .c ({new_AGEMA_signal_2993, new_AGEMA_signal_2992, new_AGEMA_signal_2991, ShiftRowsOutput[12]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_2_XOR_o1_U1 ( .a ({new_AGEMA_signal_5990, new_AGEMA_signal_5988, new_AGEMA_signal_5986, new_AGEMA_signal_5984}), .b ({new_AGEMA_signal_2990, new_AGEMA_signal_2989, new_AGEMA_signal_2988, SubCellInst_SboxInst_2_YY_3}), .c ({new_AGEMA_signal_3158, new_AGEMA_signal_3157, new_AGEMA_signal_3156, ShiftRowsOutput[13]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_AND2_U1 ( .a ({new_AGEMA_signal_5998, new_AGEMA_signal_5996, new_AGEMA_signal_5994, new_AGEMA_signal_5992}), .b ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, new_AGEMA_signal_2496, SubCellInst_SboxInst_3_Q2}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, new_AGEMA_signal_2691, SubCellInst_SboxInst_3_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_XOR4_U1 ( .a ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, new_AGEMA_signal_2691, SubCellInst_SboxInst_3_T1}), .b ({new_AGEMA_signal_6006, new_AGEMA_signal_6004, new_AGEMA_signal_6002, new_AGEMA_signal_6000}), .c ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, new_AGEMA_signal_2865, SubCellInst_SboxInst_3_L0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_AND4_U1 ( .a ({new_AGEMA_signal_6014, new_AGEMA_signal_6012, new_AGEMA_signal_6010, new_AGEMA_signal_6008}), .b ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, new_AGEMA_signal_2499, SubCellInst_SboxInst_3_Q7}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_2696, new_AGEMA_signal_2695, new_AGEMA_signal_2694, SubCellInst_SboxInst_3_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_XOR9_U1 ( .a ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, new_AGEMA_signal_2865, SubCellInst_SboxInst_3_L0}), .b ({new_AGEMA_signal_6030, new_AGEMA_signal_6026, new_AGEMA_signal_6022, new_AGEMA_signal_6018}), .c ({new_AGEMA_signal_2996, new_AGEMA_signal_2995, new_AGEMA_signal_2994, SubCellInst_SboxInst_3_YY_3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_XOR10_U1 ( .a ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, new_AGEMA_signal_2865, SubCellInst_SboxInst_3_L0}), .b ({new_AGEMA_signal_2696, new_AGEMA_signal_2695, new_AGEMA_signal_2694, SubCellInst_SboxInst_3_T3}), .c ({new_AGEMA_signal_2999, new_AGEMA_signal_2998, new_AGEMA_signal_2997, ShiftRowsOutput[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_3_XOR_o1_U1 ( .a ({new_AGEMA_signal_6038, new_AGEMA_signal_6036, new_AGEMA_signal_6034, new_AGEMA_signal_6032}), .b ({new_AGEMA_signal_2996, new_AGEMA_signal_2995, new_AGEMA_signal_2994, SubCellInst_SboxInst_3_YY_3}), .c ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, new_AGEMA_signal_3159, ShiftRowsOutput[1]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_AND2_U1 ( .a ({new_AGEMA_signal_6046, new_AGEMA_signal_6044, new_AGEMA_signal_6042, new_AGEMA_signal_6040}), .b ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, new_AGEMA_signal_2508, SubCellInst_SboxInst_4_Q2}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, new_AGEMA_signal_2703, SubCellInst_SboxInst_4_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_XOR4_U1 ( .a ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, new_AGEMA_signal_2703, SubCellInst_SboxInst_4_T1}), .b ({new_AGEMA_signal_6054, new_AGEMA_signal_6052, new_AGEMA_signal_6050, new_AGEMA_signal_6048}), .c ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, new_AGEMA_signal_2871, SubCellInst_SboxInst_4_L0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_AND4_U1 ( .a ({new_AGEMA_signal_6062, new_AGEMA_signal_6060, new_AGEMA_signal_6058, new_AGEMA_signal_6056}), .b ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, new_AGEMA_signal_2511, SubCellInst_SboxInst_4_Q7}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_2708, new_AGEMA_signal_2707, new_AGEMA_signal_2706, SubCellInst_SboxInst_4_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_XOR9_U1 ( .a ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, new_AGEMA_signal_2871, SubCellInst_SboxInst_4_L0}), .b ({new_AGEMA_signal_6078, new_AGEMA_signal_6074, new_AGEMA_signal_6070, new_AGEMA_signal_6066}), .c ({new_AGEMA_signal_3002, new_AGEMA_signal_3001, new_AGEMA_signal_3000, SubCellInst_SboxInst_4_YY_3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_XOR10_U1 ( .a ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, new_AGEMA_signal_2871, SubCellInst_SboxInst_4_L0}), .b ({new_AGEMA_signal_2708, new_AGEMA_signal_2707, new_AGEMA_signal_2706, SubCellInst_SboxInst_4_T3}), .c ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, new_AGEMA_signal_3003, ShiftRowsOutput[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_4_XOR_o1_U1 ( .a ({new_AGEMA_signal_6086, new_AGEMA_signal_6084, new_AGEMA_signal_6082, new_AGEMA_signal_6080}), .b ({new_AGEMA_signal_3002, new_AGEMA_signal_3001, new_AGEMA_signal_3000, SubCellInst_SboxInst_4_YY_3}), .c ({new_AGEMA_signal_3164, new_AGEMA_signal_3163, new_AGEMA_signal_3162, ShiftRowsOutput[25]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_AND2_U1 ( .a ({new_AGEMA_signal_6094, new_AGEMA_signal_6092, new_AGEMA_signal_6090, new_AGEMA_signal_6088}), .b ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, new_AGEMA_signal_2520, SubCellInst_SboxInst_5_Q2}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, new_AGEMA_signal_2715, SubCellInst_SboxInst_5_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_XOR4_U1 ( .a ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, new_AGEMA_signal_2715, SubCellInst_SboxInst_5_T1}), .b ({new_AGEMA_signal_6102, new_AGEMA_signal_6100, new_AGEMA_signal_6098, new_AGEMA_signal_6096}), .c ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, new_AGEMA_signal_2877, SubCellInst_SboxInst_5_L0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_AND4_U1 ( .a ({new_AGEMA_signal_6110, new_AGEMA_signal_6108, new_AGEMA_signal_6106, new_AGEMA_signal_6104}), .b ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, new_AGEMA_signal_2523, SubCellInst_SboxInst_5_Q7}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_2720, new_AGEMA_signal_2719, new_AGEMA_signal_2718, SubCellInst_SboxInst_5_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_XOR9_U1 ( .a ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, new_AGEMA_signal_2877, SubCellInst_SboxInst_5_L0}), .b ({new_AGEMA_signal_6126, new_AGEMA_signal_6122, new_AGEMA_signal_6118, new_AGEMA_signal_6114}), .c ({new_AGEMA_signal_3008, new_AGEMA_signal_3007, new_AGEMA_signal_3006, SubCellInst_SboxInst_5_YY_3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_XOR10_U1 ( .a ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, new_AGEMA_signal_2877, SubCellInst_SboxInst_5_L0}), .b ({new_AGEMA_signal_2720, new_AGEMA_signal_2719, new_AGEMA_signal_2718, SubCellInst_SboxInst_5_T3}), .c ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, new_AGEMA_signal_3009, ShiftRowsOutput[28]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_5_XOR_o1_U1 ( .a ({new_AGEMA_signal_6134, new_AGEMA_signal_6132, new_AGEMA_signal_6130, new_AGEMA_signal_6128}), .b ({new_AGEMA_signal_3008, new_AGEMA_signal_3007, new_AGEMA_signal_3006, SubCellInst_SboxInst_5_YY_3}), .c ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, new_AGEMA_signal_3165, ShiftRowsOutput[29]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_AND2_U1 ( .a ({new_AGEMA_signal_6142, new_AGEMA_signal_6140, new_AGEMA_signal_6138, new_AGEMA_signal_6136}), .b ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, new_AGEMA_signal_2532, SubCellInst_SboxInst_6_Q2}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, new_AGEMA_signal_2727, SubCellInst_SboxInst_6_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_XOR4_U1 ( .a ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, new_AGEMA_signal_2727, SubCellInst_SboxInst_6_T1}), .b ({new_AGEMA_signal_6150, new_AGEMA_signal_6148, new_AGEMA_signal_6146, new_AGEMA_signal_6144}), .c ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, new_AGEMA_signal_2883, SubCellInst_SboxInst_6_L0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_AND4_U1 ( .a ({new_AGEMA_signal_6158, new_AGEMA_signal_6156, new_AGEMA_signal_6154, new_AGEMA_signal_6152}), .b ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, new_AGEMA_signal_2535, SubCellInst_SboxInst_6_Q7}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_2732, new_AGEMA_signal_2731, new_AGEMA_signal_2730, SubCellInst_SboxInst_6_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_XOR9_U1 ( .a ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, new_AGEMA_signal_2883, SubCellInst_SboxInst_6_L0}), .b ({new_AGEMA_signal_6174, new_AGEMA_signal_6170, new_AGEMA_signal_6166, new_AGEMA_signal_6162}), .c ({new_AGEMA_signal_3014, new_AGEMA_signal_3013, new_AGEMA_signal_3012, SubCellInst_SboxInst_6_YY_3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_XOR10_U1 ( .a ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, new_AGEMA_signal_2883, SubCellInst_SboxInst_6_L0}), .b ({new_AGEMA_signal_2732, new_AGEMA_signal_2731, new_AGEMA_signal_2730, SubCellInst_SboxInst_6_T3}), .c ({new_AGEMA_signal_3017, new_AGEMA_signal_3016, new_AGEMA_signal_3015, ShiftRowsOutput[16]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_6_XOR_o1_U1 ( .a ({new_AGEMA_signal_6182, new_AGEMA_signal_6180, new_AGEMA_signal_6178, new_AGEMA_signal_6176}), .b ({new_AGEMA_signal_3014, new_AGEMA_signal_3013, new_AGEMA_signal_3012, SubCellInst_SboxInst_6_YY_3}), .c ({new_AGEMA_signal_3170, new_AGEMA_signal_3169, new_AGEMA_signal_3168, ShiftRowsOutput[17]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_AND2_U1 ( .a ({new_AGEMA_signal_6190, new_AGEMA_signal_6188, new_AGEMA_signal_6186, new_AGEMA_signal_6184}), .b ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, new_AGEMA_signal_2544, SubCellInst_SboxInst_7_Q2}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, new_AGEMA_signal_2739, SubCellInst_SboxInst_7_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_XOR4_U1 ( .a ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, new_AGEMA_signal_2739, SubCellInst_SboxInst_7_T1}), .b ({new_AGEMA_signal_6198, new_AGEMA_signal_6196, new_AGEMA_signal_6194, new_AGEMA_signal_6192}), .c ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, new_AGEMA_signal_2889, SubCellInst_SboxInst_7_L0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_AND4_U1 ( .a ({new_AGEMA_signal_6206, new_AGEMA_signal_6204, new_AGEMA_signal_6202, new_AGEMA_signal_6200}), .b ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, new_AGEMA_signal_2547, SubCellInst_SboxInst_7_Q7}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_2744, new_AGEMA_signal_2743, new_AGEMA_signal_2742, SubCellInst_SboxInst_7_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_XOR9_U1 ( .a ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, new_AGEMA_signal_2889, SubCellInst_SboxInst_7_L0}), .b ({new_AGEMA_signal_6222, new_AGEMA_signal_6218, new_AGEMA_signal_6214, new_AGEMA_signal_6210}), .c ({new_AGEMA_signal_3020, new_AGEMA_signal_3019, new_AGEMA_signal_3018, SubCellInst_SboxInst_7_YY_3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_XOR10_U1 ( .a ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, new_AGEMA_signal_2889, SubCellInst_SboxInst_7_L0}), .b ({new_AGEMA_signal_2744, new_AGEMA_signal_2743, new_AGEMA_signal_2742, SubCellInst_SboxInst_7_T3}), .c ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, new_AGEMA_signal_3021, ShiftRowsOutput[20]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_7_XOR_o1_U1 ( .a ({new_AGEMA_signal_6230, new_AGEMA_signal_6228, new_AGEMA_signal_6226, new_AGEMA_signal_6224}), .b ({new_AGEMA_signal_3020, new_AGEMA_signal_3019, new_AGEMA_signal_3018, SubCellInst_SboxInst_7_YY_3}), .c ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, new_AGEMA_signal_3171, SubCellOutput[29]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_AND2_U1 ( .a ({new_AGEMA_signal_6238, new_AGEMA_signal_6236, new_AGEMA_signal_6234, new_AGEMA_signal_6232}), .b ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, new_AGEMA_signal_2556, SubCellInst_SboxInst_8_Q2}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, new_AGEMA_signal_2751, SubCellInst_SboxInst_8_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_XOR4_U1 ( .a ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, new_AGEMA_signal_2751, SubCellInst_SboxInst_8_T1}), .b ({new_AGEMA_signal_6246, new_AGEMA_signal_6244, new_AGEMA_signal_6242, new_AGEMA_signal_6240}), .c ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, new_AGEMA_signal_2895, SubCellInst_SboxInst_8_L0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_AND4_U1 ( .a ({new_AGEMA_signal_6254, new_AGEMA_signal_6252, new_AGEMA_signal_6250, new_AGEMA_signal_6248}), .b ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, new_AGEMA_signal_2559, SubCellInst_SboxInst_8_Q7}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, new_AGEMA_signal_2754, SubCellInst_SboxInst_8_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_XOR9_U1 ( .a ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, new_AGEMA_signal_2895, SubCellInst_SboxInst_8_L0}), .b ({new_AGEMA_signal_6270, new_AGEMA_signal_6266, new_AGEMA_signal_6262, new_AGEMA_signal_6258}), .c ({new_AGEMA_signal_3026, new_AGEMA_signal_3025, new_AGEMA_signal_3024, SubCellInst_SboxInst_8_YY_3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_XOR10_U1 ( .a ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, new_AGEMA_signal_2895, SubCellInst_SboxInst_8_L0}), .b ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, new_AGEMA_signal_2754, SubCellInst_SboxInst_8_T3}), .c ({new_AGEMA_signal_3029, new_AGEMA_signal_3028, new_AGEMA_signal_3027, AddRoundConstantOutput[32]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_8_XOR_o1_U1 ( .a ({new_AGEMA_signal_6278, new_AGEMA_signal_6276, new_AGEMA_signal_6274, new_AGEMA_signal_6272}), .b ({new_AGEMA_signal_3026, new_AGEMA_signal_3025, new_AGEMA_signal_3024, SubCellInst_SboxInst_8_YY_3}), .c ({new_AGEMA_signal_3176, new_AGEMA_signal_3175, new_AGEMA_signal_3174, AddRoundConstantOutput[33]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_AND2_U1 ( .a ({new_AGEMA_signal_6286, new_AGEMA_signal_6284, new_AGEMA_signal_6282, new_AGEMA_signal_6280}), .b ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, new_AGEMA_signal_2568, SubCellInst_SboxInst_9_Q2}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, new_AGEMA_signal_2763, SubCellInst_SboxInst_9_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_XOR4_U1 ( .a ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, new_AGEMA_signal_2763, SubCellInst_SboxInst_9_T1}), .b ({new_AGEMA_signal_6294, new_AGEMA_signal_6292, new_AGEMA_signal_6290, new_AGEMA_signal_6288}), .c ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, new_AGEMA_signal_2901, SubCellInst_SboxInst_9_L0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_AND4_U1 ( .a ({new_AGEMA_signal_6302, new_AGEMA_signal_6300, new_AGEMA_signal_6298, new_AGEMA_signal_6296}), .b ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, new_AGEMA_signal_2571, SubCellInst_SboxInst_9_Q7}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, new_AGEMA_signal_2766, SubCellInst_SboxInst_9_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_XOR9_U1 ( .a ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, new_AGEMA_signal_2901, SubCellInst_SboxInst_9_L0}), .b ({new_AGEMA_signal_6318, new_AGEMA_signal_6314, new_AGEMA_signal_6310, new_AGEMA_signal_6306}), .c ({new_AGEMA_signal_3032, new_AGEMA_signal_3031, new_AGEMA_signal_3030, SubCellInst_SboxInst_9_YY_3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_XOR10_U1 ( .a ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, new_AGEMA_signal_2901, SubCellInst_SboxInst_9_L0}), .b ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, new_AGEMA_signal_2766, SubCellInst_SboxInst_9_T3}), .c ({new_AGEMA_signal_3035, new_AGEMA_signal_3034, new_AGEMA_signal_3033, AddRoundConstantOutput[36]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_9_XOR_o1_U1 ( .a ({new_AGEMA_signal_6326, new_AGEMA_signal_6324, new_AGEMA_signal_6322, new_AGEMA_signal_6320}), .b ({new_AGEMA_signal_3032, new_AGEMA_signal_3031, new_AGEMA_signal_3030, SubCellInst_SboxInst_9_YY_3}), .c ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, new_AGEMA_signal_3177, AddRoundConstantOutput[37]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_AND2_U1 ( .a ({new_AGEMA_signal_6334, new_AGEMA_signal_6332, new_AGEMA_signal_6330, new_AGEMA_signal_6328}), .b ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, new_AGEMA_signal_2580, SubCellInst_SboxInst_10_Q2}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, new_AGEMA_signal_2775, SubCellInst_SboxInst_10_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_XOR4_U1 ( .a ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, new_AGEMA_signal_2775, SubCellInst_SboxInst_10_T1}), .b ({new_AGEMA_signal_6342, new_AGEMA_signal_6340, new_AGEMA_signal_6338, new_AGEMA_signal_6336}), .c ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, new_AGEMA_signal_2907, SubCellInst_SboxInst_10_L0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_AND4_U1 ( .a ({new_AGEMA_signal_6350, new_AGEMA_signal_6348, new_AGEMA_signal_6346, new_AGEMA_signal_6344}), .b ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, new_AGEMA_signal_2583, SubCellInst_SboxInst_10_Q7}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, new_AGEMA_signal_2778, SubCellInst_SboxInst_10_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_XOR9_U1 ( .a ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, new_AGEMA_signal_2907, SubCellInst_SboxInst_10_L0}), .b ({new_AGEMA_signal_6366, new_AGEMA_signal_6362, new_AGEMA_signal_6358, new_AGEMA_signal_6354}), .c ({new_AGEMA_signal_3038, new_AGEMA_signal_3037, new_AGEMA_signal_3036, SubCellInst_SboxInst_10_YY_3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_XOR10_U1 ( .a ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, new_AGEMA_signal_2907, SubCellInst_SboxInst_10_L0}), .b ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, new_AGEMA_signal_2778, SubCellInst_SboxInst_10_T3}), .c ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, new_AGEMA_signal_3039, AddRoundConstantOutput[40]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_10_XOR_o1_U1 ( .a ({new_AGEMA_signal_6374, new_AGEMA_signal_6372, new_AGEMA_signal_6370, new_AGEMA_signal_6368}), .b ({new_AGEMA_signal_3038, new_AGEMA_signal_3037, new_AGEMA_signal_3036, SubCellInst_SboxInst_10_YY_3}), .c ({new_AGEMA_signal_3182, new_AGEMA_signal_3181, new_AGEMA_signal_3180, AddRoundConstantOutput[41]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_AND2_U1 ( .a ({new_AGEMA_signal_6382, new_AGEMA_signal_6380, new_AGEMA_signal_6378, new_AGEMA_signal_6376}), .b ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, new_AGEMA_signal_2592, SubCellInst_SboxInst_11_Q2}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, new_AGEMA_signal_2787, SubCellInst_SboxInst_11_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_XOR4_U1 ( .a ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, new_AGEMA_signal_2787, SubCellInst_SboxInst_11_T1}), .b ({new_AGEMA_signal_6390, new_AGEMA_signal_6388, new_AGEMA_signal_6386, new_AGEMA_signal_6384}), .c ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, new_AGEMA_signal_2913, SubCellInst_SboxInst_11_L0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_AND4_U1 ( .a ({new_AGEMA_signal_6398, new_AGEMA_signal_6396, new_AGEMA_signal_6394, new_AGEMA_signal_6392}), .b ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, new_AGEMA_signal_2595, SubCellInst_SboxInst_11_Q7}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, new_AGEMA_signal_2790, SubCellInst_SboxInst_11_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_XOR9_U1 ( .a ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, new_AGEMA_signal_2913, SubCellInst_SboxInst_11_L0}), .b ({new_AGEMA_signal_6414, new_AGEMA_signal_6410, new_AGEMA_signal_6406, new_AGEMA_signal_6402}), .c ({new_AGEMA_signal_3044, new_AGEMA_signal_3043, new_AGEMA_signal_3042, SubCellInst_SboxInst_11_YY_3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_XOR10_U1 ( .a ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, new_AGEMA_signal_2913, SubCellInst_SboxInst_11_L0}), .b ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, new_AGEMA_signal_2790, SubCellInst_SboxInst_11_T3}), .c ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, new_AGEMA_signal_3045, SubCellOutput[44]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_11_XOR_o1_U1 ( .a ({new_AGEMA_signal_6422, new_AGEMA_signal_6420, new_AGEMA_signal_6418, new_AGEMA_signal_6416}), .b ({new_AGEMA_signal_3044, new_AGEMA_signal_3043, new_AGEMA_signal_3042, SubCellInst_SboxInst_11_YY_3}), .c ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, new_AGEMA_signal_3183, SubCellOutput[45]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_AND2_U1 ( .a ({new_AGEMA_signal_6430, new_AGEMA_signal_6428, new_AGEMA_signal_6426, new_AGEMA_signal_6424}), .b ({new_AGEMA_signal_2606, new_AGEMA_signal_2605, new_AGEMA_signal_2604, SubCellInst_SboxInst_12_Q2}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, new_AGEMA_signal_2799, SubCellInst_SboxInst_12_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_XOR4_U1 ( .a ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, new_AGEMA_signal_2799, SubCellInst_SboxInst_12_T1}), .b ({new_AGEMA_signal_6438, new_AGEMA_signal_6436, new_AGEMA_signal_6434, new_AGEMA_signal_6432}), .c ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, new_AGEMA_signal_2919, SubCellInst_SboxInst_12_L0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_AND4_U1 ( .a ({new_AGEMA_signal_6446, new_AGEMA_signal_6444, new_AGEMA_signal_6442, new_AGEMA_signal_6440}), .b ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, new_AGEMA_signal_2607, SubCellInst_SboxInst_12_Q7}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_2804, new_AGEMA_signal_2803, new_AGEMA_signal_2802, SubCellInst_SboxInst_12_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_XOR9_U1 ( .a ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, new_AGEMA_signal_2919, SubCellInst_SboxInst_12_L0}), .b ({new_AGEMA_signal_6462, new_AGEMA_signal_6458, new_AGEMA_signal_6454, new_AGEMA_signal_6450}), .c ({new_AGEMA_signal_3050, new_AGEMA_signal_3049, new_AGEMA_signal_3048, SubCellInst_SboxInst_12_YY_3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_XOR10_U1 ( .a ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, new_AGEMA_signal_2919, SubCellInst_SboxInst_12_L0}), .b ({new_AGEMA_signal_2804, new_AGEMA_signal_2803, new_AGEMA_signal_2802, SubCellInst_SboxInst_12_T3}), .c ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, new_AGEMA_signal_3051, AddRoundConstantOutput[48]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_12_XOR_o1_U1 ( .a ({new_AGEMA_signal_6470, new_AGEMA_signal_6468, new_AGEMA_signal_6466, new_AGEMA_signal_6464}), .b ({new_AGEMA_signal_3050, new_AGEMA_signal_3049, new_AGEMA_signal_3048, SubCellInst_SboxInst_12_YY_3}), .c ({new_AGEMA_signal_3188, new_AGEMA_signal_3187, new_AGEMA_signal_3186, AddRoundConstantOutput[49]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_AND2_U1 ( .a ({new_AGEMA_signal_6478, new_AGEMA_signal_6476, new_AGEMA_signal_6474, new_AGEMA_signal_6472}), .b ({new_AGEMA_signal_2618, new_AGEMA_signal_2617, new_AGEMA_signal_2616, SubCellInst_SboxInst_13_Q2}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, new_AGEMA_signal_2811, SubCellInst_SboxInst_13_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_XOR4_U1 ( .a ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, new_AGEMA_signal_2811, SubCellInst_SboxInst_13_T1}), .b ({new_AGEMA_signal_6486, new_AGEMA_signal_6484, new_AGEMA_signal_6482, new_AGEMA_signal_6480}), .c ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, new_AGEMA_signal_2925, SubCellInst_SboxInst_13_L0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_AND4_U1 ( .a ({new_AGEMA_signal_6494, new_AGEMA_signal_6492, new_AGEMA_signal_6490, new_AGEMA_signal_6488}), .b ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, new_AGEMA_signal_2619, SubCellInst_SboxInst_13_Q7}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_2816, new_AGEMA_signal_2815, new_AGEMA_signal_2814, SubCellInst_SboxInst_13_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_XOR9_U1 ( .a ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, new_AGEMA_signal_2925, SubCellInst_SboxInst_13_L0}), .b ({new_AGEMA_signal_6510, new_AGEMA_signal_6506, new_AGEMA_signal_6502, new_AGEMA_signal_6498}), .c ({new_AGEMA_signal_3056, new_AGEMA_signal_3055, new_AGEMA_signal_3054, SubCellInst_SboxInst_13_YY_3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_XOR10_U1 ( .a ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, new_AGEMA_signal_2925, SubCellInst_SboxInst_13_L0}), .b ({new_AGEMA_signal_2816, new_AGEMA_signal_2815, new_AGEMA_signal_2814, SubCellInst_SboxInst_13_T3}), .c ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, new_AGEMA_signal_3057, AddRoundConstantOutput[52]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_13_XOR_o1_U1 ( .a ({new_AGEMA_signal_6518, new_AGEMA_signal_6516, new_AGEMA_signal_6514, new_AGEMA_signal_6512}), .b ({new_AGEMA_signal_3056, new_AGEMA_signal_3055, new_AGEMA_signal_3054, SubCellInst_SboxInst_13_YY_3}), .c ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, new_AGEMA_signal_3189, AddRoundConstantOutput[53]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_AND2_U1 ( .a ({new_AGEMA_signal_6526, new_AGEMA_signal_6524, new_AGEMA_signal_6522, new_AGEMA_signal_6520}), .b ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, new_AGEMA_signal_2628, SubCellInst_SboxInst_14_Q2}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, new_AGEMA_signal_2823, SubCellInst_SboxInst_14_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_XOR4_U1 ( .a ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, new_AGEMA_signal_2823, SubCellInst_SboxInst_14_T1}), .b ({new_AGEMA_signal_6534, new_AGEMA_signal_6532, new_AGEMA_signal_6530, new_AGEMA_signal_6528}), .c ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, new_AGEMA_signal_2931, SubCellInst_SboxInst_14_L0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_AND4_U1 ( .a ({new_AGEMA_signal_6542, new_AGEMA_signal_6540, new_AGEMA_signal_6538, new_AGEMA_signal_6536}), .b ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, new_AGEMA_signal_2631, SubCellInst_SboxInst_14_Q7}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_2828, new_AGEMA_signal_2827, new_AGEMA_signal_2826, SubCellInst_SboxInst_14_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_XOR9_U1 ( .a ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, new_AGEMA_signal_2931, SubCellInst_SboxInst_14_L0}), .b ({new_AGEMA_signal_6558, new_AGEMA_signal_6554, new_AGEMA_signal_6550, new_AGEMA_signal_6546}), .c ({new_AGEMA_signal_3062, new_AGEMA_signal_3061, new_AGEMA_signal_3060, SubCellInst_SboxInst_14_YY_3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_XOR10_U1 ( .a ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, new_AGEMA_signal_2931, SubCellInst_SboxInst_14_L0}), .b ({new_AGEMA_signal_2828, new_AGEMA_signal_2827, new_AGEMA_signal_2826, SubCellInst_SboxInst_14_T3}), .c ({new_AGEMA_signal_3065, new_AGEMA_signal_3064, new_AGEMA_signal_3063, AddRoundConstantOutput[56]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_14_XOR_o1_U1 ( .a ({new_AGEMA_signal_6566, new_AGEMA_signal_6564, new_AGEMA_signal_6562, new_AGEMA_signal_6560}), .b ({new_AGEMA_signal_3062, new_AGEMA_signal_3061, new_AGEMA_signal_3060, SubCellInst_SboxInst_14_YY_3}), .c ({new_AGEMA_signal_3194, new_AGEMA_signal_3193, new_AGEMA_signal_3192, AddRoundConstantOutput[57]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_AND2_U1 ( .a ({new_AGEMA_signal_6574, new_AGEMA_signal_6572, new_AGEMA_signal_6570, new_AGEMA_signal_6568}), .b ({new_AGEMA_signal_2642, new_AGEMA_signal_2641, new_AGEMA_signal_2640, SubCellInst_SboxInst_15_Q2}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, new_AGEMA_signal_2835, SubCellInst_SboxInst_15_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_XOR4_U1 ( .a ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, new_AGEMA_signal_2835, SubCellInst_SboxInst_15_T1}), .b ({new_AGEMA_signal_6582, new_AGEMA_signal_6580, new_AGEMA_signal_6578, new_AGEMA_signal_6576}), .c ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, new_AGEMA_signal_2937, SubCellInst_SboxInst_15_L0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_AND4_U1 ( .a ({new_AGEMA_signal_6590, new_AGEMA_signal_6588, new_AGEMA_signal_6586, new_AGEMA_signal_6584}), .b ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, new_AGEMA_signal_2643, SubCellInst_SboxInst_15_Q7}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_2840, new_AGEMA_signal_2839, new_AGEMA_signal_2838, SubCellInst_SboxInst_15_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_XOR9_U1 ( .a ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, new_AGEMA_signal_2937, SubCellInst_SboxInst_15_L0}), .b ({new_AGEMA_signal_6606, new_AGEMA_signal_6602, new_AGEMA_signal_6598, new_AGEMA_signal_6594}), .c ({new_AGEMA_signal_3068, new_AGEMA_signal_3067, new_AGEMA_signal_3066, SubCellInst_SboxInst_15_YY_3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_XOR10_U1 ( .a ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, new_AGEMA_signal_2937, SubCellInst_SboxInst_15_L0}), .b ({new_AGEMA_signal_2840, new_AGEMA_signal_2839, new_AGEMA_signal_2838, SubCellInst_SboxInst_15_T3}), .c ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, new_AGEMA_signal_3069, SubCellOutput[60]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) SubCellInst_SboxInst_15_XOR_o1_U1 ( .a ({new_AGEMA_signal_6614, new_AGEMA_signal_6612, new_AGEMA_signal_6610, new_AGEMA_signal_6608}), .b ({new_AGEMA_signal_3068, new_AGEMA_signal_3067, new_AGEMA_signal_3066, SubCellInst_SboxInst_15_YY_3}), .c ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, new_AGEMA_signal_3195, SubCellOutput[61]}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) AddConstXOR_U2 ( .a ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, new_AGEMA_signal_3171, SubCellOutput[29]}), .b ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, new_AGEMA_signal_3309, ShiftRowsOutput[21]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_3200, new_AGEMA_signal_3199, new_AGEMA_signal_3198, AddConstXOR_AddConstXOR_XORInst_0_0_n1}), .b ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_6618}), .c ({new_AGEMA_signal_3314, new_AGEMA_signal_3313, new_AGEMA_signal_3312, AddRoundConstantOutput[60]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, new_AGEMA_signal_3069, SubCellOutput[60]}), .c ({new_AGEMA_signal_3200, new_AGEMA_signal_3199, new_AGEMA_signal_3198, AddConstXOR_AddConstXOR_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, new_AGEMA_signal_3315, AddConstXOR_AddConstXOR_XORInst_0_1_n1}), .b ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_6622}), .c ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, new_AGEMA_signal_3513, AddRoundConstantOutput[61]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, new_AGEMA_signal_3195, SubCellOutput[61]}), .c ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, new_AGEMA_signal_3315, AddConstXOR_AddConstXOR_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_3206, new_AGEMA_signal_3205, new_AGEMA_signal_3204, AddConstXOR_AddConstXOR_XORInst_1_0_n1}), .b ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_6626}), .c ({new_AGEMA_signal_3320, new_AGEMA_signal_3319, new_AGEMA_signal_3318, AddRoundConstantOutput[44]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, new_AGEMA_signal_3045, SubCellOutput[44]}), .c ({new_AGEMA_signal_3206, new_AGEMA_signal_3205, new_AGEMA_signal_3204, AddConstXOR_AddConstXOR_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, new_AGEMA_signal_3321, AddConstXOR_AddConstXOR_XORInst_1_1_n1}), .b ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_6630}), .c ({new_AGEMA_signal_3518, new_AGEMA_signal_3517, new_AGEMA_signal_3516, AddRoundConstantOutput[45]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, new_AGEMA_signal_3183, SubCellOutput[45]}), .c ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, new_AGEMA_signal_3321, AddConstXOR_AddConstXOR_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_3212, new_AGEMA_signal_3211, new_AGEMA_signal_3210, AddRoundTweakeyXOR_XORInst_0_0_n1}), .b ({new_AGEMA_signal_6646, new_AGEMA_signal_6642, new_AGEMA_signal_6638, new_AGEMA_signal_6634}), .c ({new_AGEMA_signal_3326, new_AGEMA_signal_3325, new_AGEMA_signal_3324, ShiftRowsOutput[44]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3029, new_AGEMA_signal_3028, new_AGEMA_signal_3027, AddRoundConstantOutput[32]}), .c ({new_AGEMA_signal_3212, new_AGEMA_signal_3211, new_AGEMA_signal_3210, AddRoundTweakeyXOR_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, new_AGEMA_signal_3327, AddRoundTweakeyXOR_XORInst_0_1_n1}), .b ({new_AGEMA_signal_6662, new_AGEMA_signal_6658, new_AGEMA_signal_6654, new_AGEMA_signal_6650}), .c ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, new_AGEMA_signal_3519, ShiftRowsOutput[45]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3176, new_AGEMA_signal_3175, new_AGEMA_signal_3174, AddRoundConstantOutput[33]}), .c ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, new_AGEMA_signal_3327, AddRoundTweakeyXOR_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_3218, new_AGEMA_signal_3217, new_AGEMA_signal_3216, AddRoundTweakeyXOR_XORInst_1_0_n1}), .b ({new_AGEMA_signal_6678, new_AGEMA_signal_6674, new_AGEMA_signal_6670, new_AGEMA_signal_6666}), .c ({new_AGEMA_signal_3332, new_AGEMA_signal_3331, new_AGEMA_signal_3330, ShiftRowsOutput[32]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3035, new_AGEMA_signal_3034, new_AGEMA_signal_3033, AddRoundConstantOutput[36]}), .c ({new_AGEMA_signal_3218, new_AGEMA_signal_3217, new_AGEMA_signal_3216, AddRoundTweakeyXOR_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, new_AGEMA_signal_3333, AddRoundTweakeyXOR_XORInst_1_1_n1}), .b ({new_AGEMA_signal_6694, new_AGEMA_signal_6690, new_AGEMA_signal_6686, new_AGEMA_signal_6682}), .c ({new_AGEMA_signal_3524, new_AGEMA_signal_3523, new_AGEMA_signal_3522, ShiftRowsOutput[33]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, new_AGEMA_signal_3177, AddRoundConstantOutput[37]}), .c ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, new_AGEMA_signal_3333, AddRoundTweakeyXOR_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_3224, new_AGEMA_signal_3223, new_AGEMA_signal_3222, AddRoundTweakeyXOR_XORInst_2_0_n1}), .b ({new_AGEMA_signal_6710, new_AGEMA_signal_6706, new_AGEMA_signal_6702, new_AGEMA_signal_6698}), .c ({new_AGEMA_signal_3338, new_AGEMA_signal_3337, new_AGEMA_signal_3336, ShiftRowsOutput[36]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, new_AGEMA_signal_3039, AddRoundConstantOutput[40]}), .c ({new_AGEMA_signal_3224, new_AGEMA_signal_3223, new_AGEMA_signal_3222, AddRoundTweakeyXOR_XORInst_2_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, new_AGEMA_signal_3339, AddRoundTweakeyXOR_XORInst_2_1_n1}), .b ({new_AGEMA_signal_6726, new_AGEMA_signal_6722, new_AGEMA_signal_6718, new_AGEMA_signal_6714}), .c ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, new_AGEMA_signal_3525, ShiftRowsOutput[37]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3182, new_AGEMA_signal_3181, new_AGEMA_signal_3180, AddRoundConstantOutput[41]}), .c ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, new_AGEMA_signal_3339, AddRoundTweakeyXOR_XORInst_2_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_3530, new_AGEMA_signal_3529, new_AGEMA_signal_3528, AddRoundTweakeyXOR_XORInst_3_0_n1}), .b ({new_AGEMA_signal_6742, new_AGEMA_signal_6738, new_AGEMA_signal_6734, new_AGEMA_signal_6730}), .c ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, new_AGEMA_signal_3693, ShiftRowsOutput[40]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3320, new_AGEMA_signal_3319, new_AGEMA_signal_3318, AddRoundConstantOutput[44]}), .c ({new_AGEMA_signal_3530, new_AGEMA_signal_3529, new_AGEMA_signal_3528, AddRoundTweakeyXOR_XORInst_3_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_3698, new_AGEMA_signal_3697, new_AGEMA_signal_3696, AddRoundTweakeyXOR_XORInst_3_1_n1}), .b ({new_AGEMA_signal_6758, new_AGEMA_signal_6754, new_AGEMA_signal_6750, new_AGEMA_signal_6746}), .c ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, new_AGEMA_signal_3855, ShiftRowsOutput[41]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3518, new_AGEMA_signal_3517, new_AGEMA_signal_3516, AddRoundConstantOutput[45]}), .c ({new_AGEMA_signal_3698, new_AGEMA_signal_3697, new_AGEMA_signal_3696, AddRoundTweakeyXOR_XORInst_3_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_4_0_U2 ( .a ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, new_AGEMA_signal_3231, AddRoundTweakeyXOR_XORInst_4_0_n1}), .b ({new_AGEMA_signal_6774, new_AGEMA_signal_6770, new_AGEMA_signal_6766, new_AGEMA_signal_6762}), .c ({new_AGEMA_signal_3350, new_AGEMA_signal_3349, new_AGEMA_signal_3348, MCOutput[32]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_4_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, new_AGEMA_signal_3051, AddRoundConstantOutput[48]}), .c ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, new_AGEMA_signal_3231, AddRoundTweakeyXOR_XORInst_4_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_4_1_U2 ( .a ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, new_AGEMA_signal_3351, AddRoundTweakeyXOR_XORInst_4_1_n1}), .b ({new_AGEMA_signal_6790, new_AGEMA_signal_6786, new_AGEMA_signal_6782, new_AGEMA_signal_6778}), .c ({new_AGEMA_signal_3536, new_AGEMA_signal_3535, new_AGEMA_signal_3534, MCOutput[33]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_4_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3188, new_AGEMA_signal_3187, new_AGEMA_signal_3186, AddRoundConstantOutput[49]}), .c ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, new_AGEMA_signal_3351, AddRoundTweakeyXOR_XORInst_4_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_5_0_U2 ( .a ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, new_AGEMA_signal_3237, AddRoundTweakeyXOR_XORInst_5_0_n1}), .b ({new_AGEMA_signal_6806, new_AGEMA_signal_6802, new_AGEMA_signal_6798, new_AGEMA_signal_6794}), .c ({new_AGEMA_signal_3356, new_AGEMA_signal_3355, new_AGEMA_signal_3354, MCOutput[36]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_5_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, new_AGEMA_signal_3057, AddRoundConstantOutput[52]}), .c ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, new_AGEMA_signal_3237, AddRoundTweakeyXOR_XORInst_5_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_5_1_U2 ( .a ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, new_AGEMA_signal_3357, AddRoundTweakeyXOR_XORInst_5_1_n1}), .b ({new_AGEMA_signal_6822, new_AGEMA_signal_6818, new_AGEMA_signal_6814, new_AGEMA_signal_6810}), .c ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, new_AGEMA_signal_3537, MCOutput[37]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_5_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, new_AGEMA_signal_3189, AddRoundConstantOutput[53]}), .c ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, new_AGEMA_signal_3357, AddRoundTweakeyXOR_XORInst_5_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_6_0_U2 ( .a ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, new_AGEMA_signal_3243, AddRoundTweakeyXOR_XORInst_6_0_n1}), .b ({new_AGEMA_signal_6838, new_AGEMA_signal_6834, new_AGEMA_signal_6830, new_AGEMA_signal_6826}), .c ({new_AGEMA_signal_3362, new_AGEMA_signal_3361, new_AGEMA_signal_3360, MCOutput[40]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_6_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3065, new_AGEMA_signal_3064, new_AGEMA_signal_3063, AddRoundConstantOutput[56]}), .c ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, new_AGEMA_signal_3243, AddRoundTweakeyXOR_XORInst_6_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_6_1_U2 ( .a ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, new_AGEMA_signal_3363, AddRoundTweakeyXOR_XORInst_6_1_n1}), .b ({new_AGEMA_signal_6854, new_AGEMA_signal_6850, new_AGEMA_signal_6846, new_AGEMA_signal_6842}), .c ({new_AGEMA_signal_3542, new_AGEMA_signal_3541, new_AGEMA_signal_3540, MCOutput[41]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_6_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3194, new_AGEMA_signal_3193, new_AGEMA_signal_3192, AddRoundConstantOutput[57]}), .c ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, new_AGEMA_signal_3363, AddRoundTweakeyXOR_XORInst_6_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_7_0_U2 ( .a ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, new_AGEMA_signal_3543, AddRoundTweakeyXOR_XORInst_7_0_n1}), .b ({new_AGEMA_signal_6870, new_AGEMA_signal_6866, new_AGEMA_signal_6862, new_AGEMA_signal_6858}), .c ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, new_AGEMA_signal_3699, MCOutput[44]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_7_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3314, new_AGEMA_signal_3313, new_AGEMA_signal_3312, AddRoundConstantOutput[60]}), .c ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, new_AGEMA_signal_3543, AddRoundTweakeyXOR_XORInst_7_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_7_1_U2 ( .a ({new_AGEMA_signal_3704, new_AGEMA_signal_3703, new_AGEMA_signal_3702, AddRoundTweakeyXOR_XORInst_7_1_n1}), .b ({new_AGEMA_signal_6886, new_AGEMA_signal_6882, new_AGEMA_signal_6878, new_AGEMA_signal_6874}), .c ({new_AGEMA_signal_3860, new_AGEMA_signal_3859, new_AGEMA_signal_3858, MCOutput[45]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) AddRoundTweakeyXOR_XORInst_7_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, new_AGEMA_signal_3513, AddRoundConstantOutput[61]}), .c ({new_AGEMA_signal_3704, new_AGEMA_signal_3703, new_AGEMA_signal_3702, AddRoundTweakeyXOR_XORInst_7_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_0_0_U3 ( .a ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, new_AGEMA_signal_3549, MCInst_MCR0_XORInst_0_0_n2}), .b ({new_AGEMA_signal_3254, new_AGEMA_signal_3253, new_AGEMA_signal_3252, MCInst_MCR0_XORInst_0_0_n1}), .c ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, new_AGEMA_signal_3705, MCOutput[48]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_3017, new_AGEMA_signal_3016, new_AGEMA_signal_3015, ShiftRowsOutput[16]}), .b ({new_AGEMA_signal_2999, new_AGEMA_signal_2998, new_AGEMA_signal_2997, ShiftRowsOutput[0]}), .c ({new_AGEMA_signal_3254, new_AGEMA_signal_3253, new_AGEMA_signal_3252, MCInst_MCR0_XORInst_0_0_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3350, new_AGEMA_signal_3349, new_AGEMA_signal_3348, MCOutput[32]}), .c ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, new_AGEMA_signal_3549, MCInst_MCR0_XORInst_0_0_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_0_1_U3 ( .a ({new_AGEMA_signal_3710, new_AGEMA_signal_3709, new_AGEMA_signal_3708, MCInst_MCR0_XORInst_0_1_n2}), .b ({new_AGEMA_signal_3374, new_AGEMA_signal_3373, new_AGEMA_signal_3372, MCInst_MCR0_XORInst_0_1_n1}), .c ({new_AGEMA_signal_3863, new_AGEMA_signal_3862, new_AGEMA_signal_3861, MCOutput[49]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_3170, new_AGEMA_signal_3169, new_AGEMA_signal_3168, ShiftRowsOutput[17]}), .b ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, new_AGEMA_signal_3159, ShiftRowsOutput[1]}), .c ({new_AGEMA_signal_3374, new_AGEMA_signal_3373, new_AGEMA_signal_3372, MCInst_MCR0_XORInst_0_1_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3536, new_AGEMA_signal_3535, new_AGEMA_signal_3534, MCOutput[33]}), .c ({new_AGEMA_signal_3710, new_AGEMA_signal_3709, new_AGEMA_signal_3708, MCInst_MCR0_XORInst_0_1_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_1_0_U3 ( .a ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, new_AGEMA_signal_3555, MCInst_MCR0_XORInst_1_0_n2}), .b ({new_AGEMA_signal_3260, new_AGEMA_signal_3259, new_AGEMA_signal_3258, MCInst_MCR0_XORInst_1_0_n1}), .c ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, new_AGEMA_signal_3711, MCOutput[52]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, new_AGEMA_signal_3021, ShiftRowsOutput[20]}), .b ({new_AGEMA_signal_2981, new_AGEMA_signal_2980, new_AGEMA_signal_2979, ShiftRowsOutput[4]}), .c ({new_AGEMA_signal_3260, new_AGEMA_signal_3259, new_AGEMA_signal_3258, MCInst_MCR0_XORInst_1_0_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3356, new_AGEMA_signal_3355, new_AGEMA_signal_3354, MCOutput[36]}), .c ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, new_AGEMA_signal_3555, MCInst_MCR0_XORInst_1_0_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_1_1_U3 ( .a ({new_AGEMA_signal_3716, new_AGEMA_signal_3715, new_AGEMA_signal_3714, MCInst_MCR0_XORInst_1_1_n2}), .b ({new_AGEMA_signal_3560, new_AGEMA_signal_3559, new_AGEMA_signal_3558, MCInst_MCR0_XORInst_1_1_n1}), .c ({new_AGEMA_signal_3866, new_AGEMA_signal_3865, new_AGEMA_signal_3864, MCOutput[53]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, new_AGEMA_signal_3309, ShiftRowsOutput[21]}), .b ({new_AGEMA_signal_3152, new_AGEMA_signal_3151, new_AGEMA_signal_3150, ShiftRowsOutput[5]}), .c ({new_AGEMA_signal_3560, new_AGEMA_signal_3559, new_AGEMA_signal_3558, MCInst_MCR0_XORInst_1_1_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, new_AGEMA_signal_3537, MCOutput[37]}), .c ({new_AGEMA_signal_3716, new_AGEMA_signal_3715, new_AGEMA_signal_3714, MCInst_MCR0_XORInst_1_1_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_2_0_U3 ( .a ({new_AGEMA_signal_3566, new_AGEMA_signal_3565, new_AGEMA_signal_3564, MCInst_MCR0_XORInst_2_0_n2}), .b ({new_AGEMA_signal_3266, new_AGEMA_signal_3265, new_AGEMA_signal_3264, MCInst_MCR0_XORInst_2_0_n1}), .c ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, new_AGEMA_signal_3717, MCOutput[56]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, new_AGEMA_signal_3003, ShiftRowsOutput[24]}), .b ({new_AGEMA_signal_2987, new_AGEMA_signal_2986, new_AGEMA_signal_2985, ShiftRowsOutput[8]}), .c ({new_AGEMA_signal_3266, new_AGEMA_signal_3265, new_AGEMA_signal_3264, MCInst_MCR0_XORInst_2_0_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3362, new_AGEMA_signal_3361, new_AGEMA_signal_3360, MCOutput[40]}), .c ({new_AGEMA_signal_3566, new_AGEMA_signal_3565, new_AGEMA_signal_3564, MCInst_MCR0_XORInst_2_0_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_2_1_U3 ( .a ({new_AGEMA_signal_3722, new_AGEMA_signal_3721, new_AGEMA_signal_3720, MCInst_MCR0_XORInst_2_1_n2}), .b ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, new_AGEMA_signal_3387, MCInst_MCR0_XORInst_2_1_n1}), .c ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, new_AGEMA_signal_3867, MCOutput[57]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_3164, new_AGEMA_signal_3163, new_AGEMA_signal_3162, ShiftRowsOutput[25]}), .b ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, new_AGEMA_signal_3153, ShiftRowsOutput[9]}), .c ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, new_AGEMA_signal_3387, MCInst_MCR0_XORInst_2_1_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3542, new_AGEMA_signal_3541, new_AGEMA_signal_3540, MCOutput[41]}), .c ({new_AGEMA_signal_3722, new_AGEMA_signal_3721, new_AGEMA_signal_3720, MCInst_MCR0_XORInst_2_1_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_3_0_U3 ( .a ({new_AGEMA_signal_3872, new_AGEMA_signal_3871, new_AGEMA_signal_3870, MCInst_MCR0_XORInst_3_0_n2}), .b ({new_AGEMA_signal_3272, new_AGEMA_signal_3271, new_AGEMA_signal_3270, MCInst_MCR0_XORInst_3_0_n1}), .c ({new_AGEMA_signal_3986, new_AGEMA_signal_3985, new_AGEMA_signal_3984, MCOutput[60]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, new_AGEMA_signal_3009, ShiftRowsOutput[28]}), .b ({new_AGEMA_signal_2993, new_AGEMA_signal_2992, new_AGEMA_signal_2991, ShiftRowsOutput[12]}), .c ({new_AGEMA_signal_3272, new_AGEMA_signal_3271, new_AGEMA_signal_3270, MCInst_MCR0_XORInst_3_0_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, new_AGEMA_signal_3699, MCOutput[44]}), .c ({new_AGEMA_signal_3872, new_AGEMA_signal_3871, new_AGEMA_signal_3870, MCInst_MCR0_XORInst_3_0_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_3_1_U3 ( .a ({new_AGEMA_signal_3989, new_AGEMA_signal_3988, new_AGEMA_signal_3987, MCInst_MCR0_XORInst_3_1_n2}), .b ({new_AGEMA_signal_3398, new_AGEMA_signal_3397, new_AGEMA_signal_3396, MCInst_MCR0_XORInst_3_1_n1}), .c ({new_AGEMA_signal_4022, new_AGEMA_signal_4021, new_AGEMA_signal_4020, MCOutput[61]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, new_AGEMA_signal_3165, ShiftRowsOutput[29]}), .b ({new_AGEMA_signal_3158, new_AGEMA_signal_3157, new_AGEMA_signal_3156, ShiftRowsOutput[13]}), .c ({new_AGEMA_signal_3398, new_AGEMA_signal_3397, new_AGEMA_signal_3396, MCInst_MCR0_XORInst_3_1_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR0_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3860, new_AGEMA_signal_3859, new_AGEMA_signal_3858, MCOutput[45]}), .c ({new_AGEMA_signal_3989, new_AGEMA_signal_3988, new_AGEMA_signal_3987, MCInst_MCR0_XORInst_3_1_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, new_AGEMA_signal_3573, MCInst_MCR2_XORInst_0_0_n1}), .b ({new_AGEMA_signal_3017, new_AGEMA_signal_3016, new_AGEMA_signal_3015, ShiftRowsOutput[16]}), .c ({new_AGEMA_signal_3731, new_AGEMA_signal_3730, new_AGEMA_signal_3729, MCOutput[16]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3332, new_AGEMA_signal_3331, new_AGEMA_signal_3330, ShiftRowsOutput[32]}), .c ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, new_AGEMA_signal_3573, MCInst_MCR2_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_3734, new_AGEMA_signal_3733, new_AGEMA_signal_3732, MCInst_MCR2_XORInst_0_1_n1}), .b ({new_AGEMA_signal_3170, new_AGEMA_signal_3169, new_AGEMA_signal_3168, ShiftRowsOutput[17]}), .c ({new_AGEMA_signal_3878, new_AGEMA_signal_3877, new_AGEMA_signal_3876, MCOutput[17]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3524, new_AGEMA_signal_3523, new_AGEMA_signal_3522, ShiftRowsOutput[33]}), .c ({new_AGEMA_signal_3734, new_AGEMA_signal_3733, new_AGEMA_signal_3732, MCInst_MCR2_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, new_AGEMA_signal_3579, MCInst_MCR2_XORInst_1_0_n1}), .b ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, new_AGEMA_signal_3021, ShiftRowsOutput[20]}), .c ({new_AGEMA_signal_3737, new_AGEMA_signal_3736, new_AGEMA_signal_3735, MCOutput[20]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3338, new_AGEMA_signal_3337, new_AGEMA_signal_3336, ShiftRowsOutput[36]}), .c ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, new_AGEMA_signal_3579, MCInst_MCR2_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_3740, new_AGEMA_signal_3739, new_AGEMA_signal_3738, MCInst_MCR2_XORInst_1_1_n1}), .b ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, new_AGEMA_signal_3309, ShiftRowsOutput[21]}), .c ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, new_AGEMA_signal_3879, MCOutput[21]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, new_AGEMA_signal_3525, ShiftRowsOutput[37]}), .c ({new_AGEMA_signal_3740, new_AGEMA_signal_3739, new_AGEMA_signal_3738, MCInst_MCR2_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_3884, new_AGEMA_signal_3883, new_AGEMA_signal_3882, MCInst_MCR2_XORInst_2_0_n1}), .b ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, new_AGEMA_signal_3003, ShiftRowsOutput[24]}), .c ({new_AGEMA_signal_3992, new_AGEMA_signal_3991, new_AGEMA_signal_3990, MCOutput[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, new_AGEMA_signal_3693, ShiftRowsOutput[40]}), .c ({new_AGEMA_signal_3884, new_AGEMA_signal_3883, new_AGEMA_signal_3882, MCInst_MCR2_XORInst_2_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_3995, new_AGEMA_signal_3994, new_AGEMA_signal_3993, MCInst_MCR2_XORInst_2_1_n1}), .b ({new_AGEMA_signal_3164, new_AGEMA_signal_3163, new_AGEMA_signal_3162, ShiftRowsOutput[25]}), .c ({new_AGEMA_signal_4025, new_AGEMA_signal_4024, new_AGEMA_signal_4023, MCOutput[25]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, new_AGEMA_signal_3855, ShiftRowsOutput[41]}), .c ({new_AGEMA_signal_3995, new_AGEMA_signal_3994, new_AGEMA_signal_3993, MCInst_MCR2_XORInst_2_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_3590, new_AGEMA_signal_3589, new_AGEMA_signal_3588, MCInst_MCR2_XORInst_3_0_n1}), .b ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, new_AGEMA_signal_3009, ShiftRowsOutput[28]}), .c ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, new_AGEMA_signal_3747, MCOutput[28]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3326, new_AGEMA_signal_3325, new_AGEMA_signal_3324, ShiftRowsOutput[44]}), .c ({new_AGEMA_signal_3590, new_AGEMA_signal_3589, new_AGEMA_signal_3588, MCInst_MCR2_XORInst_3_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_3752, new_AGEMA_signal_3751, new_AGEMA_signal_3750, MCInst_MCR2_XORInst_3_1_n1}), .b ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, new_AGEMA_signal_3165, ShiftRowsOutput[29]}), .c ({new_AGEMA_signal_3890, new_AGEMA_signal_3889, new_AGEMA_signal_3888, MCOutput[29]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR2_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, new_AGEMA_signal_3519, ShiftRowsOutput[45]}), .c ({new_AGEMA_signal_3752, new_AGEMA_signal_3751, new_AGEMA_signal_3750, MCInst_MCR2_XORInst_3_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_3596, new_AGEMA_signal_3595, new_AGEMA_signal_3594, MCInst_MCR3_XORInst_0_0_n1}), .b ({new_AGEMA_signal_3017, new_AGEMA_signal_3016, new_AGEMA_signal_3015, ShiftRowsOutput[16]}), .c ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, new_AGEMA_signal_3753, MCOutput[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3350, new_AGEMA_signal_3349, new_AGEMA_signal_3348, MCOutput[32]}), .c ({new_AGEMA_signal_3596, new_AGEMA_signal_3595, new_AGEMA_signal_3594, MCInst_MCR3_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_3758, new_AGEMA_signal_3757, new_AGEMA_signal_3756, MCInst_MCR3_XORInst_0_1_n1}), .b ({new_AGEMA_signal_3170, new_AGEMA_signal_3169, new_AGEMA_signal_3168, ShiftRowsOutput[17]}), .c ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, new_AGEMA_signal_3891, MCOutput[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3536, new_AGEMA_signal_3535, new_AGEMA_signal_3534, MCOutput[33]}), .c ({new_AGEMA_signal_3758, new_AGEMA_signal_3757, new_AGEMA_signal_3756, MCInst_MCR3_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_3602, new_AGEMA_signal_3601, new_AGEMA_signal_3600, MCInst_MCR3_XORInst_1_0_n1}), .b ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, new_AGEMA_signal_3021, ShiftRowsOutput[20]}), .c ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, new_AGEMA_signal_3759, MCOutput[4]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3356, new_AGEMA_signal_3355, new_AGEMA_signal_3354, MCOutput[36]}), .c ({new_AGEMA_signal_3602, new_AGEMA_signal_3601, new_AGEMA_signal_3600, MCInst_MCR3_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_3764, new_AGEMA_signal_3763, new_AGEMA_signal_3762, MCInst_MCR3_XORInst_1_1_n1}), .b ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, new_AGEMA_signal_3309, ShiftRowsOutput[21]}), .c ({new_AGEMA_signal_3896, new_AGEMA_signal_3895, new_AGEMA_signal_3894, MCOutput[5]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, new_AGEMA_signal_3537, MCOutput[37]}), .c ({new_AGEMA_signal_3764, new_AGEMA_signal_3763, new_AGEMA_signal_3762, MCInst_MCR3_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_3608, new_AGEMA_signal_3607, new_AGEMA_signal_3606, MCInst_MCR3_XORInst_2_0_n1}), .b ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, new_AGEMA_signal_3003, ShiftRowsOutput[24]}), .c ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, new_AGEMA_signal_3765, MCOutput[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3362, new_AGEMA_signal_3361, new_AGEMA_signal_3360, MCOutput[40]}), .c ({new_AGEMA_signal_3608, new_AGEMA_signal_3607, new_AGEMA_signal_3606, MCInst_MCR3_XORInst_2_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_3770, new_AGEMA_signal_3769, new_AGEMA_signal_3768, MCInst_MCR3_XORInst_2_1_n1}), .b ({new_AGEMA_signal_3164, new_AGEMA_signal_3163, new_AGEMA_signal_3162, ShiftRowsOutput[25]}), .c ({new_AGEMA_signal_3899, new_AGEMA_signal_3898, new_AGEMA_signal_3897, MCOutput[9]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3542, new_AGEMA_signal_3541, new_AGEMA_signal_3540, MCOutput[41]}), .c ({new_AGEMA_signal_3770, new_AGEMA_signal_3769, new_AGEMA_signal_3768, MCInst_MCR3_XORInst_2_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_3902, new_AGEMA_signal_3901, new_AGEMA_signal_3900, MCInst_MCR3_XORInst_3_0_n1}), .b ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, new_AGEMA_signal_3009, ShiftRowsOutput[28]}), .c ({new_AGEMA_signal_3998, new_AGEMA_signal_3997, new_AGEMA_signal_3996, MCOutput[12]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, new_AGEMA_signal_3699, MCOutput[44]}), .c ({new_AGEMA_signal_3902, new_AGEMA_signal_3901, new_AGEMA_signal_3900, MCInst_MCR3_XORInst_3_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_4001, new_AGEMA_signal_4000, new_AGEMA_signal_3999, MCInst_MCR3_XORInst_3_1_n1}), .b ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, new_AGEMA_signal_3165, ShiftRowsOutput[29]}), .c ({new_AGEMA_signal_4028, new_AGEMA_signal_4027, new_AGEMA_signal_4026, MCOutput[13]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) MCInst_MCR3_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3860, new_AGEMA_signal_3859, new_AGEMA_signal_3858, MCOutput[45]}), .c ({new_AGEMA_signal_4001, new_AGEMA_signal_4000, new_AGEMA_signal_3999, MCInst_MCR3_XORInst_3_1_n1}) ) ;
    buf_clk new_AGEMA_reg_buffer_1903 ( .C (clk), .D (new_AGEMA_signal_5333), .Q (new_AGEMA_signal_5334) ) ;
    buf_clk new_AGEMA_reg_buffer_1907 ( .C (clk), .D (new_AGEMA_signal_5337), .Q (new_AGEMA_signal_5338) ) ;
    buf_clk new_AGEMA_reg_buffer_1911 ( .C (clk), .D (new_AGEMA_signal_5341), .Q (new_AGEMA_signal_5342) ) ;
    buf_clk new_AGEMA_reg_buffer_1915 ( .C (clk), .D (new_AGEMA_signal_5345), .Q (new_AGEMA_signal_5346) ) ;
    buf_clk new_AGEMA_reg_buffer_1919 ( .C (clk), .D (new_AGEMA_signal_5349), .Q (new_AGEMA_signal_5350) ) ;
    buf_clk new_AGEMA_reg_buffer_1923 ( .C (clk), .D (new_AGEMA_signal_5353), .Q (new_AGEMA_signal_5354) ) ;
    buf_clk new_AGEMA_reg_buffer_1927 ( .C (clk), .D (new_AGEMA_signal_5357), .Q (new_AGEMA_signal_5358) ) ;
    buf_clk new_AGEMA_reg_buffer_1931 ( .C (clk), .D (new_AGEMA_signal_5361), .Q (new_AGEMA_signal_5362) ) ;
    buf_clk new_AGEMA_reg_buffer_1935 ( .C (clk), .D (new_AGEMA_signal_5365), .Q (new_AGEMA_signal_5366) ) ;
    buf_clk new_AGEMA_reg_buffer_1939 ( .C (clk), .D (new_AGEMA_signal_5369), .Q (new_AGEMA_signal_5370) ) ;
    buf_clk new_AGEMA_reg_buffer_1943 ( .C (clk), .D (new_AGEMA_signal_5373), .Q (new_AGEMA_signal_5374) ) ;
    buf_clk new_AGEMA_reg_buffer_1947 ( .C (clk), .D (new_AGEMA_signal_5377), .Q (new_AGEMA_signal_5378) ) ;
    buf_clk new_AGEMA_reg_buffer_1951 ( .C (clk), .D (new_AGEMA_signal_5381), .Q (new_AGEMA_signal_5382) ) ;
    buf_clk new_AGEMA_reg_buffer_1955 ( .C (clk), .D (new_AGEMA_signal_5385), .Q (new_AGEMA_signal_5386) ) ;
    buf_clk new_AGEMA_reg_buffer_1959 ( .C (clk), .D (new_AGEMA_signal_5389), .Q (new_AGEMA_signal_5390) ) ;
    buf_clk new_AGEMA_reg_buffer_1963 ( .C (clk), .D (new_AGEMA_signal_5393), .Q (new_AGEMA_signal_5394) ) ;
    buf_clk new_AGEMA_reg_buffer_1967 ( .C (clk), .D (new_AGEMA_signal_5397), .Q (new_AGEMA_signal_5398) ) ;
    buf_clk new_AGEMA_reg_buffer_1971 ( .C (clk), .D (new_AGEMA_signal_5401), .Q (new_AGEMA_signal_5402) ) ;
    buf_clk new_AGEMA_reg_buffer_1975 ( .C (clk), .D (new_AGEMA_signal_5405), .Q (new_AGEMA_signal_5406) ) ;
    buf_clk new_AGEMA_reg_buffer_1979 ( .C (clk), .D (new_AGEMA_signal_5409), .Q (new_AGEMA_signal_5410) ) ;
    buf_clk new_AGEMA_reg_buffer_1983 ( .C (clk), .D (new_AGEMA_signal_5413), .Q (new_AGEMA_signal_5414) ) ;
    buf_clk new_AGEMA_reg_buffer_1987 ( .C (clk), .D (new_AGEMA_signal_5417), .Q (new_AGEMA_signal_5418) ) ;
    buf_clk new_AGEMA_reg_buffer_1991 ( .C (clk), .D (new_AGEMA_signal_5421), .Q (new_AGEMA_signal_5422) ) ;
    buf_clk new_AGEMA_reg_buffer_1995 ( .C (clk), .D (new_AGEMA_signal_5425), .Q (new_AGEMA_signal_5426) ) ;
    buf_clk new_AGEMA_reg_buffer_1999 ( .C (clk), .D (new_AGEMA_signal_5429), .Q (new_AGEMA_signal_5430) ) ;
    buf_clk new_AGEMA_reg_buffer_2003 ( .C (clk), .D (new_AGEMA_signal_5433), .Q (new_AGEMA_signal_5434) ) ;
    buf_clk new_AGEMA_reg_buffer_2007 ( .C (clk), .D (new_AGEMA_signal_5437), .Q (new_AGEMA_signal_5438) ) ;
    buf_clk new_AGEMA_reg_buffer_2011 ( .C (clk), .D (new_AGEMA_signal_5441), .Q (new_AGEMA_signal_5442) ) ;
    buf_clk new_AGEMA_reg_buffer_2015 ( .C (clk), .D (new_AGEMA_signal_5445), .Q (new_AGEMA_signal_5446) ) ;
    buf_clk new_AGEMA_reg_buffer_2019 ( .C (clk), .D (new_AGEMA_signal_5449), .Q (new_AGEMA_signal_5450) ) ;
    buf_clk new_AGEMA_reg_buffer_2023 ( .C (clk), .D (new_AGEMA_signal_5453), .Q (new_AGEMA_signal_5454) ) ;
    buf_clk new_AGEMA_reg_buffer_2027 ( .C (clk), .D (new_AGEMA_signal_5457), .Q (new_AGEMA_signal_5458) ) ;
    buf_clk new_AGEMA_reg_buffer_2031 ( .C (clk), .D (new_AGEMA_signal_5461), .Q (new_AGEMA_signal_5462) ) ;
    buf_clk new_AGEMA_reg_buffer_2035 ( .C (clk), .D (new_AGEMA_signal_5465), .Q (new_AGEMA_signal_5466) ) ;
    buf_clk new_AGEMA_reg_buffer_2039 ( .C (clk), .D (new_AGEMA_signal_5469), .Q (new_AGEMA_signal_5470) ) ;
    buf_clk new_AGEMA_reg_buffer_2043 ( .C (clk), .D (new_AGEMA_signal_5473), .Q (new_AGEMA_signal_5474) ) ;
    buf_clk new_AGEMA_reg_buffer_2047 ( .C (clk), .D (new_AGEMA_signal_5477), .Q (new_AGEMA_signal_5478) ) ;
    buf_clk new_AGEMA_reg_buffer_2051 ( .C (clk), .D (new_AGEMA_signal_5481), .Q (new_AGEMA_signal_5482) ) ;
    buf_clk new_AGEMA_reg_buffer_2055 ( .C (clk), .D (new_AGEMA_signal_5485), .Q (new_AGEMA_signal_5486) ) ;
    buf_clk new_AGEMA_reg_buffer_2059 ( .C (clk), .D (new_AGEMA_signal_5489), .Q (new_AGEMA_signal_5490) ) ;
    buf_clk new_AGEMA_reg_buffer_2063 ( .C (clk), .D (new_AGEMA_signal_5493), .Q (new_AGEMA_signal_5494) ) ;
    buf_clk new_AGEMA_reg_buffer_2067 ( .C (clk), .D (new_AGEMA_signal_5497), .Q (new_AGEMA_signal_5498) ) ;
    buf_clk new_AGEMA_reg_buffer_2071 ( .C (clk), .D (new_AGEMA_signal_5501), .Q (new_AGEMA_signal_5502) ) ;
    buf_clk new_AGEMA_reg_buffer_2075 ( .C (clk), .D (new_AGEMA_signal_5505), .Q (new_AGEMA_signal_5506) ) ;
    buf_clk new_AGEMA_reg_buffer_2079 ( .C (clk), .D (new_AGEMA_signal_5509), .Q (new_AGEMA_signal_5510) ) ;
    buf_clk new_AGEMA_reg_buffer_2083 ( .C (clk), .D (new_AGEMA_signal_5513), .Q (new_AGEMA_signal_5514) ) ;
    buf_clk new_AGEMA_reg_buffer_2087 ( .C (clk), .D (new_AGEMA_signal_5517), .Q (new_AGEMA_signal_5518) ) ;
    buf_clk new_AGEMA_reg_buffer_2091 ( .C (clk), .D (new_AGEMA_signal_5521), .Q (new_AGEMA_signal_5522) ) ;
    buf_clk new_AGEMA_reg_buffer_2095 ( .C (clk), .D (new_AGEMA_signal_5525), .Q (new_AGEMA_signal_5526) ) ;
    buf_clk new_AGEMA_reg_buffer_2099 ( .C (clk), .D (new_AGEMA_signal_5529), .Q (new_AGEMA_signal_5530) ) ;
    buf_clk new_AGEMA_reg_buffer_2103 ( .C (clk), .D (new_AGEMA_signal_5533), .Q (new_AGEMA_signal_5534) ) ;
    buf_clk new_AGEMA_reg_buffer_2107 ( .C (clk), .D (new_AGEMA_signal_5537), .Q (new_AGEMA_signal_5538) ) ;
    buf_clk new_AGEMA_reg_buffer_2111 ( .C (clk), .D (new_AGEMA_signal_5541), .Q (new_AGEMA_signal_5542) ) ;
    buf_clk new_AGEMA_reg_buffer_2115 ( .C (clk), .D (new_AGEMA_signal_5545), .Q (new_AGEMA_signal_5546) ) ;
    buf_clk new_AGEMA_reg_buffer_2119 ( .C (clk), .D (new_AGEMA_signal_5549), .Q (new_AGEMA_signal_5550) ) ;
    buf_clk new_AGEMA_reg_buffer_2123 ( .C (clk), .D (new_AGEMA_signal_5553), .Q (new_AGEMA_signal_5554) ) ;
    buf_clk new_AGEMA_reg_buffer_2127 ( .C (clk), .D (new_AGEMA_signal_5557), .Q (new_AGEMA_signal_5558) ) ;
    buf_clk new_AGEMA_reg_buffer_2131 ( .C (clk), .D (new_AGEMA_signal_5561), .Q (new_AGEMA_signal_5562) ) ;
    buf_clk new_AGEMA_reg_buffer_2135 ( .C (clk), .D (new_AGEMA_signal_5565), .Q (new_AGEMA_signal_5566) ) ;
    buf_clk new_AGEMA_reg_buffer_2139 ( .C (clk), .D (new_AGEMA_signal_5569), .Q (new_AGEMA_signal_5570) ) ;
    buf_clk new_AGEMA_reg_buffer_2143 ( .C (clk), .D (new_AGEMA_signal_5573), .Q (new_AGEMA_signal_5574) ) ;
    buf_clk new_AGEMA_reg_buffer_2147 ( .C (clk), .D (new_AGEMA_signal_5577), .Q (new_AGEMA_signal_5578) ) ;
    buf_clk new_AGEMA_reg_buffer_2151 ( .C (clk), .D (new_AGEMA_signal_5581), .Q (new_AGEMA_signal_5582) ) ;
    buf_clk new_AGEMA_reg_buffer_2155 ( .C (clk), .D (new_AGEMA_signal_5585), .Q (new_AGEMA_signal_5586) ) ;
    buf_clk new_AGEMA_reg_buffer_2159 ( .C (clk), .D (new_AGEMA_signal_5589), .Q (new_AGEMA_signal_5590) ) ;
    buf_clk new_AGEMA_reg_buffer_2163 ( .C (clk), .D (new_AGEMA_signal_5593), .Q (new_AGEMA_signal_5594) ) ;
    buf_clk new_AGEMA_reg_buffer_2167 ( .C (clk), .D (new_AGEMA_signal_5597), .Q (new_AGEMA_signal_5598) ) ;
    buf_clk new_AGEMA_reg_buffer_2171 ( .C (clk), .D (new_AGEMA_signal_5601), .Q (new_AGEMA_signal_5602) ) ;
    buf_clk new_AGEMA_reg_buffer_2175 ( .C (clk), .D (new_AGEMA_signal_5605), .Q (new_AGEMA_signal_5606) ) ;
    buf_clk new_AGEMA_reg_buffer_2179 ( .C (clk), .D (new_AGEMA_signal_5609), .Q (new_AGEMA_signal_5610) ) ;
    buf_clk new_AGEMA_reg_buffer_2183 ( .C (clk), .D (new_AGEMA_signal_5613), .Q (new_AGEMA_signal_5614) ) ;
    buf_clk new_AGEMA_reg_buffer_2187 ( .C (clk), .D (new_AGEMA_signal_5617), .Q (new_AGEMA_signal_5618) ) ;
    buf_clk new_AGEMA_reg_buffer_2191 ( .C (clk), .D (new_AGEMA_signal_5621), .Q (new_AGEMA_signal_5622) ) ;
    buf_clk new_AGEMA_reg_buffer_2195 ( .C (clk), .D (new_AGEMA_signal_5625), .Q (new_AGEMA_signal_5626) ) ;
    buf_clk new_AGEMA_reg_buffer_2199 ( .C (clk), .D (new_AGEMA_signal_5629), .Q (new_AGEMA_signal_5630) ) ;
    buf_clk new_AGEMA_reg_buffer_2203 ( .C (clk), .D (new_AGEMA_signal_5633), .Q (new_AGEMA_signal_5634) ) ;
    buf_clk new_AGEMA_reg_buffer_2207 ( .C (clk), .D (new_AGEMA_signal_5637), .Q (new_AGEMA_signal_5638) ) ;
    buf_clk new_AGEMA_reg_buffer_2211 ( .C (clk), .D (new_AGEMA_signal_5641), .Q (new_AGEMA_signal_5642) ) ;
    buf_clk new_AGEMA_reg_buffer_2215 ( .C (clk), .D (new_AGEMA_signal_5645), .Q (new_AGEMA_signal_5646) ) ;
    buf_clk new_AGEMA_reg_buffer_2219 ( .C (clk), .D (new_AGEMA_signal_5649), .Q (new_AGEMA_signal_5650) ) ;
    buf_clk new_AGEMA_reg_buffer_2223 ( .C (clk), .D (new_AGEMA_signal_5653), .Q (new_AGEMA_signal_5654) ) ;
    buf_clk new_AGEMA_reg_buffer_2227 ( .C (clk), .D (new_AGEMA_signal_5657), .Q (new_AGEMA_signal_5658) ) ;
    buf_clk new_AGEMA_reg_buffer_2231 ( .C (clk), .D (new_AGEMA_signal_5661), .Q (new_AGEMA_signal_5662) ) ;
    buf_clk new_AGEMA_reg_buffer_2235 ( .C (clk), .D (new_AGEMA_signal_5665), .Q (new_AGEMA_signal_5666) ) ;
    buf_clk new_AGEMA_reg_buffer_2239 ( .C (clk), .D (new_AGEMA_signal_5669), .Q (new_AGEMA_signal_5670) ) ;
    buf_clk new_AGEMA_reg_buffer_2243 ( .C (clk), .D (new_AGEMA_signal_5673), .Q (new_AGEMA_signal_5674) ) ;
    buf_clk new_AGEMA_reg_buffer_2247 ( .C (clk), .D (new_AGEMA_signal_5677), .Q (new_AGEMA_signal_5678) ) ;
    buf_clk new_AGEMA_reg_buffer_2251 ( .C (clk), .D (new_AGEMA_signal_5681), .Q (new_AGEMA_signal_5682) ) ;
    buf_clk new_AGEMA_reg_buffer_2255 ( .C (clk), .D (new_AGEMA_signal_5685), .Q (new_AGEMA_signal_5686) ) ;
    buf_clk new_AGEMA_reg_buffer_2259 ( .C (clk), .D (new_AGEMA_signal_5689), .Q (new_AGEMA_signal_5690) ) ;
    buf_clk new_AGEMA_reg_buffer_2263 ( .C (clk), .D (new_AGEMA_signal_5693), .Q (new_AGEMA_signal_5694) ) ;
    buf_clk new_AGEMA_reg_buffer_2267 ( .C (clk), .D (new_AGEMA_signal_5697), .Q (new_AGEMA_signal_5698) ) ;
    buf_clk new_AGEMA_reg_buffer_2271 ( .C (clk), .D (new_AGEMA_signal_5701), .Q (new_AGEMA_signal_5702) ) ;
    buf_clk new_AGEMA_reg_buffer_2275 ( .C (clk), .D (new_AGEMA_signal_5705), .Q (new_AGEMA_signal_5706) ) ;
    buf_clk new_AGEMA_reg_buffer_2279 ( .C (clk), .D (new_AGEMA_signal_5709), .Q (new_AGEMA_signal_5710) ) ;
    buf_clk new_AGEMA_reg_buffer_2283 ( .C (clk), .D (new_AGEMA_signal_5713), .Q (new_AGEMA_signal_5714) ) ;
    buf_clk new_AGEMA_reg_buffer_2287 ( .C (clk), .D (new_AGEMA_signal_5717), .Q (new_AGEMA_signal_5718) ) ;
    buf_clk new_AGEMA_reg_buffer_2291 ( .C (clk), .D (new_AGEMA_signal_5721), .Q (new_AGEMA_signal_5722) ) ;
    buf_clk new_AGEMA_reg_buffer_2295 ( .C (clk), .D (new_AGEMA_signal_5725), .Q (new_AGEMA_signal_5726) ) ;
    buf_clk new_AGEMA_reg_buffer_2299 ( .C (clk), .D (new_AGEMA_signal_5729), .Q (new_AGEMA_signal_5730) ) ;
    buf_clk new_AGEMA_reg_buffer_2303 ( .C (clk), .D (new_AGEMA_signal_5733), .Q (new_AGEMA_signal_5734) ) ;
    buf_clk new_AGEMA_reg_buffer_2307 ( .C (clk), .D (new_AGEMA_signal_5737), .Q (new_AGEMA_signal_5738) ) ;
    buf_clk new_AGEMA_reg_buffer_2311 ( .C (clk), .D (new_AGEMA_signal_5741), .Q (new_AGEMA_signal_5742) ) ;
    buf_clk new_AGEMA_reg_buffer_2315 ( .C (clk), .D (new_AGEMA_signal_5745), .Q (new_AGEMA_signal_5746) ) ;
    buf_clk new_AGEMA_reg_buffer_2319 ( .C (clk), .D (new_AGEMA_signal_5749), .Q (new_AGEMA_signal_5750) ) ;
    buf_clk new_AGEMA_reg_buffer_2323 ( .C (clk), .D (new_AGEMA_signal_5753), .Q (new_AGEMA_signal_5754) ) ;
    buf_clk new_AGEMA_reg_buffer_2327 ( .C (clk), .D (new_AGEMA_signal_5757), .Q (new_AGEMA_signal_5758) ) ;
    buf_clk new_AGEMA_reg_buffer_2331 ( .C (clk), .D (new_AGEMA_signal_5761), .Q (new_AGEMA_signal_5762) ) ;
    buf_clk new_AGEMA_reg_buffer_2335 ( .C (clk), .D (new_AGEMA_signal_5765), .Q (new_AGEMA_signal_5766) ) ;
    buf_clk new_AGEMA_reg_buffer_2339 ( .C (clk), .D (new_AGEMA_signal_5769), .Q (new_AGEMA_signal_5770) ) ;
    buf_clk new_AGEMA_reg_buffer_2343 ( .C (clk), .D (new_AGEMA_signal_5773), .Q (new_AGEMA_signal_5774) ) ;
    buf_clk new_AGEMA_reg_buffer_2347 ( .C (clk), .D (new_AGEMA_signal_5777), .Q (new_AGEMA_signal_5778) ) ;
    buf_clk new_AGEMA_reg_buffer_2351 ( .C (clk), .D (new_AGEMA_signal_5781), .Q (new_AGEMA_signal_5782) ) ;
    buf_clk new_AGEMA_reg_buffer_2355 ( .C (clk), .D (new_AGEMA_signal_5785), .Q (new_AGEMA_signal_5786) ) ;
    buf_clk new_AGEMA_reg_buffer_2359 ( .C (clk), .D (new_AGEMA_signal_5789), .Q (new_AGEMA_signal_5790) ) ;
    buf_clk new_AGEMA_reg_buffer_2363 ( .C (clk), .D (new_AGEMA_signal_5793), .Q (new_AGEMA_signal_5794) ) ;
    buf_clk new_AGEMA_reg_buffer_2367 ( .C (clk), .D (new_AGEMA_signal_5797), .Q (new_AGEMA_signal_5798) ) ;
    buf_clk new_AGEMA_reg_buffer_2371 ( .C (clk), .D (new_AGEMA_signal_5801), .Q (new_AGEMA_signal_5802) ) ;
    buf_clk new_AGEMA_reg_buffer_2375 ( .C (clk), .D (new_AGEMA_signal_5805), .Q (new_AGEMA_signal_5806) ) ;
    buf_clk new_AGEMA_reg_buffer_2379 ( .C (clk), .D (new_AGEMA_signal_5809), .Q (new_AGEMA_signal_5810) ) ;
    buf_clk new_AGEMA_reg_buffer_2383 ( .C (clk), .D (new_AGEMA_signal_5813), .Q (new_AGEMA_signal_5814) ) ;
    buf_clk new_AGEMA_reg_buffer_2387 ( .C (clk), .D (new_AGEMA_signal_5817), .Q (new_AGEMA_signal_5818) ) ;
    buf_clk new_AGEMA_reg_buffer_2391 ( .C (clk), .D (new_AGEMA_signal_5821), .Q (new_AGEMA_signal_5822) ) ;
    buf_clk new_AGEMA_reg_buffer_2395 ( .C (clk), .D (new_AGEMA_signal_5825), .Q (new_AGEMA_signal_5826) ) ;
    buf_clk new_AGEMA_reg_buffer_2399 ( .C (clk), .D (new_AGEMA_signal_5829), .Q (new_AGEMA_signal_5830) ) ;
    buf_clk new_AGEMA_reg_buffer_2403 ( .C (clk), .D (new_AGEMA_signal_5833), .Q (new_AGEMA_signal_5834) ) ;
    buf_clk new_AGEMA_reg_buffer_2407 ( .C (clk), .D (new_AGEMA_signal_5837), .Q (new_AGEMA_signal_5838) ) ;
    buf_clk new_AGEMA_reg_buffer_2411 ( .C (clk), .D (new_AGEMA_signal_5841), .Q (new_AGEMA_signal_5842) ) ;
    buf_clk new_AGEMA_reg_buffer_2415 ( .C (clk), .D (new_AGEMA_signal_5845), .Q (new_AGEMA_signal_5846) ) ;
    buf_clk new_AGEMA_reg_buffer_2425 ( .C (clk), .D (new_AGEMA_signal_5855), .Q (new_AGEMA_signal_5856) ) ;
    buf_clk new_AGEMA_reg_buffer_2427 ( .C (clk), .D (new_AGEMA_signal_5857), .Q (new_AGEMA_signal_5858) ) ;
    buf_clk new_AGEMA_reg_buffer_2429 ( .C (clk), .D (new_AGEMA_signal_5859), .Q (new_AGEMA_signal_5860) ) ;
    buf_clk new_AGEMA_reg_buffer_2431 ( .C (clk), .D (new_AGEMA_signal_5861), .Q (new_AGEMA_signal_5862) ) ;
    buf_clk new_AGEMA_reg_buffer_2443 ( .C (clk), .D (new_AGEMA_signal_5873), .Q (new_AGEMA_signal_5874) ) ;
    buf_clk new_AGEMA_reg_buffer_2447 ( .C (clk), .D (new_AGEMA_signal_5877), .Q (new_AGEMA_signal_5878) ) ;
    buf_clk new_AGEMA_reg_buffer_2451 ( .C (clk), .D (new_AGEMA_signal_5881), .Q (new_AGEMA_signal_5882) ) ;
    buf_clk new_AGEMA_reg_buffer_2455 ( .C (clk), .D (new_AGEMA_signal_5885), .Q (new_AGEMA_signal_5886) ) ;
    buf_clk new_AGEMA_reg_buffer_2457 ( .C (clk), .D (new_AGEMA_signal_5887), .Q (new_AGEMA_signal_5888) ) ;
    buf_clk new_AGEMA_reg_buffer_2459 ( .C (clk), .D (new_AGEMA_signal_5889), .Q (new_AGEMA_signal_5890) ) ;
    buf_clk new_AGEMA_reg_buffer_2461 ( .C (clk), .D (new_AGEMA_signal_5891), .Q (new_AGEMA_signal_5892) ) ;
    buf_clk new_AGEMA_reg_buffer_2463 ( .C (clk), .D (new_AGEMA_signal_5893), .Q (new_AGEMA_signal_5894) ) ;
    buf_clk new_AGEMA_reg_buffer_2473 ( .C (clk), .D (new_AGEMA_signal_5903), .Q (new_AGEMA_signal_5904) ) ;
    buf_clk new_AGEMA_reg_buffer_2475 ( .C (clk), .D (new_AGEMA_signal_5905), .Q (new_AGEMA_signal_5906) ) ;
    buf_clk new_AGEMA_reg_buffer_2477 ( .C (clk), .D (new_AGEMA_signal_5907), .Q (new_AGEMA_signal_5908) ) ;
    buf_clk new_AGEMA_reg_buffer_2479 ( .C (clk), .D (new_AGEMA_signal_5909), .Q (new_AGEMA_signal_5910) ) ;
    buf_clk new_AGEMA_reg_buffer_2491 ( .C (clk), .D (new_AGEMA_signal_5921), .Q (new_AGEMA_signal_5922) ) ;
    buf_clk new_AGEMA_reg_buffer_2495 ( .C (clk), .D (new_AGEMA_signal_5925), .Q (new_AGEMA_signal_5926) ) ;
    buf_clk new_AGEMA_reg_buffer_2499 ( .C (clk), .D (new_AGEMA_signal_5929), .Q (new_AGEMA_signal_5930) ) ;
    buf_clk new_AGEMA_reg_buffer_2503 ( .C (clk), .D (new_AGEMA_signal_5933), .Q (new_AGEMA_signal_5934) ) ;
    buf_clk new_AGEMA_reg_buffer_2505 ( .C (clk), .D (new_AGEMA_signal_5935), .Q (new_AGEMA_signal_5936) ) ;
    buf_clk new_AGEMA_reg_buffer_2507 ( .C (clk), .D (new_AGEMA_signal_5937), .Q (new_AGEMA_signal_5938) ) ;
    buf_clk new_AGEMA_reg_buffer_2509 ( .C (clk), .D (new_AGEMA_signal_5939), .Q (new_AGEMA_signal_5940) ) ;
    buf_clk new_AGEMA_reg_buffer_2511 ( .C (clk), .D (new_AGEMA_signal_5941), .Q (new_AGEMA_signal_5942) ) ;
    buf_clk new_AGEMA_reg_buffer_2521 ( .C (clk), .D (new_AGEMA_signal_5951), .Q (new_AGEMA_signal_5952) ) ;
    buf_clk new_AGEMA_reg_buffer_2523 ( .C (clk), .D (new_AGEMA_signal_5953), .Q (new_AGEMA_signal_5954) ) ;
    buf_clk new_AGEMA_reg_buffer_2525 ( .C (clk), .D (new_AGEMA_signal_5955), .Q (new_AGEMA_signal_5956) ) ;
    buf_clk new_AGEMA_reg_buffer_2527 ( .C (clk), .D (new_AGEMA_signal_5957), .Q (new_AGEMA_signal_5958) ) ;
    buf_clk new_AGEMA_reg_buffer_2539 ( .C (clk), .D (new_AGEMA_signal_5969), .Q (new_AGEMA_signal_5970) ) ;
    buf_clk new_AGEMA_reg_buffer_2543 ( .C (clk), .D (new_AGEMA_signal_5973), .Q (new_AGEMA_signal_5974) ) ;
    buf_clk new_AGEMA_reg_buffer_2547 ( .C (clk), .D (new_AGEMA_signal_5977), .Q (new_AGEMA_signal_5978) ) ;
    buf_clk new_AGEMA_reg_buffer_2551 ( .C (clk), .D (new_AGEMA_signal_5981), .Q (new_AGEMA_signal_5982) ) ;
    buf_clk new_AGEMA_reg_buffer_2553 ( .C (clk), .D (new_AGEMA_signal_5983), .Q (new_AGEMA_signal_5984) ) ;
    buf_clk new_AGEMA_reg_buffer_2555 ( .C (clk), .D (new_AGEMA_signal_5985), .Q (new_AGEMA_signal_5986) ) ;
    buf_clk new_AGEMA_reg_buffer_2557 ( .C (clk), .D (new_AGEMA_signal_5987), .Q (new_AGEMA_signal_5988) ) ;
    buf_clk new_AGEMA_reg_buffer_2559 ( .C (clk), .D (new_AGEMA_signal_5989), .Q (new_AGEMA_signal_5990) ) ;
    buf_clk new_AGEMA_reg_buffer_2569 ( .C (clk), .D (new_AGEMA_signal_5999), .Q (new_AGEMA_signal_6000) ) ;
    buf_clk new_AGEMA_reg_buffer_2571 ( .C (clk), .D (new_AGEMA_signal_6001), .Q (new_AGEMA_signal_6002) ) ;
    buf_clk new_AGEMA_reg_buffer_2573 ( .C (clk), .D (new_AGEMA_signal_6003), .Q (new_AGEMA_signal_6004) ) ;
    buf_clk new_AGEMA_reg_buffer_2575 ( .C (clk), .D (new_AGEMA_signal_6005), .Q (new_AGEMA_signal_6006) ) ;
    buf_clk new_AGEMA_reg_buffer_2587 ( .C (clk), .D (new_AGEMA_signal_6017), .Q (new_AGEMA_signal_6018) ) ;
    buf_clk new_AGEMA_reg_buffer_2591 ( .C (clk), .D (new_AGEMA_signal_6021), .Q (new_AGEMA_signal_6022) ) ;
    buf_clk new_AGEMA_reg_buffer_2595 ( .C (clk), .D (new_AGEMA_signal_6025), .Q (new_AGEMA_signal_6026) ) ;
    buf_clk new_AGEMA_reg_buffer_2599 ( .C (clk), .D (new_AGEMA_signal_6029), .Q (new_AGEMA_signal_6030) ) ;
    buf_clk new_AGEMA_reg_buffer_2601 ( .C (clk), .D (new_AGEMA_signal_6031), .Q (new_AGEMA_signal_6032) ) ;
    buf_clk new_AGEMA_reg_buffer_2603 ( .C (clk), .D (new_AGEMA_signal_6033), .Q (new_AGEMA_signal_6034) ) ;
    buf_clk new_AGEMA_reg_buffer_2605 ( .C (clk), .D (new_AGEMA_signal_6035), .Q (new_AGEMA_signal_6036) ) ;
    buf_clk new_AGEMA_reg_buffer_2607 ( .C (clk), .D (new_AGEMA_signal_6037), .Q (new_AGEMA_signal_6038) ) ;
    buf_clk new_AGEMA_reg_buffer_2617 ( .C (clk), .D (new_AGEMA_signal_6047), .Q (new_AGEMA_signal_6048) ) ;
    buf_clk new_AGEMA_reg_buffer_2619 ( .C (clk), .D (new_AGEMA_signal_6049), .Q (new_AGEMA_signal_6050) ) ;
    buf_clk new_AGEMA_reg_buffer_2621 ( .C (clk), .D (new_AGEMA_signal_6051), .Q (new_AGEMA_signal_6052) ) ;
    buf_clk new_AGEMA_reg_buffer_2623 ( .C (clk), .D (new_AGEMA_signal_6053), .Q (new_AGEMA_signal_6054) ) ;
    buf_clk new_AGEMA_reg_buffer_2635 ( .C (clk), .D (new_AGEMA_signal_6065), .Q (new_AGEMA_signal_6066) ) ;
    buf_clk new_AGEMA_reg_buffer_2639 ( .C (clk), .D (new_AGEMA_signal_6069), .Q (new_AGEMA_signal_6070) ) ;
    buf_clk new_AGEMA_reg_buffer_2643 ( .C (clk), .D (new_AGEMA_signal_6073), .Q (new_AGEMA_signal_6074) ) ;
    buf_clk new_AGEMA_reg_buffer_2647 ( .C (clk), .D (new_AGEMA_signal_6077), .Q (new_AGEMA_signal_6078) ) ;
    buf_clk new_AGEMA_reg_buffer_2649 ( .C (clk), .D (new_AGEMA_signal_6079), .Q (new_AGEMA_signal_6080) ) ;
    buf_clk new_AGEMA_reg_buffer_2651 ( .C (clk), .D (new_AGEMA_signal_6081), .Q (new_AGEMA_signal_6082) ) ;
    buf_clk new_AGEMA_reg_buffer_2653 ( .C (clk), .D (new_AGEMA_signal_6083), .Q (new_AGEMA_signal_6084) ) ;
    buf_clk new_AGEMA_reg_buffer_2655 ( .C (clk), .D (new_AGEMA_signal_6085), .Q (new_AGEMA_signal_6086) ) ;
    buf_clk new_AGEMA_reg_buffer_2665 ( .C (clk), .D (new_AGEMA_signal_6095), .Q (new_AGEMA_signal_6096) ) ;
    buf_clk new_AGEMA_reg_buffer_2667 ( .C (clk), .D (new_AGEMA_signal_6097), .Q (new_AGEMA_signal_6098) ) ;
    buf_clk new_AGEMA_reg_buffer_2669 ( .C (clk), .D (new_AGEMA_signal_6099), .Q (new_AGEMA_signal_6100) ) ;
    buf_clk new_AGEMA_reg_buffer_2671 ( .C (clk), .D (new_AGEMA_signal_6101), .Q (new_AGEMA_signal_6102) ) ;
    buf_clk new_AGEMA_reg_buffer_2683 ( .C (clk), .D (new_AGEMA_signal_6113), .Q (new_AGEMA_signal_6114) ) ;
    buf_clk new_AGEMA_reg_buffer_2687 ( .C (clk), .D (new_AGEMA_signal_6117), .Q (new_AGEMA_signal_6118) ) ;
    buf_clk new_AGEMA_reg_buffer_2691 ( .C (clk), .D (new_AGEMA_signal_6121), .Q (new_AGEMA_signal_6122) ) ;
    buf_clk new_AGEMA_reg_buffer_2695 ( .C (clk), .D (new_AGEMA_signal_6125), .Q (new_AGEMA_signal_6126) ) ;
    buf_clk new_AGEMA_reg_buffer_2697 ( .C (clk), .D (new_AGEMA_signal_6127), .Q (new_AGEMA_signal_6128) ) ;
    buf_clk new_AGEMA_reg_buffer_2699 ( .C (clk), .D (new_AGEMA_signal_6129), .Q (new_AGEMA_signal_6130) ) ;
    buf_clk new_AGEMA_reg_buffer_2701 ( .C (clk), .D (new_AGEMA_signal_6131), .Q (new_AGEMA_signal_6132) ) ;
    buf_clk new_AGEMA_reg_buffer_2703 ( .C (clk), .D (new_AGEMA_signal_6133), .Q (new_AGEMA_signal_6134) ) ;
    buf_clk new_AGEMA_reg_buffer_2713 ( .C (clk), .D (new_AGEMA_signal_6143), .Q (new_AGEMA_signal_6144) ) ;
    buf_clk new_AGEMA_reg_buffer_2715 ( .C (clk), .D (new_AGEMA_signal_6145), .Q (new_AGEMA_signal_6146) ) ;
    buf_clk new_AGEMA_reg_buffer_2717 ( .C (clk), .D (new_AGEMA_signal_6147), .Q (new_AGEMA_signal_6148) ) ;
    buf_clk new_AGEMA_reg_buffer_2719 ( .C (clk), .D (new_AGEMA_signal_6149), .Q (new_AGEMA_signal_6150) ) ;
    buf_clk new_AGEMA_reg_buffer_2731 ( .C (clk), .D (new_AGEMA_signal_6161), .Q (new_AGEMA_signal_6162) ) ;
    buf_clk new_AGEMA_reg_buffer_2735 ( .C (clk), .D (new_AGEMA_signal_6165), .Q (new_AGEMA_signal_6166) ) ;
    buf_clk new_AGEMA_reg_buffer_2739 ( .C (clk), .D (new_AGEMA_signal_6169), .Q (new_AGEMA_signal_6170) ) ;
    buf_clk new_AGEMA_reg_buffer_2743 ( .C (clk), .D (new_AGEMA_signal_6173), .Q (new_AGEMA_signal_6174) ) ;
    buf_clk new_AGEMA_reg_buffer_2745 ( .C (clk), .D (new_AGEMA_signal_6175), .Q (new_AGEMA_signal_6176) ) ;
    buf_clk new_AGEMA_reg_buffer_2747 ( .C (clk), .D (new_AGEMA_signal_6177), .Q (new_AGEMA_signal_6178) ) ;
    buf_clk new_AGEMA_reg_buffer_2749 ( .C (clk), .D (new_AGEMA_signal_6179), .Q (new_AGEMA_signal_6180) ) ;
    buf_clk new_AGEMA_reg_buffer_2751 ( .C (clk), .D (new_AGEMA_signal_6181), .Q (new_AGEMA_signal_6182) ) ;
    buf_clk new_AGEMA_reg_buffer_2761 ( .C (clk), .D (new_AGEMA_signal_6191), .Q (new_AGEMA_signal_6192) ) ;
    buf_clk new_AGEMA_reg_buffer_2763 ( .C (clk), .D (new_AGEMA_signal_6193), .Q (new_AGEMA_signal_6194) ) ;
    buf_clk new_AGEMA_reg_buffer_2765 ( .C (clk), .D (new_AGEMA_signal_6195), .Q (new_AGEMA_signal_6196) ) ;
    buf_clk new_AGEMA_reg_buffer_2767 ( .C (clk), .D (new_AGEMA_signal_6197), .Q (new_AGEMA_signal_6198) ) ;
    buf_clk new_AGEMA_reg_buffer_2779 ( .C (clk), .D (new_AGEMA_signal_6209), .Q (new_AGEMA_signal_6210) ) ;
    buf_clk new_AGEMA_reg_buffer_2783 ( .C (clk), .D (new_AGEMA_signal_6213), .Q (new_AGEMA_signal_6214) ) ;
    buf_clk new_AGEMA_reg_buffer_2787 ( .C (clk), .D (new_AGEMA_signal_6217), .Q (new_AGEMA_signal_6218) ) ;
    buf_clk new_AGEMA_reg_buffer_2791 ( .C (clk), .D (new_AGEMA_signal_6221), .Q (new_AGEMA_signal_6222) ) ;
    buf_clk new_AGEMA_reg_buffer_2793 ( .C (clk), .D (new_AGEMA_signal_6223), .Q (new_AGEMA_signal_6224) ) ;
    buf_clk new_AGEMA_reg_buffer_2795 ( .C (clk), .D (new_AGEMA_signal_6225), .Q (new_AGEMA_signal_6226) ) ;
    buf_clk new_AGEMA_reg_buffer_2797 ( .C (clk), .D (new_AGEMA_signal_6227), .Q (new_AGEMA_signal_6228) ) ;
    buf_clk new_AGEMA_reg_buffer_2799 ( .C (clk), .D (new_AGEMA_signal_6229), .Q (new_AGEMA_signal_6230) ) ;
    buf_clk new_AGEMA_reg_buffer_2809 ( .C (clk), .D (new_AGEMA_signal_6239), .Q (new_AGEMA_signal_6240) ) ;
    buf_clk new_AGEMA_reg_buffer_2811 ( .C (clk), .D (new_AGEMA_signal_6241), .Q (new_AGEMA_signal_6242) ) ;
    buf_clk new_AGEMA_reg_buffer_2813 ( .C (clk), .D (new_AGEMA_signal_6243), .Q (new_AGEMA_signal_6244) ) ;
    buf_clk new_AGEMA_reg_buffer_2815 ( .C (clk), .D (new_AGEMA_signal_6245), .Q (new_AGEMA_signal_6246) ) ;
    buf_clk new_AGEMA_reg_buffer_2827 ( .C (clk), .D (new_AGEMA_signal_6257), .Q (new_AGEMA_signal_6258) ) ;
    buf_clk new_AGEMA_reg_buffer_2831 ( .C (clk), .D (new_AGEMA_signal_6261), .Q (new_AGEMA_signal_6262) ) ;
    buf_clk new_AGEMA_reg_buffer_2835 ( .C (clk), .D (new_AGEMA_signal_6265), .Q (new_AGEMA_signal_6266) ) ;
    buf_clk new_AGEMA_reg_buffer_2839 ( .C (clk), .D (new_AGEMA_signal_6269), .Q (new_AGEMA_signal_6270) ) ;
    buf_clk new_AGEMA_reg_buffer_2841 ( .C (clk), .D (new_AGEMA_signal_6271), .Q (new_AGEMA_signal_6272) ) ;
    buf_clk new_AGEMA_reg_buffer_2843 ( .C (clk), .D (new_AGEMA_signal_6273), .Q (new_AGEMA_signal_6274) ) ;
    buf_clk new_AGEMA_reg_buffer_2845 ( .C (clk), .D (new_AGEMA_signal_6275), .Q (new_AGEMA_signal_6276) ) ;
    buf_clk new_AGEMA_reg_buffer_2847 ( .C (clk), .D (new_AGEMA_signal_6277), .Q (new_AGEMA_signal_6278) ) ;
    buf_clk new_AGEMA_reg_buffer_2857 ( .C (clk), .D (new_AGEMA_signal_6287), .Q (new_AGEMA_signal_6288) ) ;
    buf_clk new_AGEMA_reg_buffer_2859 ( .C (clk), .D (new_AGEMA_signal_6289), .Q (new_AGEMA_signal_6290) ) ;
    buf_clk new_AGEMA_reg_buffer_2861 ( .C (clk), .D (new_AGEMA_signal_6291), .Q (new_AGEMA_signal_6292) ) ;
    buf_clk new_AGEMA_reg_buffer_2863 ( .C (clk), .D (new_AGEMA_signal_6293), .Q (new_AGEMA_signal_6294) ) ;
    buf_clk new_AGEMA_reg_buffer_2875 ( .C (clk), .D (new_AGEMA_signal_6305), .Q (new_AGEMA_signal_6306) ) ;
    buf_clk new_AGEMA_reg_buffer_2879 ( .C (clk), .D (new_AGEMA_signal_6309), .Q (new_AGEMA_signal_6310) ) ;
    buf_clk new_AGEMA_reg_buffer_2883 ( .C (clk), .D (new_AGEMA_signal_6313), .Q (new_AGEMA_signal_6314) ) ;
    buf_clk new_AGEMA_reg_buffer_2887 ( .C (clk), .D (new_AGEMA_signal_6317), .Q (new_AGEMA_signal_6318) ) ;
    buf_clk new_AGEMA_reg_buffer_2889 ( .C (clk), .D (new_AGEMA_signal_6319), .Q (new_AGEMA_signal_6320) ) ;
    buf_clk new_AGEMA_reg_buffer_2891 ( .C (clk), .D (new_AGEMA_signal_6321), .Q (new_AGEMA_signal_6322) ) ;
    buf_clk new_AGEMA_reg_buffer_2893 ( .C (clk), .D (new_AGEMA_signal_6323), .Q (new_AGEMA_signal_6324) ) ;
    buf_clk new_AGEMA_reg_buffer_2895 ( .C (clk), .D (new_AGEMA_signal_6325), .Q (new_AGEMA_signal_6326) ) ;
    buf_clk new_AGEMA_reg_buffer_2905 ( .C (clk), .D (new_AGEMA_signal_6335), .Q (new_AGEMA_signal_6336) ) ;
    buf_clk new_AGEMA_reg_buffer_2907 ( .C (clk), .D (new_AGEMA_signal_6337), .Q (new_AGEMA_signal_6338) ) ;
    buf_clk new_AGEMA_reg_buffer_2909 ( .C (clk), .D (new_AGEMA_signal_6339), .Q (new_AGEMA_signal_6340) ) ;
    buf_clk new_AGEMA_reg_buffer_2911 ( .C (clk), .D (new_AGEMA_signal_6341), .Q (new_AGEMA_signal_6342) ) ;
    buf_clk new_AGEMA_reg_buffer_2923 ( .C (clk), .D (new_AGEMA_signal_6353), .Q (new_AGEMA_signal_6354) ) ;
    buf_clk new_AGEMA_reg_buffer_2927 ( .C (clk), .D (new_AGEMA_signal_6357), .Q (new_AGEMA_signal_6358) ) ;
    buf_clk new_AGEMA_reg_buffer_2931 ( .C (clk), .D (new_AGEMA_signal_6361), .Q (new_AGEMA_signal_6362) ) ;
    buf_clk new_AGEMA_reg_buffer_2935 ( .C (clk), .D (new_AGEMA_signal_6365), .Q (new_AGEMA_signal_6366) ) ;
    buf_clk new_AGEMA_reg_buffer_2937 ( .C (clk), .D (new_AGEMA_signal_6367), .Q (new_AGEMA_signal_6368) ) ;
    buf_clk new_AGEMA_reg_buffer_2939 ( .C (clk), .D (new_AGEMA_signal_6369), .Q (new_AGEMA_signal_6370) ) ;
    buf_clk new_AGEMA_reg_buffer_2941 ( .C (clk), .D (new_AGEMA_signal_6371), .Q (new_AGEMA_signal_6372) ) ;
    buf_clk new_AGEMA_reg_buffer_2943 ( .C (clk), .D (new_AGEMA_signal_6373), .Q (new_AGEMA_signal_6374) ) ;
    buf_clk new_AGEMA_reg_buffer_2953 ( .C (clk), .D (new_AGEMA_signal_6383), .Q (new_AGEMA_signal_6384) ) ;
    buf_clk new_AGEMA_reg_buffer_2955 ( .C (clk), .D (new_AGEMA_signal_6385), .Q (new_AGEMA_signal_6386) ) ;
    buf_clk new_AGEMA_reg_buffer_2957 ( .C (clk), .D (new_AGEMA_signal_6387), .Q (new_AGEMA_signal_6388) ) ;
    buf_clk new_AGEMA_reg_buffer_2959 ( .C (clk), .D (new_AGEMA_signal_6389), .Q (new_AGEMA_signal_6390) ) ;
    buf_clk new_AGEMA_reg_buffer_2971 ( .C (clk), .D (new_AGEMA_signal_6401), .Q (new_AGEMA_signal_6402) ) ;
    buf_clk new_AGEMA_reg_buffer_2975 ( .C (clk), .D (new_AGEMA_signal_6405), .Q (new_AGEMA_signal_6406) ) ;
    buf_clk new_AGEMA_reg_buffer_2979 ( .C (clk), .D (new_AGEMA_signal_6409), .Q (new_AGEMA_signal_6410) ) ;
    buf_clk new_AGEMA_reg_buffer_2983 ( .C (clk), .D (new_AGEMA_signal_6413), .Q (new_AGEMA_signal_6414) ) ;
    buf_clk new_AGEMA_reg_buffer_2985 ( .C (clk), .D (new_AGEMA_signal_6415), .Q (new_AGEMA_signal_6416) ) ;
    buf_clk new_AGEMA_reg_buffer_2987 ( .C (clk), .D (new_AGEMA_signal_6417), .Q (new_AGEMA_signal_6418) ) ;
    buf_clk new_AGEMA_reg_buffer_2989 ( .C (clk), .D (new_AGEMA_signal_6419), .Q (new_AGEMA_signal_6420) ) ;
    buf_clk new_AGEMA_reg_buffer_2991 ( .C (clk), .D (new_AGEMA_signal_6421), .Q (new_AGEMA_signal_6422) ) ;
    buf_clk new_AGEMA_reg_buffer_3001 ( .C (clk), .D (new_AGEMA_signal_6431), .Q (new_AGEMA_signal_6432) ) ;
    buf_clk new_AGEMA_reg_buffer_3003 ( .C (clk), .D (new_AGEMA_signal_6433), .Q (new_AGEMA_signal_6434) ) ;
    buf_clk new_AGEMA_reg_buffer_3005 ( .C (clk), .D (new_AGEMA_signal_6435), .Q (new_AGEMA_signal_6436) ) ;
    buf_clk new_AGEMA_reg_buffer_3007 ( .C (clk), .D (new_AGEMA_signal_6437), .Q (new_AGEMA_signal_6438) ) ;
    buf_clk new_AGEMA_reg_buffer_3019 ( .C (clk), .D (new_AGEMA_signal_6449), .Q (new_AGEMA_signal_6450) ) ;
    buf_clk new_AGEMA_reg_buffer_3023 ( .C (clk), .D (new_AGEMA_signal_6453), .Q (new_AGEMA_signal_6454) ) ;
    buf_clk new_AGEMA_reg_buffer_3027 ( .C (clk), .D (new_AGEMA_signal_6457), .Q (new_AGEMA_signal_6458) ) ;
    buf_clk new_AGEMA_reg_buffer_3031 ( .C (clk), .D (new_AGEMA_signal_6461), .Q (new_AGEMA_signal_6462) ) ;
    buf_clk new_AGEMA_reg_buffer_3033 ( .C (clk), .D (new_AGEMA_signal_6463), .Q (new_AGEMA_signal_6464) ) ;
    buf_clk new_AGEMA_reg_buffer_3035 ( .C (clk), .D (new_AGEMA_signal_6465), .Q (new_AGEMA_signal_6466) ) ;
    buf_clk new_AGEMA_reg_buffer_3037 ( .C (clk), .D (new_AGEMA_signal_6467), .Q (new_AGEMA_signal_6468) ) ;
    buf_clk new_AGEMA_reg_buffer_3039 ( .C (clk), .D (new_AGEMA_signal_6469), .Q (new_AGEMA_signal_6470) ) ;
    buf_clk new_AGEMA_reg_buffer_3049 ( .C (clk), .D (new_AGEMA_signal_6479), .Q (new_AGEMA_signal_6480) ) ;
    buf_clk new_AGEMA_reg_buffer_3051 ( .C (clk), .D (new_AGEMA_signal_6481), .Q (new_AGEMA_signal_6482) ) ;
    buf_clk new_AGEMA_reg_buffer_3053 ( .C (clk), .D (new_AGEMA_signal_6483), .Q (new_AGEMA_signal_6484) ) ;
    buf_clk new_AGEMA_reg_buffer_3055 ( .C (clk), .D (new_AGEMA_signal_6485), .Q (new_AGEMA_signal_6486) ) ;
    buf_clk new_AGEMA_reg_buffer_3067 ( .C (clk), .D (new_AGEMA_signal_6497), .Q (new_AGEMA_signal_6498) ) ;
    buf_clk new_AGEMA_reg_buffer_3071 ( .C (clk), .D (new_AGEMA_signal_6501), .Q (new_AGEMA_signal_6502) ) ;
    buf_clk new_AGEMA_reg_buffer_3075 ( .C (clk), .D (new_AGEMA_signal_6505), .Q (new_AGEMA_signal_6506) ) ;
    buf_clk new_AGEMA_reg_buffer_3079 ( .C (clk), .D (new_AGEMA_signal_6509), .Q (new_AGEMA_signal_6510) ) ;
    buf_clk new_AGEMA_reg_buffer_3081 ( .C (clk), .D (new_AGEMA_signal_6511), .Q (new_AGEMA_signal_6512) ) ;
    buf_clk new_AGEMA_reg_buffer_3083 ( .C (clk), .D (new_AGEMA_signal_6513), .Q (new_AGEMA_signal_6514) ) ;
    buf_clk new_AGEMA_reg_buffer_3085 ( .C (clk), .D (new_AGEMA_signal_6515), .Q (new_AGEMA_signal_6516) ) ;
    buf_clk new_AGEMA_reg_buffer_3087 ( .C (clk), .D (new_AGEMA_signal_6517), .Q (new_AGEMA_signal_6518) ) ;
    buf_clk new_AGEMA_reg_buffer_3097 ( .C (clk), .D (new_AGEMA_signal_6527), .Q (new_AGEMA_signal_6528) ) ;
    buf_clk new_AGEMA_reg_buffer_3099 ( .C (clk), .D (new_AGEMA_signal_6529), .Q (new_AGEMA_signal_6530) ) ;
    buf_clk new_AGEMA_reg_buffer_3101 ( .C (clk), .D (new_AGEMA_signal_6531), .Q (new_AGEMA_signal_6532) ) ;
    buf_clk new_AGEMA_reg_buffer_3103 ( .C (clk), .D (new_AGEMA_signal_6533), .Q (new_AGEMA_signal_6534) ) ;
    buf_clk new_AGEMA_reg_buffer_3115 ( .C (clk), .D (new_AGEMA_signal_6545), .Q (new_AGEMA_signal_6546) ) ;
    buf_clk new_AGEMA_reg_buffer_3119 ( .C (clk), .D (new_AGEMA_signal_6549), .Q (new_AGEMA_signal_6550) ) ;
    buf_clk new_AGEMA_reg_buffer_3123 ( .C (clk), .D (new_AGEMA_signal_6553), .Q (new_AGEMA_signal_6554) ) ;
    buf_clk new_AGEMA_reg_buffer_3127 ( .C (clk), .D (new_AGEMA_signal_6557), .Q (new_AGEMA_signal_6558) ) ;
    buf_clk new_AGEMA_reg_buffer_3129 ( .C (clk), .D (new_AGEMA_signal_6559), .Q (new_AGEMA_signal_6560) ) ;
    buf_clk new_AGEMA_reg_buffer_3131 ( .C (clk), .D (new_AGEMA_signal_6561), .Q (new_AGEMA_signal_6562) ) ;
    buf_clk new_AGEMA_reg_buffer_3133 ( .C (clk), .D (new_AGEMA_signal_6563), .Q (new_AGEMA_signal_6564) ) ;
    buf_clk new_AGEMA_reg_buffer_3135 ( .C (clk), .D (new_AGEMA_signal_6565), .Q (new_AGEMA_signal_6566) ) ;
    buf_clk new_AGEMA_reg_buffer_3145 ( .C (clk), .D (new_AGEMA_signal_6575), .Q (new_AGEMA_signal_6576) ) ;
    buf_clk new_AGEMA_reg_buffer_3147 ( .C (clk), .D (new_AGEMA_signal_6577), .Q (new_AGEMA_signal_6578) ) ;
    buf_clk new_AGEMA_reg_buffer_3149 ( .C (clk), .D (new_AGEMA_signal_6579), .Q (new_AGEMA_signal_6580) ) ;
    buf_clk new_AGEMA_reg_buffer_3151 ( .C (clk), .D (new_AGEMA_signal_6581), .Q (new_AGEMA_signal_6582) ) ;
    buf_clk new_AGEMA_reg_buffer_3163 ( .C (clk), .D (new_AGEMA_signal_6593), .Q (new_AGEMA_signal_6594) ) ;
    buf_clk new_AGEMA_reg_buffer_3167 ( .C (clk), .D (new_AGEMA_signal_6597), .Q (new_AGEMA_signal_6598) ) ;
    buf_clk new_AGEMA_reg_buffer_3171 ( .C (clk), .D (new_AGEMA_signal_6601), .Q (new_AGEMA_signal_6602) ) ;
    buf_clk new_AGEMA_reg_buffer_3175 ( .C (clk), .D (new_AGEMA_signal_6605), .Q (new_AGEMA_signal_6606) ) ;
    buf_clk new_AGEMA_reg_buffer_3177 ( .C (clk), .D (new_AGEMA_signal_6607), .Q (new_AGEMA_signal_6608) ) ;
    buf_clk new_AGEMA_reg_buffer_3179 ( .C (clk), .D (new_AGEMA_signal_6609), .Q (new_AGEMA_signal_6610) ) ;
    buf_clk new_AGEMA_reg_buffer_3181 ( .C (clk), .D (new_AGEMA_signal_6611), .Q (new_AGEMA_signal_6612) ) ;
    buf_clk new_AGEMA_reg_buffer_3183 ( .C (clk), .D (new_AGEMA_signal_6613), .Q (new_AGEMA_signal_6614) ) ;
    buf_clk new_AGEMA_reg_buffer_3187 ( .C (clk), .D (new_AGEMA_signal_6617), .Q (new_AGEMA_signal_6618) ) ;
    buf_clk new_AGEMA_reg_buffer_3191 ( .C (clk), .D (new_AGEMA_signal_6621), .Q (new_AGEMA_signal_6622) ) ;
    buf_clk new_AGEMA_reg_buffer_3195 ( .C (clk), .D (new_AGEMA_signal_6625), .Q (new_AGEMA_signal_6626) ) ;
    buf_clk new_AGEMA_reg_buffer_3199 ( .C (clk), .D (new_AGEMA_signal_6629), .Q (new_AGEMA_signal_6630) ) ;
    buf_clk new_AGEMA_reg_buffer_3203 ( .C (clk), .D (new_AGEMA_signal_6633), .Q (new_AGEMA_signal_6634) ) ;
    buf_clk new_AGEMA_reg_buffer_3207 ( .C (clk), .D (new_AGEMA_signal_6637), .Q (new_AGEMA_signal_6638) ) ;
    buf_clk new_AGEMA_reg_buffer_3211 ( .C (clk), .D (new_AGEMA_signal_6641), .Q (new_AGEMA_signal_6642) ) ;
    buf_clk new_AGEMA_reg_buffer_3215 ( .C (clk), .D (new_AGEMA_signal_6645), .Q (new_AGEMA_signal_6646) ) ;
    buf_clk new_AGEMA_reg_buffer_3219 ( .C (clk), .D (new_AGEMA_signal_6649), .Q (new_AGEMA_signal_6650) ) ;
    buf_clk new_AGEMA_reg_buffer_3223 ( .C (clk), .D (new_AGEMA_signal_6653), .Q (new_AGEMA_signal_6654) ) ;
    buf_clk new_AGEMA_reg_buffer_3227 ( .C (clk), .D (new_AGEMA_signal_6657), .Q (new_AGEMA_signal_6658) ) ;
    buf_clk new_AGEMA_reg_buffer_3231 ( .C (clk), .D (new_AGEMA_signal_6661), .Q (new_AGEMA_signal_6662) ) ;
    buf_clk new_AGEMA_reg_buffer_3235 ( .C (clk), .D (new_AGEMA_signal_6665), .Q (new_AGEMA_signal_6666) ) ;
    buf_clk new_AGEMA_reg_buffer_3239 ( .C (clk), .D (new_AGEMA_signal_6669), .Q (new_AGEMA_signal_6670) ) ;
    buf_clk new_AGEMA_reg_buffer_3243 ( .C (clk), .D (new_AGEMA_signal_6673), .Q (new_AGEMA_signal_6674) ) ;
    buf_clk new_AGEMA_reg_buffer_3247 ( .C (clk), .D (new_AGEMA_signal_6677), .Q (new_AGEMA_signal_6678) ) ;
    buf_clk new_AGEMA_reg_buffer_3251 ( .C (clk), .D (new_AGEMA_signal_6681), .Q (new_AGEMA_signal_6682) ) ;
    buf_clk new_AGEMA_reg_buffer_3255 ( .C (clk), .D (new_AGEMA_signal_6685), .Q (new_AGEMA_signal_6686) ) ;
    buf_clk new_AGEMA_reg_buffer_3259 ( .C (clk), .D (new_AGEMA_signal_6689), .Q (new_AGEMA_signal_6690) ) ;
    buf_clk new_AGEMA_reg_buffer_3263 ( .C (clk), .D (new_AGEMA_signal_6693), .Q (new_AGEMA_signal_6694) ) ;
    buf_clk new_AGEMA_reg_buffer_3267 ( .C (clk), .D (new_AGEMA_signal_6697), .Q (new_AGEMA_signal_6698) ) ;
    buf_clk new_AGEMA_reg_buffer_3271 ( .C (clk), .D (new_AGEMA_signal_6701), .Q (new_AGEMA_signal_6702) ) ;
    buf_clk new_AGEMA_reg_buffer_3275 ( .C (clk), .D (new_AGEMA_signal_6705), .Q (new_AGEMA_signal_6706) ) ;
    buf_clk new_AGEMA_reg_buffer_3279 ( .C (clk), .D (new_AGEMA_signal_6709), .Q (new_AGEMA_signal_6710) ) ;
    buf_clk new_AGEMA_reg_buffer_3283 ( .C (clk), .D (new_AGEMA_signal_6713), .Q (new_AGEMA_signal_6714) ) ;
    buf_clk new_AGEMA_reg_buffer_3287 ( .C (clk), .D (new_AGEMA_signal_6717), .Q (new_AGEMA_signal_6718) ) ;
    buf_clk new_AGEMA_reg_buffer_3291 ( .C (clk), .D (new_AGEMA_signal_6721), .Q (new_AGEMA_signal_6722) ) ;
    buf_clk new_AGEMA_reg_buffer_3295 ( .C (clk), .D (new_AGEMA_signal_6725), .Q (new_AGEMA_signal_6726) ) ;
    buf_clk new_AGEMA_reg_buffer_3299 ( .C (clk), .D (new_AGEMA_signal_6729), .Q (new_AGEMA_signal_6730) ) ;
    buf_clk new_AGEMA_reg_buffer_3303 ( .C (clk), .D (new_AGEMA_signal_6733), .Q (new_AGEMA_signal_6734) ) ;
    buf_clk new_AGEMA_reg_buffer_3307 ( .C (clk), .D (new_AGEMA_signal_6737), .Q (new_AGEMA_signal_6738) ) ;
    buf_clk new_AGEMA_reg_buffer_3311 ( .C (clk), .D (new_AGEMA_signal_6741), .Q (new_AGEMA_signal_6742) ) ;
    buf_clk new_AGEMA_reg_buffer_3315 ( .C (clk), .D (new_AGEMA_signal_6745), .Q (new_AGEMA_signal_6746) ) ;
    buf_clk new_AGEMA_reg_buffer_3319 ( .C (clk), .D (new_AGEMA_signal_6749), .Q (new_AGEMA_signal_6750) ) ;
    buf_clk new_AGEMA_reg_buffer_3323 ( .C (clk), .D (new_AGEMA_signal_6753), .Q (new_AGEMA_signal_6754) ) ;
    buf_clk new_AGEMA_reg_buffer_3327 ( .C (clk), .D (new_AGEMA_signal_6757), .Q (new_AGEMA_signal_6758) ) ;
    buf_clk new_AGEMA_reg_buffer_3331 ( .C (clk), .D (new_AGEMA_signal_6761), .Q (new_AGEMA_signal_6762) ) ;
    buf_clk new_AGEMA_reg_buffer_3335 ( .C (clk), .D (new_AGEMA_signal_6765), .Q (new_AGEMA_signal_6766) ) ;
    buf_clk new_AGEMA_reg_buffer_3339 ( .C (clk), .D (new_AGEMA_signal_6769), .Q (new_AGEMA_signal_6770) ) ;
    buf_clk new_AGEMA_reg_buffer_3343 ( .C (clk), .D (new_AGEMA_signal_6773), .Q (new_AGEMA_signal_6774) ) ;
    buf_clk new_AGEMA_reg_buffer_3347 ( .C (clk), .D (new_AGEMA_signal_6777), .Q (new_AGEMA_signal_6778) ) ;
    buf_clk new_AGEMA_reg_buffer_3351 ( .C (clk), .D (new_AGEMA_signal_6781), .Q (new_AGEMA_signal_6782) ) ;
    buf_clk new_AGEMA_reg_buffer_3355 ( .C (clk), .D (new_AGEMA_signal_6785), .Q (new_AGEMA_signal_6786) ) ;
    buf_clk new_AGEMA_reg_buffer_3359 ( .C (clk), .D (new_AGEMA_signal_6789), .Q (new_AGEMA_signal_6790) ) ;
    buf_clk new_AGEMA_reg_buffer_3363 ( .C (clk), .D (new_AGEMA_signal_6793), .Q (new_AGEMA_signal_6794) ) ;
    buf_clk new_AGEMA_reg_buffer_3367 ( .C (clk), .D (new_AGEMA_signal_6797), .Q (new_AGEMA_signal_6798) ) ;
    buf_clk new_AGEMA_reg_buffer_3371 ( .C (clk), .D (new_AGEMA_signal_6801), .Q (new_AGEMA_signal_6802) ) ;
    buf_clk new_AGEMA_reg_buffer_3375 ( .C (clk), .D (new_AGEMA_signal_6805), .Q (new_AGEMA_signal_6806) ) ;
    buf_clk new_AGEMA_reg_buffer_3379 ( .C (clk), .D (new_AGEMA_signal_6809), .Q (new_AGEMA_signal_6810) ) ;
    buf_clk new_AGEMA_reg_buffer_3383 ( .C (clk), .D (new_AGEMA_signal_6813), .Q (new_AGEMA_signal_6814) ) ;
    buf_clk new_AGEMA_reg_buffer_3387 ( .C (clk), .D (new_AGEMA_signal_6817), .Q (new_AGEMA_signal_6818) ) ;
    buf_clk new_AGEMA_reg_buffer_3391 ( .C (clk), .D (new_AGEMA_signal_6821), .Q (new_AGEMA_signal_6822) ) ;
    buf_clk new_AGEMA_reg_buffer_3395 ( .C (clk), .D (new_AGEMA_signal_6825), .Q (new_AGEMA_signal_6826) ) ;
    buf_clk new_AGEMA_reg_buffer_3399 ( .C (clk), .D (new_AGEMA_signal_6829), .Q (new_AGEMA_signal_6830) ) ;
    buf_clk new_AGEMA_reg_buffer_3403 ( .C (clk), .D (new_AGEMA_signal_6833), .Q (new_AGEMA_signal_6834) ) ;
    buf_clk new_AGEMA_reg_buffer_3407 ( .C (clk), .D (new_AGEMA_signal_6837), .Q (new_AGEMA_signal_6838) ) ;
    buf_clk new_AGEMA_reg_buffer_3411 ( .C (clk), .D (new_AGEMA_signal_6841), .Q (new_AGEMA_signal_6842) ) ;
    buf_clk new_AGEMA_reg_buffer_3415 ( .C (clk), .D (new_AGEMA_signal_6845), .Q (new_AGEMA_signal_6846) ) ;
    buf_clk new_AGEMA_reg_buffer_3419 ( .C (clk), .D (new_AGEMA_signal_6849), .Q (new_AGEMA_signal_6850) ) ;
    buf_clk new_AGEMA_reg_buffer_3423 ( .C (clk), .D (new_AGEMA_signal_6853), .Q (new_AGEMA_signal_6854) ) ;
    buf_clk new_AGEMA_reg_buffer_3427 ( .C (clk), .D (new_AGEMA_signal_6857), .Q (new_AGEMA_signal_6858) ) ;
    buf_clk new_AGEMA_reg_buffer_3431 ( .C (clk), .D (new_AGEMA_signal_6861), .Q (new_AGEMA_signal_6862) ) ;
    buf_clk new_AGEMA_reg_buffer_3435 ( .C (clk), .D (new_AGEMA_signal_6865), .Q (new_AGEMA_signal_6866) ) ;
    buf_clk new_AGEMA_reg_buffer_3439 ( .C (clk), .D (new_AGEMA_signal_6869), .Q (new_AGEMA_signal_6870) ) ;
    buf_clk new_AGEMA_reg_buffer_3443 ( .C (clk), .D (new_AGEMA_signal_6873), .Q (new_AGEMA_signal_6874) ) ;
    buf_clk new_AGEMA_reg_buffer_3447 ( .C (clk), .D (new_AGEMA_signal_6877), .Q (new_AGEMA_signal_6878) ) ;
    buf_clk new_AGEMA_reg_buffer_3451 ( .C (clk), .D (new_AGEMA_signal_6881), .Q (new_AGEMA_signal_6882) ) ;
    buf_clk new_AGEMA_reg_buffer_3455 ( .C (clk), .D (new_AGEMA_signal_6885), .Q (new_AGEMA_signal_6886) ) ;
    buf_clk new_AGEMA_reg_buffer_3457 ( .C (clk), .D (new_AGEMA_signal_6887), .Q (new_AGEMA_signal_6888) ) ;
    buf_clk new_AGEMA_reg_buffer_3459 ( .C (clk), .D (new_AGEMA_signal_6889), .Q (new_AGEMA_signal_6890) ) ;
    buf_clk new_AGEMA_reg_buffer_3461 ( .C (clk), .D (new_AGEMA_signal_6891), .Q (new_AGEMA_signal_6892) ) ;
    buf_clk new_AGEMA_reg_buffer_3463 ( .C (clk), .D (new_AGEMA_signal_6893), .Q (new_AGEMA_signal_6894) ) ;
    buf_clk new_AGEMA_reg_buffer_3465 ( .C (clk), .D (new_AGEMA_signal_6895), .Q (new_AGEMA_signal_6896) ) ;
    buf_clk new_AGEMA_reg_buffer_3467 ( .C (clk), .D (new_AGEMA_signal_6897), .Q (new_AGEMA_signal_6898) ) ;
    buf_clk new_AGEMA_reg_buffer_3469 ( .C (clk), .D (new_AGEMA_signal_6899), .Q (new_AGEMA_signal_6900) ) ;
    buf_clk new_AGEMA_reg_buffer_3471 ( .C (clk), .D (new_AGEMA_signal_6901), .Q (new_AGEMA_signal_6902) ) ;
    buf_clk new_AGEMA_reg_buffer_3473 ( .C (clk), .D (new_AGEMA_signal_6903), .Q (new_AGEMA_signal_6904) ) ;
    buf_clk new_AGEMA_reg_buffer_3475 ( .C (clk), .D (new_AGEMA_signal_6905), .Q (new_AGEMA_signal_6906) ) ;
    buf_clk new_AGEMA_reg_buffer_3477 ( .C (clk), .D (new_AGEMA_signal_6907), .Q (new_AGEMA_signal_6908) ) ;
    buf_clk new_AGEMA_reg_buffer_3479 ( .C (clk), .D (new_AGEMA_signal_6909), .Q (new_AGEMA_signal_6910) ) ;
    buf_clk new_AGEMA_reg_buffer_3481 ( .C (clk), .D (new_AGEMA_signal_6911), .Q (new_AGEMA_signal_6912) ) ;
    buf_clk new_AGEMA_reg_buffer_3483 ( .C (clk), .D (new_AGEMA_signal_6913), .Q (new_AGEMA_signal_6914) ) ;
    buf_clk new_AGEMA_reg_buffer_3485 ( .C (clk), .D (new_AGEMA_signal_6915), .Q (new_AGEMA_signal_6916) ) ;
    buf_clk new_AGEMA_reg_buffer_3487 ( .C (clk), .D (new_AGEMA_signal_6917), .Q (new_AGEMA_signal_6918) ) ;
    buf_clk new_AGEMA_reg_buffer_3489 ( .C (clk), .D (new_AGEMA_signal_6919), .Q (new_AGEMA_signal_6920) ) ;
    buf_clk new_AGEMA_reg_buffer_3491 ( .C (clk), .D (new_AGEMA_signal_6921), .Q (new_AGEMA_signal_6922) ) ;
    buf_clk new_AGEMA_reg_buffer_3493 ( .C (clk), .D (new_AGEMA_signal_6923), .Q (new_AGEMA_signal_6924) ) ;
    buf_clk new_AGEMA_reg_buffer_3495 ( .C (clk), .D (new_AGEMA_signal_6925), .Q (new_AGEMA_signal_6926) ) ;
    buf_clk new_AGEMA_reg_buffer_3497 ( .C (clk), .D (new_AGEMA_signal_6927), .Q (new_AGEMA_signal_6928) ) ;
    buf_clk new_AGEMA_reg_buffer_3499 ( .C (clk), .D (new_AGEMA_signal_6929), .Q (new_AGEMA_signal_6930) ) ;
    buf_clk new_AGEMA_reg_buffer_3501 ( .C (clk), .D (new_AGEMA_signal_6931), .Q (new_AGEMA_signal_6932) ) ;
    buf_clk new_AGEMA_reg_buffer_3503 ( .C (clk), .D (new_AGEMA_signal_6933), .Q (new_AGEMA_signal_6934) ) ;
    buf_clk new_AGEMA_reg_buffer_3505 ( .C (clk), .D (new_AGEMA_signal_6935), .Q (new_AGEMA_signal_6936) ) ;
    buf_clk new_AGEMA_reg_buffer_3507 ( .C (clk), .D (new_AGEMA_signal_6937), .Q (new_AGEMA_signal_6938) ) ;
    buf_clk new_AGEMA_reg_buffer_3509 ( .C (clk), .D (new_AGEMA_signal_6939), .Q (new_AGEMA_signal_6940) ) ;
    buf_clk new_AGEMA_reg_buffer_3511 ( .C (clk), .D (new_AGEMA_signal_6941), .Q (new_AGEMA_signal_6942) ) ;
    buf_clk new_AGEMA_reg_buffer_3513 ( .C (clk), .D (new_AGEMA_signal_6943), .Q (new_AGEMA_signal_6944) ) ;
    buf_clk new_AGEMA_reg_buffer_3515 ( .C (clk), .D (new_AGEMA_signal_6945), .Q (new_AGEMA_signal_6946) ) ;
    buf_clk new_AGEMA_reg_buffer_3517 ( .C (clk), .D (new_AGEMA_signal_6947), .Q (new_AGEMA_signal_6948) ) ;
    buf_clk new_AGEMA_reg_buffer_3519 ( .C (clk), .D (new_AGEMA_signal_6949), .Q (new_AGEMA_signal_6950) ) ;
    buf_clk new_AGEMA_reg_buffer_3521 ( .C (clk), .D (new_AGEMA_signal_6951), .Q (new_AGEMA_signal_6952) ) ;
    buf_clk new_AGEMA_reg_buffer_3523 ( .C (clk), .D (new_AGEMA_signal_6953), .Q (new_AGEMA_signal_6954) ) ;
    buf_clk new_AGEMA_reg_buffer_3525 ( .C (clk), .D (new_AGEMA_signal_6955), .Q (new_AGEMA_signal_6956) ) ;
    buf_clk new_AGEMA_reg_buffer_3527 ( .C (clk), .D (new_AGEMA_signal_6957), .Q (new_AGEMA_signal_6958) ) ;
    buf_clk new_AGEMA_reg_buffer_3529 ( .C (clk), .D (new_AGEMA_signal_6959), .Q (new_AGEMA_signal_6960) ) ;
    buf_clk new_AGEMA_reg_buffer_3531 ( .C (clk), .D (new_AGEMA_signal_6961), .Q (new_AGEMA_signal_6962) ) ;
    buf_clk new_AGEMA_reg_buffer_3533 ( .C (clk), .D (new_AGEMA_signal_6963), .Q (new_AGEMA_signal_6964) ) ;
    buf_clk new_AGEMA_reg_buffer_3535 ( .C (clk), .D (new_AGEMA_signal_6965), .Q (new_AGEMA_signal_6966) ) ;
    buf_clk new_AGEMA_reg_buffer_3537 ( .C (clk), .D (new_AGEMA_signal_6967), .Q (new_AGEMA_signal_6968) ) ;
    buf_clk new_AGEMA_reg_buffer_3539 ( .C (clk), .D (new_AGEMA_signal_6969), .Q (new_AGEMA_signal_6970) ) ;
    buf_clk new_AGEMA_reg_buffer_3541 ( .C (clk), .D (new_AGEMA_signal_6971), .Q (new_AGEMA_signal_6972) ) ;
    buf_clk new_AGEMA_reg_buffer_3543 ( .C (clk), .D (new_AGEMA_signal_6973), .Q (new_AGEMA_signal_6974) ) ;
    buf_clk new_AGEMA_reg_buffer_3545 ( .C (clk), .D (new_AGEMA_signal_6975), .Q (new_AGEMA_signal_6976) ) ;
    buf_clk new_AGEMA_reg_buffer_3547 ( .C (clk), .D (new_AGEMA_signal_6977), .Q (new_AGEMA_signal_6978) ) ;
    buf_clk new_AGEMA_reg_buffer_3549 ( .C (clk), .D (new_AGEMA_signal_6979), .Q (new_AGEMA_signal_6980) ) ;
    buf_clk new_AGEMA_reg_buffer_3551 ( .C (clk), .D (new_AGEMA_signal_6981), .Q (new_AGEMA_signal_6982) ) ;
    buf_clk new_AGEMA_reg_buffer_3553 ( .C (clk), .D (new_AGEMA_signal_6983), .Q (new_AGEMA_signal_6984) ) ;
    buf_clk new_AGEMA_reg_buffer_3555 ( .C (clk), .D (new_AGEMA_signal_6985), .Q (new_AGEMA_signal_6986) ) ;
    buf_clk new_AGEMA_reg_buffer_3557 ( .C (clk), .D (new_AGEMA_signal_6987), .Q (new_AGEMA_signal_6988) ) ;
    buf_clk new_AGEMA_reg_buffer_3559 ( .C (clk), .D (new_AGEMA_signal_6989), .Q (new_AGEMA_signal_6990) ) ;
    buf_clk new_AGEMA_reg_buffer_3561 ( .C (clk), .D (new_AGEMA_signal_6991), .Q (new_AGEMA_signal_6992) ) ;
    buf_clk new_AGEMA_reg_buffer_3563 ( .C (clk), .D (new_AGEMA_signal_6993), .Q (new_AGEMA_signal_6994) ) ;
    buf_clk new_AGEMA_reg_buffer_3565 ( .C (clk), .D (new_AGEMA_signal_6995), .Q (new_AGEMA_signal_6996) ) ;
    buf_clk new_AGEMA_reg_buffer_3567 ( .C (clk), .D (new_AGEMA_signal_6997), .Q (new_AGEMA_signal_6998) ) ;
    buf_clk new_AGEMA_reg_buffer_3569 ( .C (clk), .D (new_AGEMA_signal_6999), .Q (new_AGEMA_signal_7000) ) ;
    buf_clk new_AGEMA_reg_buffer_3571 ( .C (clk), .D (new_AGEMA_signal_7001), .Q (new_AGEMA_signal_7002) ) ;
    buf_clk new_AGEMA_reg_buffer_3573 ( .C (clk), .D (new_AGEMA_signal_7003), .Q (new_AGEMA_signal_7004) ) ;
    buf_clk new_AGEMA_reg_buffer_3575 ( .C (clk), .D (new_AGEMA_signal_7005), .Q (new_AGEMA_signal_7006) ) ;
    buf_clk new_AGEMA_reg_buffer_3577 ( .C (clk), .D (new_AGEMA_signal_7007), .Q (new_AGEMA_signal_7008) ) ;
    buf_clk new_AGEMA_reg_buffer_3579 ( .C (clk), .D (new_AGEMA_signal_7009), .Q (new_AGEMA_signal_7010) ) ;
    buf_clk new_AGEMA_reg_buffer_3581 ( .C (clk), .D (new_AGEMA_signal_7011), .Q (new_AGEMA_signal_7012) ) ;
    buf_clk new_AGEMA_reg_buffer_3583 ( .C (clk), .D (new_AGEMA_signal_7013), .Q (new_AGEMA_signal_7014) ) ;
    buf_clk new_AGEMA_reg_buffer_3585 ( .C (clk), .D (new_AGEMA_signal_7015), .Q (new_AGEMA_signal_7016) ) ;
    buf_clk new_AGEMA_reg_buffer_3587 ( .C (clk), .D (new_AGEMA_signal_7017), .Q (new_AGEMA_signal_7018) ) ;
    buf_clk new_AGEMA_reg_buffer_3589 ( .C (clk), .D (new_AGEMA_signal_7019), .Q (new_AGEMA_signal_7020) ) ;
    buf_clk new_AGEMA_reg_buffer_3591 ( .C (clk), .D (new_AGEMA_signal_7021), .Q (new_AGEMA_signal_7022) ) ;
    buf_clk new_AGEMA_reg_buffer_3593 ( .C (clk), .D (new_AGEMA_signal_7023), .Q (new_AGEMA_signal_7024) ) ;
    buf_clk new_AGEMA_reg_buffer_3595 ( .C (clk), .D (new_AGEMA_signal_7025), .Q (new_AGEMA_signal_7026) ) ;
    buf_clk new_AGEMA_reg_buffer_3597 ( .C (clk), .D (new_AGEMA_signal_7027), .Q (new_AGEMA_signal_7028) ) ;
    buf_clk new_AGEMA_reg_buffer_3599 ( .C (clk), .D (new_AGEMA_signal_7029), .Q (new_AGEMA_signal_7030) ) ;
    buf_clk new_AGEMA_reg_buffer_3601 ( .C (clk), .D (new_AGEMA_signal_7031), .Q (new_AGEMA_signal_7032) ) ;
    buf_clk new_AGEMA_reg_buffer_3603 ( .C (clk), .D (new_AGEMA_signal_7033), .Q (new_AGEMA_signal_7034) ) ;
    buf_clk new_AGEMA_reg_buffer_3605 ( .C (clk), .D (new_AGEMA_signal_7035), .Q (new_AGEMA_signal_7036) ) ;
    buf_clk new_AGEMA_reg_buffer_3607 ( .C (clk), .D (new_AGEMA_signal_7037), .Q (new_AGEMA_signal_7038) ) ;
    buf_clk new_AGEMA_reg_buffer_3609 ( .C (clk), .D (new_AGEMA_signal_7039), .Q (new_AGEMA_signal_7040) ) ;
    buf_clk new_AGEMA_reg_buffer_3611 ( .C (clk), .D (new_AGEMA_signal_7041), .Q (new_AGEMA_signal_7042) ) ;
    buf_clk new_AGEMA_reg_buffer_3613 ( .C (clk), .D (new_AGEMA_signal_7043), .Q (new_AGEMA_signal_7044) ) ;
    buf_clk new_AGEMA_reg_buffer_3615 ( .C (clk), .D (new_AGEMA_signal_7045), .Q (new_AGEMA_signal_7046) ) ;
    buf_clk new_AGEMA_reg_buffer_3617 ( .C (clk), .D (new_AGEMA_signal_7047), .Q (new_AGEMA_signal_7048) ) ;
    buf_clk new_AGEMA_reg_buffer_3619 ( .C (clk), .D (new_AGEMA_signal_7049), .Q (new_AGEMA_signal_7050) ) ;
    buf_clk new_AGEMA_reg_buffer_3621 ( .C (clk), .D (new_AGEMA_signal_7051), .Q (new_AGEMA_signal_7052) ) ;
    buf_clk new_AGEMA_reg_buffer_3623 ( .C (clk), .D (new_AGEMA_signal_7053), .Q (new_AGEMA_signal_7054) ) ;
    buf_clk new_AGEMA_reg_buffer_3625 ( .C (clk), .D (new_AGEMA_signal_7055), .Q (new_AGEMA_signal_7056) ) ;
    buf_clk new_AGEMA_reg_buffer_3627 ( .C (clk), .D (new_AGEMA_signal_7057), .Q (new_AGEMA_signal_7058) ) ;
    buf_clk new_AGEMA_reg_buffer_3629 ( .C (clk), .D (new_AGEMA_signal_7059), .Q (new_AGEMA_signal_7060) ) ;
    buf_clk new_AGEMA_reg_buffer_3631 ( .C (clk), .D (new_AGEMA_signal_7061), .Q (new_AGEMA_signal_7062) ) ;
    buf_clk new_AGEMA_reg_buffer_3633 ( .C (clk), .D (new_AGEMA_signal_7063), .Q (new_AGEMA_signal_7064) ) ;
    buf_clk new_AGEMA_reg_buffer_3635 ( .C (clk), .D (new_AGEMA_signal_7065), .Q (new_AGEMA_signal_7066) ) ;
    buf_clk new_AGEMA_reg_buffer_3637 ( .C (clk), .D (new_AGEMA_signal_7067), .Q (new_AGEMA_signal_7068) ) ;
    buf_clk new_AGEMA_reg_buffer_3639 ( .C (clk), .D (new_AGEMA_signal_7069), .Q (new_AGEMA_signal_7070) ) ;
    buf_clk new_AGEMA_reg_buffer_3641 ( .C (clk), .D (new_AGEMA_signal_7071), .Q (new_AGEMA_signal_7072) ) ;
    buf_clk new_AGEMA_reg_buffer_3643 ( .C (clk), .D (new_AGEMA_signal_7073), .Q (new_AGEMA_signal_7074) ) ;
    buf_clk new_AGEMA_reg_buffer_3645 ( .C (clk), .D (new_AGEMA_signal_7075), .Q (new_AGEMA_signal_7076) ) ;
    buf_clk new_AGEMA_reg_buffer_3647 ( .C (clk), .D (new_AGEMA_signal_7077), .Q (new_AGEMA_signal_7078) ) ;
    buf_clk new_AGEMA_reg_buffer_3649 ( .C (clk), .D (new_AGEMA_signal_7079), .Q (new_AGEMA_signal_7080) ) ;
    buf_clk new_AGEMA_reg_buffer_3651 ( .C (clk), .D (new_AGEMA_signal_7081), .Q (new_AGEMA_signal_7082) ) ;
    buf_clk new_AGEMA_reg_buffer_3653 ( .C (clk), .D (new_AGEMA_signal_7083), .Q (new_AGEMA_signal_7084) ) ;
    buf_clk new_AGEMA_reg_buffer_3655 ( .C (clk), .D (new_AGEMA_signal_7085), .Q (new_AGEMA_signal_7086) ) ;
    buf_clk new_AGEMA_reg_buffer_3657 ( .C (clk), .D (new_AGEMA_signal_7087), .Q (new_AGEMA_signal_7088) ) ;
    buf_clk new_AGEMA_reg_buffer_3659 ( .C (clk), .D (new_AGEMA_signal_7089), .Q (new_AGEMA_signal_7090) ) ;
    buf_clk new_AGEMA_reg_buffer_3661 ( .C (clk), .D (new_AGEMA_signal_7091), .Q (new_AGEMA_signal_7092) ) ;
    buf_clk new_AGEMA_reg_buffer_3663 ( .C (clk), .D (new_AGEMA_signal_7093), .Q (new_AGEMA_signal_7094) ) ;
    buf_clk new_AGEMA_reg_buffer_3665 ( .C (clk), .D (new_AGEMA_signal_7095), .Q (new_AGEMA_signal_7096) ) ;
    buf_clk new_AGEMA_reg_buffer_3667 ( .C (clk), .D (new_AGEMA_signal_7097), .Q (new_AGEMA_signal_7098) ) ;
    buf_clk new_AGEMA_reg_buffer_3669 ( .C (clk), .D (new_AGEMA_signal_7099), .Q (new_AGEMA_signal_7100) ) ;
    buf_clk new_AGEMA_reg_buffer_3671 ( .C (clk), .D (new_AGEMA_signal_7101), .Q (new_AGEMA_signal_7102) ) ;
    buf_clk new_AGEMA_reg_buffer_3673 ( .C (clk), .D (new_AGEMA_signal_7103), .Q (new_AGEMA_signal_7104) ) ;
    buf_clk new_AGEMA_reg_buffer_3675 ( .C (clk), .D (new_AGEMA_signal_7105), .Q (new_AGEMA_signal_7106) ) ;
    buf_clk new_AGEMA_reg_buffer_3677 ( .C (clk), .D (new_AGEMA_signal_7107), .Q (new_AGEMA_signal_7108) ) ;
    buf_clk new_AGEMA_reg_buffer_3679 ( .C (clk), .D (new_AGEMA_signal_7109), .Q (new_AGEMA_signal_7110) ) ;
    buf_clk new_AGEMA_reg_buffer_3681 ( .C (clk), .D (new_AGEMA_signal_7111), .Q (new_AGEMA_signal_7112) ) ;
    buf_clk new_AGEMA_reg_buffer_3683 ( .C (clk), .D (new_AGEMA_signal_7113), .Q (new_AGEMA_signal_7114) ) ;
    buf_clk new_AGEMA_reg_buffer_3685 ( .C (clk), .D (new_AGEMA_signal_7115), .Q (new_AGEMA_signal_7116) ) ;
    buf_clk new_AGEMA_reg_buffer_3687 ( .C (clk), .D (new_AGEMA_signal_7117), .Q (new_AGEMA_signal_7118) ) ;
    buf_clk new_AGEMA_reg_buffer_3689 ( .C (clk), .D (new_AGEMA_signal_7119), .Q (new_AGEMA_signal_7120) ) ;
    buf_clk new_AGEMA_reg_buffer_3691 ( .C (clk), .D (new_AGEMA_signal_7121), .Q (new_AGEMA_signal_7122) ) ;
    buf_clk new_AGEMA_reg_buffer_3693 ( .C (clk), .D (new_AGEMA_signal_7123), .Q (new_AGEMA_signal_7124) ) ;
    buf_clk new_AGEMA_reg_buffer_3695 ( .C (clk), .D (new_AGEMA_signal_7125), .Q (new_AGEMA_signal_7126) ) ;
    buf_clk new_AGEMA_reg_buffer_3697 ( .C (clk), .D (new_AGEMA_signal_7127), .Q (new_AGEMA_signal_7128) ) ;
    buf_clk new_AGEMA_reg_buffer_3699 ( .C (clk), .D (new_AGEMA_signal_7129), .Q (new_AGEMA_signal_7130) ) ;
    buf_clk new_AGEMA_reg_buffer_3701 ( .C (clk), .D (new_AGEMA_signal_7131), .Q (new_AGEMA_signal_7132) ) ;
    buf_clk new_AGEMA_reg_buffer_3703 ( .C (clk), .D (new_AGEMA_signal_7133), .Q (new_AGEMA_signal_7134) ) ;
    buf_clk new_AGEMA_reg_buffer_3705 ( .C (clk), .D (new_AGEMA_signal_7135), .Q (new_AGEMA_signal_7136) ) ;
    buf_clk new_AGEMA_reg_buffer_3707 ( .C (clk), .D (new_AGEMA_signal_7137), .Q (new_AGEMA_signal_7138) ) ;
    buf_clk new_AGEMA_reg_buffer_3709 ( .C (clk), .D (new_AGEMA_signal_7139), .Q (new_AGEMA_signal_7140) ) ;
    buf_clk new_AGEMA_reg_buffer_3711 ( .C (clk), .D (new_AGEMA_signal_7141), .Q (new_AGEMA_signal_7142) ) ;
    buf_clk new_AGEMA_reg_buffer_3715 ( .C (clk), .D (new_AGEMA_signal_7145), .Q (new_AGEMA_signal_7146) ) ;
    buf_clk new_AGEMA_reg_buffer_3719 ( .C (clk), .D (new_AGEMA_signal_7149), .Q (new_AGEMA_signal_7150) ) ;
    buf_clk new_AGEMA_reg_buffer_3723 ( .C (clk), .D (new_AGEMA_signal_7153), .Q (new_AGEMA_signal_7154) ) ;
    buf_clk new_AGEMA_reg_buffer_3727 ( .C (clk), .D (new_AGEMA_signal_7157), .Q (new_AGEMA_signal_7158) ) ;
    buf_clk new_AGEMA_reg_buffer_3731 ( .C (clk), .D (new_AGEMA_signal_7161), .Q (new_AGEMA_signal_7162) ) ;
    buf_clk new_AGEMA_reg_buffer_3735 ( .C (clk), .D (new_AGEMA_signal_7165), .Q (new_AGEMA_signal_7166) ) ;
    buf_clk new_AGEMA_reg_buffer_3739 ( .C (clk), .D (new_AGEMA_signal_7169), .Q (new_AGEMA_signal_7170) ) ;
    buf_clk new_AGEMA_reg_buffer_3743 ( .C (clk), .D (new_AGEMA_signal_7173), .Q (new_AGEMA_signal_7174) ) ;
    buf_clk new_AGEMA_reg_buffer_3747 ( .C (clk), .D (new_AGEMA_signal_7177), .Q (new_AGEMA_signal_7178) ) ;
    buf_clk new_AGEMA_reg_buffer_3751 ( .C (clk), .D (new_AGEMA_signal_7181), .Q (new_AGEMA_signal_7182) ) ;
    buf_clk new_AGEMA_reg_buffer_3755 ( .C (clk), .D (new_AGEMA_signal_7185), .Q (new_AGEMA_signal_7186) ) ;
    buf_clk new_AGEMA_reg_buffer_3759 ( .C (clk), .D (new_AGEMA_signal_7189), .Q (new_AGEMA_signal_7190) ) ;
    buf_clk new_AGEMA_reg_buffer_3763 ( .C (clk), .D (new_AGEMA_signal_7193), .Q (new_AGEMA_signal_7194) ) ;
    buf_clk new_AGEMA_reg_buffer_3767 ( .C (clk), .D (new_AGEMA_signal_7197), .Q (new_AGEMA_signal_7198) ) ;
    buf_clk new_AGEMA_reg_buffer_3771 ( .C (clk), .D (new_AGEMA_signal_7201), .Q (new_AGEMA_signal_7202) ) ;
    buf_clk new_AGEMA_reg_buffer_3775 ( .C (clk), .D (new_AGEMA_signal_7205), .Q (new_AGEMA_signal_7206) ) ;
    buf_clk new_AGEMA_reg_buffer_3779 ( .C (clk), .D (new_AGEMA_signal_7209), .Q (new_AGEMA_signal_7210) ) ;
    buf_clk new_AGEMA_reg_buffer_3783 ( .C (clk), .D (new_AGEMA_signal_7213), .Q (new_AGEMA_signal_7214) ) ;
    buf_clk new_AGEMA_reg_buffer_3787 ( .C (clk), .D (new_AGEMA_signal_7217), .Q (new_AGEMA_signal_7218) ) ;
    buf_clk new_AGEMA_reg_buffer_3791 ( .C (clk), .D (new_AGEMA_signal_7221), .Q (new_AGEMA_signal_7222) ) ;
    buf_clk new_AGEMA_reg_buffer_3795 ( .C (clk), .D (new_AGEMA_signal_7225), .Q (new_AGEMA_signal_7226) ) ;
    buf_clk new_AGEMA_reg_buffer_3799 ( .C (clk), .D (new_AGEMA_signal_7229), .Q (new_AGEMA_signal_7230) ) ;
    buf_clk new_AGEMA_reg_buffer_3803 ( .C (clk), .D (new_AGEMA_signal_7233), .Q (new_AGEMA_signal_7234) ) ;
    buf_clk new_AGEMA_reg_buffer_3807 ( .C (clk), .D (new_AGEMA_signal_7237), .Q (new_AGEMA_signal_7238) ) ;
    buf_clk new_AGEMA_reg_buffer_3811 ( .C (clk), .D (new_AGEMA_signal_7241), .Q (new_AGEMA_signal_7242) ) ;
    buf_clk new_AGEMA_reg_buffer_3815 ( .C (clk), .D (new_AGEMA_signal_7245), .Q (new_AGEMA_signal_7246) ) ;
    buf_clk new_AGEMA_reg_buffer_3819 ( .C (clk), .D (new_AGEMA_signal_7249), .Q (new_AGEMA_signal_7250) ) ;
    buf_clk new_AGEMA_reg_buffer_3823 ( .C (clk), .D (new_AGEMA_signal_7253), .Q (new_AGEMA_signal_7254) ) ;
    buf_clk new_AGEMA_reg_buffer_3827 ( .C (clk), .D (new_AGEMA_signal_7257), .Q (new_AGEMA_signal_7258) ) ;
    buf_clk new_AGEMA_reg_buffer_3831 ( .C (clk), .D (new_AGEMA_signal_7261), .Q (new_AGEMA_signal_7262) ) ;
    buf_clk new_AGEMA_reg_buffer_3835 ( .C (clk), .D (new_AGEMA_signal_7265), .Q (new_AGEMA_signal_7266) ) ;
    buf_clk new_AGEMA_reg_buffer_3839 ( .C (clk), .D (new_AGEMA_signal_7269), .Q (new_AGEMA_signal_7270) ) ;
    buf_clk new_AGEMA_reg_buffer_3843 ( .C (clk), .D (new_AGEMA_signal_7273), .Q (new_AGEMA_signal_7274) ) ;
    buf_clk new_AGEMA_reg_buffer_3847 ( .C (clk), .D (new_AGEMA_signal_7277), .Q (new_AGEMA_signal_7278) ) ;
    buf_clk new_AGEMA_reg_buffer_3851 ( .C (clk), .D (new_AGEMA_signal_7281), .Q (new_AGEMA_signal_7282) ) ;
    buf_clk new_AGEMA_reg_buffer_3855 ( .C (clk), .D (new_AGEMA_signal_7285), .Q (new_AGEMA_signal_7286) ) ;
    buf_clk new_AGEMA_reg_buffer_3859 ( .C (clk), .D (new_AGEMA_signal_7289), .Q (new_AGEMA_signal_7290) ) ;
    buf_clk new_AGEMA_reg_buffer_3863 ( .C (clk), .D (new_AGEMA_signal_7293), .Q (new_AGEMA_signal_7294) ) ;
    buf_clk new_AGEMA_reg_buffer_3867 ( .C (clk), .D (new_AGEMA_signal_7297), .Q (new_AGEMA_signal_7298) ) ;
    buf_clk new_AGEMA_reg_buffer_3871 ( .C (clk), .D (new_AGEMA_signal_7301), .Q (new_AGEMA_signal_7302) ) ;
    buf_clk new_AGEMA_reg_buffer_3875 ( .C (clk), .D (new_AGEMA_signal_7305), .Q (new_AGEMA_signal_7306) ) ;
    buf_clk new_AGEMA_reg_buffer_3879 ( .C (clk), .D (new_AGEMA_signal_7309), .Q (new_AGEMA_signal_7310) ) ;
    buf_clk new_AGEMA_reg_buffer_3883 ( .C (clk), .D (new_AGEMA_signal_7313), .Q (new_AGEMA_signal_7314) ) ;
    buf_clk new_AGEMA_reg_buffer_3887 ( .C (clk), .D (new_AGEMA_signal_7317), .Q (new_AGEMA_signal_7318) ) ;
    buf_clk new_AGEMA_reg_buffer_3891 ( .C (clk), .D (new_AGEMA_signal_7321), .Q (new_AGEMA_signal_7322) ) ;
    buf_clk new_AGEMA_reg_buffer_3895 ( .C (clk), .D (new_AGEMA_signal_7325), .Q (new_AGEMA_signal_7326) ) ;
    buf_clk new_AGEMA_reg_buffer_3899 ( .C (clk), .D (new_AGEMA_signal_7329), .Q (new_AGEMA_signal_7330) ) ;
    buf_clk new_AGEMA_reg_buffer_3903 ( .C (clk), .D (new_AGEMA_signal_7333), .Q (new_AGEMA_signal_7334) ) ;
    buf_clk new_AGEMA_reg_buffer_3907 ( .C (clk), .D (new_AGEMA_signal_7337), .Q (new_AGEMA_signal_7338) ) ;
    buf_clk new_AGEMA_reg_buffer_3911 ( .C (clk), .D (new_AGEMA_signal_7341), .Q (new_AGEMA_signal_7342) ) ;
    buf_clk new_AGEMA_reg_buffer_3915 ( .C (clk), .D (new_AGEMA_signal_7345), .Q (new_AGEMA_signal_7346) ) ;
    buf_clk new_AGEMA_reg_buffer_3919 ( .C (clk), .D (new_AGEMA_signal_7349), .Q (new_AGEMA_signal_7350) ) ;
    buf_clk new_AGEMA_reg_buffer_3923 ( .C (clk), .D (new_AGEMA_signal_7353), .Q (new_AGEMA_signal_7354) ) ;
    buf_clk new_AGEMA_reg_buffer_3927 ( .C (clk), .D (new_AGEMA_signal_7357), .Q (new_AGEMA_signal_7358) ) ;
    buf_clk new_AGEMA_reg_buffer_3931 ( .C (clk), .D (new_AGEMA_signal_7361), .Q (new_AGEMA_signal_7362) ) ;
    buf_clk new_AGEMA_reg_buffer_3935 ( .C (clk), .D (new_AGEMA_signal_7365), .Q (new_AGEMA_signal_7366) ) ;
    buf_clk new_AGEMA_reg_buffer_3939 ( .C (clk), .D (new_AGEMA_signal_7369), .Q (new_AGEMA_signal_7370) ) ;
    buf_clk new_AGEMA_reg_buffer_3943 ( .C (clk), .D (new_AGEMA_signal_7373), .Q (new_AGEMA_signal_7374) ) ;
    buf_clk new_AGEMA_reg_buffer_3947 ( .C (clk), .D (new_AGEMA_signal_7377), .Q (new_AGEMA_signal_7378) ) ;
    buf_clk new_AGEMA_reg_buffer_3951 ( .C (clk), .D (new_AGEMA_signal_7381), .Q (new_AGEMA_signal_7382) ) ;
    buf_clk new_AGEMA_reg_buffer_3955 ( .C (clk), .D (new_AGEMA_signal_7385), .Q (new_AGEMA_signal_7386) ) ;
    buf_clk new_AGEMA_reg_buffer_3959 ( .C (clk), .D (new_AGEMA_signal_7389), .Q (new_AGEMA_signal_7390) ) ;
    buf_clk new_AGEMA_reg_buffer_3963 ( .C (clk), .D (new_AGEMA_signal_7393), .Q (new_AGEMA_signal_7394) ) ;
    buf_clk new_AGEMA_reg_buffer_3967 ( .C (clk), .D (new_AGEMA_signal_7397), .Q (new_AGEMA_signal_7398) ) ;
    buf_clk new_AGEMA_reg_buffer_3971 ( .C (clk), .D (new_AGEMA_signal_7401), .Q (new_AGEMA_signal_7402) ) ;
    buf_clk new_AGEMA_reg_buffer_3975 ( .C (clk), .D (new_AGEMA_signal_7405), .Q (new_AGEMA_signal_7406) ) ;
    buf_clk new_AGEMA_reg_buffer_3979 ( .C (clk), .D (new_AGEMA_signal_7409), .Q (new_AGEMA_signal_7410) ) ;
    buf_clk new_AGEMA_reg_buffer_3983 ( .C (clk), .D (new_AGEMA_signal_7413), .Q (new_AGEMA_signal_7414) ) ;
    buf_clk new_AGEMA_reg_buffer_3987 ( .C (clk), .D (new_AGEMA_signal_7417), .Q (new_AGEMA_signal_7418) ) ;
    buf_clk new_AGEMA_reg_buffer_3991 ( .C (clk), .D (new_AGEMA_signal_7421), .Q (new_AGEMA_signal_7422) ) ;
    buf_clk new_AGEMA_reg_buffer_3995 ( .C (clk), .D (new_AGEMA_signal_7425), .Q (new_AGEMA_signal_7426) ) ;
    buf_clk new_AGEMA_reg_buffer_3999 ( .C (clk), .D (new_AGEMA_signal_7429), .Q (new_AGEMA_signal_7430) ) ;
    buf_clk new_AGEMA_reg_buffer_4003 ( .C (clk), .D (new_AGEMA_signal_7433), .Q (new_AGEMA_signal_7434) ) ;
    buf_clk new_AGEMA_reg_buffer_4007 ( .C (clk), .D (new_AGEMA_signal_7437), .Q (new_AGEMA_signal_7438) ) ;
    buf_clk new_AGEMA_reg_buffer_4011 ( .C (clk), .D (new_AGEMA_signal_7441), .Q (new_AGEMA_signal_7442) ) ;
    buf_clk new_AGEMA_reg_buffer_4015 ( .C (clk), .D (new_AGEMA_signal_7445), .Q (new_AGEMA_signal_7446) ) ;
    buf_clk new_AGEMA_reg_buffer_4019 ( .C (clk), .D (new_AGEMA_signal_7449), .Q (new_AGEMA_signal_7450) ) ;
    buf_clk new_AGEMA_reg_buffer_4023 ( .C (clk), .D (new_AGEMA_signal_7453), .Q (new_AGEMA_signal_7454) ) ;
    buf_clk new_AGEMA_reg_buffer_4027 ( .C (clk), .D (new_AGEMA_signal_7457), .Q (new_AGEMA_signal_7458) ) ;
    buf_clk new_AGEMA_reg_buffer_4031 ( .C (clk), .D (new_AGEMA_signal_7461), .Q (new_AGEMA_signal_7462) ) ;
    buf_clk new_AGEMA_reg_buffer_4035 ( .C (clk), .D (new_AGEMA_signal_7465), .Q (new_AGEMA_signal_7466) ) ;
    buf_clk new_AGEMA_reg_buffer_4039 ( .C (clk), .D (new_AGEMA_signal_7469), .Q (new_AGEMA_signal_7470) ) ;
    buf_clk new_AGEMA_reg_buffer_4043 ( .C (clk), .D (new_AGEMA_signal_7473), .Q (new_AGEMA_signal_7474) ) ;
    buf_clk new_AGEMA_reg_buffer_4047 ( .C (clk), .D (new_AGEMA_signal_7477), .Q (new_AGEMA_signal_7478) ) ;
    buf_clk new_AGEMA_reg_buffer_4051 ( .C (clk), .D (new_AGEMA_signal_7481), .Q (new_AGEMA_signal_7482) ) ;
    buf_clk new_AGEMA_reg_buffer_4055 ( .C (clk), .D (new_AGEMA_signal_7485), .Q (new_AGEMA_signal_7486) ) ;
    buf_clk new_AGEMA_reg_buffer_4059 ( .C (clk), .D (new_AGEMA_signal_7489), .Q (new_AGEMA_signal_7490) ) ;
    buf_clk new_AGEMA_reg_buffer_4063 ( .C (clk), .D (new_AGEMA_signal_7493), .Q (new_AGEMA_signal_7494) ) ;
    buf_clk new_AGEMA_reg_buffer_4067 ( .C (clk), .D (new_AGEMA_signal_7497), .Q (new_AGEMA_signal_7498) ) ;
    buf_clk new_AGEMA_reg_buffer_4071 ( .C (clk), .D (new_AGEMA_signal_7501), .Q (new_AGEMA_signal_7502) ) ;
    buf_clk new_AGEMA_reg_buffer_4075 ( .C (clk), .D (new_AGEMA_signal_7505), .Q (new_AGEMA_signal_7506) ) ;
    buf_clk new_AGEMA_reg_buffer_4079 ( .C (clk), .D (new_AGEMA_signal_7509), .Q (new_AGEMA_signal_7510) ) ;
    buf_clk new_AGEMA_reg_buffer_4083 ( .C (clk), .D (new_AGEMA_signal_7513), .Q (new_AGEMA_signal_7514) ) ;
    buf_clk new_AGEMA_reg_buffer_4087 ( .C (clk), .D (new_AGEMA_signal_7517), .Q (new_AGEMA_signal_7518) ) ;
    buf_clk new_AGEMA_reg_buffer_4091 ( .C (clk), .D (new_AGEMA_signal_7521), .Q (new_AGEMA_signal_7522) ) ;
    buf_clk new_AGEMA_reg_buffer_4095 ( .C (clk), .D (new_AGEMA_signal_7525), .Q (new_AGEMA_signal_7526) ) ;
    buf_clk new_AGEMA_reg_buffer_4099 ( .C (clk), .D (new_AGEMA_signal_7529), .Q (new_AGEMA_signal_7530) ) ;
    buf_clk new_AGEMA_reg_buffer_4103 ( .C (clk), .D (new_AGEMA_signal_7533), .Q (new_AGEMA_signal_7534) ) ;
    buf_clk new_AGEMA_reg_buffer_4107 ( .C (clk), .D (new_AGEMA_signal_7537), .Q (new_AGEMA_signal_7538) ) ;
    buf_clk new_AGEMA_reg_buffer_4111 ( .C (clk), .D (new_AGEMA_signal_7541), .Q (new_AGEMA_signal_7542) ) ;
    buf_clk new_AGEMA_reg_buffer_4115 ( .C (clk), .D (new_AGEMA_signal_7545), .Q (new_AGEMA_signal_7546) ) ;
    buf_clk new_AGEMA_reg_buffer_4119 ( .C (clk), .D (new_AGEMA_signal_7549), .Q (new_AGEMA_signal_7550) ) ;
    buf_clk new_AGEMA_reg_buffer_4123 ( .C (clk), .D (new_AGEMA_signal_7553), .Q (new_AGEMA_signal_7554) ) ;
    buf_clk new_AGEMA_reg_buffer_4127 ( .C (clk), .D (new_AGEMA_signal_7557), .Q (new_AGEMA_signal_7558) ) ;
    buf_clk new_AGEMA_reg_buffer_4131 ( .C (clk), .D (new_AGEMA_signal_7561), .Q (new_AGEMA_signal_7562) ) ;
    buf_clk new_AGEMA_reg_buffer_4135 ( .C (clk), .D (new_AGEMA_signal_7565), .Q (new_AGEMA_signal_7566) ) ;
    buf_clk new_AGEMA_reg_buffer_4139 ( .C (clk), .D (new_AGEMA_signal_7569), .Q (new_AGEMA_signal_7570) ) ;
    buf_clk new_AGEMA_reg_buffer_4143 ( .C (clk), .D (new_AGEMA_signal_7573), .Q (new_AGEMA_signal_7574) ) ;
    buf_clk new_AGEMA_reg_buffer_4147 ( .C (clk), .D (new_AGEMA_signal_7577), .Q (new_AGEMA_signal_7578) ) ;
    buf_clk new_AGEMA_reg_buffer_4151 ( .C (clk), .D (new_AGEMA_signal_7581), .Q (new_AGEMA_signal_7582) ) ;
    buf_clk new_AGEMA_reg_buffer_4155 ( .C (clk), .D (new_AGEMA_signal_7585), .Q (new_AGEMA_signal_7586) ) ;
    buf_clk new_AGEMA_reg_buffer_4159 ( .C (clk), .D (new_AGEMA_signal_7589), .Q (new_AGEMA_signal_7590) ) ;
    buf_clk new_AGEMA_reg_buffer_4163 ( .C (clk), .D (new_AGEMA_signal_7593), .Q (new_AGEMA_signal_7594) ) ;
    buf_clk new_AGEMA_reg_buffer_4167 ( .C (clk), .D (new_AGEMA_signal_7597), .Q (new_AGEMA_signal_7598) ) ;
    buf_clk new_AGEMA_reg_buffer_4171 ( .C (clk), .D (new_AGEMA_signal_7601), .Q (new_AGEMA_signal_7602) ) ;
    buf_clk new_AGEMA_reg_buffer_4175 ( .C (clk), .D (new_AGEMA_signal_7605), .Q (new_AGEMA_signal_7606) ) ;
    buf_clk new_AGEMA_reg_buffer_4179 ( .C (clk), .D (new_AGEMA_signal_7609), .Q (new_AGEMA_signal_7610) ) ;
    buf_clk new_AGEMA_reg_buffer_4183 ( .C (clk), .D (new_AGEMA_signal_7613), .Q (new_AGEMA_signal_7614) ) ;
    buf_clk new_AGEMA_reg_buffer_4187 ( .C (clk), .D (new_AGEMA_signal_7617), .Q (new_AGEMA_signal_7618) ) ;
    buf_clk new_AGEMA_reg_buffer_4191 ( .C (clk), .D (new_AGEMA_signal_7621), .Q (new_AGEMA_signal_7622) ) ;
    buf_clk new_AGEMA_reg_buffer_4195 ( .C (clk), .D (new_AGEMA_signal_7625), .Q (new_AGEMA_signal_7626) ) ;
    buf_clk new_AGEMA_reg_buffer_4199 ( .C (clk), .D (new_AGEMA_signal_7629), .Q (new_AGEMA_signal_7630) ) ;
    buf_clk new_AGEMA_reg_buffer_4203 ( .C (clk), .D (new_AGEMA_signal_7633), .Q (new_AGEMA_signal_7634) ) ;
    buf_clk new_AGEMA_reg_buffer_4207 ( .C (clk), .D (new_AGEMA_signal_7637), .Q (new_AGEMA_signal_7638) ) ;
    buf_clk new_AGEMA_reg_buffer_4211 ( .C (clk), .D (new_AGEMA_signal_7641), .Q (new_AGEMA_signal_7642) ) ;
    buf_clk new_AGEMA_reg_buffer_4215 ( .C (clk), .D (new_AGEMA_signal_7645), .Q (new_AGEMA_signal_7646) ) ;
    buf_clk new_AGEMA_reg_buffer_4219 ( .C (clk), .D (new_AGEMA_signal_7649), .Q (new_AGEMA_signal_7650) ) ;
    buf_clk new_AGEMA_reg_buffer_4223 ( .C (clk), .D (new_AGEMA_signal_7653), .Q (new_AGEMA_signal_7654) ) ;
    buf_clk new_AGEMA_reg_buffer_4227 ( .C (clk), .D (new_AGEMA_signal_7657), .Q (new_AGEMA_signal_7658) ) ;
    buf_clk new_AGEMA_reg_buffer_4231 ( .C (clk), .D (new_AGEMA_signal_7661), .Q (new_AGEMA_signal_7662) ) ;
    buf_clk new_AGEMA_reg_buffer_4235 ( .C (clk), .D (new_AGEMA_signal_7665), .Q (new_AGEMA_signal_7666) ) ;
    buf_clk new_AGEMA_reg_buffer_4239 ( .C (clk), .D (new_AGEMA_signal_7669), .Q (new_AGEMA_signal_7670) ) ;
    buf_clk new_AGEMA_reg_buffer_4243 ( .C (clk), .D (new_AGEMA_signal_7673), .Q (new_AGEMA_signal_7674) ) ;
    buf_clk new_AGEMA_reg_buffer_4247 ( .C (clk), .D (new_AGEMA_signal_7677), .Q (new_AGEMA_signal_7678) ) ;
    buf_clk new_AGEMA_reg_buffer_4251 ( .C (clk), .D (new_AGEMA_signal_7681), .Q (new_AGEMA_signal_7682) ) ;
    buf_clk new_AGEMA_reg_buffer_4255 ( .C (clk), .D (new_AGEMA_signal_7685), .Q (new_AGEMA_signal_7686) ) ;
    buf_clk new_AGEMA_reg_buffer_4259 ( .C (clk), .D (new_AGEMA_signal_7689), .Q (new_AGEMA_signal_7690) ) ;
    buf_clk new_AGEMA_reg_buffer_4263 ( .C (clk), .D (new_AGEMA_signal_7693), .Q (new_AGEMA_signal_7694) ) ;
    buf_clk new_AGEMA_reg_buffer_4267 ( .C (clk), .D (new_AGEMA_signal_7697), .Q (new_AGEMA_signal_7698) ) ;
    buf_clk new_AGEMA_reg_buffer_4271 ( .C (clk), .D (new_AGEMA_signal_7701), .Q (new_AGEMA_signal_7702) ) ;
    buf_clk new_AGEMA_reg_buffer_4275 ( .C (clk), .D (new_AGEMA_signal_7705), .Q (new_AGEMA_signal_7706) ) ;
    buf_clk new_AGEMA_reg_buffer_4279 ( .C (clk), .D (new_AGEMA_signal_7709), .Q (new_AGEMA_signal_7710) ) ;
    buf_clk new_AGEMA_reg_buffer_4283 ( .C (clk), .D (new_AGEMA_signal_7713), .Q (new_AGEMA_signal_7714) ) ;
    buf_clk new_AGEMA_reg_buffer_4287 ( .C (clk), .D (new_AGEMA_signal_7717), .Q (new_AGEMA_signal_7718) ) ;
    buf_clk new_AGEMA_reg_buffer_4291 ( .C (clk), .D (new_AGEMA_signal_7721), .Q (new_AGEMA_signal_7722) ) ;
    buf_clk new_AGEMA_reg_buffer_4295 ( .C (clk), .D (new_AGEMA_signal_7725), .Q (new_AGEMA_signal_7726) ) ;
    buf_clk new_AGEMA_reg_buffer_4299 ( .C (clk), .D (new_AGEMA_signal_7729), .Q (new_AGEMA_signal_7730) ) ;
    buf_clk new_AGEMA_reg_buffer_4303 ( .C (clk), .D (new_AGEMA_signal_7733), .Q (new_AGEMA_signal_7734) ) ;
    buf_clk new_AGEMA_reg_buffer_4307 ( .C (clk), .D (new_AGEMA_signal_7737), .Q (new_AGEMA_signal_7738) ) ;
    buf_clk new_AGEMA_reg_buffer_4311 ( .C (clk), .D (new_AGEMA_signal_7741), .Q (new_AGEMA_signal_7742) ) ;
    buf_clk new_AGEMA_reg_buffer_4315 ( .C (clk), .D (new_AGEMA_signal_7745), .Q (new_AGEMA_signal_7746) ) ;
    buf_clk new_AGEMA_reg_buffer_4319 ( .C (clk), .D (new_AGEMA_signal_7749), .Q (new_AGEMA_signal_7750) ) ;
    buf_clk new_AGEMA_reg_buffer_4323 ( .C (clk), .D (new_AGEMA_signal_7753), .Q (new_AGEMA_signal_7754) ) ;
    buf_clk new_AGEMA_reg_buffer_4327 ( .C (clk), .D (new_AGEMA_signal_7757), .Q (new_AGEMA_signal_7758) ) ;
    buf_clk new_AGEMA_reg_buffer_4331 ( .C (clk), .D (new_AGEMA_signal_7761), .Q (new_AGEMA_signal_7762) ) ;
    buf_clk new_AGEMA_reg_buffer_4335 ( .C (clk), .D (new_AGEMA_signal_7765), .Q (new_AGEMA_signal_7766) ) ;
    buf_clk new_AGEMA_reg_buffer_4339 ( .C (clk), .D (new_AGEMA_signal_7769), .Q (new_AGEMA_signal_7770) ) ;
    buf_clk new_AGEMA_reg_buffer_4343 ( .C (clk), .D (new_AGEMA_signal_7773), .Q (new_AGEMA_signal_7774) ) ;
    buf_clk new_AGEMA_reg_buffer_4347 ( .C (clk), .D (new_AGEMA_signal_7777), .Q (new_AGEMA_signal_7778) ) ;
    buf_clk new_AGEMA_reg_buffer_4351 ( .C (clk), .D (new_AGEMA_signal_7781), .Q (new_AGEMA_signal_7782) ) ;
    buf_clk new_AGEMA_reg_buffer_4355 ( .C (clk), .D (new_AGEMA_signal_7785), .Q (new_AGEMA_signal_7786) ) ;
    buf_clk new_AGEMA_reg_buffer_4359 ( .C (clk), .D (new_AGEMA_signal_7789), .Q (new_AGEMA_signal_7790) ) ;
    buf_clk new_AGEMA_reg_buffer_4363 ( .C (clk), .D (new_AGEMA_signal_7793), .Q (new_AGEMA_signal_7794) ) ;
    buf_clk new_AGEMA_reg_buffer_4367 ( .C (clk), .D (new_AGEMA_signal_7797), .Q (new_AGEMA_signal_7798) ) ;
    buf_clk new_AGEMA_reg_buffer_4371 ( .C (clk), .D (new_AGEMA_signal_7801), .Q (new_AGEMA_signal_7802) ) ;
    buf_clk new_AGEMA_reg_buffer_4375 ( .C (clk), .D (new_AGEMA_signal_7805), .Q (new_AGEMA_signal_7806) ) ;
    buf_clk new_AGEMA_reg_buffer_4379 ( .C (clk), .D (new_AGEMA_signal_7809), .Q (new_AGEMA_signal_7810) ) ;
    buf_clk new_AGEMA_reg_buffer_4383 ( .C (clk), .D (new_AGEMA_signal_7813), .Q (new_AGEMA_signal_7814) ) ;
    buf_clk new_AGEMA_reg_buffer_4387 ( .C (clk), .D (new_AGEMA_signal_7817), .Q (new_AGEMA_signal_7818) ) ;
    buf_clk new_AGEMA_reg_buffer_4391 ( .C (clk), .D (new_AGEMA_signal_7821), .Q (new_AGEMA_signal_7822) ) ;
    buf_clk new_AGEMA_reg_buffer_4395 ( .C (clk), .D (new_AGEMA_signal_7825), .Q (new_AGEMA_signal_7826) ) ;
    buf_clk new_AGEMA_reg_buffer_4399 ( .C (clk), .D (new_AGEMA_signal_7829), .Q (new_AGEMA_signal_7830) ) ;
    buf_clk new_AGEMA_reg_buffer_4403 ( .C (clk), .D (new_AGEMA_signal_7833), .Q (new_AGEMA_signal_7834) ) ;
    buf_clk new_AGEMA_reg_buffer_4407 ( .C (clk), .D (new_AGEMA_signal_7837), .Q (new_AGEMA_signal_7838) ) ;
    buf_clk new_AGEMA_reg_buffer_4411 ( .C (clk), .D (new_AGEMA_signal_7841), .Q (new_AGEMA_signal_7842) ) ;
    buf_clk new_AGEMA_reg_buffer_4415 ( .C (clk), .D (new_AGEMA_signal_7845), .Q (new_AGEMA_signal_7846) ) ;
    buf_clk new_AGEMA_reg_buffer_4419 ( .C (clk), .D (new_AGEMA_signal_7849), .Q (new_AGEMA_signal_7850) ) ;
    buf_clk new_AGEMA_reg_buffer_4423 ( .C (clk), .D (new_AGEMA_signal_7853), .Q (new_AGEMA_signal_7854) ) ;
    buf_clk new_AGEMA_reg_buffer_4427 ( .C (clk), .D (new_AGEMA_signal_7857), .Q (new_AGEMA_signal_7858) ) ;
    buf_clk new_AGEMA_reg_buffer_4431 ( .C (clk), .D (new_AGEMA_signal_7861), .Q (new_AGEMA_signal_7862) ) ;
    buf_clk new_AGEMA_reg_buffer_4435 ( .C (clk), .D (new_AGEMA_signal_7865), .Q (new_AGEMA_signal_7866) ) ;
    buf_clk new_AGEMA_reg_buffer_4439 ( .C (clk), .D (new_AGEMA_signal_7869), .Q (new_AGEMA_signal_7870) ) ;
    buf_clk new_AGEMA_reg_buffer_4443 ( .C (clk), .D (new_AGEMA_signal_7873), .Q (new_AGEMA_signal_7874) ) ;
    buf_clk new_AGEMA_reg_buffer_4447 ( .C (clk), .D (new_AGEMA_signal_7877), .Q (new_AGEMA_signal_7878) ) ;
    buf_clk new_AGEMA_reg_buffer_4451 ( .C (clk), .D (new_AGEMA_signal_7881), .Q (new_AGEMA_signal_7882) ) ;
    buf_clk new_AGEMA_reg_buffer_4455 ( .C (clk), .D (new_AGEMA_signal_7885), .Q (new_AGEMA_signal_7886) ) ;
    buf_clk new_AGEMA_reg_buffer_4459 ( .C (clk), .D (new_AGEMA_signal_7889), .Q (new_AGEMA_signal_7890) ) ;
    buf_clk new_AGEMA_reg_buffer_4463 ( .C (clk), .D (new_AGEMA_signal_7893), .Q (new_AGEMA_signal_7894) ) ;
    buf_clk new_AGEMA_reg_buffer_4467 ( .C (clk), .D (new_AGEMA_signal_7897), .Q (new_AGEMA_signal_7898) ) ;
    buf_clk new_AGEMA_reg_buffer_4471 ( .C (clk), .D (new_AGEMA_signal_7901), .Q (new_AGEMA_signal_7902) ) ;
    buf_clk new_AGEMA_reg_buffer_4475 ( .C (clk), .D (new_AGEMA_signal_7905), .Q (new_AGEMA_signal_7906) ) ;
    buf_clk new_AGEMA_reg_buffer_4479 ( .C (clk), .D (new_AGEMA_signal_7909), .Q (new_AGEMA_signal_7910) ) ;
    buf_clk new_AGEMA_reg_buffer_4483 ( .C (clk), .D (new_AGEMA_signal_7913), .Q (new_AGEMA_signal_7914) ) ;
    buf_clk new_AGEMA_reg_buffer_4487 ( .C (clk), .D (new_AGEMA_signal_7917), .Q (new_AGEMA_signal_7918) ) ;
    buf_clk new_AGEMA_reg_buffer_4491 ( .C (clk), .D (new_AGEMA_signal_7921), .Q (new_AGEMA_signal_7922) ) ;
    buf_clk new_AGEMA_reg_buffer_4495 ( .C (clk), .D (new_AGEMA_signal_7925), .Q (new_AGEMA_signal_7926) ) ;
    buf_clk new_AGEMA_reg_buffer_4499 ( .C (clk), .D (new_AGEMA_signal_7929), .Q (new_AGEMA_signal_7930) ) ;
    buf_clk new_AGEMA_reg_buffer_4503 ( .C (clk), .D (new_AGEMA_signal_7933), .Q (new_AGEMA_signal_7934) ) ;
    buf_clk new_AGEMA_reg_buffer_4507 ( .C (clk), .D (new_AGEMA_signal_7937), .Q (new_AGEMA_signal_7938) ) ;
    buf_clk new_AGEMA_reg_buffer_4511 ( .C (clk), .D (new_AGEMA_signal_7941), .Q (new_AGEMA_signal_7942) ) ;
    buf_clk new_AGEMA_reg_buffer_4515 ( .C (clk), .D (new_AGEMA_signal_7945), .Q (new_AGEMA_signal_7946) ) ;
    buf_clk new_AGEMA_reg_buffer_4519 ( .C (clk), .D (new_AGEMA_signal_7949), .Q (new_AGEMA_signal_7950) ) ;
    buf_clk new_AGEMA_reg_buffer_4523 ( .C (clk), .D (new_AGEMA_signal_7953), .Q (new_AGEMA_signal_7954) ) ;
    buf_clk new_AGEMA_reg_buffer_4527 ( .C (clk), .D (new_AGEMA_signal_7957), .Q (new_AGEMA_signal_7958) ) ;
    buf_clk new_AGEMA_reg_buffer_4531 ( .C (clk), .D (new_AGEMA_signal_7961), .Q (new_AGEMA_signal_7962) ) ;
    buf_clk new_AGEMA_reg_buffer_4535 ( .C (clk), .D (new_AGEMA_signal_7965), .Q (new_AGEMA_signal_7966) ) ;
    buf_clk new_AGEMA_reg_buffer_4539 ( .C (clk), .D (new_AGEMA_signal_7969), .Q (new_AGEMA_signal_7970) ) ;
    buf_clk new_AGEMA_reg_buffer_4543 ( .C (clk), .D (new_AGEMA_signal_7973), .Q (new_AGEMA_signal_7974) ) ;
    buf_clk new_AGEMA_reg_buffer_4547 ( .C (clk), .D (new_AGEMA_signal_7977), .Q (new_AGEMA_signal_7978) ) ;
    buf_clk new_AGEMA_reg_buffer_4551 ( .C (clk), .D (new_AGEMA_signal_7981), .Q (new_AGEMA_signal_7982) ) ;
    buf_clk new_AGEMA_reg_buffer_4555 ( .C (clk), .D (new_AGEMA_signal_7985), .Q (new_AGEMA_signal_7986) ) ;
    buf_clk new_AGEMA_reg_buffer_4559 ( .C (clk), .D (new_AGEMA_signal_7989), .Q (new_AGEMA_signal_7990) ) ;
    buf_clk new_AGEMA_reg_buffer_4563 ( .C (clk), .D (new_AGEMA_signal_7993), .Q (new_AGEMA_signal_7994) ) ;
    buf_clk new_AGEMA_reg_buffer_4567 ( .C (clk), .D (new_AGEMA_signal_7997), .Q (new_AGEMA_signal_7998) ) ;
    buf_clk new_AGEMA_reg_buffer_4571 ( .C (clk), .D (new_AGEMA_signal_8001), .Q (new_AGEMA_signal_8002) ) ;
    buf_clk new_AGEMA_reg_buffer_4575 ( .C (clk), .D (new_AGEMA_signal_8005), .Q (new_AGEMA_signal_8006) ) ;
    buf_clk new_AGEMA_reg_buffer_4579 ( .C (clk), .D (new_AGEMA_signal_8009), .Q (new_AGEMA_signal_8010) ) ;
    buf_clk new_AGEMA_reg_buffer_4583 ( .C (clk), .D (new_AGEMA_signal_8013), .Q (new_AGEMA_signal_8014) ) ;
    buf_clk new_AGEMA_reg_buffer_4587 ( .C (clk), .D (new_AGEMA_signal_8017), .Q (new_AGEMA_signal_8018) ) ;
    buf_clk new_AGEMA_reg_buffer_4591 ( .C (clk), .D (new_AGEMA_signal_8021), .Q (new_AGEMA_signal_8022) ) ;
    buf_clk new_AGEMA_reg_buffer_4595 ( .C (clk), .D (new_AGEMA_signal_8025), .Q (new_AGEMA_signal_8026) ) ;
    buf_clk new_AGEMA_reg_buffer_4599 ( .C (clk), .D (new_AGEMA_signal_8029), .Q (new_AGEMA_signal_8030) ) ;
    buf_clk new_AGEMA_reg_buffer_4603 ( .C (clk), .D (new_AGEMA_signal_8033), .Q (new_AGEMA_signal_8034) ) ;
    buf_clk new_AGEMA_reg_buffer_4607 ( .C (clk), .D (new_AGEMA_signal_8037), .Q (new_AGEMA_signal_8038) ) ;
    buf_clk new_AGEMA_reg_buffer_4611 ( .C (clk), .D (new_AGEMA_signal_8041), .Q (new_AGEMA_signal_8042) ) ;
    buf_clk new_AGEMA_reg_buffer_4615 ( .C (clk), .D (new_AGEMA_signal_8045), .Q (new_AGEMA_signal_8046) ) ;
    buf_clk new_AGEMA_reg_buffer_4619 ( .C (clk), .D (new_AGEMA_signal_8049), .Q (new_AGEMA_signal_8050) ) ;
    buf_clk new_AGEMA_reg_buffer_4623 ( .C (clk), .D (new_AGEMA_signal_8053), .Q (new_AGEMA_signal_8054) ) ;
    buf_clk new_AGEMA_reg_buffer_4627 ( .C (clk), .D (new_AGEMA_signal_8057), .Q (new_AGEMA_signal_8058) ) ;
    buf_clk new_AGEMA_reg_buffer_4631 ( .C (clk), .D (new_AGEMA_signal_8061), .Q (new_AGEMA_signal_8062) ) ;
    buf_clk new_AGEMA_reg_buffer_4635 ( .C (clk), .D (new_AGEMA_signal_8065), .Q (new_AGEMA_signal_8066) ) ;
    buf_clk new_AGEMA_reg_buffer_4639 ( .C (clk), .D (new_AGEMA_signal_8069), .Q (new_AGEMA_signal_8070) ) ;
    buf_clk new_AGEMA_reg_buffer_4643 ( .C (clk), .D (new_AGEMA_signal_8073), .Q (new_AGEMA_signal_8074) ) ;
    buf_clk new_AGEMA_reg_buffer_4647 ( .C (clk), .D (new_AGEMA_signal_8077), .Q (new_AGEMA_signal_8078) ) ;
    buf_clk new_AGEMA_reg_buffer_4651 ( .C (clk), .D (new_AGEMA_signal_8081), .Q (new_AGEMA_signal_8082) ) ;
    buf_clk new_AGEMA_reg_buffer_4655 ( .C (clk), .D (new_AGEMA_signal_8085), .Q (new_AGEMA_signal_8086) ) ;
    buf_clk new_AGEMA_reg_buffer_4659 ( .C (clk), .D (new_AGEMA_signal_8089), .Q (new_AGEMA_signal_8090) ) ;
    buf_clk new_AGEMA_reg_buffer_4663 ( .C (clk), .D (new_AGEMA_signal_8093), .Q (new_AGEMA_signal_8094) ) ;
    buf_clk new_AGEMA_reg_buffer_4667 ( .C (clk), .D (new_AGEMA_signal_8097), .Q (new_AGEMA_signal_8098) ) ;
    buf_clk new_AGEMA_reg_buffer_4671 ( .C (clk), .D (new_AGEMA_signal_8101), .Q (new_AGEMA_signal_8102) ) ;
    buf_clk new_AGEMA_reg_buffer_4675 ( .C (clk), .D (new_AGEMA_signal_8105), .Q (new_AGEMA_signal_8106) ) ;
    buf_clk new_AGEMA_reg_buffer_4679 ( .C (clk), .D (new_AGEMA_signal_8109), .Q (new_AGEMA_signal_8110) ) ;
    buf_clk new_AGEMA_reg_buffer_4683 ( .C (clk), .D (new_AGEMA_signal_8113), .Q (new_AGEMA_signal_8114) ) ;
    buf_clk new_AGEMA_reg_buffer_4687 ( .C (clk), .D (new_AGEMA_signal_8117), .Q (new_AGEMA_signal_8118) ) ;
    buf_clk new_AGEMA_reg_buffer_4691 ( .C (clk), .D (new_AGEMA_signal_8121), .Q (new_AGEMA_signal_8122) ) ;
    buf_clk new_AGEMA_reg_buffer_4695 ( .C (clk), .D (new_AGEMA_signal_8125), .Q (new_AGEMA_signal_8126) ) ;
    buf_clk new_AGEMA_reg_buffer_4699 ( .C (clk), .D (new_AGEMA_signal_8129), .Q (new_AGEMA_signal_8130) ) ;
    buf_clk new_AGEMA_reg_buffer_4703 ( .C (clk), .D (new_AGEMA_signal_8133), .Q (new_AGEMA_signal_8134) ) ;
    buf_clk new_AGEMA_reg_buffer_4707 ( .C (clk), .D (new_AGEMA_signal_8137), .Q (new_AGEMA_signal_8138) ) ;
    buf_clk new_AGEMA_reg_buffer_4711 ( .C (clk), .D (new_AGEMA_signal_8141), .Q (new_AGEMA_signal_8142) ) ;
    buf_clk new_AGEMA_reg_buffer_4715 ( .C (clk), .D (new_AGEMA_signal_8145), .Q (new_AGEMA_signal_8146) ) ;
    buf_clk new_AGEMA_reg_buffer_4719 ( .C (clk), .D (new_AGEMA_signal_8149), .Q (new_AGEMA_signal_8150) ) ;
    buf_clk new_AGEMA_reg_buffer_4723 ( .C (clk), .D (new_AGEMA_signal_8153), .Q (new_AGEMA_signal_8154) ) ;
    buf_clk new_AGEMA_reg_buffer_4727 ( .C (clk), .D (new_AGEMA_signal_8157), .Q (new_AGEMA_signal_8158) ) ;
    buf_clk new_AGEMA_reg_buffer_4731 ( .C (clk), .D (new_AGEMA_signal_8161), .Q (new_AGEMA_signal_8162) ) ;
    buf_clk new_AGEMA_reg_buffer_4735 ( .C (clk), .D (new_AGEMA_signal_8165), .Q (new_AGEMA_signal_8166) ) ;
    buf_clk new_AGEMA_reg_buffer_4739 ( .C (clk), .D (new_AGEMA_signal_8169), .Q (new_AGEMA_signal_8170) ) ;
    buf_clk new_AGEMA_reg_buffer_4743 ( .C (clk), .D (new_AGEMA_signal_8173), .Q (new_AGEMA_signal_8174) ) ;
    buf_clk new_AGEMA_reg_buffer_4747 ( .C (clk), .D (new_AGEMA_signal_8177), .Q (new_AGEMA_signal_8178) ) ;
    buf_clk new_AGEMA_reg_buffer_4751 ( .C (clk), .D (new_AGEMA_signal_8181), .Q (new_AGEMA_signal_8182) ) ;
    buf_clk new_AGEMA_reg_buffer_4755 ( .C (clk), .D (new_AGEMA_signal_8185), .Q (new_AGEMA_signal_8186) ) ;
    buf_clk new_AGEMA_reg_buffer_4759 ( .C (clk), .D (new_AGEMA_signal_8189), .Q (new_AGEMA_signal_8190) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_63__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6894, new_AGEMA_signal_6892, new_AGEMA_signal_6890, new_AGEMA_signal_6888}), .Q ({Ciphertext_s3[63], Ciphertext_s2[63], Ciphertext_s1[63], Ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_62__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6902, new_AGEMA_signal_6900, new_AGEMA_signal_6898, new_AGEMA_signal_6896}), .Q ({Ciphertext_s3[62], Ciphertext_s2[62], Ciphertext_s1[62], Ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_61__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4046, new_AGEMA_signal_4045, new_AGEMA_signal_4044, StateRegInput[61]}), .Q ({Ciphertext_s3[61], Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_60__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4019, new_AGEMA_signal_4018, new_AGEMA_signal_4017, StateRegInput[60]}), .Q ({Ciphertext_s3[60], Ciphertext_s2[60], Ciphertext_s1[60], Ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_59__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6910, new_AGEMA_signal_6908, new_AGEMA_signal_6906, new_AGEMA_signal_6904}), .Q ({Ciphertext_s3[59], Ciphertext_s2[59], Ciphertext_s1[59], Ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_58__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6918, new_AGEMA_signal_6916, new_AGEMA_signal_6914, new_AGEMA_signal_6912}), .Q ({Ciphertext_s3[58], Ciphertext_s2[58], Ciphertext_s1[58], Ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_57__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3977, new_AGEMA_signal_3976, new_AGEMA_signal_3975, StateRegInput[57]}), .Q ({Ciphertext_s3[57], Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_56__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3848, new_AGEMA_signal_3847, new_AGEMA_signal_3846, StateRegInput[56]}), .Q ({Ciphertext_s3[56], Ciphertext_s2[56], Ciphertext_s1[56], Ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_55__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6926, new_AGEMA_signal_6924, new_AGEMA_signal_6922, new_AGEMA_signal_6920}), .Q ({Ciphertext_s3[55], Ciphertext_s2[55], Ciphertext_s1[55], Ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_54__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6934, new_AGEMA_signal_6932, new_AGEMA_signal_6930, new_AGEMA_signal_6928}), .Q ({Ciphertext_s3[54], Ciphertext_s2[54], Ciphertext_s1[54], Ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_53__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3971, new_AGEMA_signal_3970, new_AGEMA_signal_3969, StateRegInput[53]}), .Q ({Ciphertext_s3[53], Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_52__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3842, new_AGEMA_signal_3841, new_AGEMA_signal_3840, StateRegInput[52]}), .Q ({Ciphertext_s3[52], Ciphertext_s2[52], Ciphertext_s1[52], Ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_51__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6942, new_AGEMA_signal_6940, new_AGEMA_signal_6938, new_AGEMA_signal_6936}), .Q ({Ciphertext_s3[51], Ciphertext_s2[51], Ciphertext_s1[51], Ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_50__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6950, new_AGEMA_signal_6948, new_AGEMA_signal_6946, new_AGEMA_signal_6944}), .Q ({Ciphertext_s3[50], Ciphertext_s2[50], Ciphertext_s1[50], Ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_49__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3965, new_AGEMA_signal_3964, new_AGEMA_signal_3963, StateRegInput[49]}), .Q ({Ciphertext_s3[49], Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_48__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3836, new_AGEMA_signal_3835, new_AGEMA_signal_3834, StateRegInput[48]}), .Q ({Ciphertext_s3[48], Ciphertext_s2[48], Ciphertext_s1[48], Ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_47__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6958, new_AGEMA_signal_6956, new_AGEMA_signal_6954, new_AGEMA_signal_6952}), .Q ({Ciphertext_s3[47], Ciphertext_s2[47], Ciphertext_s1[47], Ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_46__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6966, new_AGEMA_signal_6964, new_AGEMA_signal_6962, new_AGEMA_signal_6960}), .Q ({Ciphertext_s3[46], Ciphertext_s2[46], Ciphertext_s1[46], Ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_45__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, new_AGEMA_signal_3957, StateRegInput[45]}), .Q ({Ciphertext_s3[45], Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_44__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3830, new_AGEMA_signal_3829, new_AGEMA_signal_3828, StateRegInput[44]}), .Q ({Ciphertext_s3[44], Ciphertext_s2[44], Ciphertext_s1[44], Ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_43__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6974, new_AGEMA_signal_6972, new_AGEMA_signal_6970, new_AGEMA_signal_6968}), .Q ({Ciphertext_s3[43], Ciphertext_s2[43], Ciphertext_s1[43], Ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_42__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6982, new_AGEMA_signal_6980, new_AGEMA_signal_6978, new_AGEMA_signal_6976}), .Q ({Ciphertext_s3[42], Ciphertext_s2[42], Ciphertext_s1[42], Ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_41__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3668, new_AGEMA_signal_3667, new_AGEMA_signal_3666, StateRegInput[41]}), .Q ({Ciphertext_s3[41], Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_40__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3488, new_AGEMA_signal_3487, new_AGEMA_signal_3486, StateRegInput[40]}), .Q ({Ciphertext_s3[40], Ciphertext_s2[40], Ciphertext_s1[40], Ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_39__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6990, new_AGEMA_signal_6988, new_AGEMA_signal_6986, new_AGEMA_signal_6984}), .Q ({Ciphertext_s3[39], Ciphertext_s2[39], Ciphertext_s1[39], Ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_38__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6998, new_AGEMA_signal_6996, new_AGEMA_signal_6994, new_AGEMA_signal_6992}), .Q ({Ciphertext_s3[38], Ciphertext_s2[38], Ciphertext_s1[38], Ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_37__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3662, new_AGEMA_signal_3661, new_AGEMA_signal_3660, StateRegInput[37]}), .Q ({Ciphertext_s3[37], Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_36__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3482, new_AGEMA_signal_3481, new_AGEMA_signal_3480, StateRegInput[36]}), .Q ({Ciphertext_s3[36], Ciphertext_s2[36], Ciphertext_s1[36], Ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_35__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7006, new_AGEMA_signal_7004, new_AGEMA_signal_7002, new_AGEMA_signal_7000}), .Q ({Ciphertext_s3[35], Ciphertext_s2[35], Ciphertext_s1[35], Ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_34__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7014, new_AGEMA_signal_7012, new_AGEMA_signal_7010, new_AGEMA_signal_7008}), .Q ({Ciphertext_s3[34], Ciphertext_s2[34], Ciphertext_s1[34], Ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_33__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3656, new_AGEMA_signal_3655, new_AGEMA_signal_3654, StateRegInput[33]}), .Q ({Ciphertext_s3[33], Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_32__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3476, new_AGEMA_signal_3475, new_AGEMA_signal_3474, StateRegInput[32]}), .Q ({Ciphertext_s3[32], Ciphertext_s2[32], Ciphertext_s1[32], Ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_31__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7022, new_AGEMA_signal_7020, new_AGEMA_signal_7018, new_AGEMA_signal_7016}), .Q ({Ciphertext_s3[31], Ciphertext_s2[31], Ciphertext_s1[31], Ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_30__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7030, new_AGEMA_signal_7028, new_AGEMA_signal_7026, new_AGEMA_signal_7024}), .Q ({Ciphertext_s3[30], Ciphertext_s2[30], Ciphertext_s1[30], Ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_29__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3953, new_AGEMA_signal_3952, new_AGEMA_signal_3951, StateRegInput[29]}), .Q ({Ciphertext_s3[29], Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_28__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3824, new_AGEMA_signal_3823, new_AGEMA_signal_3822, StateRegInput[28]}), .Q ({Ciphertext_s3[28], Ciphertext_s2[28], Ciphertext_s1[28], Ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_27__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7038, new_AGEMA_signal_7036, new_AGEMA_signal_7034, new_AGEMA_signal_7032}), .Q ({Ciphertext_s3[27], Ciphertext_s2[27], Ciphertext_s1[27], Ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_26__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7046, new_AGEMA_signal_7044, new_AGEMA_signal_7042, new_AGEMA_signal_7040}), .Q ({Ciphertext_s3[26], Ciphertext_s2[26], Ciphertext_s1[26], Ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_25__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4040, new_AGEMA_signal_4039, new_AGEMA_signal_4038, StateRegInput[25]}), .Q ({Ciphertext_s3[25], Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_24__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4013, new_AGEMA_signal_4012, new_AGEMA_signal_4011, StateRegInput[24]}), .Q ({Ciphertext_s3[24], Ciphertext_s2[24], Ciphertext_s1[24], Ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_23__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7054, new_AGEMA_signal_7052, new_AGEMA_signal_7050, new_AGEMA_signal_7048}), .Q ({Ciphertext_s3[23], Ciphertext_s2[23], Ciphertext_s1[23], Ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_22__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7062, new_AGEMA_signal_7060, new_AGEMA_signal_7058, new_AGEMA_signal_7056}), .Q ({Ciphertext_s3[22], Ciphertext_s2[22], Ciphertext_s1[22], Ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_21__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3941, new_AGEMA_signal_3940, new_AGEMA_signal_3939, StateRegInput[21]}), .Q ({Ciphertext_s3[21], Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_20__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3812, new_AGEMA_signal_3811, new_AGEMA_signal_3810, StateRegInput[20]}), .Q ({Ciphertext_s3[20], Ciphertext_s2[20], Ciphertext_s1[20], Ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_19__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7070, new_AGEMA_signal_7068, new_AGEMA_signal_7066, new_AGEMA_signal_7064}), .Q ({Ciphertext_s3[19], Ciphertext_s2[19], Ciphertext_s1[19], Ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_18__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7078, new_AGEMA_signal_7076, new_AGEMA_signal_7074, new_AGEMA_signal_7072}), .Q ({Ciphertext_s3[18], Ciphertext_s2[18], Ciphertext_s1[18], Ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_17__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3935, new_AGEMA_signal_3934, new_AGEMA_signal_3933, StateRegInput[17]}), .Q ({Ciphertext_s3[17], Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_16__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3806, new_AGEMA_signal_3805, new_AGEMA_signal_3804, StateRegInput[16]}), .Q ({Ciphertext_s3[16], Ciphertext_s2[16], Ciphertext_s1[16], Ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_15__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7086, new_AGEMA_signal_7084, new_AGEMA_signal_7082, new_AGEMA_signal_7080}), .Q ({Ciphertext_s3[15], Ciphertext_s2[15], Ciphertext_s1[15], Ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_14__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7094, new_AGEMA_signal_7092, new_AGEMA_signal_7090, new_AGEMA_signal_7088}), .Q ({Ciphertext_s3[14], Ciphertext_s2[14], Ciphertext_s1[14], Ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_13__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4034, new_AGEMA_signal_4033, new_AGEMA_signal_4032, StateRegInput[13]}), .Q ({Ciphertext_s3[13], Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_12__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4007, new_AGEMA_signal_4006, new_AGEMA_signal_4005, StateRegInput[12]}), .Q ({Ciphertext_s3[12], Ciphertext_s2[12], Ciphertext_s1[12], Ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_11__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7102, new_AGEMA_signal_7100, new_AGEMA_signal_7098, new_AGEMA_signal_7096}), .Q ({Ciphertext_s3[11], Ciphertext_s2[11], Ciphertext_s1[11], Ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_10__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7110, new_AGEMA_signal_7108, new_AGEMA_signal_7106, new_AGEMA_signal_7104}), .Q ({Ciphertext_s3[10], Ciphertext_s2[10], Ciphertext_s1[10], Ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_9__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3923, new_AGEMA_signal_3922, new_AGEMA_signal_3921, StateRegInput[9]}), .Q ({Ciphertext_s3[9], Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_8__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3794, new_AGEMA_signal_3793, new_AGEMA_signal_3792, StateRegInput[8]}), .Q ({Ciphertext_s3[8], Ciphertext_s2[8], Ciphertext_s1[8], Ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_7__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7118, new_AGEMA_signal_7116, new_AGEMA_signal_7114, new_AGEMA_signal_7112}), .Q ({Ciphertext_s3[7], Ciphertext_s2[7], Ciphertext_s1[7], Ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_6__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7126, new_AGEMA_signal_7124, new_AGEMA_signal_7122, new_AGEMA_signal_7120}), .Q ({Ciphertext_s3[6], Ciphertext_s2[6], Ciphertext_s1[6], Ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_5__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3917, new_AGEMA_signal_3916, new_AGEMA_signal_3915, StateRegInput[5]}), .Q ({Ciphertext_s3[5], Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_4__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3788, new_AGEMA_signal_3787, new_AGEMA_signal_3786, StateRegInput[4]}), .Q ({Ciphertext_s3[4], Ciphertext_s2[4], Ciphertext_s1[4], Ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7134, new_AGEMA_signal_7132, new_AGEMA_signal_7130, new_AGEMA_signal_7128}), .Q ({Ciphertext_s3[3], Ciphertext_s2[3], Ciphertext_s1[3], Ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7142, new_AGEMA_signal_7140, new_AGEMA_signal_7138, new_AGEMA_signal_7136}), .Q ({Ciphertext_s3[2], Ciphertext_s2[2], Ciphertext_s1[2], Ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3911, new_AGEMA_signal_3910, new_AGEMA_signal_3909, StateRegInput[1]}), .Q ({Ciphertext_s3[1], Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) StateReg_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3782, new_AGEMA_signal_3781, new_AGEMA_signal_3780, StateRegInput[0]}), .Q ({Ciphertext_s3[0], Ciphertext_s2[0], Ciphertext_s1[0], Ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7158, new_AGEMA_signal_7154, new_AGEMA_signal_7150, new_AGEMA_signal_7146}), .Q ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, new_AGEMA_signal_1731, TweakeyGeneration_key_Feedback[31]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7174, new_AGEMA_signal_7170, new_AGEMA_signal_7166, new_AGEMA_signal_7162}), .Q ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, new_AGEMA_signal_1722, TweakeyGeneration_key_Feedback[30]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7190, new_AGEMA_signal_7186, new_AGEMA_signal_7182, new_AGEMA_signal_7178}), .Q ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, new_AGEMA_signal_1713, TweakeyGeneration_key_Feedback[29]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7206, new_AGEMA_signal_7202, new_AGEMA_signal_7198, new_AGEMA_signal_7194}), .Q ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, new_AGEMA_signal_1704, TweakeyGeneration_key_Feedback[28]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7222, new_AGEMA_signal_7218, new_AGEMA_signal_7214, new_AGEMA_signal_7210}), .Q ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, new_AGEMA_signal_1695, TweakeyGeneration_key_Feedback[27]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7238, new_AGEMA_signal_7234, new_AGEMA_signal_7230, new_AGEMA_signal_7226}), .Q ({new_AGEMA_signal_1688, new_AGEMA_signal_1687, new_AGEMA_signal_1686, TweakeyGeneration_key_Feedback[26]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7254, new_AGEMA_signal_7250, new_AGEMA_signal_7246, new_AGEMA_signal_7242}), .Q ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, new_AGEMA_signal_1677, TweakeyGeneration_key_Feedback[25]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7270, new_AGEMA_signal_7266, new_AGEMA_signal_7262, new_AGEMA_signal_7258}), .Q ({new_AGEMA_signal_1670, new_AGEMA_signal_1669, new_AGEMA_signal_1668, TweakeyGeneration_key_Feedback[24]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7286, new_AGEMA_signal_7282, new_AGEMA_signal_7278, new_AGEMA_signal_7274}), .Q ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, new_AGEMA_signal_1659, TweakeyGeneration_key_Feedback[23]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7302, new_AGEMA_signal_7298, new_AGEMA_signal_7294, new_AGEMA_signal_7290}), .Q ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, new_AGEMA_signal_1650, TweakeyGeneration_key_Feedback[22]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7318, new_AGEMA_signal_7314, new_AGEMA_signal_7310, new_AGEMA_signal_7306}), .Q ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, TweakeyGeneration_key_Feedback[21]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7334, new_AGEMA_signal_7330, new_AGEMA_signal_7326, new_AGEMA_signal_7322}), .Q ({new_AGEMA_signal_1634, new_AGEMA_signal_1633, new_AGEMA_signal_1632, TweakeyGeneration_key_Feedback[20]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7350, new_AGEMA_signal_7346, new_AGEMA_signal_7342, new_AGEMA_signal_7338}), .Q ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, TweakeyGeneration_key_Feedback[19]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7366, new_AGEMA_signal_7362, new_AGEMA_signal_7358, new_AGEMA_signal_7354}), .Q ({new_AGEMA_signal_1616, new_AGEMA_signal_1615, new_AGEMA_signal_1614, TweakeyGeneration_key_Feedback[18]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7382, new_AGEMA_signal_7378, new_AGEMA_signal_7374, new_AGEMA_signal_7370}), .Q ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, TweakeyGeneration_key_Feedback[17]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7398, new_AGEMA_signal_7394, new_AGEMA_signal_7390, new_AGEMA_signal_7386}), .Q ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, new_AGEMA_signal_1596, TweakeyGeneration_key_Feedback[16]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7414, new_AGEMA_signal_7410, new_AGEMA_signal_7406, new_AGEMA_signal_7402}), .Q ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, new_AGEMA_signal_1587, TweakeyGeneration_key_Feedback[15]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7430, new_AGEMA_signal_7426, new_AGEMA_signal_7422, new_AGEMA_signal_7418}), .Q ({new_AGEMA_signal_1580, new_AGEMA_signal_1579, new_AGEMA_signal_1578, TweakeyGeneration_key_Feedback[14]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7446, new_AGEMA_signal_7442, new_AGEMA_signal_7438, new_AGEMA_signal_7434}), .Q ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, new_AGEMA_signal_1569, TweakeyGeneration_key_Feedback[13]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7462, new_AGEMA_signal_7458, new_AGEMA_signal_7454, new_AGEMA_signal_7450}), .Q ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, TweakeyGeneration_key_Feedback[12]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7478, new_AGEMA_signal_7474, new_AGEMA_signal_7470, new_AGEMA_signal_7466}), .Q ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, new_AGEMA_signal_1551, TweakeyGeneration_key_Feedback[11]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7494, new_AGEMA_signal_7490, new_AGEMA_signal_7486, new_AGEMA_signal_7482}), .Q ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, new_AGEMA_signal_1542, TweakeyGeneration_key_Feedback[10]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7510, new_AGEMA_signal_7506, new_AGEMA_signal_7502, new_AGEMA_signal_7498}), .Q ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, new_AGEMA_signal_1533, TweakeyGeneration_key_Feedback[9]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7526, new_AGEMA_signal_7522, new_AGEMA_signal_7518, new_AGEMA_signal_7514}), .Q ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, new_AGEMA_signal_1524, TweakeyGeneration_key_Feedback[8]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7542, new_AGEMA_signal_7538, new_AGEMA_signal_7534, new_AGEMA_signal_7530}), .Q ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, TweakeyGeneration_key_Feedback[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7558, new_AGEMA_signal_7554, new_AGEMA_signal_7550, new_AGEMA_signal_7546}), .Q ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, new_AGEMA_signal_1506, TweakeyGeneration_key_Feedback[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7574, new_AGEMA_signal_7570, new_AGEMA_signal_7566, new_AGEMA_signal_7562}), .Q ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, new_AGEMA_signal_1497, TweakeyGeneration_key_Feedback[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7590, new_AGEMA_signal_7586, new_AGEMA_signal_7582, new_AGEMA_signal_7578}), .Q ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, new_AGEMA_signal_1488, TweakeyGeneration_key_Feedback[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7606, new_AGEMA_signal_7602, new_AGEMA_signal_7598, new_AGEMA_signal_7594}), .Q ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, new_AGEMA_signal_1479, TweakeyGeneration_key_Feedback[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7622, new_AGEMA_signal_7618, new_AGEMA_signal_7614, new_AGEMA_signal_7610}), .Q ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, new_AGEMA_signal_1470, TweakeyGeneration_key_Feedback[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7638, new_AGEMA_signal_7634, new_AGEMA_signal_7630, new_AGEMA_signal_7626}), .Q ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, new_AGEMA_signal_1461, TweakeyGeneration_key_Feedback[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7654, new_AGEMA_signal_7650, new_AGEMA_signal_7646, new_AGEMA_signal_7642}), .Q ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, new_AGEMA_signal_1452, TweakeyGeneration_key_Feedback[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7670, new_AGEMA_signal_7666, new_AGEMA_signal_7662, new_AGEMA_signal_7658}), .Q ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, new_AGEMA_signal_1947, TweakeyGeneration_key_Feedback[55]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7686, new_AGEMA_signal_7682, new_AGEMA_signal_7678, new_AGEMA_signal_7674}), .Q ({new_AGEMA_signal_1940, new_AGEMA_signal_1939, new_AGEMA_signal_1938, TweakeyGeneration_key_Feedback[54]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7702, new_AGEMA_signal_7698, new_AGEMA_signal_7694, new_AGEMA_signal_7690}), .Q ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, new_AGEMA_signal_1929, TweakeyGeneration_key_Feedback[53]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7718, new_AGEMA_signal_7714, new_AGEMA_signal_7710, new_AGEMA_signal_7706}), .Q ({new_AGEMA_signal_1922, new_AGEMA_signal_1921, new_AGEMA_signal_1920, TweakeyGeneration_key_Feedback[52]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7734, new_AGEMA_signal_7730, new_AGEMA_signal_7726, new_AGEMA_signal_7722}), .Q ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, new_AGEMA_signal_2019, TweakeyGeneration_key_Feedback[63]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7750, new_AGEMA_signal_7746, new_AGEMA_signal_7742, new_AGEMA_signal_7738}), .Q ({new_AGEMA_signal_2012, new_AGEMA_signal_2011, new_AGEMA_signal_2010, TweakeyGeneration_key_Feedback[62]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7766, new_AGEMA_signal_7762, new_AGEMA_signal_7758, new_AGEMA_signal_7754}), .Q ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, new_AGEMA_signal_2001, TweakeyGeneration_key_Feedback[61]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7782, new_AGEMA_signal_7778, new_AGEMA_signal_7774, new_AGEMA_signal_7770}), .Q ({new_AGEMA_signal_1994, new_AGEMA_signal_1993, new_AGEMA_signal_1992, TweakeyGeneration_key_Feedback[60]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7798, new_AGEMA_signal_7794, new_AGEMA_signal_7790, new_AGEMA_signal_7786}), .Q ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, new_AGEMA_signal_1875, TweakeyGeneration_key_Feedback[47]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7814, new_AGEMA_signal_7810, new_AGEMA_signal_7806, new_AGEMA_signal_7802}), .Q ({new_AGEMA_signal_1868, new_AGEMA_signal_1867, new_AGEMA_signal_1866, TweakeyGeneration_key_Feedback[46]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7830, new_AGEMA_signal_7826, new_AGEMA_signal_7822, new_AGEMA_signal_7818}), .Q ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, new_AGEMA_signal_1857, TweakeyGeneration_key_Feedback[45]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7846, new_AGEMA_signal_7842, new_AGEMA_signal_7838, new_AGEMA_signal_7834}), .Q ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, new_AGEMA_signal_1848, TweakeyGeneration_key_Feedback[44]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7862, new_AGEMA_signal_7858, new_AGEMA_signal_7854, new_AGEMA_signal_7850}), .Q ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, new_AGEMA_signal_1767, TweakeyGeneration_key_Feedback[35]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7878, new_AGEMA_signal_7874, new_AGEMA_signal_7870, new_AGEMA_signal_7866}), .Q ({new_AGEMA_signal_1760, new_AGEMA_signal_1759, new_AGEMA_signal_1758, TweakeyGeneration_key_Feedback[34]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7894, new_AGEMA_signal_7890, new_AGEMA_signal_7886, new_AGEMA_signal_7882}), .Q ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, new_AGEMA_signal_1749, TweakeyGeneration_key_Feedback[33]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7910, new_AGEMA_signal_7906, new_AGEMA_signal_7902, new_AGEMA_signal_7898}), .Q ({new_AGEMA_signal_1742, new_AGEMA_signal_1741, new_AGEMA_signal_1740, TweakeyGeneration_key_Feedback[32]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7926, new_AGEMA_signal_7922, new_AGEMA_signal_7918, new_AGEMA_signal_7914}), .Q ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, new_AGEMA_signal_1803, TweakeyGeneration_key_Feedback[39]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7942, new_AGEMA_signal_7938, new_AGEMA_signal_7934, new_AGEMA_signal_7930}), .Q ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, new_AGEMA_signal_1794, TweakeyGeneration_key_Feedback[38]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7958, new_AGEMA_signal_7954, new_AGEMA_signal_7950, new_AGEMA_signal_7946}), .Q ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, new_AGEMA_signal_1785, TweakeyGeneration_key_Feedback[37]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7974, new_AGEMA_signal_7970, new_AGEMA_signal_7966, new_AGEMA_signal_7962}), .Q ({new_AGEMA_signal_1778, new_AGEMA_signal_1777, new_AGEMA_signal_1776, TweakeyGeneration_key_Feedback[36]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7990, new_AGEMA_signal_7986, new_AGEMA_signal_7982, new_AGEMA_signal_7978}), .Q ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, new_AGEMA_signal_1911, TweakeyGeneration_key_Feedback[51]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8006, new_AGEMA_signal_8002, new_AGEMA_signal_7998, new_AGEMA_signal_7994}), .Q ({new_AGEMA_signal_1904, new_AGEMA_signal_1903, new_AGEMA_signal_1902, TweakeyGeneration_key_Feedback[50]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8022, new_AGEMA_signal_8018, new_AGEMA_signal_8014, new_AGEMA_signal_8010}), .Q ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, new_AGEMA_signal_1893, TweakeyGeneration_key_Feedback[49]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8038, new_AGEMA_signal_8034, new_AGEMA_signal_8030, new_AGEMA_signal_8026}), .Q ({new_AGEMA_signal_1886, new_AGEMA_signal_1885, new_AGEMA_signal_1884, TweakeyGeneration_key_Feedback[48]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8054, new_AGEMA_signal_8050, new_AGEMA_signal_8046, new_AGEMA_signal_8042}), .Q ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, new_AGEMA_signal_1839, TweakeyGeneration_key_Feedback[43]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8070, new_AGEMA_signal_8066, new_AGEMA_signal_8062, new_AGEMA_signal_8058}), .Q ({new_AGEMA_signal_1832, new_AGEMA_signal_1831, new_AGEMA_signal_1830, TweakeyGeneration_key_Feedback[42]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8086, new_AGEMA_signal_8082, new_AGEMA_signal_8078, new_AGEMA_signal_8074}), .Q ({new_AGEMA_signal_1823, new_AGEMA_signal_1822, new_AGEMA_signal_1821, TweakeyGeneration_key_Feedback[41]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8102, new_AGEMA_signal_8098, new_AGEMA_signal_8094, new_AGEMA_signal_8090}), .Q ({new_AGEMA_signal_1814, new_AGEMA_signal_1813, new_AGEMA_signal_1812, TweakeyGeneration_key_Feedback[40]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8118, new_AGEMA_signal_8114, new_AGEMA_signal_8110, new_AGEMA_signal_8106}), .Q ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, new_AGEMA_signal_1983, TweakeyGeneration_key_Feedback[59]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8134, new_AGEMA_signal_8130, new_AGEMA_signal_8126, new_AGEMA_signal_8122}), .Q ({new_AGEMA_signal_1976, new_AGEMA_signal_1975, new_AGEMA_signal_1974, TweakeyGeneration_key_Feedback[58]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8150, new_AGEMA_signal_8146, new_AGEMA_signal_8142, new_AGEMA_signal_8138}), .Q ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, new_AGEMA_signal_1965, TweakeyGeneration_key_Feedback[57]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8166, new_AGEMA_signal_8162, new_AGEMA_signal_8158, new_AGEMA_signal_8154}), .Q ({new_AGEMA_signal_1958, new_AGEMA_signal_1957, new_AGEMA_signal_1956, TweakeyGeneration_key_Feedback[56]}) ) ;
    DFF_X1 FSMReg_s_current_state_reg_5__FF_FF ( .CK (clk), .D (new_AGEMA_signal_8170), .Q (FSM[5]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_4__FF_FF ( .CK (clk), .D (new_AGEMA_signal_8174), .Q (FSM[4]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_3__FF_FF ( .CK (clk), .D (new_AGEMA_signal_8178), .Q (FSMUpdate[4]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_2__FF_FF ( .CK (clk), .D (new_AGEMA_signal_8182), .Q (FSMUpdate[3]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_1__FF_FF ( .CK (clk), .D (new_AGEMA_signal_8186), .Q (FSM[1]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_0__FF_FF ( .CK (clk), .D (new_AGEMA_signal_8190), .Q (FSMUpdate[1]), .QN () ) ;
endmodule
