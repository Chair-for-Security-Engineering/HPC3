////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module Midori64 in file /AGEMA/Designs/Midori_round_based/AGEMA/Midori64.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module Midori64_HPC2_ClockGating_d3 (DataIn_s0, key_s0, clk, reset, enc_dec, key_s1, key_s2, key_s3, DataIn_s1, DataIn_s2, DataIn_s3, Fresh, DataOut_s0, done, DataOut_s1, DataOut_s2, DataOut_s3, Synch);
    input [63:0] DataIn_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input enc_dec ;
    input [127:0] key_s1 ;
    input [127:0] key_s2 ;
    input [127:0] key_s3 ;
    input [63:0] DataIn_s1 ;
    input [63:0] DataIn_s2 ;
    input [63:0] DataIn_s3 ;
    input [1535:0] Fresh ;
    output [63:0] DataOut_s0 ;
    output done ;
    output [63:0] DataOut_s1 ;
    output [63:0] DataOut_s2 ;
    output [63:0] DataOut_s3 ;
    output Synch ;
    wire controller_n2 ;
    wire controller_n1 ;
    wire controller_roundCounter_n13 ;
    wire controller_roundCounter_n12 ;
    wire controller_roundCounter_n11 ;
    wire controller_roundCounter_n10 ;
    wire controller_roundCounter_n9 ;
    wire controller_roundCounter_n8 ;
    wire controller_roundCounter_n7 ;
    wire controller_roundCounter_n5 ;
    wire controller_roundCounter_n4 ;
    wire controller_roundCounter_n3 ;
    wire controller_roundCounter_n2 ;
    wire controller_roundCounter_n1 ;
    wire controller_roundCounter_N10 ;
    wire controller_roundCounter_n6 ;
    wire controller_roundCounter_N8 ;
    wire controller_roundCounter_N7 ;
    wire Midori_rounds_n16 ;
    wire Midori_rounds_n15 ;
    wire Midori_rounds_n14 ;
    wire Midori_rounds_n13 ;
    wire Midori_rounds_n12 ;
    wire Midori_rounds_n11 ;
    wire Midori_rounds_n10 ;
    wire Midori_rounds_n9 ;
    wire Midori_rounds_n8 ;
    wire Midori_rounds_n7 ;
    wire Midori_rounds_n6 ;
    wire Midori_rounds_n5 ;
    wire Midori_rounds_n4 ;
    wire Midori_rounds_n3 ;
    wire Midori_rounds_n2 ;
    wire Midori_rounds_n1 ;
    wire Midori_rounds_SelectedKey_0_ ;
    wire Midori_rounds_SelectedKey_1_ ;
    wire Midori_rounds_SelectedKey_2_ ;
    wire Midori_rounds_SelectedKey_3_ ;
    wire Midori_rounds_SelectedKey_4_ ;
    wire Midori_rounds_SelectedKey_5_ ;
    wire Midori_rounds_SelectedKey_6_ ;
    wire Midori_rounds_SelectedKey_7_ ;
    wire Midori_rounds_SelectedKey_8_ ;
    wire Midori_rounds_SelectedKey_9_ ;
    wire Midori_rounds_SelectedKey_10_ ;
    wire Midori_rounds_SelectedKey_11_ ;
    wire Midori_rounds_SelectedKey_12_ ;
    wire Midori_rounds_SelectedKey_13_ ;
    wire Midori_rounds_SelectedKey_14_ ;
    wire Midori_rounds_SelectedKey_15_ ;
    wire Midori_rounds_SelectedKey_16_ ;
    wire Midori_rounds_SelectedKey_17_ ;
    wire Midori_rounds_SelectedKey_18_ ;
    wire Midori_rounds_SelectedKey_19_ ;
    wire Midori_rounds_SelectedKey_20_ ;
    wire Midori_rounds_SelectedKey_21_ ;
    wire Midori_rounds_SelectedKey_22_ ;
    wire Midori_rounds_SelectedKey_23_ ;
    wire Midori_rounds_SelectedKey_24_ ;
    wire Midori_rounds_SelectedKey_25_ ;
    wire Midori_rounds_SelectedKey_26_ ;
    wire Midori_rounds_SelectedKey_27_ ;
    wire Midori_rounds_SelectedKey_28_ ;
    wire Midori_rounds_SelectedKey_29_ ;
    wire Midori_rounds_SelectedKey_30_ ;
    wire Midori_rounds_SelectedKey_31_ ;
    wire Midori_rounds_SelectedKey_32_ ;
    wire Midori_rounds_SelectedKey_33_ ;
    wire Midori_rounds_SelectedKey_34_ ;
    wire Midori_rounds_SelectedKey_35_ ;
    wire Midori_rounds_SelectedKey_36_ ;
    wire Midori_rounds_SelectedKey_37_ ;
    wire Midori_rounds_SelectedKey_38_ ;
    wire Midori_rounds_SelectedKey_39_ ;
    wire Midori_rounds_SelectedKey_40_ ;
    wire Midori_rounds_SelectedKey_41_ ;
    wire Midori_rounds_SelectedKey_42_ ;
    wire Midori_rounds_SelectedKey_43_ ;
    wire Midori_rounds_SelectedKey_44_ ;
    wire Midori_rounds_SelectedKey_45_ ;
    wire Midori_rounds_SelectedKey_46_ ;
    wire Midori_rounds_SelectedKey_47_ ;
    wire Midori_rounds_SelectedKey_48_ ;
    wire Midori_rounds_SelectedKey_49_ ;
    wire Midori_rounds_SelectedKey_50_ ;
    wire Midori_rounds_SelectedKey_51_ ;
    wire Midori_rounds_SelectedKey_52_ ;
    wire Midori_rounds_SelectedKey_53_ ;
    wire Midori_rounds_SelectedKey_54_ ;
    wire Midori_rounds_SelectedKey_55_ ;
    wire Midori_rounds_SelectedKey_56_ ;
    wire Midori_rounds_SelectedKey_57_ ;
    wire Midori_rounds_SelectedKey_58_ ;
    wire Midori_rounds_SelectedKey_59_ ;
    wire Midori_rounds_SelectedKey_60_ ;
    wire Midori_rounds_SelectedKey_61_ ;
    wire Midori_rounds_SelectedKey_62_ ;
    wire Midori_rounds_SelectedKey_63_ ;
    wire Midori_rounds_constant_MUX_n217 ;
    wire Midori_rounds_constant_MUX_n216 ;
    wire Midori_rounds_constant_MUX_n215 ;
    wire Midori_rounds_constant_MUX_n214 ;
    wire Midori_rounds_constant_MUX_n213 ;
    wire Midori_rounds_constant_MUX_n212 ;
    wire Midori_rounds_constant_MUX_n211 ;
    wire Midori_rounds_constant_MUX_n210 ;
    wire Midori_rounds_constant_MUX_n209 ;
    wire Midori_rounds_constant_MUX_n208 ;
    wire Midori_rounds_constant_MUX_n207 ;
    wire Midori_rounds_constant_MUX_n206 ;
    wire Midori_rounds_constant_MUX_n205 ;
    wire Midori_rounds_constant_MUX_n204 ;
    wire Midori_rounds_constant_MUX_n203 ;
    wire Midori_rounds_constant_MUX_n202 ;
    wire Midori_rounds_constant_MUX_n201 ;
    wire Midori_rounds_constant_MUX_n200 ;
    wire Midori_rounds_constant_MUX_n199 ;
    wire Midori_rounds_constant_MUX_n198 ;
    wire Midori_rounds_constant_MUX_n197 ;
    wire Midori_rounds_constant_MUX_n196 ;
    wire Midori_rounds_constant_MUX_n195 ;
    wire Midori_rounds_constant_MUX_n194 ;
    wire Midori_rounds_constant_MUX_n193 ;
    wire Midori_rounds_constant_MUX_n192 ;
    wire Midori_rounds_constant_MUX_n191 ;
    wire Midori_rounds_constant_MUX_n190 ;
    wire Midori_rounds_constant_MUX_n189 ;
    wire Midori_rounds_constant_MUX_n188 ;
    wire Midori_rounds_constant_MUX_n187 ;
    wire Midori_rounds_constant_MUX_n186 ;
    wire Midori_rounds_constant_MUX_n185 ;
    wire Midori_rounds_constant_MUX_n184 ;
    wire Midori_rounds_constant_MUX_n183 ;
    wire Midori_rounds_constant_MUX_n182 ;
    wire Midori_rounds_constant_MUX_n181 ;
    wire Midori_rounds_constant_MUX_n180 ;
    wire Midori_rounds_constant_MUX_n179 ;
    wire Midori_rounds_constant_MUX_n178 ;
    wire Midori_rounds_constant_MUX_n177 ;
    wire Midori_rounds_constant_MUX_n176 ;
    wire Midori_rounds_constant_MUX_n175 ;
    wire Midori_rounds_constant_MUX_n174 ;
    wire Midori_rounds_constant_MUX_n173 ;
    wire Midori_rounds_constant_MUX_n172 ;
    wire Midori_rounds_constant_MUX_n171 ;
    wire Midori_rounds_constant_MUX_n170 ;
    wire Midori_rounds_constant_MUX_n169 ;
    wire Midori_rounds_constant_MUX_n168 ;
    wire Midori_rounds_constant_MUX_n167 ;
    wire Midori_rounds_constant_MUX_n166 ;
    wire Midori_rounds_constant_MUX_n165 ;
    wire Midori_rounds_constant_MUX_n164 ;
    wire Midori_rounds_constant_MUX_n163 ;
    wire Midori_rounds_constant_MUX_n162 ;
    wire Midori_rounds_constant_MUX_n161 ;
    wire Midori_rounds_constant_MUX_n160 ;
    wire Midori_rounds_constant_MUX_n159 ;
    wire Midori_rounds_constant_MUX_n158 ;
    wire Midori_rounds_constant_MUX_n157 ;
    wire Midori_rounds_constant_MUX_n156 ;
    wire Midori_rounds_constant_MUX_n155 ;
    wire Midori_rounds_constant_MUX_n154 ;
    wire Midori_rounds_constant_MUX_n153 ;
    wire Midori_rounds_constant_MUX_n152 ;
    wire Midori_rounds_constant_MUX_n151 ;
    wire Midori_rounds_constant_MUX_n150 ;
    wire Midori_rounds_constant_MUX_n149 ;
    wire Midori_rounds_constant_MUX_n148 ;
    wire Midori_rounds_constant_MUX_n147 ;
    wire Midori_rounds_constant_MUX_n146 ;
    wire Midori_rounds_constant_MUX_n145 ;
    wire Midori_rounds_constant_MUX_n144 ;
    wire Midori_rounds_constant_MUX_n143 ;
    wire Midori_rounds_constant_MUX_n142 ;
    wire Midori_rounds_constant_MUX_n141 ;
    wire Midori_rounds_constant_MUX_n140 ;
    wire Midori_rounds_constant_MUX_n139 ;
    wire Midori_rounds_constant_MUX_n138 ;
    wire Midori_rounds_constant_MUX_n137 ;
    wire Midori_rounds_constant_MUX_n136 ;
    wire Midori_rounds_constant_MUX_n135 ;
    wire Midori_rounds_constant_MUX_n134 ;
    wire Midori_rounds_constant_MUX_n133 ;
    wire Midori_rounds_constant_MUX_n132 ;
    wire Midori_rounds_constant_MUX_n131 ;
    wire Midori_rounds_constant_MUX_n130 ;
    wire Midori_rounds_constant_MUX_n129 ;
    wire Midori_rounds_constant_MUX_n128 ;
    wire Midori_rounds_MUXInst_n11 ;
    wire Midori_rounds_MUXInst_n10 ;
    wire Midori_rounds_MUXInst_n9 ;
    wire Midori_rounds_MUXInst_n8 ;
    wire Midori_rounds_roundResult_Reg_SFF_0_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_1_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_2_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_3_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_4_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_5_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_6_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_7_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_8_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_9_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_10_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_11_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_12_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_13_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_14_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_15_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_16_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_17_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_18_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_19_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_20_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_21_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_22_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_23_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_24_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_25_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_26_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_27_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_28_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_29_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_30_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_31_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_32_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_33_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_34_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_35_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_36_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_37_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_38_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_39_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_40_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_41_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_42_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_43_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_44_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_45_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_46_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_47_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_48_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_49_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_50_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_51_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_52_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_53_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_54_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_55_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_56_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_57_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_58_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_59_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_60_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_61_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_62_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_63_DQ ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n1 ;
    wire Midori_rounds_mul_MC1_n8 ;
    wire Midori_rounds_mul_MC1_n7 ;
    wire Midori_rounds_mul_MC1_n6 ;
    wire Midori_rounds_mul_MC1_n5 ;
    wire Midori_rounds_mul_MC1_n4 ;
    wire Midori_rounds_mul_MC1_n3 ;
    wire Midori_rounds_mul_MC1_n2 ;
    wire Midori_rounds_mul_MC1_n1 ;
    wire Midori_rounds_mul_MC2_n8 ;
    wire Midori_rounds_mul_MC2_n7 ;
    wire Midori_rounds_mul_MC2_n6 ;
    wire Midori_rounds_mul_MC2_n5 ;
    wire Midori_rounds_mul_MC2_n4 ;
    wire Midori_rounds_mul_MC2_n3 ;
    wire Midori_rounds_mul_MC2_n2 ;
    wire Midori_rounds_mul_MC2_n1 ;
    wire Midori_rounds_mul_MC3_n8 ;
    wire Midori_rounds_mul_MC3_n7 ;
    wire Midori_rounds_mul_MC3_n6 ;
    wire Midori_rounds_mul_MC3_n5 ;
    wire Midori_rounds_mul_MC3_n4 ;
    wire Midori_rounds_mul_MC3_n3 ;
    wire Midori_rounds_mul_MC3_n2 ;
    wire Midori_rounds_mul_MC3_n1 ;
    wire Midori_rounds_mul_MC4_n8 ;
    wire Midori_rounds_mul_MC4_n7 ;
    wire Midori_rounds_mul_MC4_n6 ;
    wire Midori_rounds_mul_MC4_n5 ;
    wire Midori_rounds_mul_MC4_n4 ;
    wire Midori_rounds_mul_MC4_n3 ;
    wire Midori_rounds_mul_MC4_n2 ;
    wire Midori_rounds_mul_MC4_n1 ;
    wire [63:0] wk ;
    wire [3:0] round_Signal ;
    wire [63:0] Midori_add_Result_Start ;
    wire [63:0] Midori_rounds_mul_ResultXORkey ;
    wire [63:0] Midori_rounds_SR_Inv_Result ;
    wire [63:0] Midori_rounds_mul_input ;
    wire [63:0] Midori_rounds_sub_ResultXORkey ;
    wire [63:0] Midori_rounds_SR_Result ;
    wire [63:0] Midori_rounds_roundReg_out ;
    wire [63:0] Midori_rounds_round_Result ;
    wire [15:0] Midori_rounds_round_Constant ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4235 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4282 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4290 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4308 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4318 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4325 ;
    wire new_AGEMA_signal_4326 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4336 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4354 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4361 ;
    wire new_AGEMA_signal_4362 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4372 ;
    wire new_AGEMA_signal_4373 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4378 ;
    wire new_AGEMA_signal_4379 ;
    wire new_AGEMA_signal_4380 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4382 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4497 ;
    wire new_AGEMA_signal_4498 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5195 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U64 ( .a ({key_s3[73], key_s2[73], key_s1[73], key_s0[73]}), .b ({key_s3[9], key_s2[9], key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_1464, new_AGEMA_signal_1463, new_AGEMA_signal_1462, wk[9]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U63 ( .a ({key_s3[72], key_s2[72], key_s1[72], key_s0[72]}), .b ({key_s3[8], key_s2[8], key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, new_AGEMA_signal_1471, wk[8]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U62 ( .a ({key_s3[71], key_s2[71], key_s1[71], key_s0[71]}), .b ({key_s3[7], key_s2[7], key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_1482, new_AGEMA_signal_1481, new_AGEMA_signal_1480, wk[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U61 ( .a ({key_s3[6], key_s2[6], key_s1[6], key_s0[6]}), .b ({key_s3[70], key_s2[70], key_s1[70], key_s0[70]}), .c ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, new_AGEMA_signal_1489, wk[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U60 ( .a ({key_s3[127], key_s2[127], key_s1[127], key_s0[127]}), .b ({key_s3[63], key_s2[63], key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_1500, new_AGEMA_signal_1499, new_AGEMA_signal_1498, wk[63]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U59 ( .a ({key_s3[126], key_s2[126], key_s1[126], key_s0[126]}), .b ({key_s3[62], key_s2[62], key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, new_AGEMA_signal_1507, wk[62]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U58 ( .a ({key_s3[125], key_s2[125], key_s1[125], key_s0[125]}), .b ({key_s3[61], key_s2[61], key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_1518, new_AGEMA_signal_1517, new_AGEMA_signal_1516, wk[61]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U57 ( .a ({key_s3[124], key_s2[124], key_s1[124], key_s0[124]}), .b ({key_s3[60], key_s2[60], key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, new_AGEMA_signal_1525, wk[60]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U56 ( .a ({key_s3[5], key_s2[5], key_s1[5], key_s0[5]}), .b ({key_s3[69], key_s2[69], key_s1[69], key_s0[69]}), .c ({new_AGEMA_signal_1536, new_AGEMA_signal_1535, new_AGEMA_signal_1534, wk[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U55 ( .a ({key_s3[123], key_s2[123], key_s1[123], key_s0[123]}), .b ({key_s3[59], key_s2[59], key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, new_AGEMA_signal_1543, wk[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U54 ( .a ({key_s3[122], key_s2[122], key_s1[122], key_s0[122]}), .b ({key_s3[58], key_s2[58], key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_1554, new_AGEMA_signal_1553, new_AGEMA_signal_1552, wk[58]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U53 ( .a ({key_s3[121], key_s2[121], key_s1[121], key_s0[121]}), .b ({key_s3[57], key_s2[57], key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_1563, new_AGEMA_signal_1562, new_AGEMA_signal_1561, wk[57]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U52 ( .a ({key_s3[120], key_s2[120], key_s1[120], key_s0[120]}), .b ({key_s3[56], key_s2[56], key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, new_AGEMA_signal_1570, wk[56]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U51 ( .a ({key_s3[119], key_s2[119], key_s1[119], key_s0[119]}), .b ({key_s3[55], key_s2[55], key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, new_AGEMA_signal_1579, wk[55]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U50 ( .a ({key_s3[118], key_s2[118], key_s1[118], key_s0[118]}), .b ({key_s3[54], key_s2[54], key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_1590, new_AGEMA_signal_1589, new_AGEMA_signal_1588, wk[54]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U49 ( .a ({key_s3[117], key_s2[117], key_s1[117], key_s0[117]}), .b ({key_s3[53], key_s2[53], key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, new_AGEMA_signal_1597, wk[53]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U48 ( .a ({key_s3[116], key_s2[116], key_s1[116], key_s0[116]}), .b ({key_s3[52], key_s2[52], key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, new_AGEMA_signal_1606, wk[52]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U47 ( .a ({key_s3[115], key_s2[115], key_s1[115], key_s0[115]}), .b ({key_s3[51], key_s2[51], key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, new_AGEMA_signal_1615, wk[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U46 ( .a ({key_s3[114], key_s2[114], key_s1[114], key_s0[114]}), .b ({key_s3[50], key_s2[50], key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_1626, new_AGEMA_signal_1625, new_AGEMA_signal_1624, wk[50]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U45 ( .a ({key_s3[4], key_s2[4], key_s1[4], key_s0[4]}), .b ({key_s3[68], key_s2[68], key_s1[68], key_s0[68]}), .c ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, new_AGEMA_signal_1633, wk[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U44 ( .a ({key_s3[113], key_s2[113], key_s1[113], key_s0[113]}), .b ({key_s3[49], key_s2[49], key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_1644, new_AGEMA_signal_1643, new_AGEMA_signal_1642, wk[49]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U43 ( .a ({key_s3[112], key_s2[112], key_s1[112], key_s0[112]}), .b ({key_s3[48], key_s2[48], key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, new_AGEMA_signal_1651, wk[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U42 ( .a ({key_s3[111], key_s2[111], key_s1[111], key_s0[111]}), .b ({key_s3[47], key_s2[47], key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_1662, new_AGEMA_signal_1661, new_AGEMA_signal_1660, wk[47]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U41 ( .a ({key_s3[110], key_s2[110], key_s1[110], key_s0[110]}), .b ({key_s3[46], key_s2[46], key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, new_AGEMA_signal_1669, wk[46]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U40 ( .a ({key_s3[109], key_s2[109], key_s1[109], key_s0[109]}), .b ({key_s3[45], key_s2[45], key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_1680, new_AGEMA_signal_1679, new_AGEMA_signal_1678, wk[45]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U39 ( .a ({key_s3[108], key_s2[108], key_s1[108], key_s0[108]}), .b ({key_s3[44], key_s2[44], key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, new_AGEMA_signal_1687, wk[44]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U38 ( .a ({key_s3[107], key_s2[107], key_s1[107], key_s0[107]}), .b ({key_s3[43], key_s2[43], key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, new_AGEMA_signal_1696, wk[43]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U37 ( .a ({key_s3[106], key_s2[106], key_s1[106], key_s0[106]}), .b ({key_s3[42], key_s2[42], key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, new_AGEMA_signal_1705, wk[42]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U36 ( .a ({key_s3[105], key_s2[105], key_s1[105], key_s0[105]}), .b ({key_s3[41], key_s2[41], key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_1716, new_AGEMA_signal_1715, new_AGEMA_signal_1714, wk[41]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U35 ( .a ({key_s3[104], key_s2[104], key_s1[104], key_s0[104]}), .b ({key_s3[40], key_s2[40], key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, new_AGEMA_signal_1723, wk[40]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U34 ( .a ({key_s3[3], key_s2[3], key_s1[3], key_s0[3]}), .b ({key_s3[67], key_s2[67], key_s1[67], key_s0[67]}), .c ({new_AGEMA_signal_1734, new_AGEMA_signal_1733, new_AGEMA_signal_1732, wk[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U33 ( .a ({key_s3[103], key_s2[103], key_s1[103], key_s0[103]}), .b ({key_s3[39], key_s2[39], key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, new_AGEMA_signal_1741, wk[39]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U32 ( .a ({key_s3[102], key_s2[102], key_s1[102], key_s0[102]}), .b ({key_s3[38], key_s2[38], key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_1752, new_AGEMA_signal_1751, new_AGEMA_signal_1750, wk[38]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U31 ( .a ({key_s3[101], key_s2[101], key_s1[101], key_s0[101]}), .b ({key_s3[37], key_s2[37], key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, new_AGEMA_signal_1759, wk[37]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U30 ( .a ({key_s3[100], key_s2[100], key_s1[100], key_s0[100]}), .b ({key_s3[36], key_s2[36], key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, new_AGEMA_signal_1768, wk[36]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U29 ( .a ({key_s3[35], key_s2[35], key_s1[35], key_s0[35]}), .b ({key_s3[99], key_s2[99], key_s1[99], key_s0[99]}), .c ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, new_AGEMA_signal_1777, wk[35]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U28 ( .a ({key_s3[34], key_s2[34], key_s1[34], key_s0[34]}), .b ({key_s3[98], key_s2[98], key_s1[98], key_s0[98]}), .c ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, new_AGEMA_signal_1786, wk[34]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U27 ( .a ({key_s3[33], key_s2[33], key_s1[33], key_s0[33]}), .b ({key_s3[97], key_s2[97], key_s1[97], key_s0[97]}), .c ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, new_AGEMA_signal_1795, wk[33]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U26 ( .a ({key_s3[32], key_s2[32], key_s1[32], key_s0[32]}), .b ({key_s3[96], key_s2[96], key_s1[96], key_s0[96]}), .c ({new_AGEMA_signal_1806, new_AGEMA_signal_1805, new_AGEMA_signal_1804, wk[32]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U25 ( .a ({key_s3[31], key_s2[31], key_s1[31], key_s0[31]}), .b ({key_s3[95], key_s2[95], key_s1[95], key_s0[95]}), .c ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, new_AGEMA_signal_1813, wk[31]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U24 ( .a ({key_s3[30], key_s2[30], key_s1[30], key_s0[30]}), .b ({key_s3[94], key_s2[94], key_s1[94], key_s0[94]}), .c ({new_AGEMA_signal_1824, new_AGEMA_signal_1823, new_AGEMA_signal_1822, wk[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U23 ( .a ({key_s3[2], key_s2[2], key_s1[2], key_s0[2]}), .b ({key_s3[66], key_s2[66], key_s1[66], key_s0[66]}), .c ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, new_AGEMA_signal_1831, wk[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U22 ( .a ({key_s3[29], key_s2[29], key_s1[29], key_s0[29]}), .b ({key_s3[93], key_s2[93], key_s1[93], key_s0[93]}), .c ({new_AGEMA_signal_1842, new_AGEMA_signal_1841, new_AGEMA_signal_1840, wk[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U21 ( .a ({key_s3[28], key_s2[28], key_s1[28], key_s0[28]}), .b ({key_s3[92], key_s2[92], key_s1[92], key_s0[92]}), .c ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, new_AGEMA_signal_1849, wk[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U20 ( .a ({key_s3[27], key_s2[27], key_s1[27], key_s0[27]}), .b ({key_s3[91], key_s2[91], key_s1[91], key_s0[91]}), .c ({new_AGEMA_signal_1860, new_AGEMA_signal_1859, new_AGEMA_signal_1858, wk[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U19 ( .a ({key_s3[26], key_s2[26], key_s1[26], key_s0[26]}), .b ({key_s3[90], key_s2[90], key_s1[90], key_s0[90]}), .c ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, new_AGEMA_signal_1867, wk[26]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U18 ( .a ({key_s3[25], key_s2[25], key_s1[25], key_s0[25]}), .b ({key_s3[89], key_s2[89], key_s1[89], key_s0[89]}), .c ({new_AGEMA_signal_1878, new_AGEMA_signal_1877, new_AGEMA_signal_1876, wk[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U17 ( .a ({key_s3[24], key_s2[24], key_s1[24], key_s0[24]}), .b ({key_s3[88], key_s2[88], key_s1[88], key_s0[88]}), .c ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, new_AGEMA_signal_1885, wk[24]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U16 ( .a ({key_s3[23], key_s2[23], key_s1[23], key_s0[23]}), .b ({key_s3[87], key_s2[87], key_s1[87], key_s0[87]}), .c ({new_AGEMA_signal_1896, new_AGEMA_signal_1895, new_AGEMA_signal_1894, wk[23]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U15 ( .a ({key_s3[22], key_s2[22], key_s1[22], key_s0[22]}), .b ({key_s3[86], key_s2[86], key_s1[86], key_s0[86]}), .c ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, new_AGEMA_signal_1903, wk[22]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U14 ( .a ({key_s3[21], key_s2[21], key_s1[21], key_s0[21]}), .b ({key_s3[85], key_s2[85], key_s1[85], key_s0[85]}), .c ({new_AGEMA_signal_1914, new_AGEMA_signal_1913, new_AGEMA_signal_1912, wk[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U13 ( .a ({key_s3[20], key_s2[20], key_s1[20], key_s0[20]}), .b ({key_s3[84], key_s2[84], key_s1[84], key_s0[84]}), .c ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, new_AGEMA_signal_1921, wk[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U12 ( .a ({key_s3[1], key_s2[1], key_s1[1], key_s0[1]}), .b ({key_s3[65], key_s2[65], key_s1[65], key_s0[65]}), .c ({new_AGEMA_signal_1932, new_AGEMA_signal_1931, new_AGEMA_signal_1930, wk[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U11 ( .a ({key_s3[19], key_s2[19], key_s1[19], key_s0[19]}), .b ({key_s3[83], key_s2[83], key_s1[83], key_s0[83]}), .c ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, new_AGEMA_signal_1939, wk[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U10 ( .a ({key_s3[18], key_s2[18], key_s1[18], key_s0[18]}), .b ({key_s3[82], key_s2[82], key_s1[82], key_s0[82]}), .c ({new_AGEMA_signal_1950, new_AGEMA_signal_1949, new_AGEMA_signal_1948, wk[18]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U9 ( .a ({key_s3[17], key_s2[17], key_s1[17], key_s0[17]}), .b ({key_s3[81], key_s2[81], key_s1[81], key_s0[81]}), .c ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, new_AGEMA_signal_1957, wk[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U8 ( .a ({key_s3[16], key_s2[16], key_s1[16], key_s0[16]}), .b ({key_s3[80], key_s2[80], key_s1[80], key_s0[80]}), .c ({new_AGEMA_signal_1968, new_AGEMA_signal_1967, new_AGEMA_signal_1966, wk[16]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U7 ( .a ({key_s3[15], key_s2[15], key_s1[15], key_s0[15]}), .b ({key_s3[79], key_s2[79], key_s1[79], key_s0[79]}), .c ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, new_AGEMA_signal_1975, wk[15]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U6 ( .a ({key_s3[14], key_s2[14], key_s1[14], key_s0[14]}), .b ({key_s3[78], key_s2[78], key_s1[78], key_s0[78]}), .c ({new_AGEMA_signal_1986, new_AGEMA_signal_1985, new_AGEMA_signal_1984, wk[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U5 ( .a ({key_s3[13], key_s2[13], key_s1[13], key_s0[13]}), .b ({key_s3[77], key_s2[77], key_s1[77], key_s0[77]}), .c ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, new_AGEMA_signal_1993, wk[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U4 ( .a ({key_s3[12], key_s2[12], key_s1[12], key_s0[12]}), .b ({key_s3[76], key_s2[76], key_s1[76], key_s0[76]}), .c ({new_AGEMA_signal_2004, new_AGEMA_signal_2003, new_AGEMA_signal_2002, wk[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U3 ( .a ({key_s3[11], key_s2[11], key_s1[11], key_s0[11]}), .b ({key_s3[75], key_s2[75], key_s1[75], key_s0[75]}), .c ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, new_AGEMA_signal_2011, wk[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U2 ( .a ({key_s3[10], key_s2[10], key_s1[10], key_s0[10]}), .b ({key_s3[74], key_s2[74], key_s1[74], key_s0[74]}), .c ({new_AGEMA_signal_2022, new_AGEMA_signal_2021, new_AGEMA_signal_2020, wk[10]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) keys_U1 ( .a ({key_s3[0], key_s2[0], key_s1[0], key_s0[0]}), .b ({key_s3[64], key_s2[64], key_s1[64], key_s0[64]}), .c ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, new_AGEMA_signal_2029, wk[0]}) ) ;
    NOR2_X1 controller_U3 ( .A1 (controller_n2), .A2 (controller_n1), .ZN (done) ) ;
    NAND2_X1 controller_U2 ( .A1 (round_Signal[0]), .A2 (round_Signal[1]), .ZN (controller_n1) ) ;
    NAND2_X1 controller_U1 ( .A1 (round_Signal[2]), .A2 (round_Signal[3]), .ZN (controller_n2) ) ;
    INV_X1 controller_roundCounter_U14 ( .A (controller_roundCounter_n13), .ZN (controller_roundCounter_n2) ) ;
    MUX2_X1 controller_roundCounter_U13 ( .S (controller_roundCounter_n6), .A (controller_roundCounter_n12), .B (controller_roundCounter_n11), .Z (controller_roundCounter_n13) ) ;
    NOR2_X1 controller_roundCounter_U12 ( .A1 (reset), .A2 (controller_roundCounter_n10), .ZN (controller_roundCounter_N8) ) ;
    XNOR2_X1 controller_roundCounter_U11 ( .A (round_Signal[0]), .B (round_Signal[1]), .ZN (controller_roundCounter_n10) ) ;
    MUX2_X1 controller_roundCounter_U10 ( .S (round_Signal[3]), .A (controller_roundCounter_n9), .B (controller_roundCounter_n8), .Z (controller_roundCounter_N10) ) ;
    NAND2_X1 controller_roundCounter_U9 ( .A1 (controller_roundCounter_n12), .A2 (controller_roundCounter_n7), .ZN (controller_roundCounter_n8) ) ;
    NAND2_X1 controller_roundCounter_U8 ( .A1 (controller_roundCounter_n6), .A2 (controller_roundCounter_n3), .ZN (controller_roundCounter_n7) ) ;
    NOR2_X1 controller_roundCounter_U7 ( .A1 (controller_roundCounter_n5), .A2 (controller_roundCounter_N7), .ZN (controller_roundCounter_n12) ) ;
    NOR2_X1 controller_roundCounter_U6 ( .A1 (round_Signal[1]), .A2 (reset), .ZN (controller_roundCounter_n5) ) ;
    NOR2_X1 controller_roundCounter_U5 ( .A1 (controller_roundCounter_n6), .A2 (controller_roundCounter_n11), .ZN (controller_roundCounter_n9) ) ;
    NAND2_X1 controller_roundCounter_U4 ( .A1 (round_Signal[1]), .A2 (controller_roundCounter_n4), .ZN (controller_roundCounter_n11) ) ;
    NOR2_X1 controller_roundCounter_U3 ( .A1 (reset), .A2 (controller_roundCounter_n1), .ZN (controller_roundCounter_n4) ) ;
    NOR2_X1 controller_roundCounter_U2 ( .A1 (reset), .A2 (round_Signal[0]), .ZN (controller_roundCounter_N7) ) ;
    INV_X1 controller_roundCounter_U1 ( .A (reset), .ZN (controller_roundCounter_n3) ) ;
    INV_X1 controller_roundCounter_count_reg_0__U1 ( .A (round_Signal[0]), .ZN (controller_roundCounter_n1) ) ;
    INV_X1 controller_roundCounter_count_reg_2__U1 ( .A (round_Signal[2]), .ZN (controller_roundCounter_n6) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U64 ( .a ({new_AGEMA_signal_1464, new_AGEMA_signal_1463, new_AGEMA_signal_1462, wk[9]}), .b ({DataIn_s3[9], DataIn_s2[9], DataIn_s1[9], DataIn_s0[9]}), .c ({new_AGEMA_signal_2460, new_AGEMA_signal_2459, new_AGEMA_signal_2458, Midori_add_Result_Start[9]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U63 ( .a ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, new_AGEMA_signal_1471, wk[8]}), .b ({DataIn_s3[8], DataIn_s2[8], DataIn_s1[8], DataIn_s0[8]}), .c ({new_AGEMA_signal_2466, new_AGEMA_signal_2465, new_AGEMA_signal_2464, Midori_add_Result_Start[8]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U62 ( .a ({new_AGEMA_signal_1482, new_AGEMA_signal_1481, new_AGEMA_signal_1480, wk[7]}), .b ({DataIn_s3[7], DataIn_s2[7], DataIn_s1[7], DataIn_s0[7]}), .c ({new_AGEMA_signal_2472, new_AGEMA_signal_2471, new_AGEMA_signal_2470, Midori_add_Result_Start[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U61 ( .a ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, new_AGEMA_signal_1489, wk[6]}), .b ({DataIn_s3[6], DataIn_s2[6], DataIn_s1[6], DataIn_s0[6]}), .c ({new_AGEMA_signal_2478, new_AGEMA_signal_2477, new_AGEMA_signal_2476, Midori_add_Result_Start[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U60 ( .a ({new_AGEMA_signal_1500, new_AGEMA_signal_1499, new_AGEMA_signal_1498, wk[63]}), .b ({DataIn_s3[63], DataIn_s2[63], DataIn_s1[63], DataIn_s0[63]}), .c ({new_AGEMA_signal_2484, new_AGEMA_signal_2483, new_AGEMA_signal_2482, Midori_add_Result_Start[63]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U59 ( .a ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, new_AGEMA_signal_1507, wk[62]}), .b ({DataIn_s3[62], DataIn_s2[62], DataIn_s1[62], DataIn_s0[62]}), .c ({new_AGEMA_signal_2490, new_AGEMA_signal_2489, new_AGEMA_signal_2488, Midori_add_Result_Start[62]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U58 ( .a ({new_AGEMA_signal_1518, new_AGEMA_signal_1517, new_AGEMA_signal_1516, wk[61]}), .b ({DataIn_s3[61], DataIn_s2[61], DataIn_s1[61], DataIn_s0[61]}), .c ({new_AGEMA_signal_2496, new_AGEMA_signal_2495, new_AGEMA_signal_2494, Midori_add_Result_Start[61]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U57 ( .a ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, new_AGEMA_signal_1525, wk[60]}), .b ({DataIn_s3[60], DataIn_s2[60], DataIn_s1[60], DataIn_s0[60]}), .c ({new_AGEMA_signal_2502, new_AGEMA_signal_2501, new_AGEMA_signal_2500, Midori_add_Result_Start[60]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U56 ( .a ({new_AGEMA_signal_1536, new_AGEMA_signal_1535, new_AGEMA_signal_1534, wk[5]}), .b ({DataIn_s3[5], DataIn_s2[5], DataIn_s1[5], DataIn_s0[5]}), .c ({new_AGEMA_signal_2508, new_AGEMA_signal_2507, new_AGEMA_signal_2506, Midori_add_Result_Start[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U55 ( .a ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, new_AGEMA_signal_1543, wk[59]}), .b ({DataIn_s3[59], DataIn_s2[59], DataIn_s1[59], DataIn_s0[59]}), .c ({new_AGEMA_signal_2514, new_AGEMA_signal_2513, new_AGEMA_signal_2512, Midori_add_Result_Start[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U54 ( .a ({new_AGEMA_signal_1554, new_AGEMA_signal_1553, new_AGEMA_signal_1552, wk[58]}), .b ({DataIn_s3[58], DataIn_s2[58], DataIn_s1[58], DataIn_s0[58]}), .c ({new_AGEMA_signal_2520, new_AGEMA_signal_2519, new_AGEMA_signal_2518, Midori_add_Result_Start[58]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U53 ( .a ({new_AGEMA_signal_1563, new_AGEMA_signal_1562, new_AGEMA_signal_1561, wk[57]}), .b ({DataIn_s3[57], DataIn_s2[57], DataIn_s1[57], DataIn_s0[57]}), .c ({new_AGEMA_signal_2526, new_AGEMA_signal_2525, new_AGEMA_signal_2524, Midori_add_Result_Start[57]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U52 ( .a ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, new_AGEMA_signal_1570, wk[56]}), .b ({DataIn_s3[56], DataIn_s2[56], DataIn_s1[56], DataIn_s0[56]}), .c ({new_AGEMA_signal_2532, new_AGEMA_signal_2531, new_AGEMA_signal_2530, Midori_add_Result_Start[56]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U51 ( .a ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, new_AGEMA_signal_1579, wk[55]}), .b ({DataIn_s3[55], DataIn_s2[55], DataIn_s1[55], DataIn_s0[55]}), .c ({new_AGEMA_signal_2538, new_AGEMA_signal_2537, new_AGEMA_signal_2536, Midori_add_Result_Start[55]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U50 ( .a ({new_AGEMA_signal_1590, new_AGEMA_signal_1589, new_AGEMA_signal_1588, wk[54]}), .b ({DataIn_s3[54], DataIn_s2[54], DataIn_s1[54], DataIn_s0[54]}), .c ({new_AGEMA_signal_2544, new_AGEMA_signal_2543, new_AGEMA_signal_2542, Midori_add_Result_Start[54]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U49 ( .a ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, new_AGEMA_signal_1597, wk[53]}), .b ({DataIn_s3[53], DataIn_s2[53], DataIn_s1[53], DataIn_s0[53]}), .c ({new_AGEMA_signal_2550, new_AGEMA_signal_2549, new_AGEMA_signal_2548, Midori_add_Result_Start[53]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U48 ( .a ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, new_AGEMA_signal_1606, wk[52]}), .b ({DataIn_s3[52], DataIn_s2[52], DataIn_s1[52], DataIn_s0[52]}), .c ({new_AGEMA_signal_2556, new_AGEMA_signal_2555, new_AGEMA_signal_2554, Midori_add_Result_Start[52]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U47 ( .a ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, new_AGEMA_signal_1615, wk[51]}), .b ({DataIn_s3[51], DataIn_s2[51], DataIn_s1[51], DataIn_s0[51]}), .c ({new_AGEMA_signal_2562, new_AGEMA_signal_2561, new_AGEMA_signal_2560, Midori_add_Result_Start[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U46 ( .a ({new_AGEMA_signal_1626, new_AGEMA_signal_1625, new_AGEMA_signal_1624, wk[50]}), .b ({DataIn_s3[50], DataIn_s2[50], DataIn_s1[50], DataIn_s0[50]}), .c ({new_AGEMA_signal_2568, new_AGEMA_signal_2567, new_AGEMA_signal_2566, Midori_add_Result_Start[50]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U45 ( .a ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, new_AGEMA_signal_1633, wk[4]}), .b ({DataIn_s3[4], DataIn_s2[4], DataIn_s1[4], DataIn_s0[4]}), .c ({new_AGEMA_signal_2574, new_AGEMA_signal_2573, new_AGEMA_signal_2572, Midori_add_Result_Start[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U44 ( .a ({new_AGEMA_signal_1644, new_AGEMA_signal_1643, new_AGEMA_signal_1642, wk[49]}), .b ({DataIn_s3[49], DataIn_s2[49], DataIn_s1[49], DataIn_s0[49]}), .c ({new_AGEMA_signal_2580, new_AGEMA_signal_2579, new_AGEMA_signal_2578, Midori_add_Result_Start[49]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U43 ( .a ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, new_AGEMA_signal_1651, wk[48]}), .b ({DataIn_s3[48], DataIn_s2[48], DataIn_s1[48], DataIn_s0[48]}), .c ({new_AGEMA_signal_2586, new_AGEMA_signal_2585, new_AGEMA_signal_2584, Midori_add_Result_Start[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U42 ( .a ({new_AGEMA_signal_1662, new_AGEMA_signal_1661, new_AGEMA_signal_1660, wk[47]}), .b ({DataIn_s3[47], DataIn_s2[47], DataIn_s1[47], DataIn_s0[47]}), .c ({new_AGEMA_signal_2592, new_AGEMA_signal_2591, new_AGEMA_signal_2590, Midori_add_Result_Start[47]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U41 ( .a ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, new_AGEMA_signal_1669, wk[46]}), .b ({DataIn_s3[46], DataIn_s2[46], DataIn_s1[46], DataIn_s0[46]}), .c ({new_AGEMA_signal_2598, new_AGEMA_signal_2597, new_AGEMA_signal_2596, Midori_add_Result_Start[46]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U40 ( .a ({new_AGEMA_signal_1680, new_AGEMA_signal_1679, new_AGEMA_signal_1678, wk[45]}), .b ({DataIn_s3[45], DataIn_s2[45], DataIn_s1[45], DataIn_s0[45]}), .c ({new_AGEMA_signal_2604, new_AGEMA_signal_2603, new_AGEMA_signal_2602, Midori_add_Result_Start[45]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U39 ( .a ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, new_AGEMA_signal_1687, wk[44]}), .b ({DataIn_s3[44], DataIn_s2[44], DataIn_s1[44], DataIn_s0[44]}), .c ({new_AGEMA_signal_2610, new_AGEMA_signal_2609, new_AGEMA_signal_2608, Midori_add_Result_Start[44]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U38 ( .a ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, new_AGEMA_signal_1696, wk[43]}), .b ({DataIn_s3[43], DataIn_s2[43], DataIn_s1[43], DataIn_s0[43]}), .c ({new_AGEMA_signal_2616, new_AGEMA_signal_2615, new_AGEMA_signal_2614, Midori_add_Result_Start[43]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U37 ( .a ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, new_AGEMA_signal_1705, wk[42]}), .b ({DataIn_s3[42], DataIn_s2[42], DataIn_s1[42], DataIn_s0[42]}), .c ({new_AGEMA_signal_2622, new_AGEMA_signal_2621, new_AGEMA_signal_2620, Midori_add_Result_Start[42]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U36 ( .a ({new_AGEMA_signal_1716, new_AGEMA_signal_1715, new_AGEMA_signal_1714, wk[41]}), .b ({DataIn_s3[41], DataIn_s2[41], DataIn_s1[41], DataIn_s0[41]}), .c ({new_AGEMA_signal_2628, new_AGEMA_signal_2627, new_AGEMA_signal_2626, Midori_add_Result_Start[41]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U35 ( .a ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, new_AGEMA_signal_1723, wk[40]}), .b ({DataIn_s3[40], DataIn_s2[40], DataIn_s1[40], DataIn_s0[40]}), .c ({new_AGEMA_signal_2634, new_AGEMA_signal_2633, new_AGEMA_signal_2632, Midori_add_Result_Start[40]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U34 ( .a ({new_AGEMA_signal_1734, new_AGEMA_signal_1733, new_AGEMA_signal_1732, wk[3]}), .b ({DataIn_s3[3], DataIn_s2[3], DataIn_s1[3], DataIn_s0[3]}), .c ({new_AGEMA_signal_2640, new_AGEMA_signal_2639, new_AGEMA_signal_2638, Midori_add_Result_Start[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U33 ( .a ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, new_AGEMA_signal_1741, wk[39]}), .b ({DataIn_s3[39], DataIn_s2[39], DataIn_s1[39], DataIn_s0[39]}), .c ({new_AGEMA_signal_2646, new_AGEMA_signal_2645, new_AGEMA_signal_2644, Midori_add_Result_Start[39]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U32 ( .a ({new_AGEMA_signal_1752, new_AGEMA_signal_1751, new_AGEMA_signal_1750, wk[38]}), .b ({DataIn_s3[38], DataIn_s2[38], DataIn_s1[38], DataIn_s0[38]}), .c ({new_AGEMA_signal_2652, new_AGEMA_signal_2651, new_AGEMA_signal_2650, Midori_add_Result_Start[38]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U31 ( .a ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, new_AGEMA_signal_1759, wk[37]}), .b ({DataIn_s3[37], DataIn_s2[37], DataIn_s1[37], DataIn_s0[37]}), .c ({new_AGEMA_signal_2658, new_AGEMA_signal_2657, new_AGEMA_signal_2656, Midori_add_Result_Start[37]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U30 ( .a ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, new_AGEMA_signal_1768, wk[36]}), .b ({DataIn_s3[36], DataIn_s2[36], DataIn_s1[36], DataIn_s0[36]}), .c ({new_AGEMA_signal_2664, new_AGEMA_signal_2663, new_AGEMA_signal_2662, Midori_add_Result_Start[36]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U29 ( .a ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, new_AGEMA_signal_1777, wk[35]}), .b ({DataIn_s3[35], DataIn_s2[35], DataIn_s1[35], DataIn_s0[35]}), .c ({new_AGEMA_signal_2670, new_AGEMA_signal_2669, new_AGEMA_signal_2668, Midori_add_Result_Start[35]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U28 ( .a ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, new_AGEMA_signal_1786, wk[34]}), .b ({DataIn_s3[34], DataIn_s2[34], DataIn_s1[34], DataIn_s0[34]}), .c ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, new_AGEMA_signal_2674, Midori_add_Result_Start[34]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U27 ( .a ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, new_AGEMA_signal_1795, wk[33]}), .b ({DataIn_s3[33], DataIn_s2[33], DataIn_s1[33], DataIn_s0[33]}), .c ({new_AGEMA_signal_2682, new_AGEMA_signal_2681, new_AGEMA_signal_2680, Midori_add_Result_Start[33]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U26 ( .a ({new_AGEMA_signal_1806, new_AGEMA_signal_1805, new_AGEMA_signal_1804, wk[32]}), .b ({DataIn_s3[32], DataIn_s2[32], DataIn_s1[32], DataIn_s0[32]}), .c ({new_AGEMA_signal_2688, new_AGEMA_signal_2687, new_AGEMA_signal_2686, Midori_add_Result_Start[32]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U25 ( .a ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, new_AGEMA_signal_1813, wk[31]}), .b ({DataIn_s3[31], DataIn_s2[31], DataIn_s1[31], DataIn_s0[31]}), .c ({new_AGEMA_signal_2694, new_AGEMA_signal_2693, new_AGEMA_signal_2692, Midori_add_Result_Start[31]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U24 ( .a ({new_AGEMA_signal_1824, new_AGEMA_signal_1823, new_AGEMA_signal_1822, wk[30]}), .b ({DataIn_s3[30], DataIn_s2[30], DataIn_s1[30], DataIn_s0[30]}), .c ({new_AGEMA_signal_2700, new_AGEMA_signal_2699, new_AGEMA_signal_2698, Midori_add_Result_Start[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U23 ( .a ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, new_AGEMA_signal_1831, wk[2]}), .b ({DataIn_s3[2], DataIn_s2[2], DataIn_s1[2], DataIn_s0[2]}), .c ({new_AGEMA_signal_2706, new_AGEMA_signal_2705, new_AGEMA_signal_2704, Midori_add_Result_Start[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U22 ( .a ({new_AGEMA_signal_1842, new_AGEMA_signal_1841, new_AGEMA_signal_1840, wk[29]}), .b ({DataIn_s3[29], DataIn_s2[29], DataIn_s1[29], DataIn_s0[29]}), .c ({new_AGEMA_signal_2712, new_AGEMA_signal_2711, new_AGEMA_signal_2710, Midori_add_Result_Start[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U21 ( .a ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, new_AGEMA_signal_1849, wk[28]}), .b ({DataIn_s3[28], DataIn_s2[28], DataIn_s1[28], DataIn_s0[28]}), .c ({new_AGEMA_signal_2718, new_AGEMA_signal_2717, new_AGEMA_signal_2716, Midori_add_Result_Start[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U20 ( .a ({new_AGEMA_signal_1860, new_AGEMA_signal_1859, new_AGEMA_signal_1858, wk[27]}), .b ({DataIn_s3[27], DataIn_s2[27], DataIn_s1[27], DataIn_s0[27]}), .c ({new_AGEMA_signal_2724, new_AGEMA_signal_2723, new_AGEMA_signal_2722, Midori_add_Result_Start[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U19 ( .a ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, new_AGEMA_signal_1867, wk[26]}), .b ({DataIn_s3[26], DataIn_s2[26], DataIn_s1[26], DataIn_s0[26]}), .c ({new_AGEMA_signal_2730, new_AGEMA_signal_2729, new_AGEMA_signal_2728, Midori_add_Result_Start[26]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U18 ( .a ({new_AGEMA_signal_1878, new_AGEMA_signal_1877, new_AGEMA_signal_1876, wk[25]}), .b ({DataIn_s3[25], DataIn_s2[25], DataIn_s1[25], DataIn_s0[25]}), .c ({new_AGEMA_signal_2736, new_AGEMA_signal_2735, new_AGEMA_signal_2734, Midori_add_Result_Start[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U17 ( .a ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, new_AGEMA_signal_1885, wk[24]}), .b ({DataIn_s3[24], DataIn_s2[24], DataIn_s1[24], DataIn_s0[24]}), .c ({new_AGEMA_signal_2742, new_AGEMA_signal_2741, new_AGEMA_signal_2740, Midori_add_Result_Start[24]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U16 ( .a ({new_AGEMA_signal_1896, new_AGEMA_signal_1895, new_AGEMA_signal_1894, wk[23]}), .b ({DataIn_s3[23], DataIn_s2[23], DataIn_s1[23], DataIn_s0[23]}), .c ({new_AGEMA_signal_2748, new_AGEMA_signal_2747, new_AGEMA_signal_2746, Midori_add_Result_Start[23]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U15 ( .a ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, new_AGEMA_signal_1903, wk[22]}), .b ({DataIn_s3[22], DataIn_s2[22], DataIn_s1[22], DataIn_s0[22]}), .c ({new_AGEMA_signal_2754, new_AGEMA_signal_2753, new_AGEMA_signal_2752, Midori_add_Result_Start[22]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U14 ( .a ({new_AGEMA_signal_1914, new_AGEMA_signal_1913, new_AGEMA_signal_1912, wk[21]}), .b ({DataIn_s3[21], DataIn_s2[21], DataIn_s1[21], DataIn_s0[21]}), .c ({new_AGEMA_signal_2760, new_AGEMA_signal_2759, new_AGEMA_signal_2758, Midori_add_Result_Start[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U13 ( .a ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, new_AGEMA_signal_1921, wk[20]}), .b ({DataIn_s3[20], DataIn_s2[20], DataIn_s1[20], DataIn_s0[20]}), .c ({new_AGEMA_signal_2766, new_AGEMA_signal_2765, new_AGEMA_signal_2764, Midori_add_Result_Start[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U12 ( .a ({new_AGEMA_signal_1932, new_AGEMA_signal_1931, new_AGEMA_signal_1930, wk[1]}), .b ({DataIn_s3[1], DataIn_s2[1], DataIn_s1[1], DataIn_s0[1]}), .c ({new_AGEMA_signal_2772, new_AGEMA_signal_2771, new_AGEMA_signal_2770, Midori_add_Result_Start[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U11 ( .a ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, new_AGEMA_signal_1939, wk[19]}), .b ({DataIn_s3[19], DataIn_s2[19], DataIn_s1[19], DataIn_s0[19]}), .c ({new_AGEMA_signal_2778, new_AGEMA_signal_2777, new_AGEMA_signal_2776, Midori_add_Result_Start[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U10 ( .a ({new_AGEMA_signal_1950, new_AGEMA_signal_1949, new_AGEMA_signal_1948, wk[18]}), .b ({DataIn_s3[18], DataIn_s2[18], DataIn_s1[18], DataIn_s0[18]}), .c ({new_AGEMA_signal_2784, new_AGEMA_signal_2783, new_AGEMA_signal_2782, Midori_add_Result_Start[18]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U9 ( .a ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, new_AGEMA_signal_1957, wk[17]}), .b ({DataIn_s3[17], DataIn_s2[17], DataIn_s1[17], DataIn_s0[17]}), .c ({new_AGEMA_signal_2790, new_AGEMA_signal_2789, new_AGEMA_signal_2788, Midori_add_Result_Start[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U8 ( .a ({new_AGEMA_signal_1968, new_AGEMA_signal_1967, new_AGEMA_signal_1966, wk[16]}), .b ({DataIn_s3[16], DataIn_s2[16], DataIn_s1[16], DataIn_s0[16]}), .c ({new_AGEMA_signal_2796, new_AGEMA_signal_2795, new_AGEMA_signal_2794, Midori_add_Result_Start[16]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U7 ( .a ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, new_AGEMA_signal_1975, wk[15]}), .b ({DataIn_s3[15], DataIn_s2[15], DataIn_s1[15], DataIn_s0[15]}), .c ({new_AGEMA_signal_2802, new_AGEMA_signal_2801, new_AGEMA_signal_2800, Midori_add_Result_Start[15]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U6 ( .a ({new_AGEMA_signal_1986, new_AGEMA_signal_1985, new_AGEMA_signal_1984, wk[14]}), .b ({DataIn_s3[14], DataIn_s2[14], DataIn_s1[14], DataIn_s0[14]}), .c ({new_AGEMA_signal_2808, new_AGEMA_signal_2807, new_AGEMA_signal_2806, Midori_add_Result_Start[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U5 ( .a ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, new_AGEMA_signal_1993, wk[13]}), .b ({DataIn_s3[13], DataIn_s2[13], DataIn_s1[13], DataIn_s0[13]}), .c ({new_AGEMA_signal_2814, new_AGEMA_signal_2813, new_AGEMA_signal_2812, Midori_add_Result_Start[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U4 ( .a ({new_AGEMA_signal_2004, new_AGEMA_signal_2003, new_AGEMA_signal_2002, wk[12]}), .b ({DataIn_s3[12], DataIn_s2[12], DataIn_s1[12], DataIn_s0[12]}), .c ({new_AGEMA_signal_2820, new_AGEMA_signal_2819, new_AGEMA_signal_2818, Midori_add_Result_Start[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U3 ( .a ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, new_AGEMA_signal_2011, wk[11]}), .b ({DataIn_s3[11], DataIn_s2[11], DataIn_s1[11], DataIn_s0[11]}), .c ({new_AGEMA_signal_2826, new_AGEMA_signal_2825, new_AGEMA_signal_2824, Midori_add_Result_Start[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U2 ( .a ({new_AGEMA_signal_2022, new_AGEMA_signal_2021, new_AGEMA_signal_2020, wk[10]}), .b ({DataIn_s3[10], DataIn_s2[10], DataIn_s1[10], DataIn_s0[10]}), .c ({new_AGEMA_signal_2832, new_AGEMA_signal_2831, new_AGEMA_signal_2830, Midori_add_Result_Start[10]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U1 ( .a ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, new_AGEMA_signal_2029, wk[0]}), .b ({DataIn_s3[0], DataIn_s2[0], DataIn_s1[0], DataIn_s0[0]}), .c ({new_AGEMA_signal_2838, new_AGEMA_signal_2837, new_AGEMA_signal_2836, Midori_add_Result_Start[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U78 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, new_AGEMA_signal_2047, Midori_rounds_SelectedKey_8_}), .b ({1'b0, 1'b0, 1'b0, Midori_rounds_round_Constant[2]}), .c ({new_AGEMA_signal_4413, new_AGEMA_signal_4412, new_AGEMA_signal_4411, Midori_rounds_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U71 ( .a ({new_AGEMA_signal_3270, new_AGEMA_signal_3269, new_AGEMA_signal_3268, Midori_rounds_SelectedKey_60_}), .b ({1'b0, 1'b0, 1'b0, Midori_rounds_round_Constant[15]}), .c ({new_AGEMA_signal_4578, new_AGEMA_signal_4577, new_AGEMA_signal_4576, Midori_rounds_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U65 ( .a ({new_AGEMA_signal_3258, new_AGEMA_signal_3257, new_AGEMA_signal_3256, Midori_rounds_SelectedKey_56_}), .b ({1'b0, 1'b0, 1'b0, Midori_rounds_round_Constant[14]}), .c ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, new_AGEMA_signal_4579, Midori_rounds_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U60 ( .a ({new_AGEMA_signal_3246, new_AGEMA_signal_3245, new_AGEMA_signal_3244, Midori_rounds_SelectedKey_52_}), .b ({1'b0, 1'b0, 1'b0, Midori_rounds_round_Constant[13]}), .c ({new_AGEMA_signal_4584, new_AGEMA_signal_4583, new_AGEMA_signal_4582, Midori_rounds_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U56 ( .a ({new_AGEMA_signal_2046, new_AGEMA_signal_2045, new_AGEMA_signal_2044, Midori_rounds_SelectedKey_4_}), .b ({1'b0, 1'b0, 1'b0, Midori_rounds_round_Constant[1]}), .c ({new_AGEMA_signal_4587, new_AGEMA_signal_4586, new_AGEMA_signal_4585, Midori_rounds_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U53 ( .a ({new_AGEMA_signal_3234, new_AGEMA_signal_3233, new_AGEMA_signal_3232, Midori_rounds_SelectedKey_48_}), .b ({1'b0, 1'b0, 1'b0, Midori_rounds_round_Constant[12]}), .c ({new_AGEMA_signal_4944, new_AGEMA_signal_4943, new_AGEMA_signal_4942, Midori_rounds_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U48 ( .a ({new_AGEMA_signal_3222, new_AGEMA_signal_3221, new_AGEMA_signal_3220, Midori_rounds_SelectedKey_44_}), .b ({1'b0, 1'b0, 1'b0, Midori_rounds_round_Constant[11]}), .c ({new_AGEMA_signal_4470, new_AGEMA_signal_4469, new_AGEMA_signal_4468, Midori_rounds_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U43 ( .a ({new_AGEMA_signal_3210, new_AGEMA_signal_3209, new_AGEMA_signal_3208, Midori_rounds_SelectedKey_40_}), .b ({1'b0, 1'b0, 1'b0, Midori_rounds_round_Constant[10]}), .c ({new_AGEMA_signal_4590, new_AGEMA_signal_4589, new_AGEMA_signal_4588, Midori_rounds_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U37 ( .a ({new_AGEMA_signal_3198, new_AGEMA_signal_3197, new_AGEMA_signal_3196, Midori_rounds_SelectedKey_36_}), .b ({1'b0, 1'b0, 1'b0, Midori_rounds_round_Constant[9]}), .c ({new_AGEMA_signal_4494, new_AGEMA_signal_4493, new_AGEMA_signal_4492, Midori_rounds_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U32 ( .a ({new_AGEMA_signal_3186, new_AGEMA_signal_3185, new_AGEMA_signal_3184, Midori_rounds_SelectedKey_32_}), .b ({1'b0, 1'b0, 1'b0, Midori_rounds_round_Constant[8]}), .c ({new_AGEMA_signal_4593, new_AGEMA_signal_4592, new_AGEMA_signal_4591, Midori_rounds_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U26 ( .a ({new_AGEMA_signal_3174, new_AGEMA_signal_3173, new_AGEMA_signal_3172, Midori_rounds_SelectedKey_28_}), .b ({1'b0, 1'b0, 1'b0, Midori_rounds_round_Constant[7]}), .c ({new_AGEMA_signal_4782, new_AGEMA_signal_4781, new_AGEMA_signal_4780, Midori_rounds_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U21 ( .a ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, new_AGEMA_signal_3163, Midori_rounds_SelectedKey_24_}), .b ({1'b0, 1'b0, 1'b0, Midori_rounds_round_Constant[6]}), .c ({new_AGEMA_signal_4596, new_AGEMA_signal_4595, new_AGEMA_signal_4594, Midori_rounds_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U16 ( .a ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, new_AGEMA_signal_3151, Midori_rounds_SelectedKey_20_}), .b ({1'b0, 1'b0, 1'b0, Midori_rounds_round_Constant[5]}), .c ({new_AGEMA_signal_4536, new_AGEMA_signal_4535, new_AGEMA_signal_4534, Midori_rounds_n4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U10 ( .a ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, new_AGEMA_signal_3139, Midori_rounds_SelectedKey_16_}), .b ({1'b0, 1'b0, 1'b0, Midori_rounds_round_Constant[4]}), .c ({new_AGEMA_signal_4599, new_AGEMA_signal_4598, new_AGEMA_signal_4597, Midori_rounds_n3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U5 ( .a ({new_AGEMA_signal_3138, new_AGEMA_signal_3137, new_AGEMA_signal_3136, Midori_rounds_SelectedKey_12_}), .b ({1'b0, 1'b0, 1'b0, Midori_rounds_round_Constant[3]}), .c ({new_AGEMA_signal_4602, new_AGEMA_signal_4601, new_AGEMA_signal_4600, Midori_rounds_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U1 ( .a ({new_AGEMA_signal_2034, new_AGEMA_signal_2033, new_AGEMA_signal_2032, Midori_rounds_SelectedKey_0_}), .b ({1'b0, 1'b0, 1'b0, Midori_rounds_round_Constant[0]}), .c ({new_AGEMA_signal_4605, new_AGEMA_signal_4604, new_AGEMA_signal_4603, Midori_rounds_n1}) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U106 ( .A1 (Midori_rounds_constant_MUX_n217), .A2 (Midori_rounds_constant_MUX_n216), .ZN (Midori_rounds_round_Constant[9]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U105 ( .A1 (Midori_rounds_constant_MUX_n215), .A2 (Midori_rounds_constant_MUX_n214), .ZN (Midori_rounds_constant_MUX_n217) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U104 ( .A1 (Midori_rounds_constant_MUX_n213), .A2 (Midori_rounds_constant_MUX_n212), .ZN (Midori_rounds_constant_MUX_n214) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U103 ( .A1 (Midori_rounds_constant_MUX_n211), .A2 (Midori_rounds_constant_MUX_n210), .ZN (Midori_rounds_round_Constant[8]) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U102 ( .A1 (Midori_rounds_constant_MUX_n209), .A2 (Midori_rounds_constant_MUX_n208), .ZN (Midori_rounds_round_Constant[7]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U101 ( .A1 (Midori_rounds_round_Constant[11]), .A2 (Midori_rounds_constant_MUX_n207), .ZN (Midori_rounds_constant_MUX_n208) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U100 ( .A1 (Midori_rounds_constant_MUX_n206), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n207) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U99 ( .A1 (Midori_rounds_constant_MUX_n204), .A2 (Midori_rounds_constant_MUX_n203), .ZN (Midori_rounds_constant_MUX_n206) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U98 ( .A1 (Midori_rounds_constant_MUX_n202), .A2 (Midori_rounds_constant_MUX_n201), .ZN (Midori_rounds_round_Constant[6]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U97 ( .A1 (Midori_rounds_constant_MUX_n200), .A2 (Midori_rounds_constant_MUX_n199), .ZN (Midori_rounds_constant_MUX_n201) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U96 ( .A1 (Midori_rounds_constant_MUX_n198), .A2 (Midori_rounds_constant_MUX_n197), .ZN (Midori_rounds_round_Constant[5]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U95 ( .A1 (Midori_rounds_constant_MUX_n212), .A2 (Midori_rounds_constant_MUX_n196), .ZN (Midori_rounds_constant_MUX_n197) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U94 ( .A1 (Midori_rounds_constant_MUX_n195), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n196) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U93 ( .A1 (Midori_rounds_constant_MUX_n194), .A2 (Midori_rounds_constant_MUX_n195), .ZN (Midori_rounds_round_Constant[4]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U92 ( .A1 (Midori_rounds_constant_MUX_n193), .A2 (Midori_rounds_constant_MUX_n192), .ZN (Midori_rounds_constant_MUX_n195) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U91 ( .A1 (Midori_rounds_constant_MUX_n191), .A2 (Midori_rounds_constant_MUX_n190), .ZN (Midori_rounds_round_Constant[3]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U90 ( .A1 (Midori_rounds_constant_MUX_n215), .A2 (Midori_rounds_constant_MUX_n189), .ZN (Midori_rounds_constant_MUX_n191) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U89 ( .A1 (Midori_rounds_constant_MUX_n188), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n189) ) ;
    INV_X1 Midori_rounds_constant_MUX_U88 ( .A (Midori_rounds_constant_MUX_n187), .ZN (Midori_rounds_constant_MUX_n188) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U87 ( .A1 (Midori_rounds_constant_MUX_n215), .A2 (Midori_rounds_constant_MUX_n186), .ZN (Midori_rounds_round_Constant[2]) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U86 ( .A1 (Midori_rounds_constant_MUX_n202), .A2 (Midori_rounds_constant_MUX_n185), .ZN (Midori_rounds_constant_MUX_n186) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U85 ( .A1 (Midori_rounds_constant_MUX_n184), .A2 (Midori_rounds_constant_MUX_n212), .ZN (Midori_rounds_constant_MUX_n202) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U84 ( .A1 (Midori_rounds_constant_MUX_n183), .A2 (Midori_rounds_constant_MUX_n210), .ZN (Midori_rounds_constant_MUX_n215) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U83 ( .A1 (Midori_rounds_constant_MUX_n182), .A2 (Midori_rounds_constant_MUX_n181), .ZN (Midori_rounds_round_Constant[1]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U82 ( .A1 (Midori_rounds_constant_MUX_n187), .A2 (Midori_rounds_constant_MUX_n180), .ZN (Midori_rounds_constant_MUX_n181) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U81 ( .A1 (Midori_rounds_constant_MUX_n212), .A2 (Midori_rounds_constant_MUX_n204), .ZN (Midori_rounds_constant_MUX_n180) ) ;
    INV_X1 Midori_rounds_constant_MUX_U80 ( .A (Midori_rounds_constant_MUX_n183), .ZN (Midori_rounds_constant_MUX_n204) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U79 ( .A1 (Midori_rounds_constant_MUX_n179), .A2 (Midori_rounds_constant_MUX_n178), .ZN (Midori_rounds_constant_MUX_n183) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U78 ( .A1 (Midori_rounds_constant_MUX_n177), .A2 (Midori_rounds_constant_MUX_n176), .ZN (Midori_rounds_constant_MUX_n178) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U77 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n175), .ZN (Midori_rounds_constant_MUX_n212) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U76 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n174), .B (Midori_rounds_constant_MUX_n173), .Z (Midori_rounds_constant_MUX_n175) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U75 ( .A1 (Midori_rounds_constant_MUX_n172), .A2 (Midori_rounds_constant_MUX_n171), .ZN (Midori_rounds_round_Constant[15]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U74 ( .A1 (Midori_rounds_constant_MUX_n200), .A2 (Midori_rounds_constant_MUX_n187), .ZN (Midori_rounds_constant_MUX_n172) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U73 ( .A1 (Midori_rounds_constant_MUX_n170), .A2 (Midori_rounds_constant_MUX_n194), .ZN (Midori_rounds_round_Constant[14]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U72 ( .A1 (Midori_rounds_constant_MUX_n169), .A2 (Midori_rounds_constant_MUX_n168), .ZN (Midori_rounds_constant_MUX_n194) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U71 ( .A1 (Midori_rounds_constant_MUX_n216), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n168) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U70 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n167), .ZN (Midori_rounds_constant_MUX_n205) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U69 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n166), .B (Midori_rounds_constant_MUX_n165), .Z (Midori_rounds_constant_MUX_n167) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U68 ( .A1 (Midori_rounds_constant_MUX_n185), .A2 (Midori_rounds_constant_MUX_n164), .ZN (Midori_rounds_round_Constant[13]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U67 ( .A1 (Midori_rounds_constant_MUX_n163), .A2 (Midori_rounds_constant_MUX_n162), .ZN (Midori_rounds_constant_MUX_n164) ) ;
    INV_X1 Midori_rounds_constant_MUX_U66 ( .A (Midori_rounds_constant_MUX_n170), .ZN (Midori_rounds_constant_MUX_n162) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U65 ( .A1 (Midori_rounds_constant_MUX_n161), .A2 (Midori_rounds_constant_MUX_n192), .ZN (Midori_rounds_constant_MUX_n185) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U64 ( .A1 (Midori_rounds_constant_MUX_n160), .A2 (Midori_rounds_constant_MUX_n190), .ZN (Midori_rounds_round_Constant[12]) ) ;
    INV_X1 Midori_rounds_constant_MUX_U63 ( .A (Midori_rounds_constant_MUX_n184), .ZN (Midori_rounds_constant_MUX_n190) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U62 ( .A1 (Midori_rounds_constant_MUX_n203), .A2 (Midori_rounds_constant_MUX_n159), .ZN (Midori_rounds_constant_MUX_n160) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U61 ( .A1 (Midori_rounds_constant_MUX_n211), .A2 (Midori_rounds_constant_MUX_n170), .ZN (Midori_rounds_constant_MUX_n159) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U60 ( .A1 (Midori_rounds_constant_MUX_n193), .A2 (Midori_rounds_constant_MUX_n169), .ZN (Midori_rounds_constant_MUX_n211) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U59 ( .A1 (Midori_rounds_constant_MUX_n198), .A2 (Midori_rounds_constant_MUX_n158), .ZN (Midori_rounds_constant_MUX_n169) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U58 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n157), .ZN (Midori_rounds_constant_MUX_n158) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U57 ( .A1 (Midori_rounds_constant_MUX_n165), .A2 (Midori_rounds_constant_MUX_n177), .ZN (Midori_rounds_constant_MUX_n157) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U56 ( .A1 (Midori_rounds_constant_MUX_n200), .A2 (Midori_rounds_constant_MUX_n156), .ZN (Midori_rounds_constant_MUX_n198) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U55 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n155), .ZN (Midori_rounds_constant_MUX_n156) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U54 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n176), .B (Midori_rounds_constant_MUX_n166), .Z (Midori_rounds_constant_MUX_n155) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U53 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n154), .ZN (Midori_rounds_constant_MUX_n200) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U52 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n174), .B (Midori_rounds_constant_MUX_n153), .Z (Midori_rounds_constant_MUX_n154) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U51 ( .A1 (Midori_rounds_constant_MUX_n199), .A2 (Midori_rounds_constant_MUX_n213), .ZN (Midori_rounds_round_Constant[11]) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U50 ( .A1 (Midori_rounds_constant_MUX_n170), .A2 (Midori_rounds_constant_MUX_n210), .ZN (Midori_rounds_constant_MUX_n199) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U49 ( .A1 (Midori_rounds_constant_MUX_n152), .A2 (Midori_rounds_constant_MUX_n151), .ZN (Midori_rounds_constant_MUX_n210) ) ;
    AND2_X1 Midori_rounds_constant_MUX_U48 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (round_Signal[2]), .ZN (Midori_rounds_constant_MUX_n151) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U47 ( .A1 (Midori_rounds_constant_MUX_n150), .A2 (Midori_rounds_constant_MUX_n187), .ZN (Midori_rounds_constant_MUX_n170) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U46 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n149), .ZN (Midori_rounds_constant_MUX_n187) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U45 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n165), .B (Midori_rounds_constant_MUX_n166), .Z (Midori_rounds_constant_MUX_n149) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U44 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n148), .ZN (Midori_rounds_constant_MUX_n150) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U43 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n153), .B (Midori_rounds_constant_MUX_n174), .Z (Midori_rounds_constant_MUX_n148) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U42 ( .A1 (Midori_rounds_constant_MUX_n147), .A2 (Midori_rounds_constant_MUX_n171), .ZN (Midori_rounds_round_Constant[10]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U41 ( .A1 (Midori_rounds_constant_MUX_n146), .A2 (Midori_rounds_constant_MUX_n213), .ZN (Midori_rounds_constant_MUX_n171) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U40 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n145), .ZN (Midori_rounds_constant_MUX_n213) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U39 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n165), .B (Midori_rounds_constant_MUX_n177), .Z (Midori_rounds_constant_MUX_n145) ) ;
    INV_X1 Midori_rounds_constant_MUX_U38 ( .A (Midori_rounds_constant_MUX_n144), .ZN (Midori_rounds_constant_MUX_n146) ) ;
    INV_X1 Midori_rounds_constant_MUX_U37 ( .A (Midori_rounds_constant_MUX_n193), .ZN (Midori_rounds_constant_MUX_n147) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U36 ( .A1 (Midori_rounds_constant_MUX_n182), .A2 (Midori_rounds_constant_MUX_n144), .ZN (Midori_rounds_round_Constant[0]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U35 ( .A1 (Midori_rounds_constant_MUX_n203), .A2 (Midori_rounds_constant_MUX_n192), .ZN (Midori_rounds_constant_MUX_n144) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U34 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n143), .ZN (Midori_rounds_constant_MUX_n192) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U33 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n173), .B (Midori_rounds_constant_MUX_n174), .Z (Midori_rounds_constant_MUX_n143) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U32 ( .A1 (Midori_rounds_constant_MUX_n142), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n174) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U31 ( .A1 (Midori_rounds_constant_MUX_n140), .A2 (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n173) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U30 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n139), .ZN (Midori_rounds_constant_MUX_n203) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U29 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n166), .B (Midori_rounds_constant_MUX_n176), .Z (Midori_rounds_constant_MUX_n139) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U28 ( .A1 (enc_dec), .A2 (Midori_rounds_constant_MUX_n152), .ZN (Midori_rounds_constant_MUX_n176) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U27 ( .A1 (round_Signal[3]), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n152) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U26 ( .A1 (Midori_rounds_constant_MUX_n138), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n166) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U25 ( .A1 (Midori_rounds_constant_MUX_n184), .A2 (Midori_rounds_constant_MUX_n137), .ZN (Midori_rounds_constant_MUX_n182) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U24 ( .A1 (Midori_rounds_constant_MUX_n209), .A2 (Midori_rounds_constant_MUX_n216), .ZN (Midori_rounds_constant_MUX_n137) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U23 ( .A1 (Midori_rounds_constant_MUX_n163), .A2 (Midori_rounds_constant_MUX_n136), .ZN (Midori_rounds_constant_MUX_n216) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U22 ( .A1 (Midori_rounds_constant_MUX_n140), .A2 (Midori_rounds_constant_MUX_n142), .ZN (Midori_rounds_constant_MUX_n136) ) ;
    AND2_X1 Midori_rounds_constant_MUX_U21 ( .A1 (round_Signal[1]), .A2 (Midori_rounds_constant_MUX_n179), .ZN (Midori_rounds_constant_MUX_n163) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U20 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (round_Signal[2]), .ZN (Midori_rounds_constant_MUX_n179) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U19 ( .A1 (Midori_rounds_constant_MUX_n193), .A2 (Midori_rounds_constant_MUX_n161), .ZN (Midori_rounds_constant_MUX_n209) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U18 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n135), .ZN (Midori_rounds_constant_MUX_n161) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U17 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n177), .B (Midori_rounds_constant_MUX_n165), .Z (Midori_rounds_constant_MUX_n135) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U16 ( .A1 (enc_dec), .A2 (Midori_rounds_constant_MUX_n134), .ZN (Midori_rounds_constant_MUX_n165) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U15 ( .A1 (round_Signal[3]), .A2 (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n134) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U14 ( .A1 (round_Signal[1]), .A2 (Midori_rounds_constant_MUX_n138), .ZN (Midori_rounds_constant_MUX_n177) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U13 ( .A1 (enc_dec), .A2 (Midori_rounds_constant_MUX_n133), .ZN (Midori_rounds_constant_MUX_n138) ) ;
    INV_X1 Midori_rounds_constant_MUX_U12 ( .A (round_Signal[3]), .ZN (Midori_rounds_constant_MUX_n133) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U11 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n132), .ZN (Midori_rounds_constant_MUX_n193) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U10 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n153), .B (Midori_rounds_constant_MUX_n131), .Z (Midori_rounds_constant_MUX_n132) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U9 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n130), .ZN (Midori_rounds_constant_MUX_n184) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U8 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n131), .B (Midori_rounds_constant_MUX_n153), .Z (Midori_rounds_constant_MUX_n130) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U7 ( .A1 (Midori_rounds_constant_MUX_n140), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n153) ) ;
    INV_X1 Midori_rounds_constant_MUX_U6 ( .A (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n141) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U5 ( .A1 (enc_dec), .A2 (round_Signal[3]), .ZN (Midori_rounds_constant_MUX_n140) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U4 ( .A1 (Midori_rounds_constant_MUX_n142), .A2 (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n131) ) ;
    AND2_X1 Midori_rounds_constant_MUX_U3 ( .A1 (enc_dec), .A2 (round_Signal[3]), .ZN (Midori_rounds_constant_MUX_n142) ) ;
    INV_X1 Midori_rounds_constant_MUX_U2 ( .A (Midori_rounds_constant_MUX_n129), .ZN (Midori_rounds_constant_MUX_n128) ) ;
    INV_X1 Midori_rounds_constant_MUX_U1 ( .A (round_Signal[0]), .ZN (Midori_rounds_constant_MUX_n129) ) ;
    INV_X1 Midori_rounds_MUXInst_U4 ( .A (round_Signal[0]), .ZN (Midori_rounds_MUXInst_n11) ) ;
    INV_X1 Midori_rounds_MUXInst_U3 ( .A (Midori_rounds_MUXInst_n11), .ZN (Midori_rounds_MUXInst_n8) ) ;
    INV_X1 Midori_rounds_MUXInst_U2 ( .A (Midori_rounds_MUXInst_n11), .ZN (Midori_rounds_MUXInst_n9) ) ;
    INV_X1 Midori_rounds_MUXInst_U1 ( .A (Midori_rounds_MUXInst_n11), .ZN (Midori_rounds_MUXInst_n10) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_0_U1 ( .s (round_Signal[0]), .b ({key_s3[64], key_s2[64], key_s1[64], key_s0[64]}), .a ({key_s3[0], key_s2[0], key_s1[0], key_s0[0]}), .c ({new_AGEMA_signal_2034, new_AGEMA_signal_2033, new_AGEMA_signal_2032, Midori_rounds_SelectedKey_0_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_1_U1 ( .s (round_Signal[0]), .b ({key_s3[65], key_s2[65], key_s1[65], key_s0[65]}), .a ({key_s3[1], key_s2[1], key_s1[1], key_s0[1]}), .c ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, new_AGEMA_signal_2035, Midori_rounds_SelectedKey_1_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_2_U1 ( .s (round_Signal[0]), .b ({key_s3[66], key_s2[66], key_s1[66], key_s0[66]}), .a ({key_s3[2], key_s2[2], key_s1[2], key_s0[2]}), .c ({new_AGEMA_signal_2040, new_AGEMA_signal_2039, new_AGEMA_signal_2038, Midori_rounds_SelectedKey_2_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_3_U1 ( .s (round_Signal[0]), .b ({key_s3[67], key_s2[67], key_s1[67], key_s0[67]}), .a ({key_s3[3], key_s2[3], key_s1[3], key_s0[3]}), .c ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, new_AGEMA_signal_2041, Midori_rounds_SelectedKey_3_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_4_U1 ( .s (round_Signal[0]), .b ({key_s3[68], key_s2[68], key_s1[68], key_s0[68]}), .a ({key_s3[4], key_s2[4], key_s1[4], key_s0[4]}), .c ({new_AGEMA_signal_2046, new_AGEMA_signal_2045, new_AGEMA_signal_2044, Midori_rounds_SelectedKey_4_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_5_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s3[69], key_s2[69], key_s1[69], key_s0[69]}), .a ({key_s3[5], key_s2[5], key_s1[5], key_s0[5]}), .c ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, new_AGEMA_signal_3127, Midori_rounds_SelectedKey_5_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_6_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[70], key_s2[70], key_s1[70], key_s0[70]}), .a ({key_s3[6], key_s2[6], key_s1[6], key_s0[6]}), .c ({new_AGEMA_signal_3132, new_AGEMA_signal_3131, new_AGEMA_signal_3130, Midori_rounds_SelectedKey_6_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_7_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s3[71], key_s2[71], key_s1[71], key_s0[71]}), .a ({key_s3[7], key_s2[7], key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, new_AGEMA_signal_3133, Midori_rounds_SelectedKey_7_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_8_U1 ( .s (round_Signal[0]), .b ({key_s3[72], key_s2[72], key_s1[72], key_s0[72]}), .a ({key_s3[8], key_s2[8], key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, new_AGEMA_signal_2047, Midori_rounds_SelectedKey_8_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_9_U1 ( .s (round_Signal[0]), .b ({key_s3[73], key_s2[73], key_s1[73], key_s0[73]}), .a ({key_s3[9], key_s2[9], key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_2052, new_AGEMA_signal_2051, new_AGEMA_signal_2050, Midori_rounds_SelectedKey_9_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_10_U1 ( .s (round_Signal[0]), .b ({key_s3[74], key_s2[74], key_s1[74], key_s0[74]}), .a ({key_s3[10], key_s2[10], key_s1[10], key_s0[10]}), .c ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, new_AGEMA_signal_2053, Midori_rounds_SelectedKey_10_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_11_U1 ( .s (round_Signal[0]), .b ({key_s3[75], key_s2[75], key_s1[75], key_s0[75]}), .a ({key_s3[11], key_s2[11], key_s1[11], key_s0[11]}), .c ({new_AGEMA_signal_2058, new_AGEMA_signal_2057, new_AGEMA_signal_2056, Midori_rounds_SelectedKey_11_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_12_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s3[76], key_s2[76], key_s1[76], key_s0[76]}), .a ({key_s3[12], key_s2[12], key_s1[12], key_s0[12]}), .c ({new_AGEMA_signal_3138, new_AGEMA_signal_3137, new_AGEMA_signal_3136, Midori_rounds_SelectedKey_12_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_13_U1 ( .s (round_Signal[0]), .b ({key_s3[77], key_s2[77], key_s1[77], key_s0[77]}), .a ({key_s3[13], key_s2[13], key_s1[13], key_s0[13]}), .c ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, new_AGEMA_signal_2059, Midori_rounds_SelectedKey_13_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_14_U1 ( .s (round_Signal[0]), .b ({key_s3[78], key_s2[78], key_s1[78], key_s0[78]}), .a ({key_s3[14], key_s2[14], key_s1[14], key_s0[14]}), .c ({new_AGEMA_signal_2064, new_AGEMA_signal_2063, new_AGEMA_signal_2062, Midori_rounds_SelectedKey_14_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_15_U1 ( .s (round_Signal[0]), .b ({key_s3[79], key_s2[79], key_s1[79], key_s0[79]}), .a ({key_s3[15], key_s2[15], key_s1[15], key_s0[15]}), .c ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, new_AGEMA_signal_2065, Midori_rounds_SelectedKey_15_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_16_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[80], key_s2[80], key_s1[80], key_s0[80]}), .a ({key_s3[16], key_s2[16], key_s1[16], key_s0[16]}), .c ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, new_AGEMA_signal_3139, Midori_rounds_SelectedKey_16_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_17_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s3[81], key_s2[81], key_s1[81], key_s0[81]}), .a ({key_s3[17], key_s2[17], key_s1[17], key_s0[17]}), .c ({new_AGEMA_signal_3144, new_AGEMA_signal_3143, new_AGEMA_signal_3142, Midori_rounds_SelectedKey_17_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_18_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[82], key_s2[82], key_s1[82], key_s0[82]}), .a ({key_s3[18], key_s2[18], key_s1[18], key_s0[18]}), .c ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, new_AGEMA_signal_3145, Midori_rounds_SelectedKey_18_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_19_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[83], key_s2[83], key_s1[83], key_s0[83]}), .a ({key_s3[19], key_s2[19], key_s1[19], key_s0[19]}), .c ({new_AGEMA_signal_3150, new_AGEMA_signal_3149, new_AGEMA_signal_3148, Midori_rounds_SelectedKey_19_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_20_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[84], key_s2[84], key_s1[84], key_s0[84]}), .a ({key_s3[20], key_s2[20], key_s1[20], key_s0[20]}), .c ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, new_AGEMA_signal_3151, Midori_rounds_SelectedKey_20_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_21_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[85], key_s2[85], key_s1[85], key_s0[85]}), .a ({key_s3[21], key_s2[21], key_s1[21], key_s0[21]}), .c ({new_AGEMA_signal_3156, new_AGEMA_signal_3155, new_AGEMA_signal_3154, Midori_rounds_SelectedKey_21_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_22_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s3[86], key_s2[86], key_s1[86], key_s0[86]}), .a ({key_s3[22], key_s2[22], key_s1[22], key_s0[22]}), .c ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, new_AGEMA_signal_3157, Midori_rounds_SelectedKey_22_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_23_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s3[87], key_s2[87], key_s1[87], key_s0[87]}), .a ({key_s3[23], key_s2[23], key_s1[23], key_s0[23]}), .c ({new_AGEMA_signal_3162, new_AGEMA_signal_3161, new_AGEMA_signal_3160, Midori_rounds_SelectedKey_23_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_24_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[88], key_s2[88], key_s1[88], key_s0[88]}), .a ({key_s3[24], key_s2[24], key_s1[24], key_s0[24]}), .c ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, new_AGEMA_signal_3163, Midori_rounds_SelectedKey_24_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_25_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s3[89], key_s2[89], key_s1[89], key_s0[89]}), .a ({key_s3[25], key_s2[25], key_s1[25], key_s0[25]}), .c ({new_AGEMA_signal_3168, new_AGEMA_signal_3167, new_AGEMA_signal_3166, Midori_rounds_SelectedKey_25_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_26_U1 ( .s (round_Signal[0]), .b ({key_s3[90], key_s2[90], key_s1[90], key_s0[90]}), .a ({key_s3[26], key_s2[26], key_s1[26], key_s0[26]}), .c ({new_AGEMA_signal_2070, new_AGEMA_signal_2069, new_AGEMA_signal_2068, Midori_rounds_SelectedKey_26_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_27_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[91], key_s2[91], key_s1[91], key_s0[91]}), .a ({key_s3[27], key_s2[27], key_s1[27], key_s0[27]}), .c ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, new_AGEMA_signal_3169, Midori_rounds_SelectedKey_27_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_28_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[92], key_s2[92], key_s1[92], key_s0[92]}), .a ({key_s3[28], key_s2[28], key_s1[28], key_s0[28]}), .c ({new_AGEMA_signal_3174, new_AGEMA_signal_3173, new_AGEMA_signal_3172, Midori_rounds_SelectedKey_28_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_29_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[93], key_s2[93], key_s1[93], key_s0[93]}), .a ({key_s3[29], key_s2[29], key_s1[29], key_s0[29]}), .c ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, new_AGEMA_signal_3175, Midori_rounds_SelectedKey_29_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_30_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[94], key_s2[94], key_s1[94], key_s0[94]}), .a ({key_s3[30], key_s2[30], key_s1[30], key_s0[30]}), .c ({new_AGEMA_signal_3180, new_AGEMA_signal_3179, new_AGEMA_signal_3178, Midori_rounds_SelectedKey_30_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_31_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[95], key_s2[95], key_s1[95], key_s0[95]}), .a ({key_s3[31], key_s2[31], key_s1[31], key_s0[31]}), .c ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, new_AGEMA_signal_3181, Midori_rounds_SelectedKey_31_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_32_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[96], key_s2[96], key_s1[96], key_s0[96]}), .a ({key_s3[32], key_s2[32], key_s1[32], key_s0[32]}), .c ({new_AGEMA_signal_3186, new_AGEMA_signal_3185, new_AGEMA_signal_3184, Midori_rounds_SelectedKey_32_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_33_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[97], key_s2[97], key_s1[97], key_s0[97]}), .a ({key_s3[33], key_s2[33], key_s1[33], key_s0[33]}), .c ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, new_AGEMA_signal_3187, Midori_rounds_SelectedKey_33_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_34_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[98], key_s2[98], key_s1[98], key_s0[98]}), .a ({key_s3[34], key_s2[34], key_s1[34], key_s0[34]}), .c ({new_AGEMA_signal_3192, new_AGEMA_signal_3191, new_AGEMA_signal_3190, Midori_rounds_SelectedKey_34_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_35_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[99], key_s2[99], key_s1[99], key_s0[99]}), .a ({key_s3[35], key_s2[35], key_s1[35], key_s0[35]}), .c ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, new_AGEMA_signal_3193, Midori_rounds_SelectedKey_35_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_36_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[100], key_s2[100], key_s1[100], key_s0[100]}), .a ({key_s3[36], key_s2[36], key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_3198, new_AGEMA_signal_3197, new_AGEMA_signal_3196, Midori_rounds_SelectedKey_36_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_37_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[101], key_s2[101], key_s1[101], key_s0[101]}), .a ({key_s3[37], key_s2[37], key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, new_AGEMA_signal_3199, Midori_rounds_SelectedKey_37_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_38_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[102], key_s2[102], key_s1[102], key_s0[102]}), .a ({key_s3[38], key_s2[38], key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_3204, new_AGEMA_signal_3203, new_AGEMA_signal_3202, Midori_rounds_SelectedKey_38_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_39_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s3[103], key_s2[103], key_s1[103], key_s0[103]}), .a ({key_s3[39], key_s2[39], key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, new_AGEMA_signal_3205, Midori_rounds_SelectedKey_39_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_40_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s3[104], key_s2[104], key_s1[104], key_s0[104]}), .a ({key_s3[40], key_s2[40], key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_3210, new_AGEMA_signal_3209, new_AGEMA_signal_3208, Midori_rounds_SelectedKey_40_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_41_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s3[105], key_s2[105], key_s1[105], key_s0[105]}), .a ({key_s3[41], key_s2[41], key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, new_AGEMA_signal_3211, Midori_rounds_SelectedKey_41_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_42_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s3[106], key_s2[106], key_s1[106], key_s0[106]}), .a ({key_s3[42], key_s2[42], key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_3216, new_AGEMA_signal_3215, new_AGEMA_signal_3214, Midori_rounds_SelectedKey_42_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_43_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s3[107], key_s2[107], key_s1[107], key_s0[107]}), .a ({key_s3[43], key_s2[43], key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, new_AGEMA_signal_3217, Midori_rounds_SelectedKey_43_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_44_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s3[108], key_s2[108], key_s1[108], key_s0[108]}), .a ({key_s3[44], key_s2[44], key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_3222, new_AGEMA_signal_3221, new_AGEMA_signal_3220, Midori_rounds_SelectedKey_44_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_45_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s3[109], key_s2[109], key_s1[109], key_s0[109]}), .a ({key_s3[45], key_s2[45], key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, new_AGEMA_signal_3223, Midori_rounds_SelectedKey_45_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_46_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s3[110], key_s2[110], key_s1[110], key_s0[110]}), .a ({key_s3[46], key_s2[46], key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_3228, new_AGEMA_signal_3227, new_AGEMA_signal_3226, Midori_rounds_SelectedKey_46_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_47_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s3[111], key_s2[111], key_s1[111], key_s0[111]}), .a ({key_s3[47], key_s2[47], key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, new_AGEMA_signal_3229, Midori_rounds_SelectedKey_47_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_48_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s3[112], key_s2[112], key_s1[112], key_s0[112]}), .a ({key_s3[48], key_s2[48], key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_3234, new_AGEMA_signal_3233, new_AGEMA_signal_3232, Midori_rounds_SelectedKey_48_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_49_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s3[113], key_s2[113], key_s1[113], key_s0[113]}), .a ({key_s3[49], key_s2[49], key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, new_AGEMA_signal_3235, Midori_rounds_SelectedKey_49_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_50_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s3[114], key_s2[114], key_s1[114], key_s0[114]}), .a ({key_s3[50], key_s2[50], key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_3240, new_AGEMA_signal_3239, new_AGEMA_signal_3238, Midori_rounds_SelectedKey_50_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_51_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s3[115], key_s2[115], key_s1[115], key_s0[115]}), .a ({key_s3[51], key_s2[51], key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, new_AGEMA_signal_3241, Midori_rounds_SelectedKey_51_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_52_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s3[116], key_s2[116], key_s1[116], key_s0[116]}), .a ({key_s3[52], key_s2[52], key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_3246, new_AGEMA_signal_3245, new_AGEMA_signal_3244, Midori_rounds_SelectedKey_52_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_53_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s3[117], key_s2[117], key_s1[117], key_s0[117]}), .a ({key_s3[53], key_s2[53], key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, new_AGEMA_signal_3247, Midori_rounds_SelectedKey_53_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_54_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s3[118], key_s2[118], key_s1[118], key_s0[118]}), .a ({key_s3[54], key_s2[54], key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_3252, new_AGEMA_signal_3251, new_AGEMA_signal_3250, Midori_rounds_SelectedKey_54_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_55_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s3[119], key_s2[119], key_s1[119], key_s0[119]}), .a ({key_s3[55], key_s2[55], key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, new_AGEMA_signal_3253, Midori_rounds_SelectedKey_55_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_56_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s3[120], key_s2[120], key_s1[120], key_s0[120]}), .a ({key_s3[56], key_s2[56], key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_3258, new_AGEMA_signal_3257, new_AGEMA_signal_3256, Midori_rounds_SelectedKey_56_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_57_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s3[121], key_s2[121], key_s1[121], key_s0[121]}), .a ({key_s3[57], key_s2[57], key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, new_AGEMA_signal_3259, Midori_rounds_SelectedKey_57_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_58_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s3[122], key_s2[122], key_s1[122], key_s0[122]}), .a ({key_s3[58], key_s2[58], key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_3264, new_AGEMA_signal_3263, new_AGEMA_signal_3262, Midori_rounds_SelectedKey_58_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_59_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s3[123], key_s2[123], key_s1[123], key_s0[123]}), .a ({key_s3[59], key_s2[59], key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, new_AGEMA_signal_3265, Midori_rounds_SelectedKey_59_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_60_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s3[124], key_s2[124], key_s1[124], key_s0[124]}), .a ({key_s3[60], key_s2[60], key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_3270, new_AGEMA_signal_3269, new_AGEMA_signal_3268, Midori_rounds_SelectedKey_60_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_61_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s3[125], key_s2[125], key_s1[125], key_s0[125]}), .a ({key_s3[61], key_s2[61], key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, new_AGEMA_signal_3271, Midori_rounds_SelectedKey_61_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_62_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s3[126], key_s2[126], key_s1[126], key_s0[126]}), .a ({key_s3[62], key_s2[62], key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_3276, new_AGEMA_signal_3275, new_AGEMA_signal_3274, Midori_rounds_SelectedKey_62_}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_63_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s3[127], key_s2[127], key_s1[127], key_s0[127]}), .a ({key_s3[63], key_s2[63], key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, new_AGEMA_signal_3277, Midori_rounds_SelectedKey_63_}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U4 ( .a ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, new_AGEMA_signal_2071, Midori_rounds_roundReg_out[0]}), .b ({new_AGEMA_signal_2088, new_AGEMA_signal_2087, new_AGEMA_signal_2086, Midori_rounds_sub_sBox_PRINCE_0_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U2 ( .a ({new_AGEMA_signal_2076, new_AGEMA_signal_2075, new_AGEMA_signal_2074, Midori_rounds_roundReg_out[3]}), .b ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, new_AGEMA_signal_2089, Midori_rounds_sub_sBox_PRINCE_0_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U1 ( .a ({new_AGEMA_signal_2082, new_AGEMA_signal_2081, new_AGEMA_signal_2080, Midori_rounds_roundReg_out[2]}), .b ({new_AGEMA_signal_2094, new_AGEMA_signal_2093, new_AGEMA_signal_2092, Midori_rounds_sub_sBox_PRINCE_0_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U4 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, new_AGEMA_signal_2095, Midori_rounds_roundReg_out[4]}), .b ({new_AGEMA_signal_2112, new_AGEMA_signal_2111, new_AGEMA_signal_2110, Midori_rounds_sub_sBox_PRINCE_1_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U2 ( .a ({new_AGEMA_signal_2100, new_AGEMA_signal_2099, new_AGEMA_signal_2098, Midori_rounds_roundReg_out[7]}), .b ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, new_AGEMA_signal_2113, Midori_rounds_sub_sBox_PRINCE_1_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U1 ( .a ({new_AGEMA_signal_2106, new_AGEMA_signal_2105, new_AGEMA_signal_2104, Midori_rounds_roundReg_out[6]}), .b ({new_AGEMA_signal_2118, new_AGEMA_signal_2117, new_AGEMA_signal_2116, Midori_rounds_sub_sBox_PRINCE_1_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U4 ( .a ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, new_AGEMA_signal_2119, Midori_rounds_roundReg_out[8]}), .b ({new_AGEMA_signal_2136, new_AGEMA_signal_2135, new_AGEMA_signal_2134, Midori_rounds_sub_sBox_PRINCE_2_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U2 ( .a ({new_AGEMA_signal_2124, new_AGEMA_signal_2123, new_AGEMA_signal_2122, Midori_rounds_roundReg_out[11]}), .b ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, new_AGEMA_signal_2137, Midori_rounds_sub_sBox_PRINCE_2_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U1 ( .a ({new_AGEMA_signal_2130, new_AGEMA_signal_2129, new_AGEMA_signal_2128, Midori_rounds_roundReg_out[10]}), .b ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, new_AGEMA_signal_2140, Midori_rounds_sub_sBox_PRINCE_2_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U4 ( .a ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, new_AGEMA_signal_2143, Midori_rounds_roundReg_out[12]}), .b ({new_AGEMA_signal_2160, new_AGEMA_signal_2159, new_AGEMA_signal_2158, Midori_rounds_sub_sBox_PRINCE_3_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U2 ( .a ({new_AGEMA_signal_2148, new_AGEMA_signal_2147, new_AGEMA_signal_2146, Midori_rounds_roundReg_out[15]}), .b ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, new_AGEMA_signal_2161, Midori_rounds_sub_sBox_PRINCE_3_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U1 ( .a ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, new_AGEMA_signal_2152, Midori_rounds_roundReg_out[14]}), .b ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, new_AGEMA_signal_2164, Midori_rounds_sub_sBox_PRINCE_3_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U4 ( .a ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, new_AGEMA_signal_2167, Midori_rounds_roundReg_out[16]}), .b ({new_AGEMA_signal_2184, new_AGEMA_signal_2183, new_AGEMA_signal_2182, Midori_rounds_sub_sBox_PRINCE_4_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U2 ( .a ({new_AGEMA_signal_2172, new_AGEMA_signal_2171, new_AGEMA_signal_2170, Midori_rounds_roundReg_out[19]}), .b ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, new_AGEMA_signal_2185, Midori_rounds_sub_sBox_PRINCE_4_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U1 ( .a ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, new_AGEMA_signal_2176, Midori_rounds_roundReg_out[18]}), .b ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, new_AGEMA_signal_2188, Midori_rounds_sub_sBox_PRINCE_4_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U4 ( .a ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, new_AGEMA_signal_2191, Midori_rounds_roundReg_out[20]}), .b ({new_AGEMA_signal_2208, new_AGEMA_signal_2207, new_AGEMA_signal_2206, Midori_rounds_sub_sBox_PRINCE_5_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U2 ( .a ({new_AGEMA_signal_2196, new_AGEMA_signal_2195, new_AGEMA_signal_2194, Midori_rounds_roundReg_out[23]}), .b ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, new_AGEMA_signal_2209, Midori_rounds_sub_sBox_PRINCE_5_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U1 ( .a ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, new_AGEMA_signal_2200, Midori_rounds_roundReg_out[22]}), .b ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, new_AGEMA_signal_2212, Midori_rounds_sub_sBox_PRINCE_5_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U4 ( .a ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, new_AGEMA_signal_2215, Midori_rounds_roundReg_out[24]}), .b ({new_AGEMA_signal_2232, new_AGEMA_signal_2231, new_AGEMA_signal_2230, Midori_rounds_sub_sBox_PRINCE_6_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U2 ( .a ({new_AGEMA_signal_2220, new_AGEMA_signal_2219, new_AGEMA_signal_2218, Midori_rounds_roundReg_out[27]}), .b ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, new_AGEMA_signal_2233, Midori_rounds_sub_sBox_PRINCE_6_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U1 ( .a ({new_AGEMA_signal_2226, new_AGEMA_signal_2225, new_AGEMA_signal_2224, Midori_rounds_roundReg_out[26]}), .b ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, new_AGEMA_signal_2236, Midori_rounds_sub_sBox_PRINCE_6_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U4 ( .a ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, new_AGEMA_signal_2239, Midori_rounds_roundReg_out[28]}), .b ({new_AGEMA_signal_2256, new_AGEMA_signal_2255, new_AGEMA_signal_2254, Midori_rounds_sub_sBox_PRINCE_7_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U2 ( .a ({new_AGEMA_signal_2244, new_AGEMA_signal_2243, new_AGEMA_signal_2242, Midori_rounds_roundReg_out[31]}), .b ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, new_AGEMA_signal_2257, Midori_rounds_sub_sBox_PRINCE_7_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U1 ( .a ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, new_AGEMA_signal_2248, Midori_rounds_roundReg_out[30]}), .b ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, new_AGEMA_signal_2260, Midori_rounds_sub_sBox_PRINCE_7_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U4 ( .a ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, new_AGEMA_signal_2263, Midori_rounds_roundReg_out[32]}), .b ({new_AGEMA_signal_2280, new_AGEMA_signal_2279, new_AGEMA_signal_2278, Midori_rounds_sub_sBox_PRINCE_8_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U2 ( .a ({new_AGEMA_signal_2268, new_AGEMA_signal_2267, new_AGEMA_signal_2266, Midori_rounds_roundReg_out[35]}), .b ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, new_AGEMA_signal_2281, Midori_rounds_sub_sBox_PRINCE_8_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U1 ( .a ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, new_AGEMA_signal_2272, Midori_rounds_roundReg_out[34]}), .b ({new_AGEMA_signal_2286, new_AGEMA_signal_2285, new_AGEMA_signal_2284, Midori_rounds_sub_sBox_PRINCE_8_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U4 ( .a ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, new_AGEMA_signal_2287, Midori_rounds_roundReg_out[36]}), .b ({new_AGEMA_signal_2304, new_AGEMA_signal_2303, new_AGEMA_signal_2302, Midori_rounds_sub_sBox_PRINCE_9_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U2 ( .a ({new_AGEMA_signal_2292, new_AGEMA_signal_2291, new_AGEMA_signal_2290, Midori_rounds_roundReg_out[39]}), .b ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, new_AGEMA_signal_2305, Midori_rounds_sub_sBox_PRINCE_9_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U1 ( .a ({new_AGEMA_signal_2298, new_AGEMA_signal_2297, new_AGEMA_signal_2296, Midori_rounds_roundReg_out[38]}), .b ({new_AGEMA_signal_2310, new_AGEMA_signal_2309, new_AGEMA_signal_2308, Midori_rounds_sub_sBox_PRINCE_9_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U4 ( .a ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, new_AGEMA_signal_2311, Midori_rounds_roundReg_out[40]}), .b ({new_AGEMA_signal_2328, new_AGEMA_signal_2327, new_AGEMA_signal_2326, Midori_rounds_sub_sBox_PRINCE_10_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U2 ( .a ({new_AGEMA_signal_2316, new_AGEMA_signal_2315, new_AGEMA_signal_2314, Midori_rounds_roundReg_out[43]}), .b ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, new_AGEMA_signal_2329, Midori_rounds_sub_sBox_PRINCE_10_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U1 ( .a ({new_AGEMA_signal_2322, new_AGEMA_signal_2321, new_AGEMA_signal_2320, Midori_rounds_roundReg_out[42]}), .b ({new_AGEMA_signal_2334, new_AGEMA_signal_2333, new_AGEMA_signal_2332, Midori_rounds_sub_sBox_PRINCE_10_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U4 ( .a ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, new_AGEMA_signal_2335, Midori_rounds_roundReg_out[44]}), .b ({new_AGEMA_signal_2352, new_AGEMA_signal_2351, new_AGEMA_signal_2350, Midori_rounds_sub_sBox_PRINCE_11_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U2 ( .a ({new_AGEMA_signal_2340, new_AGEMA_signal_2339, new_AGEMA_signal_2338, Midori_rounds_roundReg_out[47]}), .b ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, new_AGEMA_signal_2353, Midori_rounds_sub_sBox_PRINCE_11_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U1 ( .a ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, new_AGEMA_signal_2344, Midori_rounds_roundReg_out[46]}), .b ({new_AGEMA_signal_2358, new_AGEMA_signal_2357, new_AGEMA_signal_2356, Midori_rounds_sub_sBox_PRINCE_11_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U4 ( .a ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, new_AGEMA_signal_2359, Midori_rounds_roundReg_out[48]}), .b ({new_AGEMA_signal_2376, new_AGEMA_signal_2375, new_AGEMA_signal_2374, Midori_rounds_sub_sBox_PRINCE_12_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U2 ( .a ({new_AGEMA_signal_2364, new_AGEMA_signal_2363, new_AGEMA_signal_2362, Midori_rounds_roundReg_out[51]}), .b ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, new_AGEMA_signal_2377, Midori_rounds_sub_sBox_PRINCE_12_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U1 ( .a ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, new_AGEMA_signal_2368, Midori_rounds_roundReg_out[50]}), .b ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, new_AGEMA_signal_2380, Midori_rounds_sub_sBox_PRINCE_12_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U4 ( .a ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, new_AGEMA_signal_2383, Midori_rounds_roundReg_out[52]}), .b ({new_AGEMA_signal_2400, new_AGEMA_signal_2399, new_AGEMA_signal_2398, Midori_rounds_sub_sBox_PRINCE_13_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U2 ( .a ({new_AGEMA_signal_2388, new_AGEMA_signal_2387, new_AGEMA_signal_2386, Midori_rounds_roundReg_out[55]}), .b ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, new_AGEMA_signal_2401, Midori_rounds_sub_sBox_PRINCE_13_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U1 ( .a ({new_AGEMA_signal_2394, new_AGEMA_signal_2393, new_AGEMA_signal_2392, Midori_rounds_roundReg_out[54]}), .b ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, new_AGEMA_signal_2404, Midori_rounds_sub_sBox_PRINCE_13_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U4 ( .a ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, new_AGEMA_signal_2407, Midori_rounds_roundReg_out[56]}), .b ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, new_AGEMA_signal_2422, Midori_rounds_sub_sBox_PRINCE_14_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U2 ( .a ({new_AGEMA_signal_2412, new_AGEMA_signal_2411, new_AGEMA_signal_2410, Midori_rounds_roundReg_out[59]}), .b ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, new_AGEMA_signal_2425, Midori_rounds_sub_sBox_PRINCE_14_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U1 ( .a ({new_AGEMA_signal_2418, new_AGEMA_signal_2417, new_AGEMA_signal_2416, Midori_rounds_roundReg_out[58]}), .b ({new_AGEMA_signal_2430, new_AGEMA_signal_2429, new_AGEMA_signal_2428, Midori_rounds_sub_sBox_PRINCE_14_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U4 ( .a ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, new_AGEMA_signal_2431, Midori_rounds_roundReg_out[60]}), .b ({new_AGEMA_signal_2448, new_AGEMA_signal_2447, new_AGEMA_signal_2446, Midori_rounds_sub_sBox_PRINCE_15_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U2 ( .a ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, new_AGEMA_signal_2434, Midori_rounds_roundReg_out[63]}), .b ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, new_AGEMA_signal_2449, Midori_rounds_sub_sBox_PRINCE_15_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U1 ( .a ({new_AGEMA_signal_2442, new_AGEMA_signal_2441, new_AGEMA_signal_2440, Midori_rounds_roundReg_out[62]}), .b ({new_AGEMA_signal_2454, new_AGEMA_signal_2453, new_AGEMA_signal_2452, Midori_rounds_sub_sBox_PRINCE_15_n9}) ) ;
    ClockGatingController #(9) ClockGatingInst ( .clk (clk), .rst (reset), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U14 ( .a ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, new_AGEMA_signal_2071, Midori_rounds_roundReg_out[0]}), .b ({new_AGEMA_signal_2076, new_AGEMA_signal_2075, new_AGEMA_signal_2074, Midori_rounds_roundReg_out[3]}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, new_AGEMA_signal_2077, Midori_rounds_sub_sBox_PRINCE_0_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U13 ( .a ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, new_AGEMA_signal_2089, Midori_rounds_sub_sBox_PRINCE_0_n8}), .b ({new_AGEMA_signal_2088, new_AGEMA_signal_2087, new_AGEMA_signal_2086, Midori_rounds_sub_sBox_PRINCE_0_n7}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_2844, new_AGEMA_signal_2843, new_AGEMA_signal_2842, Midori_rounds_sub_sBox_PRINCE_0_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U10 ( .a ({new_AGEMA_signal_2076, new_AGEMA_signal_2075, new_AGEMA_signal_2074, Midori_rounds_roundReg_out[3]}), .b ({new_AGEMA_signal_2094, new_AGEMA_signal_2093, new_AGEMA_signal_2092, Midori_rounds_sub_sBox_PRINCE_0_n9}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, new_AGEMA_signal_2845, Midori_rounds_sub_sBox_PRINCE_0_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U9 ( .a ({new_AGEMA_signal_2082, new_AGEMA_signal_2081, new_AGEMA_signal_2080, Midori_rounds_roundReg_out[2]}), .b ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, new_AGEMA_signal_2089, Midori_rounds_sub_sBox_PRINCE_0_n8}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_2850, new_AGEMA_signal_2849, new_AGEMA_signal_2848, Midori_rounds_sub_sBox_PRINCE_0_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U5 ( .a ({new_AGEMA_signal_2082, new_AGEMA_signal_2081, new_AGEMA_signal_2080, Midori_rounds_roundReg_out[2]}), .b ({new_AGEMA_signal_2076, new_AGEMA_signal_2075, new_AGEMA_signal_2074, Midori_rounds_roundReg_out[3]}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, new_AGEMA_signal_2083, Midori_rounds_sub_sBox_PRINCE_0_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U3 ( .a ({new_AGEMA_signal_2094, new_AGEMA_signal_2093, new_AGEMA_signal_2092, Midori_rounds_sub_sBox_PRINCE_0_n9}), .b ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, new_AGEMA_signal_2089, Midori_rounds_sub_sBox_PRINCE_0_n8}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_2856, new_AGEMA_signal_2855, new_AGEMA_signal_2854, Midori_rounds_sub_sBox_PRINCE_0_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U14 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, new_AGEMA_signal_2095, Midori_rounds_roundReg_out[4]}), .b ({new_AGEMA_signal_2100, new_AGEMA_signal_2099, new_AGEMA_signal_2098, Midori_rounds_roundReg_out[7]}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, new_AGEMA_signal_2101, Midori_rounds_sub_sBox_PRINCE_1_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U13 ( .a ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, new_AGEMA_signal_2113, Midori_rounds_sub_sBox_PRINCE_1_n8}), .b ({new_AGEMA_signal_2112, new_AGEMA_signal_2111, new_AGEMA_signal_2110, Midori_rounds_sub_sBox_PRINCE_1_n7}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_2862, new_AGEMA_signal_2861, new_AGEMA_signal_2860, Midori_rounds_sub_sBox_PRINCE_1_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U10 ( .a ({new_AGEMA_signal_2100, new_AGEMA_signal_2099, new_AGEMA_signal_2098, Midori_rounds_roundReg_out[7]}), .b ({new_AGEMA_signal_2118, new_AGEMA_signal_2117, new_AGEMA_signal_2116, Midori_rounds_sub_sBox_PRINCE_1_n9}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, new_AGEMA_signal_2863, Midori_rounds_sub_sBox_PRINCE_1_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U9 ( .a ({new_AGEMA_signal_2106, new_AGEMA_signal_2105, new_AGEMA_signal_2104, Midori_rounds_roundReg_out[6]}), .b ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, new_AGEMA_signal_2113, Midori_rounds_sub_sBox_PRINCE_1_n8}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_2868, new_AGEMA_signal_2867, new_AGEMA_signal_2866, Midori_rounds_sub_sBox_PRINCE_1_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U5 ( .a ({new_AGEMA_signal_2106, new_AGEMA_signal_2105, new_AGEMA_signal_2104, Midori_rounds_roundReg_out[6]}), .b ({new_AGEMA_signal_2100, new_AGEMA_signal_2099, new_AGEMA_signal_2098, Midori_rounds_roundReg_out[7]}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, new_AGEMA_signal_2107, Midori_rounds_sub_sBox_PRINCE_1_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U3 ( .a ({new_AGEMA_signal_2118, new_AGEMA_signal_2117, new_AGEMA_signal_2116, Midori_rounds_sub_sBox_PRINCE_1_n9}), .b ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, new_AGEMA_signal_2113, Midori_rounds_sub_sBox_PRINCE_1_n8}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_2874, new_AGEMA_signal_2873, new_AGEMA_signal_2872, Midori_rounds_sub_sBox_PRINCE_1_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U14 ( .a ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, new_AGEMA_signal_2119, Midori_rounds_roundReg_out[8]}), .b ({new_AGEMA_signal_2124, new_AGEMA_signal_2123, new_AGEMA_signal_2122, Midori_rounds_roundReg_out[11]}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, new_AGEMA_signal_2125, Midori_rounds_sub_sBox_PRINCE_2_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U13 ( .a ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, new_AGEMA_signal_2137, Midori_rounds_sub_sBox_PRINCE_2_n8}), .b ({new_AGEMA_signal_2136, new_AGEMA_signal_2135, new_AGEMA_signal_2134, Midori_rounds_sub_sBox_PRINCE_2_n7}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_2880, new_AGEMA_signal_2879, new_AGEMA_signal_2878, Midori_rounds_sub_sBox_PRINCE_2_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U10 ( .a ({new_AGEMA_signal_2124, new_AGEMA_signal_2123, new_AGEMA_signal_2122, Midori_rounds_roundReg_out[11]}), .b ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, new_AGEMA_signal_2140, Midori_rounds_sub_sBox_PRINCE_2_n9}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, new_AGEMA_signal_2881, Midori_rounds_sub_sBox_PRINCE_2_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U9 ( .a ({new_AGEMA_signal_2130, new_AGEMA_signal_2129, new_AGEMA_signal_2128, Midori_rounds_roundReg_out[10]}), .b ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, new_AGEMA_signal_2137, Midori_rounds_sub_sBox_PRINCE_2_n8}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_2886, new_AGEMA_signal_2885, new_AGEMA_signal_2884, Midori_rounds_sub_sBox_PRINCE_2_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U5 ( .a ({new_AGEMA_signal_2130, new_AGEMA_signal_2129, new_AGEMA_signal_2128, Midori_rounds_roundReg_out[10]}), .b ({new_AGEMA_signal_2124, new_AGEMA_signal_2123, new_AGEMA_signal_2122, Midori_rounds_roundReg_out[11]}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, new_AGEMA_signal_2131, Midori_rounds_sub_sBox_PRINCE_2_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U3 ( .a ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, new_AGEMA_signal_2140, Midori_rounds_sub_sBox_PRINCE_2_n9}), .b ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, new_AGEMA_signal_2137, Midori_rounds_sub_sBox_PRINCE_2_n8}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_2892, new_AGEMA_signal_2891, new_AGEMA_signal_2890, Midori_rounds_sub_sBox_PRINCE_2_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U14 ( .a ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, new_AGEMA_signal_2143, Midori_rounds_roundReg_out[12]}), .b ({new_AGEMA_signal_2148, new_AGEMA_signal_2147, new_AGEMA_signal_2146, Midori_rounds_roundReg_out[15]}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, new_AGEMA_signal_2149, Midori_rounds_sub_sBox_PRINCE_3_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U13 ( .a ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, new_AGEMA_signal_2161, Midori_rounds_sub_sBox_PRINCE_3_n8}), .b ({new_AGEMA_signal_2160, new_AGEMA_signal_2159, new_AGEMA_signal_2158, Midori_rounds_sub_sBox_PRINCE_3_n7}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_2898, new_AGEMA_signal_2897, new_AGEMA_signal_2896, Midori_rounds_sub_sBox_PRINCE_3_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U10 ( .a ({new_AGEMA_signal_2148, new_AGEMA_signal_2147, new_AGEMA_signal_2146, Midori_rounds_roundReg_out[15]}), .b ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, new_AGEMA_signal_2164, Midori_rounds_sub_sBox_PRINCE_3_n9}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, new_AGEMA_signal_2899, Midori_rounds_sub_sBox_PRINCE_3_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U9 ( .a ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, new_AGEMA_signal_2152, Midori_rounds_roundReg_out[14]}), .b ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, new_AGEMA_signal_2161, Midori_rounds_sub_sBox_PRINCE_3_n8}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_2904, new_AGEMA_signal_2903, new_AGEMA_signal_2902, Midori_rounds_sub_sBox_PRINCE_3_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U5 ( .a ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, new_AGEMA_signal_2152, Midori_rounds_roundReg_out[14]}), .b ({new_AGEMA_signal_2148, new_AGEMA_signal_2147, new_AGEMA_signal_2146, Midori_rounds_roundReg_out[15]}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, new_AGEMA_signal_2155, Midori_rounds_sub_sBox_PRINCE_3_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U3 ( .a ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, new_AGEMA_signal_2164, Midori_rounds_sub_sBox_PRINCE_3_n9}), .b ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, new_AGEMA_signal_2161, Midori_rounds_sub_sBox_PRINCE_3_n8}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_2910, new_AGEMA_signal_2909, new_AGEMA_signal_2908, Midori_rounds_sub_sBox_PRINCE_3_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U14 ( .a ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, new_AGEMA_signal_2167, Midori_rounds_roundReg_out[16]}), .b ({new_AGEMA_signal_2172, new_AGEMA_signal_2171, new_AGEMA_signal_2170, Midori_rounds_roundReg_out[19]}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, new_AGEMA_signal_2173, Midori_rounds_sub_sBox_PRINCE_4_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U13 ( .a ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, new_AGEMA_signal_2185, Midori_rounds_sub_sBox_PRINCE_4_n8}), .b ({new_AGEMA_signal_2184, new_AGEMA_signal_2183, new_AGEMA_signal_2182, Midori_rounds_sub_sBox_PRINCE_4_n7}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_2916, new_AGEMA_signal_2915, new_AGEMA_signal_2914, Midori_rounds_sub_sBox_PRINCE_4_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U10 ( .a ({new_AGEMA_signal_2172, new_AGEMA_signal_2171, new_AGEMA_signal_2170, Midori_rounds_roundReg_out[19]}), .b ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, new_AGEMA_signal_2188, Midori_rounds_sub_sBox_PRINCE_4_n9}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, new_AGEMA_signal_2917, Midori_rounds_sub_sBox_PRINCE_4_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U9 ( .a ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, new_AGEMA_signal_2176, Midori_rounds_roundReg_out[18]}), .b ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, new_AGEMA_signal_2185, Midori_rounds_sub_sBox_PRINCE_4_n8}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_2922, new_AGEMA_signal_2921, new_AGEMA_signal_2920, Midori_rounds_sub_sBox_PRINCE_4_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U5 ( .a ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, new_AGEMA_signal_2176, Midori_rounds_roundReg_out[18]}), .b ({new_AGEMA_signal_2172, new_AGEMA_signal_2171, new_AGEMA_signal_2170, Midori_rounds_roundReg_out[19]}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, new_AGEMA_signal_2179, Midori_rounds_sub_sBox_PRINCE_4_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U3 ( .a ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, new_AGEMA_signal_2188, Midori_rounds_sub_sBox_PRINCE_4_n9}), .b ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, new_AGEMA_signal_2185, Midori_rounds_sub_sBox_PRINCE_4_n8}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_2928, new_AGEMA_signal_2927, new_AGEMA_signal_2926, Midori_rounds_sub_sBox_PRINCE_4_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U14 ( .a ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, new_AGEMA_signal_2191, Midori_rounds_roundReg_out[20]}), .b ({new_AGEMA_signal_2196, new_AGEMA_signal_2195, new_AGEMA_signal_2194, Midori_rounds_roundReg_out[23]}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, new_AGEMA_signal_2197, Midori_rounds_sub_sBox_PRINCE_5_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U13 ( .a ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, new_AGEMA_signal_2209, Midori_rounds_sub_sBox_PRINCE_5_n8}), .b ({new_AGEMA_signal_2208, new_AGEMA_signal_2207, new_AGEMA_signal_2206, Midori_rounds_sub_sBox_PRINCE_5_n7}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_2934, new_AGEMA_signal_2933, new_AGEMA_signal_2932, Midori_rounds_sub_sBox_PRINCE_5_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U10 ( .a ({new_AGEMA_signal_2196, new_AGEMA_signal_2195, new_AGEMA_signal_2194, Midori_rounds_roundReg_out[23]}), .b ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, new_AGEMA_signal_2212, Midori_rounds_sub_sBox_PRINCE_5_n9}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, new_AGEMA_signal_2935, Midori_rounds_sub_sBox_PRINCE_5_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U9 ( .a ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, new_AGEMA_signal_2200, Midori_rounds_roundReg_out[22]}), .b ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, new_AGEMA_signal_2209, Midori_rounds_sub_sBox_PRINCE_5_n8}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_2940, new_AGEMA_signal_2939, new_AGEMA_signal_2938, Midori_rounds_sub_sBox_PRINCE_5_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U5 ( .a ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, new_AGEMA_signal_2200, Midori_rounds_roundReg_out[22]}), .b ({new_AGEMA_signal_2196, new_AGEMA_signal_2195, new_AGEMA_signal_2194, Midori_rounds_roundReg_out[23]}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, new_AGEMA_signal_2203, Midori_rounds_sub_sBox_PRINCE_5_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U3 ( .a ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, new_AGEMA_signal_2212, Midori_rounds_sub_sBox_PRINCE_5_n9}), .b ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, new_AGEMA_signal_2209, Midori_rounds_sub_sBox_PRINCE_5_n8}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_2946, new_AGEMA_signal_2945, new_AGEMA_signal_2944, Midori_rounds_sub_sBox_PRINCE_5_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U14 ( .a ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, new_AGEMA_signal_2215, Midori_rounds_roundReg_out[24]}), .b ({new_AGEMA_signal_2220, new_AGEMA_signal_2219, new_AGEMA_signal_2218, Midori_rounds_roundReg_out[27]}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, new_AGEMA_signal_2221, Midori_rounds_sub_sBox_PRINCE_6_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U13 ( .a ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, new_AGEMA_signal_2233, Midori_rounds_sub_sBox_PRINCE_6_n8}), .b ({new_AGEMA_signal_2232, new_AGEMA_signal_2231, new_AGEMA_signal_2230, Midori_rounds_sub_sBox_PRINCE_6_n7}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_2952, new_AGEMA_signal_2951, new_AGEMA_signal_2950, Midori_rounds_sub_sBox_PRINCE_6_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U10 ( .a ({new_AGEMA_signal_2220, new_AGEMA_signal_2219, new_AGEMA_signal_2218, Midori_rounds_roundReg_out[27]}), .b ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, new_AGEMA_signal_2236, Midori_rounds_sub_sBox_PRINCE_6_n9}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, new_AGEMA_signal_2953, Midori_rounds_sub_sBox_PRINCE_6_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U9 ( .a ({new_AGEMA_signal_2226, new_AGEMA_signal_2225, new_AGEMA_signal_2224, Midori_rounds_roundReg_out[26]}), .b ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, new_AGEMA_signal_2233, Midori_rounds_sub_sBox_PRINCE_6_n8}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_2958, new_AGEMA_signal_2957, new_AGEMA_signal_2956, Midori_rounds_sub_sBox_PRINCE_6_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U5 ( .a ({new_AGEMA_signal_2226, new_AGEMA_signal_2225, new_AGEMA_signal_2224, Midori_rounds_roundReg_out[26]}), .b ({new_AGEMA_signal_2220, new_AGEMA_signal_2219, new_AGEMA_signal_2218, Midori_rounds_roundReg_out[27]}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, new_AGEMA_signal_2227, Midori_rounds_sub_sBox_PRINCE_6_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U3 ( .a ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, new_AGEMA_signal_2236, Midori_rounds_sub_sBox_PRINCE_6_n9}), .b ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, new_AGEMA_signal_2233, Midori_rounds_sub_sBox_PRINCE_6_n8}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_2964, new_AGEMA_signal_2963, new_AGEMA_signal_2962, Midori_rounds_sub_sBox_PRINCE_6_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U14 ( .a ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, new_AGEMA_signal_2239, Midori_rounds_roundReg_out[28]}), .b ({new_AGEMA_signal_2244, new_AGEMA_signal_2243, new_AGEMA_signal_2242, Midori_rounds_roundReg_out[31]}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, new_AGEMA_signal_2245, Midori_rounds_sub_sBox_PRINCE_7_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U13 ( .a ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, new_AGEMA_signal_2257, Midori_rounds_sub_sBox_PRINCE_7_n8}), .b ({new_AGEMA_signal_2256, new_AGEMA_signal_2255, new_AGEMA_signal_2254, Midori_rounds_sub_sBox_PRINCE_7_n7}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_2970, new_AGEMA_signal_2969, new_AGEMA_signal_2968, Midori_rounds_sub_sBox_PRINCE_7_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U10 ( .a ({new_AGEMA_signal_2244, new_AGEMA_signal_2243, new_AGEMA_signal_2242, Midori_rounds_roundReg_out[31]}), .b ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, new_AGEMA_signal_2260, Midori_rounds_sub_sBox_PRINCE_7_n9}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, new_AGEMA_signal_2971, Midori_rounds_sub_sBox_PRINCE_7_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U9 ( .a ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, new_AGEMA_signal_2248, Midori_rounds_roundReg_out[30]}), .b ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, new_AGEMA_signal_2257, Midori_rounds_sub_sBox_PRINCE_7_n8}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_2976, new_AGEMA_signal_2975, new_AGEMA_signal_2974, Midori_rounds_sub_sBox_PRINCE_7_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U5 ( .a ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, new_AGEMA_signal_2248, Midori_rounds_roundReg_out[30]}), .b ({new_AGEMA_signal_2244, new_AGEMA_signal_2243, new_AGEMA_signal_2242, Midori_rounds_roundReg_out[31]}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, new_AGEMA_signal_2251, Midori_rounds_sub_sBox_PRINCE_7_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U3 ( .a ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, new_AGEMA_signal_2260, Midori_rounds_sub_sBox_PRINCE_7_n9}), .b ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, new_AGEMA_signal_2257, Midori_rounds_sub_sBox_PRINCE_7_n8}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_2982, new_AGEMA_signal_2981, new_AGEMA_signal_2980, Midori_rounds_sub_sBox_PRINCE_7_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U14 ( .a ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, new_AGEMA_signal_2263, Midori_rounds_roundReg_out[32]}), .b ({new_AGEMA_signal_2268, new_AGEMA_signal_2267, new_AGEMA_signal_2266, Midori_rounds_roundReg_out[35]}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, new_AGEMA_signal_2269, Midori_rounds_sub_sBox_PRINCE_8_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U13 ( .a ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, new_AGEMA_signal_2281, Midori_rounds_sub_sBox_PRINCE_8_n8}), .b ({new_AGEMA_signal_2280, new_AGEMA_signal_2279, new_AGEMA_signal_2278, Midori_rounds_sub_sBox_PRINCE_8_n7}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_2988, new_AGEMA_signal_2987, new_AGEMA_signal_2986, Midori_rounds_sub_sBox_PRINCE_8_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U10 ( .a ({new_AGEMA_signal_2268, new_AGEMA_signal_2267, new_AGEMA_signal_2266, Midori_rounds_roundReg_out[35]}), .b ({new_AGEMA_signal_2286, new_AGEMA_signal_2285, new_AGEMA_signal_2284, Midori_rounds_sub_sBox_PRINCE_8_n9}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, new_AGEMA_signal_2989, Midori_rounds_sub_sBox_PRINCE_8_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U9 ( .a ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, new_AGEMA_signal_2272, Midori_rounds_roundReg_out[34]}), .b ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, new_AGEMA_signal_2281, Midori_rounds_sub_sBox_PRINCE_8_n8}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_2994, new_AGEMA_signal_2993, new_AGEMA_signal_2992, Midori_rounds_sub_sBox_PRINCE_8_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U5 ( .a ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, new_AGEMA_signal_2272, Midori_rounds_roundReg_out[34]}), .b ({new_AGEMA_signal_2268, new_AGEMA_signal_2267, new_AGEMA_signal_2266, Midori_rounds_roundReg_out[35]}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, new_AGEMA_signal_2275, Midori_rounds_sub_sBox_PRINCE_8_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U3 ( .a ({new_AGEMA_signal_2286, new_AGEMA_signal_2285, new_AGEMA_signal_2284, Midori_rounds_sub_sBox_PRINCE_8_n9}), .b ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, new_AGEMA_signal_2281, Midori_rounds_sub_sBox_PRINCE_8_n8}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_3000, new_AGEMA_signal_2999, new_AGEMA_signal_2998, Midori_rounds_sub_sBox_PRINCE_8_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U14 ( .a ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, new_AGEMA_signal_2287, Midori_rounds_roundReg_out[36]}), .b ({new_AGEMA_signal_2292, new_AGEMA_signal_2291, new_AGEMA_signal_2290, Midori_rounds_roundReg_out[39]}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, new_AGEMA_signal_2293, Midori_rounds_sub_sBox_PRINCE_9_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U13 ( .a ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, new_AGEMA_signal_2305, Midori_rounds_sub_sBox_PRINCE_9_n8}), .b ({new_AGEMA_signal_2304, new_AGEMA_signal_2303, new_AGEMA_signal_2302, Midori_rounds_sub_sBox_PRINCE_9_n7}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_3006, new_AGEMA_signal_3005, new_AGEMA_signal_3004, Midori_rounds_sub_sBox_PRINCE_9_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U10 ( .a ({new_AGEMA_signal_2292, new_AGEMA_signal_2291, new_AGEMA_signal_2290, Midori_rounds_roundReg_out[39]}), .b ({new_AGEMA_signal_2310, new_AGEMA_signal_2309, new_AGEMA_signal_2308, Midori_rounds_sub_sBox_PRINCE_9_n9}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_3009, new_AGEMA_signal_3008, new_AGEMA_signal_3007, Midori_rounds_sub_sBox_PRINCE_9_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U9 ( .a ({new_AGEMA_signal_2298, new_AGEMA_signal_2297, new_AGEMA_signal_2296, Midori_rounds_roundReg_out[38]}), .b ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, new_AGEMA_signal_2305, Midori_rounds_sub_sBox_PRINCE_9_n8}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_3012, new_AGEMA_signal_3011, new_AGEMA_signal_3010, Midori_rounds_sub_sBox_PRINCE_9_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U5 ( .a ({new_AGEMA_signal_2298, new_AGEMA_signal_2297, new_AGEMA_signal_2296, Midori_rounds_roundReg_out[38]}), .b ({new_AGEMA_signal_2292, new_AGEMA_signal_2291, new_AGEMA_signal_2290, Midori_rounds_roundReg_out[39]}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, new_AGEMA_signal_2299, Midori_rounds_sub_sBox_PRINCE_9_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U3 ( .a ({new_AGEMA_signal_2310, new_AGEMA_signal_2309, new_AGEMA_signal_2308, Midori_rounds_sub_sBox_PRINCE_9_n9}), .b ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, new_AGEMA_signal_2305, Midori_rounds_sub_sBox_PRINCE_9_n8}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_3018, new_AGEMA_signal_3017, new_AGEMA_signal_3016, Midori_rounds_sub_sBox_PRINCE_9_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U14 ( .a ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, new_AGEMA_signal_2311, Midori_rounds_roundReg_out[40]}), .b ({new_AGEMA_signal_2316, new_AGEMA_signal_2315, new_AGEMA_signal_2314, Midori_rounds_roundReg_out[43]}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, new_AGEMA_signal_2317, Midori_rounds_sub_sBox_PRINCE_10_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U13 ( .a ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, new_AGEMA_signal_2329, Midori_rounds_sub_sBox_PRINCE_10_n8}), .b ({new_AGEMA_signal_2328, new_AGEMA_signal_2327, new_AGEMA_signal_2326, Midori_rounds_sub_sBox_PRINCE_10_n7}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_3024, new_AGEMA_signal_3023, new_AGEMA_signal_3022, Midori_rounds_sub_sBox_PRINCE_10_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U10 ( .a ({new_AGEMA_signal_2316, new_AGEMA_signal_2315, new_AGEMA_signal_2314, Midori_rounds_roundReg_out[43]}), .b ({new_AGEMA_signal_2334, new_AGEMA_signal_2333, new_AGEMA_signal_2332, Midori_rounds_sub_sBox_PRINCE_10_n9}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, new_AGEMA_signal_3025, Midori_rounds_sub_sBox_PRINCE_10_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U9 ( .a ({new_AGEMA_signal_2322, new_AGEMA_signal_2321, new_AGEMA_signal_2320, Midori_rounds_roundReg_out[42]}), .b ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, new_AGEMA_signal_2329, Midori_rounds_sub_sBox_PRINCE_10_n8}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_3030, new_AGEMA_signal_3029, new_AGEMA_signal_3028, Midori_rounds_sub_sBox_PRINCE_10_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U5 ( .a ({new_AGEMA_signal_2322, new_AGEMA_signal_2321, new_AGEMA_signal_2320, Midori_rounds_roundReg_out[42]}), .b ({new_AGEMA_signal_2316, new_AGEMA_signal_2315, new_AGEMA_signal_2314, Midori_rounds_roundReg_out[43]}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, new_AGEMA_signal_2323, Midori_rounds_sub_sBox_PRINCE_10_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U3 ( .a ({new_AGEMA_signal_2334, new_AGEMA_signal_2333, new_AGEMA_signal_2332, Midori_rounds_sub_sBox_PRINCE_10_n9}), .b ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, new_AGEMA_signal_2329, Midori_rounds_sub_sBox_PRINCE_10_n8}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_3036, new_AGEMA_signal_3035, new_AGEMA_signal_3034, Midori_rounds_sub_sBox_PRINCE_10_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U14 ( .a ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, new_AGEMA_signal_2335, Midori_rounds_roundReg_out[44]}), .b ({new_AGEMA_signal_2340, new_AGEMA_signal_2339, new_AGEMA_signal_2338, Midori_rounds_roundReg_out[47]}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, new_AGEMA_signal_2341, Midori_rounds_sub_sBox_PRINCE_11_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U13 ( .a ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, new_AGEMA_signal_2353, Midori_rounds_sub_sBox_PRINCE_11_n8}), .b ({new_AGEMA_signal_2352, new_AGEMA_signal_2351, new_AGEMA_signal_2350, Midori_rounds_sub_sBox_PRINCE_11_n7}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_3042, new_AGEMA_signal_3041, new_AGEMA_signal_3040, Midori_rounds_sub_sBox_PRINCE_11_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U10 ( .a ({new_AGEMA_signal_2340, new_AGEMA_signal_2339, new_AGEMA_signal_2338, Midori_rounds_roundReg_out[47]}), .b ({new_AGEMA_signal_2358, new_AGEMA_signal_2357, new_AGEMA_signal_2356, Midori_rounds_sub_sBox_PRINCE_11_n9}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, new_AGEMA_signal_3043, Midori_rounds_sub_sBox_PRINCE_11_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U9 ( .a ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, new_AGEMA_signal_2344, Midori_rounds_roundReg_out[46]}), .b ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, new_AGEMA_signal_2353, Midori_rounds_sub_sBox_PRINCE_11_n8}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_3048, new_AGEMA_signal_3047, new_AGEMA_signal_3046, Midori_rounds_sub_sBox_PRINCE_11_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U5 ( .a ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, new_AGEMA_signal_2344, Midori_rounds_roundReg_out[46]}), .b ({new_AGEMA_signal_2340, new_AGEMA_signal_2339, new_AGEMA_signal_2338, Midori_rounds_roundReg_out[47]}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, new_AGEMA_signal_2347, Midori_rounds_sub_sBox_PRINCE_11_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U3 ( .a ({new_AGEMA_signal_2358, new_AGEMA_signal_2357, new_AGEMA_signal_2356, Midori_rounds_sub_sBox_PRINCE_11_n9}), .b ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, new_AGEMA_signal_2353, Midori_rounds_sub_sBox_PRINCE_11_n8}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_3054, new_AGEMA_signal_3053, new_AGEMA_signal_3052, Midori_rounds_sub_sBox_PRINCE_11_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U14 ( .a ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, new_AGEMA_signal_2359, Midori_rounds_roundReg_out[48]}), .b ({new_AGEMA_signal_2364, new_AGEMA_signal_2363, new_AGEMA_signal_2362, Midori_rounds_roundReg_out[51]}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, new_AGEMA_signal_2365, Midori_rounds_sub_sBox_PRINCE_12_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U13 ( .a ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, new_AGEMA_signal_2377, Midori_rounds_sub_sBox_PRINCE_12_n8}), .b ({new_AGEMA_signal_2376, new_AGEMA_signal_2375, new_AGEMA_signal_2374, Midori_rounds_sub_sBox_PRINCE_12_n7}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_3060, new_AGEMA_signal_3059, new_AGEMA_signal_3058, Midori_rounds_sub_sBox_PRINCE_12_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U10 ( .a ({new_AGEMA_signal_2364, new_AGEMA_signal_2363, new_AGEMA_signal_2362, Midori_rounds_roundReg_out[51]}), .b ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, new_AGEMA_signal_2380, Midori_rounds_sub_sBox_PRINCE_12_n9}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, new_AGEMA_signal_3061, Midori_rounds_sub_sBox_PRINCE_12_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U9 ( .a ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, new_AGEMA_signal_2368, Midori_rounds_roundReg_out[50]}), .b ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, new_AGEMA_signal_2377, Midori_rounds_sub_sBox_PRINCE_12_n8}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_3066, new_AGEMA_signal_3065, new_AGEMA_signal_3064, Midori_rounds_sub_sBox_PRINCE_12_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U5 ( .a ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, new_AGEMA_signal_2368, Midori_rounds_roundReg_out[50]}), .b ({new_AGEMA_signal_2364, new_AGEMA_signal_2363, new_AGEMA_signal_2362, Midori_rounds_roundReg_out[51]}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, new_AGEMA_signal_2371, Midori_rounds_sub_sBox_PRINCE_12_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U3 ( .a ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, new_AGEMA_signal_2380, Midori_rounds_sub_sBox_PRINCE_12_n9}), .b ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, new_AGEMA_signal_2377, Midori_rounds_sub_sBox_PRINCE_12_n8}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_3072, new_AGEMA_signal_3071, new_AGEMA_signal_3070, Midori_rounds_sub_sBox_PRINCE_12_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U14 ( .a ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, new_AGEMA_signal_2383, Midori_rounds_roundReg_out[52]}), .b ({new_AGEMA_signal_2388, new_AGEMA_signal_2387, new_AGEMA_signal_2386, Midori_rounds_roundReg_out[55]}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, new_AGEMA_signal_2389, Midori_rounds_sub_sBox_PRINCE_13_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U13 ( .a ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, new_AGEMA_signal_2401, Midori_rounds_sub_sBox_PRINCE_13_n8}), .b ({new_AGEMA_signal_2400, new_AGEMA_signal_2399, new_AGEMA_signal_2398, Midori_rounds_sub_sBox_PRINCE_13_n7}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_3078, new_AGEMA_signal_3077, new_AGEMA_signal_3076, Midori_rounds_sub_sBox_PRINCE_13_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U10 ( .a ({new_AGEMA_signal_2388, new_AGEMA_signal_2387, new_AGEMA_signal_2386, Midori_rounds_roundReg_out[55]}), .b ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, new_AGEMA_signal_2404, Midori_rounds_sub_sBox_PRINCE_13_n9}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, new_AGEMA_signal_3079, Midori_rounds_sub_sBox_PRINCE_13_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U9 ( .a ({new_AGEMA_signal_2394, new_AGEMA_signal_2393, new_AGEMA_signal_2392, Midori_rounds_roundReg_out[54]}), .b ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, new_AGEMA_signal_2401, Midori_rounds_sub_sBox_PRINCE_13_n8}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_3084, new_AGEMA_signal_3083, new_AGEMA_signal_3082, Midori_rounds_sub_sBox_PRINCE_13_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U5 ( .a ({new_AGEMA_signal_2394, new_AGEMA_signal_2393, new_AGEMA_signal_2392, Midori_rounds_roundReg_out[54]}), .b ({new_AGEMA_signal_2388, new_AGEMA_signal_2387, new_AGEMA_signal_2386, Midori_rounds_roundReg_out[55]}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, new_AGEMA_signal_2395, Midori_rounds_sub_sBox_PRINCE_13_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U3 ( .a ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, new_AGEMA_signal_2404, Midori_rounds_sub_sBox_PRINCE_13_n9}), .b ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, new_AGEMA_signal_2401, Midori_rounds_sub_sBox_PRINCE_13_n8}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_3090, new_AGEMA_signal_3089, new_AGEMA_signal_3088, Midori_rounds_sub_sBox_PRINCE_13_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U14 ( .a ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, new_AGEMA_signal_2407, Midori_rounds_roundReg_out[56]}), .b ({new_AGEMA_signal_2412, new_AGEMA_signal_2411, new_AGEMA_signal_2410, Midori_rounds_roundReg_out[59]}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, new_AGEMA_signal_2413, Midori_rounds_sub_sBox_PRINCE_14_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U13 ( .a ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, new_AGEMA_signal_2425, Midori_rounds_sub_sBox_PRINCE_14_n8}), .b ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, new_AGEMA_signal_2422, Midori_rounds_sub_sBox_PRINCE_14_n7}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_3096, new_AGEMA_signal_3095, new_AGEMA_signal_3094, Midori_rounds_sub_sBox_PRINCE_14_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U10 ( .a ({new_AGEMA_signal_2412, new_AGEMA_signal_2411, new_AGEMA_signal_2410, Midori_rounds_roundReg_out[59]}), .b ({new_AGEMA_signal_2430, new_AGEMA_signal_2429, new_AGEMA_signal_2428, Midori_rounds_sub_sBox_PRINCE_14_n9}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, new_AGEMA_signal_3097, Midori_rounds_sub_sBox_PRINCE_14_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U9 ( .a ({new_AGEMA_signal_2418, new_AGEMA_signal_2417, new_AGEMA_signal_2416, Midori_rounds_roundReg_out[58]}), .b ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, new_AGEMA_signal_2425, Midori_rounds_sub_sBox_PRINCE_14_n8}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_3102, new_AGEMA_signal_3101, new_AGEMA_signal_3100, Midori_rounds_sub_sBox_PRINCE_14_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U5 ( .a ({new_AGEMA_signal_2418, new_AGEMA_signal_2417, new_AGEMA_signal_2416, Midori_rounds_roundReg_out[58]}), .b ({new_AGEMA_signal_2412, new_AGEMA_signal_2411, new_AGEMA_signal_2410, Midori_rounds_roundReg_out[59]}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, new_AGEMA_signal_2419, Midori_rounds_sub_sBox_PRINCE_14_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U3 ( .a ({new_AGEMA_signal_2430, new_AGEMA_signal_2429, new_AGEMA_signal_2428, Midori_rounds_sub_sBox_PRINCE_14_n9}), .b ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, new_AGEMA_signal_2425, Midori_rounds_sub_sBox_PRINCE_14_n8}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_3108, new_AGEMA_signal_3107, new_AGEMA_signal_3106, Midori_rounds_sub_sBox_PRINCE_14_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U14 ( .a ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, new_AGEMA_signal_2431, Midori_rounds_roundReg_out[60]}), .b ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, new_AGEMA_signal_2434, Midori_rounds_roundReg_out[63]}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, new_AGEMA_signal_2437, Midori_rounds_sub_sBox_PRINCE_15_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U13 ( .a ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, new_AGEMA_signal_2449, Midori_rounds_sub_sBox_PRINCE_15_n8}), .b ({new_AGEMA_signal_2448, new_AGEMA_signal_2447, new_AGEMA_signal_2446, Midori_rounds_sub_sBox_PRINCE_15_n7}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_3114, new_AGEMA_signal_3113, new_AGEMA_signal_3112, Midori_rounds_sub_sBox_PRINCE_15_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U10 ( .a ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, new_AGEMA_signal_2434, Midori_rounds_roundReg_out[63]}), .b ({new_AGEMA_signal_2454, new_AGEMA_signal_2453, new_AGEMA_signal_2452, Midori_rounds_sub_sBox_PRINCE_15_n9}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, new_AGEMA_signal_3115, Midori_rounds_sub_sBox_PRINCE_15_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U9 ( .a ({new_AGEMA_signal_2442, new_AGEMA_signal_2441, new_AGEMA_signal_2440, Midori_rounds_roundReg_out[62]}), .b ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, new_AGEMA_signal_2449, Midori_rounds_sub_sBox_PRINCE_15_n8}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_3120, new_AGEMA_signal_3119, new_AGEMA_signal_3118, Midori_rounds_sub_sBox_PRINCE_15_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U5 ( .a ({new_AGEMA_signal_2442, new_AGEMA_signal_2441, new_AGEMA_signal_2440, Midori_rounds_roundReg_out[62]}), .b ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, new_AGEMA_signal_2434, Midori_rounds_roundReg_out[63]}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, new_AGEMA_signal_2443, Midori_rounds_sub_sBox_PRINCE_15_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U3 ( .a ({new_AGEMA_signal_2454, new_AGEMA_signal_2453, new_AGEMA_signal_2452, Midori_rounds_sub_sBox_PRINCE_15_n9}), .b ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, new_AGEMA_signal_2449, Midori_rounds_sub_sBox_PRINCE_15_n8}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_3126, new_AGEMA_signal_3125, new_AGEMA_signal_3124, Midori_rounds_sub_sBox_PRINCE_15_n13}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    or_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U18 ( .a ({new_AGEMA_signal_2856, new_AGEMA_signal_2855, new_AGEMA_signal_2854, Midori_rounds_sub_sBox_PRINCE_0_n13}), .b ({new_AGEMA_signal_3282, new_AGEMA_signal_3281, new_AGEMA_signal_3280, Midori_rounds_roundReg_out[1]}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, new_AGEMA_signal_3283, Midori_rounds_sub_sBox_PRINCE_0_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U15 ( .a ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, new_AGEMA_signal_2077, Midori_rounds_sub_sBox_PRINCE_0_n10}), .b ({new_AGEMA_signal_2094, new_AGEMA_signal_2093, new_AGEMA_signal_2092, Midori_rounds_sub_sBox_PRINCE_0_n9}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, new_AGEMA_signal_2839, Midori_rounds_sub_sBox_PRINCE_0_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U11 ( .a ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, new_AGEMA_signal_2071, Midori_rounds_roundReg_out[0]}), .b ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, new_AGEMA_signal_2845, Midori_rounds_sub_sBox_PRINCE_0_n4}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, new_AGEMA_signal_3289, Midori_rounds_sub_sBox_PRINCE_0_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U6 ( .a ({new_AGEMA_signal_2088, new_AGEMA_signal_2087, new_AGEMA_signal_2086, Midori_rounds_sub_sBox_PRINCE_0_n7}), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, new_AGEMA_signal_2083, Midori_rounds_sub_sBox_PRINCE_0_n1}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, new_AGEMA_signal_2851, Midori_rounds_sub_sBox_PRINCE_0_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U18 ( .a ({new_AGEMA_signal_2874, new_AGEMA_signal_2873, new_AGEMA_signal_2872, Midori_rounds_sub_sBox_PRINCE_1_n13}), .b ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, new_AGEMA_signal_3295, Midori_rounds_roundReg_out[5]}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_3300, new_AGEMA_signal_3299, new_AGEMA_signal_3298, Midori_rounds_sub_sBox_PRINCE_1_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U15 ( .a ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, new_AGEMA_signal_2101, Midori_rounds_sub_sBox_PRINCE_1_n10}), .b ({new_AGEMA_signal_2118, new_AGEMA_signal_2117, new_AGEMA_signal_2116, Midori_rounds_sub_sBox_PRINCE_1_n9}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, new_AGEMA_signal_2857, Midori_rounds_sub_sBox_PRINCE_1_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U11 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, new_AGEMA_signal_2095, Midori_rounds_roundReg_out[4]}), .b ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, new_AGEMA_signal_2863, Midori_rounds_sub_sBox_PRINCE_1_n4}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_3306, new_AGEMA_signal_3305, new_AGEMA_signal_3304, Midori_rounds_sub_sBox_PRINCE_1_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U6 ( .a ({new_AGEMA_signal_2112, new_AGEMA_signal_2111, new_AGEMA_signal_2110, Midori_rounds_sub_sBox_PRINCE_1_n7}), .b ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, new_AGEMA_signal_2107, Midori_rounds_sub_sBox_PRINCE_1_n1}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, new_AGEMA_signal_2869, Midori_rounds_sub_sBox_PRINCE_1_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U18 ( .a ({new_AGEMA_signal_2892, new_AGEMA_signal_2891, new_AGEMA_signal_2890, Midori_rounds_sub_sBox_PRINCE_2_n13}), .b ({new_AGEMA_signal_3312, new_AGEMA_signal_3311, new_AGEMA_signal_3310, Midori_rounds_roundReg_out[9]}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, new_AGEMA_signal_3313, Midori_rounds_sub_sBox_PRINCE_2_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U15 ( .a ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, new_AGEMA_signal_2125, Midori_rounds_sub_sBox_PRINCE_2_n10}), .b ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, new_AGEMA_signal_2140, Midori_rounds_sub_sBox_PRINCE_2_n9}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, new_AGEMA_signal_2875, Midori_rounds_sub_sBox_PRINCE_2_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U11 ( .a ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, new_AGEMA_signal_2119, Midori_rounds_roundReg_out[8]}), .b ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, new_AGEMA_signal_2881, Midori_rounds_sub_sBox_PRINCE_2_n4}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, new_AGEMA_signal_3319, Midori_rounds_sub_sBox_PRINCE_2_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U6 ( .a ({new_AGEMA_signal_2136, new_AGEMA_signal_2135, new_AGEMA_signal_2134, Midori_rounds_sub_sBox_PRINCE_2_n7}), .b ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, new_AGEMA_signal_2131, Midori_rounds_sub_sBox_PRINCE_2_n1}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, new_AGEMA_signal_2887, Midori_rounds_sub_sBox_PRINCE_2_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U18 ( .a ({new_AGEMA_signal_2910, new_AGEMA_signal_2909, new_AGEMA_signal_2908, Midori_rounds_sub_sBox_PRINCE_3_n13}), .b ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, new_AGEMA_signal_3325, Midori_rounds_roundReg_out[13]}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_3330, new_AGEMA_signal_3329, new_AGEMA_signal_3328, Midori_rounds_sub_sBox_PRINCE_3_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U15 ( .a ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, new_AGEMA_signal_2149, Midori_rounds_sub_sBox_PRINCE_3_n10}), .b ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, new_AGEMA_signal_2164, Midori_rounds_sub_sBox_PRINCE_3_n9}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, new_AGEMA_signal_2893, Midori_rounds_sub_sBox_PRINCE_3_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U11 ( .a ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, new_AGEMA_signal_2143, Midori_rounds_roundReg_out[12]}), .b ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, new_AGEMA_signal_2899, Midori_rounds_sub_sBox_PRINCE_3_n4}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_3336, new_AGEMA_signal_3335, new_AGEMA_signal_3334, Midori_rounds_sub_sBox_PRINCE_3_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U6 ( .a ({new_AGEMA_signal_2160, new_AGEMA_signal_2159, new_AGEMA_signal_2158, Midori_rounds_sub_sBox_PRINCE_3_n7}), .b ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, new_AGEMA_signal_2155, Midori_rounds_sub_sBox_PRINCE_3_n1}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, new_AGEMA_signal_2905, Midori_rounds_sub_sBox_PRINCE_3_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U18 ( .a ({new_AGEMA_signal_2928, new_AGEMA_signal_2927, new_AGEMA_signal_2926, Midori_rounds_sub_sBox_PRINCE_4_n13}), .b ({new_AGEMA_signal_3342, new_AGEMA_signal_3341, new_AGEMA_signal_3340, Midori_rounds_roundReg_out[17]}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, new_AGEMA_signal_3343, Midori_rounds_sub_sBox_PRINCE_4_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U15 ( .a ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, new_AGEMA_signal_2173, Midori_rounds_sub_sBox_PRINCE_4_n10}), .b ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, new_AGEMA_signal_2188, Midori_rounds_sub_sBox_PRINCE_4_n9}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, new_AGEMA_signal_2911, Midori_rounds_sub_sBox_PRINCE_4_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U11 ( .a ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, new_AGEMA_signal_2167, Midori_rounds_roundReg_out[16]}), .b ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, new_AGEMA_signal_2917, Midori_rounds_sub_sBox_PRINCE_4_n4}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, new_AGEMA_signal_3349, Midori_rounds_sub_sBox_PRINCE_4_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U6 ( .a ({new_AGEMA_signal_2184, new_AGEMA_signal_2183, new_AGEMA_signal_2182, Midori_rounds_sub_sBox_PRINCE_4_n7}), .b ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, new_AGEMA_signal_2179, Midori_rounds_sub_sBox_PRINCE_4_n1}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, new_AGEMA_signal_2923, Midori_rounds_sub_sBox_PRINCE_4_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U18 ( .a ({new_AGEMA_signal_2946, new_AGEMA_signal_2945, new_AGEMA_signal_2944, Midori_rounds_sub_sBox_PRINCE_5_n13}), .b ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, new_AGEMA_signal_3355, Midori_rounds_roundReg_out[21]}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_3360, new_AGEMA_signal_3359, new_AGEMA_signal_3358, Midori_rounds_sub_sBox_PRINCE_5_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U15 ( .a ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, new_AGEMA_signal_2197, Midori_rounds_sub_sBox_PRINCE_5_n10}), .b ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, new_AGEMA_signal_2212, Midori_rounds_sub_sBox_PRINCE_5_n9}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, new_AGEMA_signal_2929, Midori_rounds_sub_sBox_PRINCE_5_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U11 ( .a ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, new_AGEMA_signal_2191, Midori_rounds_roundReg_out[20]}), .b ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, new_AGEMA_signal_2935, Midori_rounds_sub_sBox_PRINCE_5_n4}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_3366, new_AGEMA_signal_3365, new_AGEMA_signal_3364, Midori_rounds_sub_sBox_PRINCE_5_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U6 ( .a ({new_AGEMA_signal_2208, new_AGEMA_signal_2207, new_AGEMA_signal_2206, Midori_rounds_sub_sBox_PRINCE_5_n7}), .b ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, new_AGEMA_signal_2203, Midori_rounds_sub_sBox_PRINCE_5_n1}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, new_AGEMA_signal_2941, Midori_rounds_sub_sBox_PRINCE_5_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U18 ( .a ({new_AGEMA_signal_2964, new_AGEMA_signal_2963, new_AGEMA_signal_2962, Midori_rounds_sub_sBox_PRINCE_6_n13}), .b ({new_AGEMA_signal_3372, new_AGEMA_signal_3371, new_AGEMA_signal_3370, Midori_rounds_roundReg_out[25]}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, new_AGEMA_signal_3373, Midori_rounds_sub_sBox_PRINCE_6_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U15 ( .a ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, new_AGEMA_signal_2221, Midori_rounds_sub_sBox_PRINCE_6_n10}), .b ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, new_AGEMA_signal_2236, Midori_rounds_sub_sBox_PRINCE_6_n9}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, new_AGEMA_signal_2947, Midori_rounds_sub_sBox_PRINCE_6_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U11 ( .a ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, new_AGEMA_signal_2215, Midori_rounds_roundReg_out[24]}), .b ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, new_AGEMA_signal_2953, Midori_rounds_sub_sBox_PRINCE_6_n4}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, new_AGEMA_signal_3379, Midori_rounds_sub_sBox_PRINCE_6_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U6 ( .a ({new_AGEMA_signal_2232, new_AGEMA_signal_2231, new_AGEMA_signal_2230, Midori_rounds_sub_sBox_PRINCE_6_n7}), .b ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, new_AGEMA_signal_2227, Midori_rounds_sub_sBox_PRINCE_6_n1}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, new_AGEMA_signal_2959, Midori_rounds_sub_sBox_PRINCE_6_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U18 ( .a ({new_AGEMA_signal_2982, new_AGEMA_signal_2981, new_AGEMA_signal_2980, Midori_rounds_sub_sBox_PRINCE_7_n13}), .b ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, new_AGEMA_signal_3385, Midori_rounds_roundReg_out[29]}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_3390, new_AGEMA_signal_3389, new_AGEMA_signal_3388, Midori_rounds_sub_sBox_PRINCE_7_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U15 ( .a ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, new_AGEMA_signal_2245, Midori_rounds_sub_sBox_PRINCE_7_n10}), .b ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, new_AGEMA_signal_2260, Midori_rounds_sub_sBox_PRINCE_7_n9}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_2967, new_AGEMA_signal_2966, new_AGEMA_signal_2965, Midori_rounds_sub_sBox_PRINCE_7_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U11 ( .a ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, new_AGEMA_signal_2239, Midori_rounds_roundReg_out[28]}), .b ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, new_AGEMA_signal_2971, Midori_rounds_sub_sBox_PRINCE_7_n4}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_3396, new_AGEMA_signal_3395, new_AGEMA_signal_3394, Midori_rounds_sub_sBox_PRINCE_7_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U6 ( .a ({new_AGEMA_signal_2256, new_AGEMA_signal_2255, new_AGEMA_signal_2254, Midori_rounds_sub_sBox_PRINCE_7_n7}), .b ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, new_AGEMA_signal_2251, Midori_rounds_sub_sBox_PRINCE_7_n1}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_2979, new_AGEMA_signal_2978, new_AGEMA_signal_2977, Midori_rounds_sub_sBox_PRINCE_7_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U18 ( .a ({new_AGEMA_signal_3000, new_AGEMA_signal_2999, new_AGEMA_signal_2998, Midori_rounds_sub_sBox_PRINCE_8_n13}), .b ({new_AGEMA_signal_3402, new_AGEMA_signal_3401, new_AGEMA_signal_3400, Midori_rounds_roundReg_out[33]}), .clk (clk), .r ({Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, new_AGEMA_signal_3403, Midori_rounds_sub_sBox_PRINCE_8_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U15 ( .a ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, new_AGEMA_signal_2269, Midori_rounds_sub_sBox_PRINCE_8_n10}), .b ({new_AGEMA_signal_2286, new_AGEMA_signal_2285, new_AGEMA_signal_2284, Midori_rounds_sub_sBox_PRINCE_8_n9}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774]}), .c ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, new_AGEMA_signal_2983, Midori_rounds_sub_sBox_PRINCE_8_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U11 ( .a ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, new_AGEMA_signal_2263, Midori_rounds_roundReg_out[32]}), .b ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, new_AGEMA_signal_2989, Midori_rounds_sub_sBox_PRINCE_8_n4}), .clk (clk), .r ({Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_3411, new_AGEMA_signal_3410, new_AGEMA_signal_3409, Midori_rounds_sub_sBox_PRINCE_8_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U6 ( .a ({new_AGEMA_signal_2280, new_AGEMA_signal_2279, new_AGEMA_signal_2278, Midori_rounds_sub_sBox_PRINCE_8_n7}), .b ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, new_AGEMA_signal_2275, Midori_rounds_sub_sBox_PRINCE_8_n1}), .clk (clk), .r ({Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786]}), .c ({new_AGEMA_signal_2997, new_AGEMA_signal_2996, new_AGEMA_signal_2995, Midori_rounds_sub_sBox_PRINCE_8_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U18 ( .a ({new_AGEMA_signal_3018, new_AGEMA_signal_3017, new_AGEMA_signal_3016, Midori_rounds_sub_sBox_PRINCE_9_n13}), .b ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, new_AGEMA_signal_3415, Midori_rounds_roundReg_out[37]}), .clk (clk), .r ({Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_3420, new_AGEMA_signal_3419, new_AGEMA_signal_3418, Midori_rounds_sub_sBox_PRINCE_9_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U15 ( .a ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, new_AGEMA_signal_2293, Midori_rounds_sub_sBox_PRINCE_9_n10}), .b ({new_AGEMA_signal_2310, new_AGEMA_signal_2309, new_AGEMA_signal_2308, Midori_rounds_sub_sBox_PRINCE_9_n9}), .clk (clk), .r ({Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798]}), .c ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, new_AGEMA_signal_3001, Midori_rounds_sub_sBox_PRINCE_9_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U11 ( .a ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, new_AGEMA_signal_2287, Midori_rounds_roundReg_out[36]}), .b ({new_AGEMA_signal_3009, new_AGEMA_signal_3008, new_AGEMA_signal_3007, Midori_rounds_sub_sBox_PRINCE_9_n4}), .clk (clk), .r ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_3426, new_AGEMA_signal_3425, new_AGEMA_signal_3424, Midori_rounds_sub_sBox_PRINCE_9_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U6 ( .a ({new_AGEMA_signal_2304, new_AGEMA_signal_2303, new_AGEMA_signal_2302, Midori_rounds_sub_sBox_PRINCE_9_n7}), .b ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, new_AGEMA_signal_2299, Midori_rounds_sub_sBox_PRINCE_9_n1}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .c ({new_AGEMA_signal_3015, new_AGEMA_signal_3014, new_AGEMA_signal_3013, Midori_rounds_sub_sBox_PRINCE_9_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U18 ( .a ({new_AGEMA_signal_3036, new_AGEMA_signal_3035, new_AGEMA_signal_3034, Midori_rounds_sub_sBox_PRINCE_10_n13}), .b ({new_AGEMA_signal_3432, new_AGEMA_signal_3431, new_AGEMA_signal_3430, Midori_rounds_roundReg_out[41]}), .clk (clk), .r ({Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .c ({new_AGEMA_signal_3435, new_AGEMA_signal_3434, new_AGEMA_signal_3433, Midori_rounds_sub_sBox_PRINCE_10_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U15 ( .a ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, new_AGEMA_signal_2317, Midori_rounds_sub_sBox_PRINCE_10_n10}), .b ({new_AGEMA_signal_2334, new_AGEMA_signal_2333, new_AGEMA_signal_2332, Midori_rounds_sub_sBox_PRINCE_10_n9}), .clk (clk), .r ({Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822]}), .c ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, new_AGEMA_signal_3019, Midori_rounds_sub_sBox_PRINCE_10_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U11 ( .a ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, new_AGEMA_signal_2311, Midori_rounds_roundReg_out[40]}), .b ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, new_AGEMA_signal_3025, Midori_rounds_sub_sBox_PRINCE_10_n4}), .clk (clk), .r ({Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828]}), .c ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, new_AGEMA_signal_3439, Midori_rounds_sub_sBox_PRINCE_10_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U6 ( .a ({new_AGEMA_signal_2328, new_AGEMA_signal_2327, new_AGEMA_signal_2326, Midori_rounds_sub_sBox_PRINCE_10_n7}), .b ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, new_AGEMA_signal_2323, Midori_rounds_sub_sBox_PRINCE_10_n1}), .clk (clk), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834]}), .c ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, new_AGEMA_signal_3031, Midori_rounds_sub_sBox_PRINCE_10_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U18 ( .a ({new_AGEMA_signal_3054, new_AGEMA_signal_3053, new_AGEMA_signal_3052, Midori_rounds_sub_sBox_PRINCE_11_n13}), .b ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, new_AGEMA_signal_3445, Midori_rounds_roundReg_out[45]}), .clk (clk), .r ({Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({new_AGEMA_signal_3450, new_AGEMA_signal_3449, new_AGEMA_signal_3448, Midori_rounds_sub_sBox_PRINCE_11_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U15 ( .a ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, new_AGEMA_signal_2341, Midori_rounds_sub_sBox_PRINCE_11_n10}), .b ({new_AGEMA_signal_2358, new_AGEMA_signal_2357, new_AGEMA_signal_2356, Midori_rounds_sub_sBox_PRINCE_11_n9}), .clk (clk), .r ({Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846]}), .c ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, new_AGEMA_signal_3037, Midori_rounds_sub_sBox_PRINCE_11_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U11 ( .a ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, new_AGEMA_signal_2335, Midori_rounds_roundReg_out[44]}), .b ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, new_AGEMA_signal_3043, Midori_rounds_sub_sBox_PRINCE_11_n4}), .clk (clk), .r ({Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852]}), .c ({new_AGEMA_signal_3456, new_AGEMA_signal_3455, new_AGEMA_signal_3454, Midori_rounds_sub_sBox_PRINCE_11_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U6 ( .a ({new_AGEMA_signal_2352, new_AGEMA_signal_2351, new_AGEMA_signal_2350, Midori_rounds_sub_sBox_PRINCE_11_n7}), .b ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, new_AGEMA_signal_2347, Midori_rounds_sub_sBox_PRINCE_11_n1}), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858]}), .c ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, new_AGEMA_signal_3049, Midori_rounds_sub_sBox_PRINCE_11_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U18 ( .a ({new_AGEMA_signal_3072, new_AGEMA_signal_3071, new_AGEMA_signal_3070, Midori_rounds_sub_sBox_PRINCE_12_n13}), .b ({new_AGEMA_signal_3462, new_AGEMA_signal_3461, new_AGEMA_signal_3460, Midori_rounds_roundReg_out[49]}), .clk (clk), .r ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .c ({new_AGEMA_signal_3465, new_AGEMA_signal_3464, new_AGEMA_signal_3463, Midori_rounds_sub_sBox_PRINCE_12_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U15 ( .a ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, new_AGEMA_signal_2365, Midori_rounds_sub_sBox_PRINCE_12_n10}), .b ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, new_AGEMA_signal_2380, Midori_rounds_sub_sBox_PRINCE_12_n9}), .clk (clk), .r ({Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .c ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, new_AGEMA_signal_3055, Midori_rounds_sub_sBox_PRINCE_12_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U11 ( .a ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, new_AGEMA_signal_2359, Midori_rounds_roundReg_out[48]}), .b ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, new_AGEMA_signal_3061, Midori_rounds_sub_sBox_PRINCE_12_n4}), .clk (clk), .r ({Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876]}), .c ({new_AGEMA_signal_3471, new_AGEMA_signal_3470, new_AGEMA_signal_3469, Midori_rounds_sub_sBox_PRINCE_12_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U6 ( .a ({new_AGEMA_signal_2376, new_AGEMA_signal_2375, new_AGEMA_signal_2374, Midori_rounds_sub_sBox_PRINCE_12_n7}), .b ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, new_AGEMA_signal_2371, Midori_rounds_sub_sBox_PRINCE_12_n1}), .clk (clk), .r ({Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882]}), .c ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, new_AGEMA_signal_3067, Midori_rounds_sub_sBox_PRINCE_12_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U18 ( .a ({new_AGEMA_signal_3090, new_AGEMA_signal_3089, new_AGEMA_signal_3088, Midori_rounds_sub_sBox_PRINCE_13_n13}), .b ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, new_AGEMA_signal_3475, Midori_rounds_roundReg_out[53]}), .clk (clk), .r ({Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888]}), .c ({new_AGEMA_signal_3480, new_AGEMA_signal_3479, new_AGEMA_signal_3478, Midori_rounds_sub_sBox_PRINCE_13_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U15 ( .a ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, new_AGEMA_signal_2389, Midori_rounds_sub_sBox_PRINCE_13_n10}), .b ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, new_AGEMA_signal_2404, Midori_rounds_sub_sBox_PRINCE_13_n9}), .clk (clk), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894]}), .c ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, new_AGEMA_signal_3073, Midori_rounds_sub_sBox_PRINCE_13_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U11 ( .a ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, new_AGEMA_signal_2383, Midori_rounds_roundReg_out[52]}), .b ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, new_AGEMA_signal_3079, Midori_rounds_sub_sBox_PRINCE_13_n4}), .clk (clk), .r ({Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({new_AGEMA_signal_3486, new_AGEMA_signal_3485, new_AGEMA_signal_3484, Midori_rounds_sub_sBox_PRINCE_13_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U6 ( .a ({new_AGEMA_signal_2400, new_AGEMA_signal_2399, new_AGEMA_signal_2398, Midori_rounds_sub_sBox_PRINCE_13_n7}), .b ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, new_AGEMA_signal_2395, Midori_rounds_sub_sBox_PRINCE_13_n1}), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906]}), .c ({new_AGEMA_signal_3087, new_AGEMA_signal_3086, new_AGEMA_signal_3085, Midori_rounds_sub_sBox_PRINCE_13_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U18 ( .a ({new_AGEMA_signal_3108, new_AGEMA_signal_3107, new_AGEMA_signal_3106, Midori_rounds_sub_sBox_PRINCE_14_n13}), .b ({new_AGEMA_signal_3492, new_AGEMA_signal_3491, new_AGEMA_signal_3490, Midori_rounds_roundReg_out[57]}), .clk (clk), .r ({Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .c ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, new_AGEMA_signal_3493, Midori_rounds_sub_sBox_PRINCE_14_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U15 ( .a ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, new_AGEMA_signal_2413, Midori_rounds_sub_sBox_PRINCE_14_n10}), .b ({new_AGEMA_signal_2430, new_AGEMA_signal_2429, new_AGEMA_signal_2428, Midori_rounds_sub_sBox_PRINCE_14_n9}), .clk (clk), .r ({Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918]}), .c ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, new_AGEMA_signal_3091, Midori_rounds_sub_sBox_PRINCE_14_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U11 ( .a ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, new_AGEMA_signal_2407, Midori_rounds_roundReg_out[56]}), .b ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, new_AGEMA_signal_3097, Midori_rounds_sub_sBox_PRINCE_14_n4}), .clk (clk), .r ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924]}), .c ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, new_AGEMA_signal_3499, Midori_rounds_sub_sBox_PRINCE_14_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U6 ( .a ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, new_AGEMA_signal_2422, Midori_rounds_sub_sBox_PRINCE_14_n7}), .b ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, new_AGEMA_signal_2419, Midori_rounds_sub_sBox_PRINCE_14_n1}), .clk (clk), .r ({Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .c ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, new_AGEMA_signal_3103, Midori_rounds_sub_sBox_PRINCE_14_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U18 ( .a ({new_AGEMA_signal_3126, new_AGEMA_signal_3125, new_AGEMA_signal_3124, Midori_rounds_sub_sBox_PRINCE_15_n13}), .b ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, new_AGEMA_signal_3505, Midori_rounds_roundReg_out[61]}), .clk (clk), .r ({Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936]}), .c ({new_AGEMA_signal_3510, new_AGEMA_signal_3509, new_AGEMA_signal_3508, Midori_rounds_sub_sBox_PRINCE_15_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U15 ( .a ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, new_AGEMA_signal_2437, Midori_rounds_sub_sBox_PRINCE_15_n10}), .b ({new_AGEMA_signal_2454, new_AGEMA_signal_2453, new_AGEMA_signal_2452, Midori_rounds_sub_sBox_PRINCE_15_n9}), .clk (clk), .r ({Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942]}), .c ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, new_AGEMA_signal_3109, Midori_rounds_sub_sBox_PRINCE_15_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U11 ( .a ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, new_AGEMA_signal_2431, Midori_rounds_roundReg_out[60]}), .b ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, new_AGEMA_signal_3115, Midori_rounds_sub_sBox_PRINCE_15_n4}), .clk (clk), .r ({Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948]}), .c ({new_AGEMA_signal_3516, new_AGEMA_signal_3515, new_AGEMA_signal_3514, Midori_rounds_sub_sBox_PRINCE_15_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U6 ( .a ({new_AGEMA_signal_2448, new_AGEMA_signal_2447, new_AGEMA_signal_2446, Midori_rounds_sub_sBox_PRINCE_15_n7}), .b ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, new_AGEMA_signal_2443, Midori_rounds_sub_sBox_PRINCE_15_n1}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954]}), .c ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, new_AGEMA_signal_3121, Midori_rounds_sub_sBox_PRINCE_15_n2}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U128 ( .a ({new_AGEMA_signal_1464, new_AGEMA_signal_1463, new_AGEMA_signal_1462, wk[9]}), .b ({new_AGEMA_signal_3552, new_AGEMA_signal_3551, new_AGEMA_signal_3550, Midori_rounds_SR_Result[9]}), .c ({DataOut_s3[9], DataOut_s2[9], DataOut_s1[9], DataOut_s0[9]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U126 ( .a ({new_AGEMA_signal_1482, new_AGEMA_signal_1481, new_AGEMA_signal_1480, wk[7]}), .b ({new_AGEMA_signal_3534, new_AGEMA_signal_3533, new_AGEMA_signal_3532, Midori_rounds_SR_Result[47]}), .c ({DataOut_s3[7], DataOut_s2[7], DataOut_s1[7], DataOut_s0[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U124 ( .a ({new_AGEMA_signal_1500, new_AGEMA_signal_1499, new_AGEMA_signal_1498, wk[63]}), .b ({new_AGEMA_signal_3702, new_AGEMA_signal_3701, new_AGEMA_signal_3700, Midori_rounds_SR_Result[63]}), .c ({DataOut_s3[63], DataOut_s2[63], DataOut_s1[63], DataOut_s0[63]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U122 ( .a ({new_AGEMA_signal_1518, new_AGEMA_signal_1517, new_AGEMA_signal_1516, wk[61]}), .b ({new_AGEMA_signal_3708, new_AGEMA_signal_3707, new_AGEMA_signal_3706, Midori_rounds_SR_Result[61]}), .c ({DataOut_s3[61], DataOut_s2[61], DataOut_s1[61], DataOut_s0[61]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U120 ( .a ({new_AGEMA_signal_1536, new_AGEMA_signal_1535, new_AGEMA_signal_1534, wk[5]}), .b ({new_AGEMA_signal_3540, new_AGEMA_signal_3539, new_AGEMA_signal_3538, Midori_rounds_SR_Result[45]}), .c ({DataOut_s3[5], DataOut_s2[5], DataOut_s1[5], DataOut_s0[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U119 ( .a ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, new_AGEMA_signal_1543, wk[59]}), .b ({new_AGEMA_signal_3690, new_AGEMA_signal_3689, new_AGEMA_signal_3688, Midori_rounds_SR_Result[35]}), .c ({DataOut_s3[59], DataOut_s2[59], DataOut_s1[59], DataOut_s0[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U117 ( .a ({new_AGEMA_signal_1563, new_AGEMA_signal_1562, new_AGEMA_signal_1561, wk[57]}), .b ({new_AGEMA_signal_3696, new_AGEMA_signal_3695, new_AGEMA_signal_3694, Midori_rounds_SR_Result[33]}), .c ({DataOut_s3[57], DataOut_s2[57], DataOut_s1[57], DataOut_s0[57]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U115 ( .a ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, new_AGEMA_signal_1579, wk[55]}), .b ({new_AGEMA_signal_3678, new_AGEMA_signal_3677, new_AGEMA_signal_3676, Midori_rounds_SR_Result[7]}), .c ({DataOut_s3[55], DataOut_s2[55], DataOut_s1[55], DataOut_s0[55]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U113 ( .a ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, new_AGEMA_signal_1597, wk[53]}), .b ({new_AGEMA_signal_3684, new_AGEMA_signal_3683, new_AGEMA_signal_3682, Midori_rounds_SR_Result[5]}), .c ({DataOut_s3[53], DataOut_s2[53], DataOut_s1[53], DataOut_s0[53]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U111 ( .a ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, new_AGEMA_signal_1615, wk[51]}), .b ({new_AGEMA_signal_3666, new_AGEMA_signal_3665, new_AGEMA_signal_3664, Midori_rounds_SR_Result[27]}), .c ({DataOut_s3[51], DataOut_s2[51], DataOut_s1[51], DataOut_s0[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U108 ( .a ({new_AGEMA_signal_1644, new_AGEMA_signal_1643, new_AGEMA_signal_1642, wk[49]}), .b ({new_AGEMA_signal_3672, new_AGEMA_signal_3671, new_AGEMA_signal_3670, Midori_rounds_SR_Result[25]}), .c ({DataOut_s3[49], DataOut_s2[49], DataOut_s1[49], DataOut_s0[49]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U106 ( .a ({new_AGEMA_signal_1662, new_AGEMA_signal_1661, new_AGEMA_signal_1660, wk[47]}), .b ({new_AGEMA_signal_3654, new_AGEMA_signal_3653, new_AGEMA_signal_3652, Midori_rounds_SR_Result[43]}), .c ({DataOut_s3[47], DataOut_s2[47], DataOut_s1[47], DataOut_s0[47]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U104 ( .a ({new_AGEMA_signal_1680, new_AGEMA_signal_1679, new_AGEMA_signal_1678, wk[45]}), .b ({new_AGEMA_signal_3660, new_AGEMA_signal_3659, new_AGEMA_signal_3658, Midori_rounds_SR_Result[41]}), .c ({DataOut_s3[45], DataOut_s2[45], DataOut_s1[45], DataOut_s0[45]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U102 ( .a ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, new_AGEMA_signal_1696, wk[43]}), .b ({new_AGEMA_signal_3642, new_AGEMA_signal_3641, new_AGEMA_signal_3640, Midori_rounds_SR_Result[55]}), .c ({DataOut_s3[43], DataOut_s2[43], DataOut_s1[43], DataOut_s0[43]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U100 ( .a ({new_AGEMA_signal_1716, new_AGEMA_signal_1715, new_AGEMA_signal_1714, wk[41]}), .b ({new_AGEMA_signal_3648, new_AGEMA_signal_3647, new_AGEMA_signal_3646, Midori_rounds_SR_Result[53]}), .c ({DataOut_s3[41], DataOut_s2[41], DataOut_s1[41], DataOut_s0[41]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U98 ( .a ({new_AGEMA_signal_1734, new_AGEMA_signal_1733, new_AGEMA_signal_1732, wk[3]}), .b ({new_AGEMA_signal_3522, new_AGEMA_signal_3521, new_AGEMA_signal_3520, Midori_rounds_SR_Result[51]}), .c ({DataOut_s3[3], DataOut_s2[3], DataOut_s1[3], DataOut_s0[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U97 ( .a ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, new_AGEMA_signal_1741, wk[39]}), .b ({new_AGEMA_signal_3630, new_AGEMA_signal_3629, new_AGEMA_signal_3628, Midori_rounds_SR_Result[19]}), .c ({DataOut_s3[39], DataOut_s2[39], DataOut_s1[39], DataOut_s0[39]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U95 ( .a ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, new_AGEMA_signal_1759, wk[37]}), .b ({new_AGEMA_signal_3636, new_AGEMA_signal_3635, new_AGEMA_signal_3634, Midori_rounds_SR_Result[17]}), .c ({DataOut_s3[37], DataOut_s2[37], DataOut_s1[37], DataOut_s0[37]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U93 ( .a ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, new_AGEMA_signal_1777, wk[35]}), .b ({new_AGEMA_signal_3618, new_AGEMA_signal_3617, new_AGEMA_signal_3616, Midori_rounds_SR_Result[15]}), .c ({DataOut_s3[35], DataOut_s2[35], DataOut_s1[35], DataOut_s0[35]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U91 ( .a ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, new_AGEMA_signal_1795, wk[33]}), .b ({new_AGEMA_signal_3624, new_AGEMA_signal_3623, new_AGEMA_signal_3622, Midori_rounds_SR_Result[13]}), .c ({DataOut_s3[33], DataOut_s2[33], DataOut_s1[33], DataOut_s0[33]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U89 ( .a ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, new_AGEMA_signal_1813, wk[31]}), .b ({new_AGEMA_signal_3606, new_AGEMA_signal_3605, new_AGEMA_signal_3604, Midori_rounds_SR_Result[3]}), .c ({DataOut_s3[31], DataOut_s2[31], DataOut_s1[31], DataOut_s0[31]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U86 ( .a ({new_AGEMA_signal_1842, new_AGEMA_signal_1841, new_AGEMA_signal_1840, wk[29]}), .b ({new_AGEMA_signal_3612, new_AGEMA_signal_3611, new_AGEMA_signal_3610, Midori_rounds_SR_Result[1]}), .c ({DataOut_s3[29], DataOut_s2[29], DataOut_s1[29], DataOut_s0[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U84 ( .a ({new_AGEMA_signal_1860, new_AGEMA_signal_1859, new_AGEMA_signal_1858, wk[27]}), .b ({new_AGEMA_signal_3594, new_AGEMA_signal_3593, new_AGEMA_signal_3592, Midori_rounds_SR_Result[31]}), .c ({DataOut_s3[27], DataOut_s2[27], DataOut_s1[27], DataOut_s0[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U82 ( .a ({new_AGEMA_signal_1878, new_AGEMA_signal_1877, new_AGEMA_signal_1876, wk[25]}), .b ({new_AGEMA_signal_3600, new_AGEMA_signal_3599, new_AGEMA_signal_3598, Midori_rounds_SR_Result[29]}), .c ({DataOut_s3[25], DataOut_s2[25], DataOut_s1[25], DataOut_s0[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U80 ( .a ({new_AGEMA_signal_1896, new_AGEMA_signal_1895, new_AGEMA_signal_1894, wk[23]}), .b ({new_AGEMA_signal_3582, new_AGEMA_signal_3581, new_AGEMA_signal_3580, Midori_rounds_SR_Result[59]}), .c ({DataOut_s3[23], DataOut_s2[23], DataOut_s1[23], DataOut_s0[23]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U78 ( .a ({new_AGEMA_signal_1914, new_AGEMA_signal_1913, new_AGEMA_signal_1912, wk[21]}), .b ({new_AGEMA_signal_3588, new_AGEMA_signal_3587, new_AGEMA_signal_3586, Midori_rounds_SR_Result[57]}), .c ({DataOut_s3[21], DataOut_s2[21], DataOut_s1[21], DataOut_s0[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U76 ( .a ({new_AGEMA_signal_1932, new_AGEMA_signal_1931, new_AGEMA_signal_1930, wk[1]}), .b ({new_AGEMA_signal_3528, new_AGEMA_signal_3527, new_AGEMA_signal_3526, Midori_rounds_SR_Result[49]}), .c ({DataOut_s3[1], DataOut_s2[1], DataOut_s1[1], DataOut_s0[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U75 ( .a ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, new_AGEMA_signal_1939, wk[19]}), .b ({new_AGEMA_signal_3570, new_AGEMA_signal_3569, new_AGEMA_signal_3568, Midori_rounds_SR_Result[39]}), .c ({DataOut_s3[19], DataOut_s2[19], DataOut_s1[19], DataOut_s0[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U73 ( .a ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, new_AGEMA_signal_1957, wk[17]}), .b ({new_AGEMA_signal_3576, new_AGEMA_signal_3575, new_AGEMA_signal_3574, Midori_rounds_SR_Result[37]}), .c ({DataOut_s3[17], DataOut_s2[17], DataOut_s1[17], DataOut_s0[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U71 ( .a ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, new_AGEMA_signal_1975, wk[15]}), .b ({new_AGEMA_signal_3558, new_AGEMA_signal_3557, new_AGEMA_signal_3556, Midori_rounds_SR_Result[23]}), .c ({DataOut_s3[15], DataOut_s2[15], DataOut_s1[15], DataOut_s0[15]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U69 ( .a ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, new_AGEMA_signal_1993, wk[13]}), .b ({new_AGEMA_signal_3564, new_AGEMA_signal_3563, new_AGEMA_signal_3562, Midori_rounds_SR_Result[21]}), .c ({DataOut_s3[13], DataOut_s2[13], DataOut_s1[13], DataOut_s0[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U67 ( .a ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, new_AGEMA_signal_2011, wk[11]}), .b ({new_AGEMA_signal_3546, new_AGEMA_signal_3545, new_AGEMA_signal_3544, Midori_rounds_SR_Result[11]}), .c ({DataOut_s3[11], DataOut_s2[11], DataOut_s1[11], DataOut_s0[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U144 ( .a ({new_AGEMA_signal_2052, new_AGEMA_signal_2051, new_AGEMA_signal_2050, Midori_rounds_SelectedKey_9_}), .b ({new_AGEMA_signal_3552, new_AGEMA_signal_3551, new_AGEMA_signal_3550, Midori_rounds_SR_Result[9]}), .c ({new_AGEMA_signal_3906, new_AGEMA_signal_3905, new_AGEMA_signal_3904, Midori_rounds_sub_ResultXORkey[9]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U142 ( .a ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, new_AGEMA_signal_3133, Midori_rounds_SelectedKey_7_}), .b ({new_AGEMA_signal_3534, new_AGEMA_signal_3533, new_AGEMA_signal_3532, Midori_rounds_SR_Result[47]}), .c ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, new_AGEMA_signal_3907, Midori_rounds_sub_ResultXORkey[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U140 ( .a ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, new_AGEMA_signal_3277, Midori_rounds_SelectedKey_63_}), .b ({new_AGEMA_signal_3702, new_AGEMA_signal_3701, new_AGEMA_signal_3700, Midori_rounds_SR_Result[63]}), .c ({new_AGEMA_signal_3915, new_AGEMA_signal_3914, new_AGEMA_signal_3913, Midori_rounds_sub_ResultXORkey[63]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U138 ( .a ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, new_AGEMA_signal_3271, Midori_rounds_SelectedKey_61_}), .b ({new_AGEMA_signal_3708, new_AGEMA_signal_3707, new_AGEMA_signal_3706, Midori_rounds_SR_Result[61]}), .c ({new_AGEMA_signal_3921, new_AGEMA_signal_3920, new_AGEMA_signal_3919, Midori_rounds_sub_ResultXORkey[61]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U136 ( .a ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, new_AGEMA_signal_3127, Midori_rounds_SelectedKey_5_}), .b ({new_AGEMA_signal_3540, new_AGEMA_signal_3539, new_AGEMA_signal_3538, Midori_rounds_SR_Result[45]}), .c ({new_AGEMA_signal_3924, new_AGEMA_signal_3923, new_AGEMA_signal_3922, Midori_rounds_sub_ResultXORkey[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U135 ( .a ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, new_AGEMA_signal_3265, Midori_rounds_SelectedKey_59_}), .b ({new_AGEMA_signal_3690, new_AGEMA_signal_3689, new_AGEMA_signal_3688, Midori_rounds_SR_Result[35]}), .c ({new_AGEMA_signal_3927, new_AGEMA_signal_3926, new_AGEMA_signal_3925, Midori_rounds_sub_ResultXORkey[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U133 ( .a ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, new_AGEMA_signal_3259, Midori_rounds_SelectedKey_57_}), .b ({new_AGEMA_signal_3696, new_AGEMA_signal_3695, new_AGEMA_signal_3694, Midori_rounds_SR_Result[33]}), .c ({new_AGEMA_signal_3933, new_AGEMA_signal_3932, new_AGEMA_signal_3931, Midori_rounds_sub_ResultXORkey[57]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U131 ( .a ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, new_AGEMA_signal_3253, Midori_rounds_SelectedKey_55_}), .b ({new_AGEMA_signal_3678, new_AGEMA_signal_3677, new_AGEMA_signal_3676, Midori_rounds_SR_Result[7]}), .c ({new_AGEMA_signal_3936, new_AGEMA_signal_3935, new_AGEMA_signal_3934, Midori_rounds_sub_ResultXORkey[55]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U129 ( .a ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, new_AGEMA_signal_3247, Midori_rounds_SelectedKey_53_}), .b ({new_AGEMA_signal_3684, new_AGEMA_signal_3683, new_AGEMA_signal_3682, Midori_rounds_SR_Result[5]}), .c ({new_AGEMA_signal_3942, new_AGEMA_signal_3941, new_AGEMA_signal_3940, Midori_rounds_sub_ResultXORkey[53]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U127 ( .a ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, new_AGEMA_signal_3241, Midori_rounds_SelectedKey_51_}), .b ({new_AGEMA_signal_3666, new_AGEMA_signal_3665, new_AGEMA_signal_3664, Midori_rounds_SR_Result[27]}), .c ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, new_AGEMA_signal_3943, Midori_rounds_sub_ResultXORkey[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U124 ( .a ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, new_AGEMA_signal_3235, Midori_rounds_SelectedKey_49_}), .b ({new_AGEMA_signal_3672, new_AGEMA_signal_3671, new_AGEMA_signal_3670, Midori_rounds_SR_Result[25]}), .c ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, new_AGEMA_signal_3949, Midori_rounds_sub_ResultXORkey[49]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U122 ( .a ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, new_AGEMA_signal_3229, Midori_rounds_SelectedKey_47_}), .b ({new_AGEMA_signal_3654, new_AGEMA_signal_3653, new_AGEMA_signal_3652, Midori_rounds_SR_Result[43]}), .c ({new_AGEMA_signal_3954, new_AGEMA_signal_3953, new_AGEMA_signal_3952, Midori_rounds_sub_ResultXORkey[47]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U120 ( .a ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, new_AGEMA_signal_3223, Midori_rounds_SelectedKey_45_}), .b ({new_AGEMA_signal_3660, new_AGEMA_signal_3659, new_AGEMA_signal_3658, Midori_rounds_SR_Result[41]}), .c ({new_AGEMA_signal_3960, new_AGEMA_signal_3959, new_AGEMA_signal_3958, Midori_rounds_sub_ResultXORkey[45]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U118 ( .a ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, new_AGEMA_signal_3217, Midori_rounds_SelectedKey_43_}), .b ({new_AGEMA_signal_3642, new_AGEMA_signal_3641, new_AGEMA_signal_3640, Midori_rounds_SR_Result[55]}), .c ({new_AGEMA_signal_3963, new_AGEMA_signal_3962, new_AGEMA_signal_3961, Midori_rounds_sub_ResultXORkey[43]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U116 ( .a ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, new_AGEMA_signal_3211, Midori_rounds_SelectedKey_41_}), .b ({new_AGEMA_signal_3648, new_AGEMA_signal_3647, new_AGEMA_signal_3646, Midori_rounds_SR_Result[53]}), .c ({new_AGEMA_signal_3969, new_AGEMA_signal_3968, new_AGEMA_signal_3967, Midori_rounds_sub_ResultXORkey[41]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U114 ( .a ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, new_AGEMA_signal_2041, Midori_rounds_SelectedKey_3_}), .b ({new_AGEMA_signal_3522, new_AGEMA_signal_3521, new_AGEMA_signal_3520, Midori_rounds_SR_Result[51]}), .c ({new_AGEMA_signal_3972, new_AGEMA_signal_3971, new_AGEMA_signal_3970, Midori_rounds_sub_ResultXORkey[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U113 ( .a ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, new_AGEMA_signal_3205, Midori_rounds_SelectedKey_39_}), .b ({new_AGEMA_signal_3630, new_AGEMA_signal_3629, new_AGEMA_signal_3628, Midori_rounds_SR_Result[19]}), .c ({new_AGEMA_signal_3975, new_AGEMA_signal_3974, new_AGEMA_signal_3973, Midori_rounds_sub_ResultXORkey[39]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U111 ( .a ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, new_AGEMA_signal_3199, Midori_rounds_SelectedKey_37_}), .b ({new_AGEMA_signal_3636, new_AGEMA_signal_3635, new_AGEMA_signal_3634, Midori_rounds_SR_Result[17]}), .c ({new_AGEMA_signal_3981, new_AGEMA_signal_3980, new_AGEMA_signal_3979, Midori_rounds_sub_ResultXORkey[37]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U109 ( .a ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, new_AGEMA_signal_3193, Midori_rounds_SelectedKey_35_}), .b ({new_AGEMA_signal_3618, new_AGEMA_signal_3617, new_AGEMA_signal_3616, Midori_rounds_SR_Result[15]}), .c ({new_AGEMA_signal_3984, new_AGEMA_signal_3983, new_AGEMA_signal_3982, Midori_rounds_sub_ResultXORkey[35]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U107 ( .a ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, new_AGEMA_signal_3187, Midori_rounds_SelectedKey_33_}), .b ({new_AGEMA_signal_3624, new_AGEMA_signal_3623, new_AGEMA_signal_3622, Midori_rounds_SR_Result[13]}), .c ({new_AGEMA_signal_3990, new_AGEMA_signal_3989, new_AGEMA_signal_3988, Midori_rounds_sub_ResultXORkey[33]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U105 ( .a ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, new_AGEMA_signal_3181, Midori_rounds_SelectedKey_31_}), .b ({new_AGEMA_signal_3606, new_AGEMA_signal_3605, new_AGEMA_signal_3604, Midori_rounds_SR_Result[3]}), .c ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, new_AGEMA_signal_3991, Midori_rounds_sub_ResultXORkey[31]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U102 ( .a ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, new_AGEMA_signal_3175, Midori_rounds_SelectedKey_29_}), .b ({new_AGEMA_signal_3612, new_AGEMA_signal_3611, new_AGEMA_signal_3610, Midori_rounds_SR_Result[1]}), .c ({new_AGEMA_signal_4002, new_AGEMA_signal_4001, new_AGEMA_signal_4000, Midori_rounds_sub_ResultXORkey[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U100 ( .a ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, new_AGEMA_signal_3169, Midori_rounds_SelectedKey_27_}), .b ({new_AGEMA_signal_3594, new_AGEMA_signal_3593, new_AGEMA_signal_3592, Midori_rounds_SR_Result[31]}), .c ({new_AGEMA_signal_4005, new_AGEMA_signal_4004, new_AGEMA_signal_4003, Midori_rounds_sub_ResultXORkey[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U98 ( .a ({new_AGEMA_signal_3168, new_AGEMA_signal_3167, new_AGEMA_signal_3166, Midori_rounds_SelectedKey_25_}), .b ({new_AGEMA_signal_3600, new_AGEMA_signal_3599, new_AGEMA_signal_3598, Midori_rounds_SR_Result[29]}), .c ({new_AGEMA_signal_4011, new_AGEMA_signal_4010, new_AGEMA_signal_4009, Midori_rounds_sub_ResultXORkey[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U96 ( .a ({new_AGEMA_signal_3162, new_AGEMA_signal_3161, new_AGEMA_signal_3160, Midori_rounds_SelectedKey_23_}), .b ({new_AGEMA_signal_3582, new_AGEMA_signal_3581, new_AGEMA_signal_3580, Midori_rounds_SR_Result[59]}), .c ({new_AGEMA_signal_4014, new_AGEMA_signal_4013, new_AGEMA_signal_4012, Midori_rounds_sub_ResultXORkey[23]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U94 ( .a ({new_AGEMA_signal_3156, new_AGEMA_signal_3155, new_AGEMA_signal_3154, Midori_rounds_SelectedKey_21_}), .b ({new_AGEMA_signal_3588, new_AGEMA_signal_3587, new_AGEMA_signal_3586, Midori_rounds_SR_Result[57]}), .c ({new_AGEMA_signal_4020, new_AGEMA_signal_4019, new_AGEMA_signal_4018, Midori_rounds_sub_ResultXORkey[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U92 ( .a ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, new_AGEMA_signal_2035, Midori_rounds_SelectedKey_1_}), .b ({new_AGEMA_signal_3528, new_AGEMA_signal_3527, new_AGEMA_signal_3526, Midori_rounds_SR_Result[49]}), .c ({new_AGEMA_signal_4023, new_AGEMA_signal_4022, new_AGEMA_signal_4021, Midori_rounds_sub_ResultXORkey[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U91 ( .a ({new_AGEMA_signal_3150, new_AGEMA_signal_3149, new_AGEMA_signal_3148, Midori_rounds_SelectedKey_19_}), .b ({new_AGEMA_signal_3570, new_AGEMA_signal_3569, new_AGEMA_signal_3568, Midori_rounds_SR_Result[39]}), .c ({new_AGEMA_signal_4026, new_AGEMA_signal_4025, new_AGEMA_signal_4024, Midori_rounds_sub_ResultXORkey[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U89 ( .a ({new_AGEMA_signal_3144, new_AGEMA_signal_3143, new_AGEMA_signal_3142, Midori_rounds_SelectedKey_17_}), .b ({new_AGEMA_signal_3576, new_AGEMA_signal_3575, new_AGEMA_signal_3574, Midori_rounds_SR_Result[37]}), .c ({new_AGEMA_signal_4032, new_AGEMA_signal_4031, new_AGEMA_signal_4030, Midori_rounds_sub_ResultXORkey[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U87 ( .a ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, new_AGEMA_signal_2065, Midori_rounds_SelectedKey_15_}), .b ({new_AGEMA_signal_3558, new_AGEMA_signal_3557, new_AGEMA_signal_3556, Midori_rounds_SR_Result[23]}), .c ({new_AGEMA_signal_4035, new_AGEMA_signal_4034, new_AGEMA_signal_4033, Midori_rounds_sub_ResultXORkey[15]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U85 ( .a ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, new_AGEMA_signal_2059, Midori_rounds_SelectedKey_13_}), .b ({new_AGEMA_signal_3564, new_AGEMA_signal_3563, new_AGEMA_signal_3562, Midori_rounds_SR_Result[21]}), .c ({new_AGEMA_signal_4041, new_AGEMA_signal_4040, new_AGEMA_signal_4039, Midori_rounds_sub_ResultXORkey[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U83 ( .a ({new_AGEMA_signal_2058, new_AGEMA_signal_2057, new_AGEMA_signal_2056, Midori_rounds_SelectedKey_11_}), .b ({new_AGEMA_signal_3546, new_AGEMA_signal_3545, new_AGEMA_signal_3544, Midori_rounds_SR_Result[11]}), .c ({new_AGEMA_signal_4044, new_AGEMA_signal_4043, new_AGEMA_signal_4042, Midori_rounds_sub_ResultXORkey[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U80 ( .a ({new_AGEMA_signal_2052, new_AGEMA_signal_2051, new_AGEMA_signal_2050, Midori_rounds_SelectedKey_9_}), .b ({new_AGEMA_signal_4374, new_AGEMA_signal_4373, new_AGEMA_signal_4372, Midori_rounds_SR_Inv_Result[9]}), .c ({new_AGEMA_signal_4410, new_AGEMA_signal_4409, new_AGEMA_signal_4408, Midori_rounds_mul_ResultXORkey[9]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U77 ( .a ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, new_AGEMA_signal_3133, Midori_rounds_SelectedKey_7_}), .b ({new_AGEMA_signal_4377, new_AGEMA_signal_4376, new_AGEMA_signal_4375, Midori_rounds_SR_Inv_Result[55]}), .c ({new_AGEMA_signal_4416, new_AGEMA_signal_4415, new_AGEMA_signal_4414, Midori_rounds_mul_ResultXORkey[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U75 ( .a ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, new_AGEMA_signal_3277, Midori_rounds_SelectedKey_63_}), .b ({new_AGEMA_signal_4287, new_AGEMA_signal_4286, new_AGEMA_signal_4285, Midori_rounds_SR_Inv_Result[63]}), .c ({new_AGEMA_signal_4422, new_AGEMA_signal_4421, new_AGEMA_signal_4420, Midori_rounds_mul_ResultXORkey[63]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U73 ( .a ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, new_AGEMA_signal_3271, Midori_rounds_SelectedKey_61_}), .b ({new_AGEMA_signal_4293, new_AGEMA_signal_4292, new_AGEMA_signal_4291, Midori_rounds_SR_Inv_Result[61]}), .c ({new_AGEMA_signal_4428, new_AGEMA_signal_4427, new_AGEMA_signal_4426, Midori_rounds_mul_ResultXORkey[61]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U70 ( .a ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, new_AGEMA_signal_3127, Midori_rounds_SelectedKey_5_}), .b ({new_AGEMA_signal_4383, new_AGEMA_signal_4382, new_AGEMA_signal_4381, Midori_rounds_SR_Inv_Result[53]}), .c ({new_AGEMA_signal_4431, new_AGEMA_signal_4430, new_AGEMA_signal_4429, Midori_rounds_mul_ResultXORkey[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U69 ( .a ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, new_AGEMA_signal_3265, Midori_rounds_SelectedKey_59_}), .b ({new_AGEMA_signal_4296, new_AGEMA_signal_4295, new_AGEMA_signal_4294, Midori_rounds_SR_Inv_Result[23]}), .c ({new_AGEMA_signal_4434, new_AGEMA_signal_4433, new_AGEMA_signal_4432, Midori_rounds_mul_ResultXORkey[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U67 ( .a ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, new_AGEMA_signal_3259, Midori_rounds_SelectedKey_57_}), .b ({new_AGEMA_signal_4266, new_AGEMA_signal_4265, new_AGEMA_signal_4264, Midori_rounds_SR_Inv_Result[21]}), .c ({new_AGEMA_signal_4440, new_AGEMA_signal_4439, new_AGEMA_signal_4438, Midori_rounds_mul_ResultXORkey[57]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U64 ( .a ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, new_AGEMA_signal_3253, Midori_rounds_SelectedKey_55_}), .b ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, new_AGEMA_signal_4267, Midori_rounds_SR_Inv_Result[43]}), .c ({new_AGEMA_signal_4443, new_AGEMA_signal_4442, new_AGEMA_signal_4441, Midori_rounds_mul_ResultXORkey[55]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U62 ( .a ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, new_AGEMA_signal_3247, Midori_rounds_SelectedKey_53_}), .b ({new_AGEMA_signal_4275, new_AGEMA_signal_4274, new_AGEMA_signal_4273, Midori_rounds_SR_Inv_Result[41]}), .c ({new_AGEMA_signal_4449, new_AGEMA_signal_4448, new_AGEMA_signal_4447, Midori_rounds_mul_ResultXORkey[53]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U59 ( .a ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, new_AGEMA_signal_3241, Midori_rounds_SelectedKey_51_}), .b ({new_AGEMA_signal_4278, new_AGEMA_signal_4277, new_AGEMA_signal_4276, Midori_rounds_SR_Inv_Result[3]}), .c ({new_AGEMA_signal_4452, new_AGEMA_signal_4451, new_AGEMA_signal_4450, Midori_rounds_mul_ResultXORkey[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U55 ( .a ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, new_AGEMA_signal_3235, Midori_rounds_SelectedKey_49_}), .b ({new_AGEMA_signal_4284, new_AGEMA_signal_4283, new_AGEMA_signal_4282, Midori_rounds_SR_Inv_Result[1]}), .c ({new_AGEMA_signal_4458, new_AGEMA_signal_4457, new_AGEMA_signal_4456, Midori_rounds_mul_ResultXORkey[49]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U52 ( .a ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, new_AGEMA_signal_3229, Midori_rounds_SelectedKey_47_}), .b ({new_AGEMA_signal_4323, new_AGEMA_signal_4322, new_AGEMA_signal_4321, Midori_rounds_SR_Inv_Result[7]}), .c ({new_AGEMA_signal_4461, new_AGEMA_signal_4460, new_AGEMA_signal_4459, Midori_rounds_mul_ResultXORkey[47]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U50 ( .a ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, new_AGEMA_signal_3223, Midori_rounds_SelectedKey_45_}), .b ({new_AGEMA_signal_4329, new_AGEMA_signal_4328, new_AGEMA_signal_4327, Midori_rounds_SR_Inv_Result[5]}), .c ({new_AGEMA_signal_4467, new_AGEMA_signal_4466, new_AGEMA_signal_4465, Midori_rounds_mul_ResultXORkey[45]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U47 ( .a ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, new_AGEMA_signal_3217, Midori_rounds_SelectedKey_43_}), .b ({new_AGEMA_signal_4332, new_AGEMA_signal_4331, new_AGEMA_signal_4330, Midori_rounds_SR_Inv_Result[47]}), .c ({new_AGEMA_signal_4473, new_AGEMA_signal_4472, new_AGEMA_signal_4471, Midori_rounds_mul_ResultXORkey[43]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U45 ( .a ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, new_AGEMA_signal_3211, Midori_rounds_SelectedKey_41_}), .b ({new_AGEMA_signal_4302, new_AGEMA_signal_4301, new_AGEMA_signal_4300, Midori_rounds_SR_Inv_Result[45]}), .c ({new_AGEMA_signal_4479, new_AGEMA_signal_4478, new_AGEMA_signal_4477, Midori_rounds_mul_ResultXORkey[41]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U42 ( .a ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, new_AGEMA_signal_2041, Midori_rounds_SelectedKey_3_}), .b ({new_AGEMA_signal_4386, new_AGEMA_signal_4385, new_AGEMA_signal_4384, Midori_rounds_SR_Inv_Result[31]}), .c ({new_AGEMA_signal_4482, new_AGEMA_signal_4481, new_AGEMA_signal_4480, Midori_rounds_mul_ResultXORkey[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U41 ( .a ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, new_AGEMA_signal_3205, Midori_rounds_SelectedKey_39_}), .b ({new_AGEMA_signal_4305, new_AGEMA_signal_4304, new_AGEMA_signal_4303, Midori_rounds_SR_Inv_Result[19]}), .c ({new_AGEMA_signal_4485, new_AGEMA_signal_4484, new_AGEMA_signal_4483, Midori_rounds_mul_ResultXORkey[39]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U39 ( .a ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, new_AGEMA_signal_3199, Midori_rounds_SelectedKey_37_}), .b ({new_AGEMA_signal_4311, new_AGEMA_signal_4310, new_AGEMA_signal_4309, Midori_rounds_SR_Inv_Result[17]}), .c ({new_AGEMA_signal_4491, new_AGEMA_signal_4490, new_AGEMA_signal_4489, Midori_rounds_mul_ResultXORkey[37]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U36 ( .a ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, new_AGEMA_signal_3193, Midori_rounds_SelectedKey_35_}), .b ({new_AGEMA_signal_4314, new_AGEMA_signal_4313, new_AGEMA_signal_4312, Midori_rounds_SR_Inv_Result[59]}), .c ({new_AGEMA_signal_4497, new_AGEMA_signal_4496, new_AGEMA_signal_4495, Midori_rounds_mul_ResultXORkey[35]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U34 ( .a ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, new_AGEMA_signal_3187, Midori_rounds_SelectedKey_33_}), .b ({new_AGEMA_signal_4320, new_AGEMA_signal_4319, new_AGEMA_signal_4318, Midori_rounds_SR_Inv_Result[57]}), .c ({new_AGEMA_signal_4503, new_AGEMA_signal_4502, new_AGEMA_signal_4501, Midori_rounds_mul_ResultXORkey[33]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U31 ( .a ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, new_AGEMA_signal_3181, Midori_rounds_SelectedKey_31_}), .b ({new_AGEMA_signal_4359, new_AGEMA_signal_4358, new_AGEMA_signal_4357, Midori_rounds_SR_Inv_Result[27]}), .c ({new_AGEMA_signal_4506, new_AGEMA_signal_4505, new_AGEMA_signal_4504, Midori_rounds_mul_ResultXORkey[31]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U28 ( .a ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, new_AGEMA_signal_3175, Midori_rounds_SelectedKey_29_}), .b ({new_AGEMA_signal_4365, new_AGEMA_signal_4364, new_AGEMA_signal_4363, Midori_rounds_SR_Inv_Result[25]}), .c ({new_AGEMA_signal_4515, new_AGEMA_signal_4514, new_AGEMA_signal_4513, Midori_rounds_mul_ResultXORkey[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U25 ( .a ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, new_AGEMA_signal_3169, Midori_rounds_SelectedKey_27_}), .b ({new_AGEMA_signal_4368, new_AGEMA_signal_4367, new_AGEMA_signal_4366, Midori_rounds_SR_Inv_Result[51]}), .c ({new_AGEMA_signal_4518, new_AGEMA_signal_4517, new_AGEMA_signal_4516, Midori_rounds_mul_ResultXORkey[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U23 ( .a ({new_AGEMA_signal_3168, new_AGEMA_signal_3167, new_AGEMA_signal_3166, Midori_rounds_SelectedKey_25_}), .b ({new_AGEMA_signal_4338, new_AGEMA_signal_4337, new_AGEMA_signal_4336, Midori_rounds_SR_Inv_Result[49]}), .c ({new_AGEMA_signal_4524, new_AGEMA_signal_4523, new_AGEMA_signal_4522, Midori_rounds_mul_ResultXORkey[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U20 ( .a ({new_AGEMA_signal_3162, new_AGEMA_signal_3161, new_AGEMA_signal_3160, Midori_rounds_SelectedKey_23_}), .b ({new_AGEMA_signal_4341, new_AGEMA_signal_4340, new_AGEMA_signal_4339, Midori_rounds_SR_Inv_Result[15]}), .c ({new_AGEMA_signal_4527, new_AGEMA_signal_4526, new_AGEMA_signal_4525, Midori_rounds_mul_ResultXORkey[23]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U18 ( .a ({new_AGEMA_signal_3156, new_AGEMA_signal_3155, new_AGEMA_signal_3154, Midori_rounds_SelectedKey_21_}), .b ({new_AGEMA_signal_4347, new_AGEMA_signal_4346, new_AGEMA_signal_4345, Midori_rounds_SR_Inv_Result[13]}), .c ({new_AGEMA_signal_4533, new_AGEMA_signal_4532, new_AGEMA_signal_4531, Midori_rounds_mul_ResultXORkey[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U15 ( .a ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, new_AGEMA_signal_2035, Midori_rounds_SelectedKey_1_}), .b ({new_AGEMA_signal_4392, new_AGEMA_signal_4391, new_AGEMA_signal_4390, Midori_rounds_SR_Inv_Result[29]}), .c ({new_AGEMA_signal_4539, new_AGEMA_signal_4538, new_AGEMA_signal_4537, Midori_rounds_mul_ResultXORkey[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U14 ( .a ({new_AGEMA_signal_3150, new_AGEMA_signal_3149, new_AGEMA_signal_3148, Midori_rounds_SelectedKey_19_}), .b ({new_AGEMA_signal_4350, new_AGEMA_signal_4349, new_AGEMA_signal_4348, Midori_rounds_SR_Inv_Result[39]}), .c ({new_AGEMA_signal_4542, new_AGEMA_signal_4541, new_AGEMA_signal_4540, Midori_rounds_mul_ResultXORkey[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U12 ( .a ({new_AGEMA_signal_3144, new_AGEMA_signal_3143, new_AGEMA_signal_3142, Midori_rounds_SelectedKey_17_}), .b ({new_AGEMA_signal_4356, new_AGEMA_signal_4355, new_AGEMA_signal_4354, Midori_rounds_SR_Inv_Result[37]}), .c ({new_AGEMA_signal_4548, new_AGEMA_signal_4547, new_AGEMA_signal_4546, Midori_rounds_mul_ResultXORkey[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U9 ( .a ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, new_AGEMA_signal_2065, Midori_rounds_SelectedKey_15_}), .b ({new_AGEMA_signal_4395, new_AGEMA_signal_4394, new_AGEMA_signal_4393, Midori_rounds_SR_Inv_Result[35]}), .c ({new_AGEMA_signal_4551, new_AGEMA_signal_4550, new_AGEMA_signal_4549, Midori_rounds_mul_ResultXORkey[15]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U7 ( .a ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, new_AGEMA_signal_2059, Midori_rounds_SelectedKey_13_}), .b ({new_AGEMA_signal_4401, new_AGEMA_signal_4400, new_AGEMA_signal_4399, Midori_rounds_SR_Inv_Result[33]}), .c ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, new_AGEMA_signal_4555, Midori_rounds_mul_ResultXORkey[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U4 ( .a ({new_AGEMA_signal_2058, new_AGEMA_signal_2057, new_AGEMA_signal_2056, Midori_rounds_SelectedKey_11_}), .b ({new_AGEMA_signal_4404, new_AGEMA_signal_4403, new_AGEMA_signal_4402, Midori_rounds_SR_Inv_Result[11]}), .c ({new_AGEMA_signal_4560, new_AGEMA_signal_4559, new_AGEMA_signal_4558, Midori_rounds_mul_ResultXORkey[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4608, new_AGEMA_signal_4607, new_AGEMA_signal_4606, Midori_rounds_round_Result[1]}), .a ({new_AGEMA_signal_2772, new_AGEMA_signal_2771, new_AGEMA_signal_2770, Midori_add_Result_Start[1]}), .c ({new_AGEMA_signal_4785, new_AGEMA_signal_4784, new_AGEMA_signal_4783, Midori_rounds_roundResult_Reg_SFF_1_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4614, new_AGEMA_signal_4613, new_AGEMA_signal_4612, Midori_rounds_round_Result[3]}), .a ({new_AGEMA_signal_2640, new_AGEMA_signal_2639, new_AGEMA_signal_2638, Midori_add_Result_Start[3]}), .c ({new_AGEMA_signal_4791, new_AGEMA_signal_4790, new_AGEMA_signal_4789, Midori_rounds_roundResult_Reg_SFF_3_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4617, new_AGEMA_signal_4616, new_AGEMA_signal_4615, Midori_rounds_round_Result[5]}), .a ({new_AGEMA_signal_2508, new_AGEMA_signal_2507, new_AGEMA_signal_2506, Midori_add_Result_Start[5]}), .c ({new_AGEMA_signal_4794, new_AGEMA_signal_4793, new_AGEMA_signal_4792, Midori_rounds_roundResult_Reg_SFF_5_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4623, new_AGEMA_signal_4622, new_AGEMA_signal_4621, Midori_rounds_round_Result[7]}), .a ({new_AGEMA_signal_2472, new_AGEMA_signal_2471, new_AGEMA_signal_2470, Midori_add_Result_Start[7]}), .c ({new_AGEMA_signal_4800, new_AGEMA_signal_4799, new_AGEMA_signal_4798, Midori_rounds_roundResult_Reg_SFF_7_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4626, new_AGEMA_signal_4625, new_AGEMA_signal_4624, Midori_rounds_round_Result[9]}), .a ({new_AGEMA_signal_2460, new_AGEMA_signal_2459, new_AGEMA_signal_2458, Midori_add_Result_Start[9]}), .c ({new_AGEMA_signal_4803, new_AGEMA_signal_4802, new_AGEMA_signal_4801, Midori_rounds_roundResult_Reg_SFF_9_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4632, new_AGEMA_signal_4631, new_AGEMA_signal_4630, Midori_rounds_round_Result[11]}), .a ({new_AGEMA_signal_2826, new_AGEMA_signal_2825, new_AGEMA_signal_2824, Midori_add_Result_Start[11]}), .c ({new_AGEMA_signal_4809, new_AGEMA_signal_4808, new_AGEMA_signal_4807, Midori_rounds_roundResult_Reg_SFF_11_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4635, new_AGEMA_signal_4634, new_AGEMA_signal_4633, Midori_rounds_round_Result[13]}), .a ({new_AGEMA_signal_2814, new_AGEMA_signal_2813, new_AGEMA_signal_2812, Midori_add_Result_Start[13]}), .c ({new_AGEMA_signal_4812, new_AGEMA_signal_4811, new_AGEMA_signal_4810, Midori_rounds_roundResult_Reg_SFF_13_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4641, new_AGEMA_signal_4640, new_AGEMA_signal_4639, Midori_rounds_round_Result[15]}), .a ({new_AGEMA_signal_2802, new_AGEMA_signal_2801, new_AGEMA_signal_2800, Midori_add_Result_Start[15]}), .c ({new_AGEMA_signal_4818, new_AGEMA_signal_4817, new_AGEMA_signal_4816, Midori_rounds_roundResult_Reg_SFF_15_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4644, new_AGEMA_signal_4643, new_AGEMA_signal_4642, Midori_rounds_round_Result[17]}), .a ({new_AGEMA_signal_2790, new_AGEMA_signal_2789, new_AGEMA_signal_2788, Midori_add_Result_Start[17]}), .c ({new_AGEMA_signal_4821, new_AGEMA_signal_4820, new_AGEMA_signal_4819, Midori_rounds_roundResult_Reg_SFF_17_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4650, new_AGEMA_signal_4649, new_AGEMA_signal_4648, Midori_rounds_round_Result[19]}), .a ({new_AGEMA_signal_2778, new_AGEMA_signal_2777, new_AGEMA_signal_2776, Midori_add_Result_Start[19]}), .c ({new_AGEMA_signal_4827, new_AGEMA_signal_4826, new_AGEMA_signal_4825, Midori_rounds_roundResult_Reg_SFF_19_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, new_AGEMA_signal_4651, Midori_rounds_round_Result[21]}), .a ({new_AGEMA_signal_2760, new_AGEMA_signal_2759, new_AGEMA_signal_2758, Midori_add_Result_Start[21]}), .c ({new_AGEMA_signal_4830, new_AGEMA_signal_4829, new_AGEMA_signal_4828, Midori_rounds_roundResult_Reg_SFF_21_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4659, new_AGEMA_signal_4658, new_AGEMA_signal_4657, Midori_rounds_round_Result[23]}), .a ({new_AGEMA_signal_2748, new_AGEMA_signal_2747, new_AGEMA_signal_2746, Midori_add_Result_Start[23]}), .c ({new_AGEMA_signal_4836, new_AGEMA_signal_4835, new_AGEMA_signal_4834, Midori_rounds_roundResult_Reg_SFF_23_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4662, new_AGEMA_signal_4661, new_AGEMA_signal_4660, Midori_rounds_round_Result[25]}), .a ({new_AGEMA_signal_2736, new_AGEMA_signal_2735, new_AGEMA_signal_2734, Midori_add_Result_Start[25]}), .c ({new_AGEMA_signal_4839, new_AGEMA_signal_4838, new_AGEMA_signal_4837, Midori_rounds_roundResult_Reg_SFF_25_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4668, new_AGEMA_signal_4667, new_AGEMA_signal_4666, Midori_rounds_round_Result[27]}), .a ({new_AGEMA_signal_2724, new_AGEMA_signal_2723, new_AGEMA_signal_2722, Midori_add_Result_Start[27]}), .c ({new_AGEMA_signal_4845, new_AGEMA_signal_4844, new_AGEMA_signal_4843, Midori_rounds_roundResult_Reg_SFF_27_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, new_AGEMA_signal_4669, Midori_rounds_round_Result[29]}), .a ({new_AGEMA_signal_2712, new_AGEMA_signal_2711, new_AGEMA_signal_2710, Midori_add_Result_Start[29]}), .c ({new_AGEMA_signal_4848, new_AGEMA_signal_4847, new_AGEMA_signal_4846, Midori_rounds_roundResult_Reg_SFF_29_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4677, new_AGEMA_signal_4676, new_AGEMA_signal_4675, Midori_rounds_round_Result[31]}), .a ({new_AGEMA_signal_2694, new_AGEMA_signal_2693, new_AGEMA_signal_2692, Midori_add_Result_Start[31]}), .c ({new_AGEMA_signal_4854, new_AGEMA_signal_4853, new_AGEMA_signal_4852, Midori_rounds_roundResult_Reg_SFF_31_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4680, new_AGEMA_signal_4679, new_AGEMA_signal_4678, Midori_rounds_round_Result[33]}), .a ({new_AGEMA_signal_2682, new_AGEMA_signal_2681, new_AGEMA_signal_2680, Midori_add_Result_Start[33]}), .c ({new_AGEMA_signal_4857, new_AGEMA_signal_4856, new_AGEMA_signal_4855, Midori_rounds_roundResult_Reg_SFF_33_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4686, new_AGEMA_signal_4685, new_AGEMA_signal_4684, Midori_rounds_round_Result[35]}), .a ({new_AGEMA_signal_2670, new_AGEMA_signal_2669, new_AGEMA_signal_2668, Midori_add_Result_Start[35]}), .c ({new_AGEMA_signal_4863, new_AGEMA_signal_4862, new_AGEMA_signal_4861, Midori_rounds_roundResult_Reg_SFF_35_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4689, new_AGEMA_signal_4688, new_AGEMA_signal_4687, Midori_rounds_round_Result[37]}), .a ({new_AGEMA_signal_2658, new_AGEMA_signal_2657, new_AGEMA_signal_2656, Midori_add_Result_Start[37]}), .c ({new_AGEMA_signal_4866, new_AGEMA_signal_4865, new_AGEMA_signal_4864, Midori_rounds_roundResult_Reg_SFF_37_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4695, new_AGEMA_signal_4694, new_AGEMA_signal_4693, Midori_rounds_round_Result[39]}), .a ({new_AGEMA_signal_2646, new_AGEMA_signal_2645, new_AGEMA_signal_2644, Midori_add_Result_Start[39]}), .c ({new_AGEMA_signal_4872, new_AGEMA_signal_4871, new_AGEMA_signal_4870, Midori_rounds_roundResult_Reg_SFF_39_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4698, new_AGEMA_signal_4697, new_AGEMA_signal_4696, Midori_rounds_round_Result[41]}), .a ({new_AGEMA_signal_2628, new_AGEMA_signal_2627, new_AGEMA_signal_2626, Midori_add_Result_Start[41]}), .c ({new_AGEMA_signal_4875, new_AGEMA_signal_4874, new_AGEMA_signal_4873, Midori_rounds_roundResult_Reg_SFF_41_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4704, new_AGEMA_signal_4703, new_AGEMA_signal_4702, Midori_rounds_round_Result[43]}), .a ({new_AGEMA_signal_2616, new_AGEMA_signal_2615, new_AGEMA_signal_2614, Midori_add_Result_Start[43]}), .c ({new_AGEMA_signal_4881, new_AGEMA_signal_4880, new_AGEMA_signal_4879, Midori_rounds_roundResult_Reg_SFF_43_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4707, new_AGEMA_signal_4706, new_AGEMA_signal_4705, Midori_rounds_round_Result[45]}), .a ({new_AGEMA_signal_2604, new_AGEMA_signal_2603, new_AGEMA_signal_2602, Midori_add_Result_Start[45]}), .c ({new_AGEMA_signal_4884, new_AGEMA_signal_4883, new_AGEMA_signal_4882, Midori_rounds_roundResult_Reg_SFF_45_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, new_AGEMA_signal_4711, Midori_rounds_round_Result[47]}), .a ({new_AGEMA_signal_2592, new_AGEMA_signal_2591, new_AGEMA_signal_2590, Midori_add_Result_Start[47]}), .c ({new_AGEMA_signal_4890, new_AGEMA_signal_4889, new_AGEMA_signal_4888, Midori_rounds_roundResult_Reg_SFF_47_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4716, new_AGEMA_signal_4715, new_AGEMA_signal_4714, Midori_rounds_round_Result[49]}), .a ({new_AGEMA_signal_2580, new_AGEMA_signal_2579, new_AGEMA_signal_2578, Midori_add_Result_Start[49]}), .c ({new_AGEMA_signal_4893, new_AGEMA_signal_4892, new_AGEMA_signal_4891, Midori_rounds_roundResult_Reg_SFF_49_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4722, new_AGEMA_signal_4721, new_AGEMA_signal_4720, Midori_rounds_round_Result[51]}), .a ({new_AGEMA_signal_2562, new_AGEMA_signal_2561, new_AGEMA_signal_2560, Midori_add_Result_Start[51]}), .c ({new_AGEMA_signal_4899, new_AGEMA_signal_4898, new_AGEMA_signal_4897, Midori_rounds_roundResult_Reg_SFF_51_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, new_AGEMA_signal_4723, Midori_rounds_round_Result[53]}), .a ({new_AGEMA_signal_2550, new_AGEMA_signal_2549, new_AGEMA_signal_2548, Midori_add_Result_Start[53]}), .c ({new_AGEMA_signal_4902, new_AGEMA_signal_4901, new_AGEMA_signal_4900, Midori_rounds_roundResult_Reg_SFF_53_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, new_AGEMA_signal_4729, Midori_rounds_round_Result[55]}), .a ({new_AGEMA_signal_2538, new_AGEMA_signal_2537, new_AGEMA_signal_2536, Midori_add_Result_Start[55]}), .c ({new_AGEMA_signal_4908, new_AGEMA_signal_4907, new_AGEMA_signal_4906, Midori_rounds_roundResult_Reg_SFF_55_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4734, new_AGEMA_signal_4733, new_AGEMA_signal_4732, Midori_rounds_round_Result[57]}), .a ({new_AGEMA_signal_2526, new_AGEMA_signal_2525, new_AGEMA_signal_2524, Midori_add_Result_Start[57]}), .c ({new_AGEMA_signal_4911, new_AGEMA_signal_4910, new_AGEMA_signal_4909, Midori_rounds_roundResult_Reg_SFF_57_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4740, new_AGEMA_signal_4739, new_AGEMA_signal_4738, Midori_rounds_round_Result[59]}), .a ({new_AGEMA_signal_2514, new_AGEMA_signal_2513, new_AGEMA_signal_2512, Midori_add_Result_Start[59]}), .c ({new_AGEMA_signal_4917, new_AGEMA_signal_4916, new_AGEMA_signal_4915, Midori_rounds_roundResult_Reg_SFF_59_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, new_AGEMA_signal_4741, Midori_rounds_round_Result[61]}), .a ({new_AGEMA_signal_2496, new_AGEMA_signal_2495, new_AGEMA_signal_2494, Midori_add_Result_Start[61]}), .c ({new_AGEMA_signal_4920, new_AGEMA_signal_4919, new_AGEMA_signal_4918, Midori_rounds_roundResult_Reg_SFF_61_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, new_AGEMA_signal_4747, Midori_rounds_round_Result[63]}), .a ({new_AGEMA_signal_2484, new_AGEMA_signal_2483, new_AGEMA_signal_2482, Midori_add_Result_Start[63]}), .c ({new_AGEMA_signal_4926, new_AGEMA_signal_4925, new_AGEMA_signal_4924, Midori_rounds_roundResult_Reg_SFF_63_DQ}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U19 ( .a ({new_AGEMA_signal_2844, new_AGEMA_signal_2843, new_AGEMA_signal_2842, Midori_rounds_sub_sBox_PRINCE_0_n15}), .b ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, new_AGEMA_signal_3283, Midori_rounds_sub_sBox_PRINCE_0_n14}), .clk (clk), .r ({Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({new_AGEMA_signal_3522, new_AGEMA_signal_3521, new_AGEMA_signal_3520, Midori_rounds_SR_Result[51]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U16 ( .a ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, new_AGEMA_signal_2839, Midori_rounds_sub_sBox_PRINCE_0_n11}), .b ({new_AGEMA_signal_3282, new_AGEMA_signal_3281, new_AGEMA_signal_3280, Midori_rounds_roundReg_out[1]}), .clk (clk), .r ({Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966]}), .c ({new_AGEMA_signal_3288, new_AGEMA_signal_3287, new_AGEMA_signal_3286, Midori_rounds_sub_sBox_PRINCE_0_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U12 ( .a ({new_AGEMA_signal_2850, new_AGEMA_signal_2849, new_AGEMA_signal_2848, Midori_rounds_sub_sBox_PRINCE_0_n6}), .b ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, new_AGEMA_signal_3289, Midori_rounds_sub_sBox_PRINCE_0_n5}), .clk (clk), .r ({Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972]}), .c ({new_AGEMA_signal_3528, new_AGEMA_signal_3527, new_AGEMA_signal_3526, Midori_rounds_SR_Result[49]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U7 ( .a ({new_AGEMA_signal_3282, new_AGEMA_signal_3281, new_AGEMA_signal_3280, Midori_rounds_roundReg_out[1]}), .b ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, new_AGEMA_signal_2851, Midori_rounds_sub_sBox_PRINCE_0_n2}), .clk (clk), .r ({Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978]}), .c ({new_AGEMA_signal_3294, new_AGEMA_signal_3293, new_AGEMA_signal_3292, Midori_rounds_sub_sBox_PRINCE_0_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U19 ( .a ({new_AGEMA_signal_2862, new_AGEMA_signal_2861, new_AGEMA_signal_2860, Midori_rounds_sub_sBox_PRINCE_1_n15}), .b ({new_AGEMA_signal_3300, new_AGEMA_signal_3299, new_AGEMA_signal_3298, Midori_rounds_sub_sBox_PRINCE_1_n14}), .clk (clk), .r ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984]}), .c ({new_AGEMA_signal_3534, new_AGEMA_signal_3533, new_AGEMA_signal_3532, Midori_rounds_SR_Result[47]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U16 ( .a ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, new_AGEMA_signal_2857, Midori_rounds_sub_sBox_PRINCE_1_n11}), .b ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, new_AGEMA_signal_3295, Midori_rounds_roundReg_out[5]}), .clk (clk), .r ({Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .c ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, new_AGEMA_signal_3301, Midori_rounds_sub_sBox_PRINCE_1_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U12 ( .a ({new_AGEMA_signal_2868, new_AGEMA_signal_2867, new_AGEMA_signal_2866, Midori_rounds_sub_sBox_PRINCE_1_n6}), .b ({new_AGEMA_signal_3306, new_AGEMA_signal_3305, new_AGEMA_signal_3304, Midori_rounds_sub_sBox_PRINCE_1_n5}), .clk (clk), .r ({Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996]}), .c ({new_AGEMA_signal_3540, new_AGEMA_signal_3539, new_AGEMA_signal_3538, Midori_rounds_SR_Result[45]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U7 ( .a ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, new_AGEMA_signal_3295, Midori_rounds_roundReg_out[5]}), .b ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, new_AGEMA_signal_2869, Midori_rounds_sub_sBox_PRINCE_1_n2}), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, new_AGEMA_signal_3307, Midori_rounds_sub_sBox_PRINCE_1_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U19 ( .a ({new_AGEMA_signal_2880, new_AGEMA_signal_2879, new_AGEMA_signal_2878, Midori_rounds_sub_sBox_PRINCE_2_n15}), .b ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, new_AGEMA_signal_3313, Midori_rounds_sub_sBox_PRINCE_2_n14}), .clk (clk), .r ({Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({new_AGEMA_signal_3546, new_AGEMA_signal_3545, new_AGEMA_signal_3544, Midori_rounds_SR_Result[11]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U16 ( .a ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, new_AGEMA_signal_2875, Midori_rounds_sub_sBox_PRINCE_2_n11}), .b ({new_AGEMA_signal_3312, new_AGEMA_signal_3311, new_AGEMA_signal_3310, Midori_rounds_roundReg_out[9]}), .clk (clk), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({new_AGEMA_signal_3318, new_AGEMA_signal_3317, new_AGEMA_signal_3316, Midori_rounds_sub_sBox_PRINCE_2_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U12 ( .a ({new_AGEMA_signal_2886, new_AGEMA_signal_2885, new_AGEMA_signal_2884, Midori_rounds_sub_sBox_PRINCE_2_n6}), .b ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, new_AGEMA_signal_3319, Midori_rounds_sub_sBox_PRINCE_2_n5}), .clk (clk), .r ({Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({new_AGEMA_signal_3552, new_AGEMA_signal_3551, new_AGEMA_signal_3550, Midori_rounds_SR_Result[9]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U7 ( .a ({new_AGEMA_signal_3312, new_AGEMA_signal_3311, new_AGEMA_signal_3310, Midori_rounds_roundReg_out[9]}), .b ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, new_AGEMA_signal_2887, Midori_rounds_sub_sBox_PRINCE_2_n2}), .clk (clk), .r ({Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({new_AGEMA_signal_3324, new_AGEMA_signal_3323, new_AGEMA_signal_3322, Midori_rounds_sub_sBox_PRINCE_2_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U19 ( .a ({new_AGEMA_signal_2898, new_AGEMA_signal_2897, new_AGEMA_signal_2896, Midori_rounds_sub_sBox_PRINCE_3_n15}), .b ({new_AGEMA_signal_3330, new_AGEMA_signal_3329, new_AGEMA_signal_3328, Midori_rounds_sub_sBox_PRINCE_3_n14}), .clk (clk), .r ({Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({new_AGEMA_signal_3558, new_AGEMA_signal_3557, new_AGEMA_signal_3556, Midori_rounds_SR_Result[23]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U16 ( .a ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, new_AGEMA_signal_2893, Midori_rounds_sub_sBox_PRINCE_3_n11}), .b ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, new_AGEMA_signal_3325, Midori_rounds_roundReg_out[13]}), .clk (clk), .r ({Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, new_AGEMA_signal_3331, Midori_rounds_sub_sBox_PRINCE_3_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U12 ( .a ({new_AGEMA_signal_2904, new_AGEMA_signal_2903, new_AGEMA_signal_2902, Midori_rounds_sub_sBox_PRINCE_3_n6}), .b ({new_AGEMA_signal_3336, new_AGEMA_signal_3335, new_AGEMA_signal_3334, Midori_rounds_sub_sBox_PRINCE_3_n5}), .clk (clk), .r ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({new_AGEMA_signal_3564, new_AGEMA_signal_3563, new_AGEMA_signal_3562, Midori_rounds_SR_Result[21]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U7 ( .a ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, new_AGEMA_signal_3325, Midori_rounds_roundReg_out[13]}), .b ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, new_AGEMA_signal_2905, Midori_rounds_sub_sBox_PRINCE_3_n2}), .clk (clk), .r ({Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, new_AGEMA_signal_3337, Midori_rounds_sub_sBox_PRINCE_3_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U19 ( .a ({new_AGEMA_signal_2916, new_AGEMA_signal_2915, new_AGEMA_signal_2914, Midori_rounds_sub_sBox_PRINCE_4_n15}), .b ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, new_AGEMA_signal_3343, Midori_rounds_sub_sBox_PRINCE_4_n14}), .clk (clk), .r ({Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({new_AGEMA_signal_3570, new_AGEMA_signal_3569, new_AGEMA_signal_3568, Midori_rounds_SR_Result[39]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U16 ( .a ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, new_AGEMA_signal_2911, Midori_rounds_sub_sBox_PRINCE_4_n11}), .b ({new_AGEMA_signal_3342, new_AGEMA_signal_3341, new_AGEMA_signal_3340, Midori_rounds_roundReg_out[17]}), .clk (clk), .r ({Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({new_AGEMA_signal_3348, new_AGEMA_signal_3347, new_AGEMA_signal_3346, Midori_rounds_sub_sBox_PRINCE_4_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U12 ( .a ({new_AGEMA_signal_2922, new_AGEMA_signal_2921, new_AGEMA_signal_2920, Midori_rounds_sub_sBox_PRINCE_4_n6}), .b ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, new_AGEMA_signal_3349, Midori_rounds_sub_sBox_PRINCE_4_n5}), .clk (clk), .r ({Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({new_AGEMA_signal_3576, new_AGEMA_signal_3575, new_AGEMA_signal_3574, Midori_rounds_SR_Result[37]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U7 ( .a ({new_AGEMA_signal_3342, new_AGEMA_signal_3341, new_AGEMA_signal_3340, Midori_rounds_roundReg_out[17]}), .b ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, new_AGEMA_signal_2923, Midori_rounds_sub_sBox_PRINCE_4_n2}), .clk (clk), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({new_AGEMA_signal_3354, new_AGEMA_signal_3353, new_AGEMA_signal_3352, Midori_rounds_sub_sBox_PRINCE_4_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U19 ( .a ({new_AGEMA_signal_2934, new_AGEMA_signal_2933, new_AGEMA_signal_2932, Midori_rounds_sub_sBox_PRINCE_5_n15}), .b ({new_AGEMA_signal_3360, new_AGEMA_signal_3359, new_AGEMA_signal_3358, Midori_rounds_sub_sBox_PRINCE_5_n14}), .clk (clk), .r ({Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({new_AGEMA_signal_3582, new_AGEMA_signal_3581, new_AGEMA_signal_3580, Midori_rounds_SR_Result[59]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U16 ( .a ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, new_AGEMA_signal_2929, Midori_rounds_sub_sBox_PRINCE_5_n11}), .b ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, new_AGEMA_signal_3355, Midori_rounds_roundReg_out[21]}), .clk (clk), .r ({Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, new_AGEMA_signal_3361, Midori_rounds_sub_sBox_PRINCE_5_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U12 ( .a ({new_AGEMA_signal_2940, new_AGEMA_signal_2939, new_AGEMA_signal_2938, Midori_rounds_sub_sBox_PRINCE_5_n6}), .b ({new_AGEMA_signal_3366, new_AGEMA_signal_3365, new_AGEMA_signal_3364, Midori_rounds_sub_sBox_PRINCE_5_n5}), .clk (clk), .r ({Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({new_AGEMA_signal_3588, new_AGEMA_signal_3587, new_AGEMA_signal_3586, Midori_rounds_SR_Result[57]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U7 ( .a ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, new_AGEMA_signal_3355, Midori_rounds_roundReg_out[21]}), .b ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, new_AGEMA_signal_2941, Midori_rounds_sub_sBox_PRINCE_5_n2}), .clk (clk), .r ({Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, new_AGEMA_signal_3367, Midori_rounds_sub_sBox_PRINCE_5_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U19 ( .a ({new_AGEMA_signal_2952, new_AGEMA_signal_2951, new_AGEMA_signal_2950, Midori_rounds_sub_sBox_PRINCE_6_n15}), .b ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, new_AGEMA_signal_3373, Midori_rounds_sub_sBox_PRINCE_6_n14}), .clk (clk), .r ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({new_AGEMA_signal_3594, new_AGEMA_signal_3593, new_AGEMA_signal_3592, Midori_rounds_SR_Result[31]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U16 ( .a ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, new_AGEMA_signal_2947, Midori_rounds_sub_sBox_PRINCE_6_n11}), .b ({new_AGEMA_signal_3372, new_AGEMA_signal_3371, new_AGEMA_signal_3370, Midori_rounds_roundReg_out[25]}), .clk (clk), .r ({Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({new_AGEMA_signal_3378, new_AGEMA_signal_3377, new_AGEMA_signal_3376, Midori_rounds_sub_sBox_PRINCE_6_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U12 ( .a ({new_AGEMA_signal_2958, new_AGEMA_signal_2957, new_AGEMA_signal_2956, Midori_rounds_sub_sBox_PRINCE_6_n6}), .b ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, new_AGEMA_signal_3379, Midori_rounds_sub_sBox_PRINCE_6_n5}), .clk (clk), .r ({Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({new_AGEMA_signal_3600, new_AGEMA_signal_3599, new_AGEMA_signal_3598, Midori_rounds_SR_Result[29]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U7 ( .a ({new_AGEMA_signal_3372, new_AGEMA_signal_3371, new_AGEMA_signal_3370, Midori_rounds_roundReg_out[25]}), .b ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, new_AGEMA_signal_2959, Midori_rounds_sub_sBox_PRINCE_6_n2}), .clk (clk), .r ({Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({new_AGEMA_signal_3384, new_AGEMA_signal_3383, new_AGEMA_signal_3382, Midori_rounds_sub_sBox_PRINCE_6_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U19 ( .a ({new_AGEMA_signal_2970, new_AGEMA_signal_2969, new_AGEMA_signal_2968, Midori_rounds_sub_sBox_PRINCE_7_n15}), .b ({new_AGEMA_signal_3390, new_AGEMA_signal_3389, new_AGEMA_signal_3388, Midori_rounds_sub_sBox_PRINCE_7_n14}), .clk (clk), .r ({Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({new_AGEMA_signal_3606, new_AGEMA_signal_3605, new_AGEMA_signal_3604, Midori_rounds_SR_Result[3]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U16 ( .a ({new_AGEMA_signal_2967, new_AGEMA_signal_2966, new_AGEMA_signal_2965, Midori_rounds_sub_sBox_PRINCE_7_n11}), .b ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, new_AGEMA_signal_3385, Midori_rounds_roundReg_out[29]}), .clk (clk), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, new_AGEMA_signal_3391, Midori_rounds_sub_sBox_PRINCE_7_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U12 ( .a ({new_AGEMA_signal_2976, new_AGEMA_signal_2975, new_AGEMA_signal_2974, Midori_rounds_sub_sBox_PRINCE_7_n6}), .b ({new_AGEMA_signal_3396, new_AGEMA_signal_3395, new_AGEMA_signal_3394, Midori_rounds_sub_sBox_PRINCE_7_n5}), .clk (clk), .r ({Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({new_AGEMA_signal_3612, new_AGEMA_signal_3611, new_AGEMA_signal_3610, Midori_rounds_SR_Result[1]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U7 ( .a ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, new_AGEMA_signal_3385, Midori_rounds_roundReg_out[29]}), .b ({new_AGEMA_signal_2979, new_AGEMA_signal_2978, new_AGEMA_signal_2977, Midori_rounds_sub_sBox_PRINCE_7_n2}), .clk (clk), .r ({Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, new_AGEMA_signal_3397, Midori_rounds_sub_sBox_PRINCE_7_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U19 ( .a ({new_AGEMA_signal_2988, new_AGEMA_signal_2987, new_AGEMA_signal_2986, Midori_rounds_sub_sBox_PRINCE_8_n15}), .b ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, new_AGEMA_signal_3403, Midori_rounds_sub_sBox_PRINCE_8_n14}), .clk (clk), .r ({Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({new_AGEMA_signal_3618, new_AGEMA_signal_3617, new_AGEMA_signal_3616, Midori_rounds_SR_Result[15]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U16 ( .a ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, new_AGEMA_signal_2983, Midori_rounds_sub_sBox_PRINCE_8_n11}), .b ({new_AGEMA_signal_3402, new_AGEMA_signal_3401, new_AGEMA_signal_3400, Midori_rounds_roundReg_out[33]}), .clk (clk), .r ({Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({new_AGEMA_signal_3408, new_AGEMA_signal_3407, new_AGEMA_signal_3406, Midori_rounds_sub_sBox_PRINCE_8_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U12 ( .a ({new_AGEMA_signal_2994, new_AGEMA_signal_2993, new_AGEMA_signal_2992, Midori_rounds_sub_sBox_PRINCE_8_n6}), .b ({new_AGEMA_signal_3411, new_AGEMA_signal_3410, new_AGEMA_signal_3409, Midori_rounds_sub_sBox_PRINCE_8_n5}), .clk (clk), .r ({Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({new_AGEMA_signal_3624, new_AGEMA_signal_3623, new_AGEMA_signal_3622, Midori_rounds_SR_Result[13]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U7 ( .a ({new_AGEMA_signal_3402, new_AGEMA_signal_3401, new_AGEMA_signal_3400, Midori_rounds_roundReg_out[33]}), .b ({new_AGEMA_signal_2997, new_AGEMA_signal_2996, new_AGEMA_signal_2995, Midori_rounds_sub_sBox_PRINCE_8_n2}), .clk (clk), .r ({Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({new_AGEMA_signal_3414, new_AGEMA_signal_3413, new_AGEMA_signal_3412, Midori_rounds_sub_sBox_PRINCE_8_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U19 ( .a ({new_AGEMA_signal_3006, new_AGEMA_signal_3005, new_AGEMA_signal_3004, Midori_rounds_sub_sBox_PRINCE_9_n15}), .b ({new_AGEMA_signal_3420, new_AGEMA_signal_3419, new_AGEMA_signal_3418, Midori_rounds_sub_sBox_PRINCE_9_n14}), .clk (clk), .r ({Fresh[1181], Fresh[1180], Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({new_AGEMA_signal_3630, new_AGEMA_signal_3629, new_AGEMA_signal_3628, Midori_rounds_SR_Result[19]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U16 ( .a ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, new_AGEMA_signal_3001, Midori_rounds_sub_sBox_PRINCE_9_n11}), .b ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, new_AGEMA_signal_3415, Midori_rounds_roundReg_out[37]}), .clk (clk), .r ({Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, new_AGEMA_signal_3421, Midori_rounds_sub_sBox_PRINCE_9_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U12 ( .a ({new_AGEMA_signal_3012, new_AGEMA_signal_3011, new_AGEMA_signal_3010, Midori_rounds_sub_sBox_PRINCE_9_n6}), .b ({new_AGEMA_signal_3426, new_AGEMA_signal_3425, new_AGEMA_signal_3424, Midori_rounds_sub_sBox_PRINCE_9_n5}), .clk (clk), .r ({Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({new_AGEMA_signal_3636, new_AGEMA_signal_3635, new_AGEMA_signal_3634, Midori_rounds_SR_Result[17]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U7 ( .a ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, new_AGEMA_signal_3415, Midori_rounds_roundReg_out[37]}), .b ({new_AGEMA_signal_3015, new_AGEMA_signal_3014, new_AGEMA_signal_3013, Midori_rounds_sub_sBox_PRINCE_9_n2}), .clk (clk), .r ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, new_AGEMA_signal_3427, Midori_rounds_sub_sBox_PRINCE_9_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U19 ( .a ({new_AGEMA_signal_3024, new_AGEMA_signal_3023, new_AGEMA_signal_3022, Midori_rounds_sub_sBox_PRINCE_10_n15}), .b ({new_AGEMA_signal_3435, new_AGEMA_signal_3434, new_AGEMA_signal_3433, Midori_rounds_sub_sBox_PRINCE_10_n14}), .clk (clk), .r ({Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({new_AGEMA_signal_3642, new_AGEMA_signal_3641, new_AGEMA_signal_3640, Midori_rounds_SR_Result[55]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U16 ( .a ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, new_AGEMA_signal_3019, Midori_rounds_sub_sBox_PRINCE_10_n11}), .b ({new_AGEMA_signal_3432, new_AGEMA_signal_3431, new_AGEMA_signal_3430, Midori_rounds_roundReg_out[41]}), .clk (clk), .r ({Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({new_AGEMA_signal_3438, new_AGEMA_signal_3437, new_AGEMA_signal_3436, Midori_rounds_sub_sBox_PRINCE_10_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U12 ( .a ({new_AGEMA_signal_3030, new_AGEMA_signal_3029, new_AGEMA_signal_3028, Midori_rounds_sub_sBox_PRINCE_10_n6}), .b ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, new_AGEMA_signal_3439, Midori_rounds_sub_sBox_PRINCE_10_n5}), .clk (clk), .r ({Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({new_AGEMA_signal_3648, new_AGEMA_signal_3647, new_AGEMA_signal_3646, Midori_rounds_SR_Result[53]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U7 ( .a ({new_AGEMA_signal_3432, new_AGEMA_signal_3431, new_AGEMA_signal_3430, Midori_rounds_roundReg_out[41]}), .b ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, new_AGEMA_signal_3031, Midori_rounds_sub_sBox_PRINCE_10_n2}), .clk (clk), .r ({Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({new_AGEMA_signal_3444, new_AGEMA_signal_3443, new_AGEMA_signal_3442, Midori_rounds_sub_sBox_PRINCE_10_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U19 ( .a ({new_AGEMA_signal_3042, new_AGEMA_signal_3041, new_AGEMA_signal_3040, Midori_rounds_sub_sBox_PRINCE_11_n15}), .b ({new_AGEMA_signal_3450, new_AGEMA_signal_3449, new_AGEMA_signal_3448, Midori_rounds_sub_sBox_PRINCE_11_n14}), .clk (clk), .r ({Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({new_AGEMA_signal_3654, new_AGEMA_signal_3653, new_AGEMA_signal_3652, Midori_rounds_SR_Result[43]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U16 ( .a ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, new_AGEMA_signal_3037, Midori_rounds_sub_sBox_PRINCE_11_n11}), .b ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, new_AGEMA_signal_3445, Midori_rounds_roundReg_out[45]}), .clk (clk), .r ({Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, new_AGEMA_signal_3451, Midori_rounds_sub_sBox_PRINCE_11_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U12 ( .a ({new_AGEMA_signal_3048, new_AGEMA_signal_3047, new_AGEMA_signal_3046, Midori_rounds_sub_sBox_PRINCE_11_n6}), .b ({new_AGEMA_signal_3456, new_AGEMA_signal_3455, new_AGEMA_signal_3454, Midori_rounds_sub_sBox_PRINCE_11_n5}), .clk (clk), .r ({Fresh[1241], Fresh[1240], Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({new_AGEMA_signal_3660, new_AGEMA_signal_3659, new_AGEMA_signal_3658, Midori_rounds_SR_Result[41]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U7 ( .a ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, new_AGEMA_signal_3445, Midori_rounds_roundReg_out[45]}), .b ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, new_AGEMA_signal_3049, Midori_rounds_sub_sBox_PRINCE_11_n2}), .clk (clk), .r ({Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242]}), .c ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, new_AGEMA_signal_3457, Midori_rounds_sub_sBox_PRINCE_11_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U19 ( .a ({new_AGEMA_signal_3060, new_AGEMA_signal_3059, new_AGEMA_signal_3058, Midori_rounds_sub_sBox_PRINCE_12_n15}), .b ({new_AGEMA_signal_3465, new_AGEMA_signal_3464, new_AGEMA_signal_3463, Midori_rounds_sub_sBox_PRINCE_12_n14}), .clk (clk), .r ({Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({new_AGEMA_signal_3666, new_AGEMA_signal_3665, new_AGEMA_signal_3664, Midori_rounds_SR_Result[27]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U16 ( .a ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, new_AGEMA_signal_3055, Midori_rounds_sub_sBox_PRINCE_12_n11}), .b ({new_AGEMA_signal_3462, new_AGEMA_signal_3461, new_AGEMA_signal_3460, Midori_rounds_roundReg_out[49]}), .clk (clk), .r ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254]}), .c ({new_AGEMA_signal_3468, new_AGEMA_signal_3467, new_AGEMA_signal_3466, Midori_rounds_sub_sBox_PRINCE_12_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U12 ( .a ({new_AGEMA_signal_3066, new_AGEMA_signal_3065, new_AGEMA_signal_3064, Midori_rounds_sub_sBox_PRINCE_12_n6}), .b ({new_AGEMA_signal_3471, new_AGEMA_signal_3470, new_AGEMA_signal_3469, Midori_rounds_sub_sBox_PRINCE_12_n5}), .clk (clk), .r ({Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({new_AGEMA_signal_3672, new_AGEMA_signal_3671, new_AGEMA_signal_3670, Midori_rounds_SR_Result[25]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U7 ( .a ({new_AGEMA_signal_3462, new_AGEMA_signal_3461, new_AGEMA_signal_3460, Midori_rounds_roundReg_out[49]}), .b ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, new_AGEMA_signal_3067, Midori_rounds_sub_sBox_PRINCE_12_n2}), .clk (clk), .r ({Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266]}), .c ({new_AGEMA_signal_3474, new_AGEMA_signal_3473, new_AGEMA_signal_3472, Midori_rounds_sub_sBox_PRINCE_12_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U19 ( .a ({new_AGEMA_signal_3078, new_AGEMA_signal_3077, new_AGEMA_signal_3076, Midori_rounds_sub_sBox_PRINCE_13_n15}), .b ({new_AGEMA_signal_3480, new_AGEMA_signal_3479, new_AGEMA_signal_3478, Midori_rounds_sub_sBox_PRINCE_13_n14}), .clk (clk), .r ({Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({new_AGEMA_signal_3678, new_AGEMA_signal_3677, new_AGEMA_signal_3676, Midori_rounds_SR_Result[7]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U16 ( .a ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, new_AGEMA_signal_3073, Midori_rounds_sub_sBox_PRINCE_13_n11}), .b ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, new_AGEMA_signal_3475, Midori_rounds_roundReg_out[53]}), .clk (clk), .r ({Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280], Fresh[1279], Fresh[1278]}), .c ({new_AGEMA_signal_3483, new_AGEMA_signal_3482, new_AGEMA_signal_3481, Midori_rounds_sub_sBox_PRINCE_13_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U12 ( .a ({new_AGEMA_signal_3084, new_AGEMA_signal_3083, new_AGEMA_signal_3082, Midori_rounds_sub_sBox_PRINCE_13_n6}), .b ({new_AGEMA_signal_3486, new_AGEMA_signal_3485, new_AGEMA_signal_3484, Midori_rounds_sub_sBox_PRINCE_13_n5}), .clk (clk), .r ({Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({new_AGEMA_signal_3684, new_AGEMA_signal_3683, new_AGEMA_signal_3682, Midori_rounds_SR_Result[5]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U7 ( .a ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, new_AGEMA_signal_3475, Midori_rounds_roundReg_out[53]}), .b ({new_AGEMA_signal_3087, new_AGEMA_signal_3086, new_AGEMA_signal_3085, Midori_rounds_sub_sBox_PRINCE_13_n2}), .clk (clk), .r ({Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, new_AGEMA_signal_3487, Midori_rounds_sub_sBox_PRINCE_13_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U19 ( .a ({new_AGEMA_signal_3096, new_AGEMA_signal_3095, new_AGEMA_signal_3094, Midori_rounds_sub_sBox_PRINCE_14_n15}), .b ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, new_AGEMA_signal_3493, Midori_rounds_sub_sBox_PRINCE_14_n14}), .clk (clk), .r ({Fresh[1301], Fresh[1300], Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({new_AGEMA_signal_3690, new_AGEMA_signal_3689, new_AGEMA_signal_3688, Midori_rounds_SR_Result[35]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U16 ( .a ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, new_AGEMA_signal_3091, Midori_rounds_sub_sBox_PRINCE_14_n11}), .b ({new_AGEMA_signal_3492, new_AGEMA_signal_3491, new_AGEMA_signal_3490, Midori_rounds_roundReg_out[57]}), .clk (clk), .r ({Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302]}), .c ({new_AGEMA_signal_3498, new_AGEMA_signal_3497, new_AGEMA_signal_3496, Midori_rounds_sub_sBox_PRINCE_14_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U12 ( .a ({new_AGEMA_signal_3102, new_AGEMA_signal_3101, new_AGEMA_signal_3100, Midori_rounds_sub_sBox_PRINCE_14_n6}), .b ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, new_AGEMA_signal_3499, Midori_rounds_sub_sBox_PRINCE_14_n5}), .clk (clk), .r ({Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({new_AGEMA_signal_3696, new_AGEMA_signal_3695, new_AGEMA_signal_3694, Midori_rounds_SR_Result[33]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U7 ( .a ({new_AGEMA_signal_3492, new_AGEMA_signal_3491, new_AGEMA_signal_3490, Midori_rounds_roundReg_out[57]}), .b ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, new_AGEMA_signal_3103, Midori_rounds_sub_sBox_PRINCE_14_n2}), .clk (clk), .r ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314]}), .c ({new_AGEMA_signal_3504, new_AGEMA_signal_3503, new_AGEMA_signal_3502, Midori_rounds_sub_sBox_PRINCE_14_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U19 ( .a ({new_AGEMA_signal_3114, new_AGEMA_signal_3113, new_AGEMA_signal_3112, Midori_rounds_sub_sBox_PRINCE_15_n15}), .b ({new_AGEMA_signal_3510, new_AGEMA_signal_3509, new_AGEMA_signal_3508, Midori_rounds_sub_sBox_PRINCE_15_n14}), .clk (clk), .r ({Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({new_AGEMA_signal_3702, new_AGEMA_signal_3701, new_AGEMA_signal_3700, Midori_rounds_SR_Result[63]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U16 ( .a ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, new_AGEMA_signal_3109, Midori_rounds_sub_sBox_PRINCE_15_n11}), .b ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, new_AGEMA_signal_3505, Midori_rounds_roundReg_out[61]}), .clk (clk), .r ({Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326]}), .c ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, new_AGEMA_signal_3511, Midori_rounds_sub_sBox_PRINCE_15_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U12 ( .a ({new_AGEMA_signal_3120, new_AGEMA_signal_3119, new_AGEMA_signal_3118, Midori_rounds_sub_sBox_PRINCE_15_n6}), .b ({new_AGEMA_signal_3516, new_AGEMA_signal_3515, new_AGEMA_signal_3514, Midori_rounds_sub_sBox_PRINCE_15_n5}), .clk (clk), .r ({Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({new_AGEMA_signal_3708, new_AGEMA_signal_3707, new_AGEMA_signal_3706, Midori_rounds_SR_Result[61]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U7 ( .a ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, new_AGEMA_signal_3505, Midori_rounds_roundReg_out[61]}), .b ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, new_AGEMA_signal_3121, Midori_rounds_sub_sBox_PRINCE_15_n2}), .clk (clk), .r ({Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340], Fresh[1339], Fresh[1338]}), .c ({new_AGEMA_signal_3519, new_AGEMA_signal_3518, new_AGEMA_signal_3517, Midori_rounds_sub_sBox_PRINCE_15_n3}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_1_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3612, new_AGEMA_signal_3611, new_AGEMA_signal_3610, Midori_rounds_SR_Result[1]}), .a ({new_AGEMA_signal_4023, new_AGEMA_signal_4022, new_AGEMA_signal_4021, Midori_rounds_sub_ResultXORkey[1]}), .c ({new_AGEMA_signal_4050, new_AGEMA_signal_4049, new_AGEMA_signal_4048, Midori_rounds_mul_input[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_3_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3606, new_AGEMA_signal_3605, new_AGEMA_signal_3604, Midori_rounds_SR_Result[3]}), .a ({new_AGEMA_signal_3972, new_AGEMA_signal_3971, new_AGEMA_signal_3970, Midori_rounds_sub_ResultXORkey[3]}), .c ({new_AGEMA_signal_4056, new_AGEMA_signal_4055, new_AGEMA_signal_4054, Midori_rounds_mul_input[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_5_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3684, new_AGEMA_signal_3683, new_AGEMA_signal_3682, Midori_rounds_SR_Result[5]}), .a ({new_AGEMA_signal_3924, new_AGEMA_signal_3923, new_AGEMA_signal_3922, Midori_rounds_sub_ResultXORkey[5]}), .c ({new_AGEMA_signal_4059, new_AGEMA_signal_4058, new_AGEMA_signal_4057, Midori_rounds_mul_input[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_7_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3678, new_AGEMA_signal_3677, new_AGEMA_signal_3676, Midori_rounds_SR_Result[7]}), .a ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, new_AGEMA_signal_3907, Midori_rounds_sub_ResultXORkey[7]}), .c ({new_AGEMA_signal_4065, new_AGEMA_signal_4064, new_AGEMA_signal_4063, Midori_rounds_mul_input[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_9_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3552, new_AGEMA_signal_3551, new_AGEMA_signal_3550, Midori_rounds_SR_Result[9]}), .a ({new_AGEMA_signal_3906, new_AGEMA_signal_3905, new_AGEMA_signal_3904, Midori_rounds_sub_ResultXORkey[9]}), .c ({new_AGEMA_signal_4068, new_AGEMA_signal_4067, new_AGEMA_signal_4066, Midori_rounds_mul_input[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_11_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3546, new_AGEMA_signal_3545, new_AGEMA_signal_3544, Midori_rounds_SR_Result[11]}), .a ({new_AGEMA_signal_4044, new_AGEMA_signal_4043, new_AGEMA_signal_4042, Midori_rounds_sub_ResultXORkey[11]}), .c ({new_AGEMA_signal_4074, new_AGEMA_signal_4073, new_AGEMA_signal_4072, Midori_rounds_mul_input[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_13_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3624, new_AGEMA_signal_3623, new_AGEMA_signal_3622, Midori_rounds_SR_Result[13]}), .a ({new_AGEMA_signal_4041, new_AGEMA_signal_4040, new_AGEMA_signal_4039, Midori_rounds_sub_ResultXORkey[13]}), .c ({new_AGEMA_signal_4077, new_AGEMA_signal_4076, new_AGEMA_signal_4075, Midori_rounds_mul_input[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_15_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3618, new_AGEMA_signal_3617, new_AGEMA_signal_3616, Midori_rounds_SR_Result[15]}), .a ({new_AGEMA_signal_4035, new_AGEMA_signal_4034, new_AGEMA_signal_4033, Midori_rounds_sub_ResultXORkey[15]}), .c ({new_AGEMA_signal_4083, new_AGEMA_signal_4082, new_AGEMA_signal_4081, Midori_rounds_mul_input[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_17_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3636, new_AGEMA_signal_3635, new_AGEMA_signal_3634, Midori_rounds_SR_Result[17]}), .a ({new_AGEMA_signal_4032, new_AGEMA_signal_4031, new_AGEMA_signal_4030, Midori_rounds_sub_ResultXORkey[17]}), .c ({new_AGEMA_signal_4086, new_AGEMA_signal_4085, new_AGEMA_signal_4084, Midori_rounds_mul_input[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_19_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3630, new_AGEMA_signal_3629, new_AGEMA_signal_3628, Midori_rounds_SR_Result[19]}), .a ({new_AGEMA_signal_4026, new_AGEMA_signal_4025, new_AGEMA_signal_4024, Midori_rounds_sub_ResultXORkey[19]}), .c ({new_AGEMA_signal_4092, new_AGEMA_signal_4091, new_AGEMA_signal_4090, Midori_rounds_mul_input[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_21_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3564, new_AGEMA_signal_3563, new_AGEMA_signal_3562, Midori_rounds_SR_Result[21]}), .a ({new_AGEMA_signal_4020, new_AGEMA_signal_4019, new_AGEMA_signal_4018, Midori_rounds_sub_ResultXORkey[21]}), .c ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, new_AGEMA_signal_4093, Midori_rounds_mul_input[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_23_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3558, new_AGEMA_signal_3557, new_AGEMA_signal_3556, Midori_rounds_SR_Result[23]}), .a ({new_AGEMA_signal_4014, new_AGEMA_signal_4013, new_AGEMA_signal_4012, Midori_rounds_sub_ResultXORkey[23]}), .c ({new_AGEMA_signal_4101, new_AGEMA_signal_4100, new_AGEMA_signal_4099, Midori_rounds_mul_input[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_25_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3672, new_AGEMA_signal_3671, new_AGEMA_signal_3670, Midori_rounds_SR_Result[25]}), .a ({new_AGEMA_signal_4011, new_AGEMA_signal_4010, new_AGEMA_signal_4009, Midori_rounds_sub_ResultXORkey[25]}), .c ({new_AGEMA_signal_4104, new_AGEMA_signal_4103, new_AGEMA_signal_4102, Midori_rounds_mul_input[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_27_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3666, new_AGEMA_signal_3665, new_AGEMA_signal_3664, Midori_rounds_SR_Result[27]}), .a ({new_AGEMA_signal_4005, new_AGEMA_signal_4004, new_AGEMA_signal_4003, Midori_rounds_sub_ResultXORkey[27]}), .c ({new_AGEMA_signal_4110, new_AGEMA_signal_4109, new_AGEMA_signal_4108, Midori_rounds_mul_input[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_29_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3600, new_AGEMA_signal_3599, new_AGEMA_signal_3598, Midori_rounds_SR_Result[29]}), .a ({new_AGEMA_signal_4002, new_AGEMA_signal_4001, new_AGEMA_signal_4000, Midori_rounds_sub_ResultXORkey[29]}), .c ({new_AGEMA_signal_4113, new_AGEMA_signal_4112, new_AGEMA_signal_4111, Midori_rounds_mul_input[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_31_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3594, new_AGEMA_signal_3593, new_AGEMA_signal_3592, Midori_rounds_SR_Result[31]}), .a ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, new_AGEMA_signal_3991, Midori_rounds_sub_ResultXORkey[31]}), .c ({new_AGEMA_signal_4119, new_AGEMA_signal_4118, new_AGEMA_signal_4117, Midori_rounds_mul_input[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_33_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3696, new_AGEMA_signal_3695, new_AGEMA_signal_3694, Midori_rounds_SR_Result[33]}), .a ({new_AGEMA_signal_3990, new_AGEMA_signal_3989, new_AGEMA_signal_3988, Midori_rounds_sub_ResultXORkey[33]}), .c ({new_AGEMA_signal_4122, new_AGEMA_signal_4121, new_AGEMA_signal_4120, Midori_rounds_mul_input[33]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_35_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3690, new_AGEMA_signal_3689, new_AGEMA_signal_3688, Midori_rounds_SR_Result[35]}), .a ({new_AGEMA_signal_3984, new_AGEMA_signal_3983, new_AGEMA_signal_3982, Midori_rounds_sub_ResultXORkey[35]}), .c ({new_AGEMA_signal_4128, new_AGEMA_signal_4127, new_AGEMA_signal_4126, Midori_rounds_mul_input[35]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_37_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3576, new_AGEMA_signal_3575, new_AGEMA_signal_3574, Midori_rounds_SR_Result[37]}), .a ({new_AGEMA_signal_3981, new_AGEMA_signal_3980, new_AGEMA_signal_3979, Midori_rounds_sub_ResultXORkey[37]}), .c ({new_AGEMA_signal_4131, new_AGEMA_signal_4130, new_AGEMA_signal_4129, Midori_rounds_mul_input[37]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_39_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3570, new_AGEMA_signal_3569, new_AGEMA_signal_3568, Midori_rounds_SR_Result[39]}), .a ({new_AGEMA_signal_3975, new_AGEMA_signal_3974, new_AGEMA_signal_3973, Midori_rounds_sub_ResultXORkey[39]}), .c ({new_AGEMA_signal_4137, new_AGEMA_signal_4136, new_AGEMA_signal_4135, Midori_rounds_mul_input[39]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_41_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3660, new_AGEMA_signal_3659, new_AGEMA_signal_3658, Midori_rounds_SR_Result[41]}), .a ({new_AGEMA_signal_3969, new_AGEMA_signal_3968, new_AGEMA_signal_3967, Midori_rounds_sub_ResultXORkey[41]}), .c ({new_AGEMA_signal_4140, new_AGEMA_signal_4139, new_AGEMA_signal_4138, Midori_rounds_mul_input[41]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_43_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3654, new_AGEMA_signal_3653, new_AGEMA_signal_3652, Midori_rounds_SR_Result[43]}), .a ({new_AGEMA_signal_3963, new_AGEMA_signal_3962, new_AGEMA_signal_3961, Midori_rounds_sub_ResultXORkey[43]}), .c ({new_AGEMA_signal_4146, new_AGEMA_signal_4145, new_AGEMA_signal_4144, Midori_rounds_mul_input[43]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_45_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3540, new_AGEMA_signal_3539, new_AGEMA_signal_3538, Midori_rounds_SR_Result[45]}), .a ({new_AGEMA_signal_3960, new_AGEMA_signal_3959, new_AGEMA_signal_3958, Midori_rounds_sub_ResultXORkey[45]}), .c ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, new_AGEMA_signal_4147, Midori_rounds_mul_input[45]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_47_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3534, new_AGEMA_signal_3533, new_AGEMA_signal_3532, Midori_rounds_SR_Result[47]}), .a ({new_AGEMA_signal_3954, new_AGEMA_signal_3953, new_AGEMA_signal_3952, Midori_rounds_sub_ResultXORkey[47]}), .c ({new_AGEMA_signal_4155, new_AGEMA_signal_4154, new_AGEMA_signal_4153, Midori_rounds_mul_input[47]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_49_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3528, new_AGEMA_signal_3527, new_AGEMA_signal_3526, Midori_rounds_SR_Result[49]}), .a ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, new_AGEMA_signal_3949, Midori_rounds_sub_ResultXORkey[49]}), .c ({new_AGEMA_signal_4158, new_AGEMA_signal_4157, new_AGEMA_signal_4156, Midori_rounds_mul_input[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_51_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3522, new_AGEMA_signal_3521, new_AGEMA_signal_3520, Midori_rounds_SR_Result[51]}), .a ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, new_AGEMA_signal_3943, Midori_rounds_sub_ResultXORkey[51]}), .c ({new_AGEMA_signal_4164, new_AGEMA_signal_4163, new_AGEMA_signal_4162, Midori_rounds_mul_input[51]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_53_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3648, new_AGEMA_signal_3647, new_AGEMA_signal_3646, Midori_rounds_SR_Result[53]}), .a ({new_AGEMA_signal_3942, new_AGEMA_signal_3941, new_AGEMA_signal_3940, Midori_rounds_sub_ResultXORkey[53]}), .c ({new_AGEMA_signal_4167, new_AGEMA_signal_4166, new_AGEMA_signal_4165, Midori_rounds_mul_input[53]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_55_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3642, new_AGEMA_signal_3641, new_AGEMA_signal_3640, Midori_rounds_SR_Result[55]}), .a ({new_AGEMA_signal_3936, new_AGEMA_signal_3935, new_AGEMA_signal_3934, Midori_rounds_sub_ResultXORkey[55]}), .c ({new_AGEMA_signal_4173, new_AGEMA_signal_4172, new_AGEMA_signal_4171, Midori_rounds_mul_input[55]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_57_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3588, new_AGEMA_signal_3587, new_AGEMA_signal_3586, Midori_rounds_SR_Result[57]}), .a ({new_AGEMA_signal_3933, new_AGEMA_signal_3932, new_AGEMA_signal_3931, Midori_rounds_sub_ResultXORkey[57]}), .c ({new_AGEMA_signal_4176, new_AGEMA_signal_4175, new_AGEMA_signal_4174, Midori_rounds_mul_input[57]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_59_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3582, new_AGEMA_signal_3581, new_AGEMA_signal_3580, Midori_rounds_SR_Result[59]}), .a ({new_AGEMA_signal_3927, new_AGEMA_signal_3926, new_AGEMA_signal_3925, Midori_rounds_sub_ResultXORkey[59]}), .c ({new_AGEMA_signal_4182, new_AGEMA_signal_4181, new_AGEMA_signal_4180, Midori_rounds_mul_input[59]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_61_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3708, new_AGEMA_signal_3707, new_AGEMA_signal_3706, Midori_rounds_SR_Result[61]}), .a ({new_AGEMA_signal_3921, new_AGEMA_signal_3920, new_AGEMA_signal_3919, Midori_rounds_sub_ResultXORkey[61]}), .c ({new_AGEMA_signal_4185, new_AGEMA_signal_4184, new_AGEMA_signal_4183, Midori_rounds_mul_input[61]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_63_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3702, new_AGEMA_signal_3701, new_AGEMA_signal_3700, Midori_rounds_SR_Result[63]}), .a ({new_AGEMA_signal_3915, new_AGEMA_signal_3914, new_AGEMA_signal_3913, Midori_rounds_sub_ResultXORkey[63]}), .c ({new_AGEMA_signal_4191, new_AGEMA_signal_4190, new_AGEMA_signal_4189, Midori_rounds_mul_input[63]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U24 ( .a ({new_AGEMA_signal_4185, new_AGEMA_signal_4184, new_AGEMA_signal_4183, Midori_rounds_mul_input[61]}), .b ({new_AGEMA_signal_4203, new_AGEMA_signal_4202, new_AGEMA_signal_4201, Midori_rounds_mul_MC1_n8}), .c ({new_AGEMA_signal_4266, new_AGEMA_signal_4265, new_AGEMA_signal_4264, Midori_rounds_SR_Inv_Result[21]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U22 ( .a ({new_AGEMA_signal_4164, new_AGEMA_signal_4163, new_AGEMA_signal_4162, Midori_rounds_mul_input[51]}), .b ({new_AGEMA_signal_4194, new_AGEMA_signal_4193, new_AGEMA_signal_4192, Midori_rounds_mul_MC1_n6}), .c ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, new_AGEMA_signal_4267, Midori_rounds_SR_Inv_Result[43]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U20 ( .a ({new_AGEMA_signal_4158, new_AGEMA_signal_4157, new_AGEMA_signal_4156, Midori_rounds_mul_input[49]}), .b ({new_AGEMA_signal_4200, new_AGEMA_signal_4199, new_AGEMA_signal_4198, Midori_rounds_mul_MC1_n4}), .c ({new_AGEMA_signal_4275, new_AGEMA_signal_4274, new_AGEMA_signal_4273, Midori_rounds_SR_Inv_Result[41]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U18 ( .a ({new_AGEMA_signal_4173, new_AGEMA_signal_4172, new_AGEMA_signal_4171, Midori_rounds_mul_input[55]}), .b ({new_AGEMA_signal_4194, new_AGEMA_signal_4193, new_AGEMA_signal_4192, Midori_rounds_mul_MC1_n6}), .c ({new_AGEMA_signal_4278, new_AGEMA_signal_4277, new_AGEMA_signal_4276, Midori_rounds_SR_Inv_Result[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U17 ( .a ({new_AGEMA_signal_4191, new_AGEMA_signal_4190, new_AGEMA_signal_4189, Midori_rounds_mul_input[63]}), .b ({new_AGEMA_signal_4182, new_AGEMA_signal_4181, new_AGEMA_signal_4180, Midori_rounds_mul_input[59]}), .c ({new_AGEMA_signal_4194, new_AGEMA_signal_4193, new_AGEMA_signal_4192, Midori_rounds_mul_MC1_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U14 ( .a ({new_AGEMA_signal_4167, new_AGEMA_signal_4166, new_AGEMA_signal_4165, Midori_rounds_mul_input[53]}), .b ({new_AGEMA_signal_4200, new_AGEMA_signal_4199, new_AGEMA_signal_4198, Midori_rounds_mul_MC1_n4}), .c ({new_AGEMA_signal_4284, new_AGEMA_signal_4283, new_AGEMA_signal_4282, Midori_rounds_SR_Inv_Result[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U13 ( .a ({new_AGEMA_signal_4176, new_AGEMA_signal_4175, new_AGEMA_signal_4174, Midori_rounds_mul_input[57]}), .b ({new_AGEMA_signal_4185, new_AGEMA_signal_4184, new_AGEMA_signal_4183, Midori_rounds_mul_input[61]}), .c ({new_AGEMA_signal_4200, new_AGEMA_signal_4199, new_AGEMA_signal_4198, Midori_rounds_mul_MC1_n4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U12 ( .a ({new_AGEMA_signal_4182, new_AGEMA_signal_4181, new_AGEMA_signal_4180, Midori_rounds_mul_input[59]}), .b ({new_AGEMA_signal_4206, new_AGEMA_signal_4205, new_AGEMA_signal_4204, Midori_rounds_mul_MC1_n2}), .c ({new_AGEMA_signal_4287, new_AGEMA_signal_4286, new_AGEMA_signal_4285, Midori_rounds_SR_Inv_Result[63]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U10 ( .a ({new_AGEMA_signal_4176, new_AGEMA_signal_4175, new_AGEMA_signal_4174, Midori_rounds_mul_input[57]}), .b ({new_AGEMA_signal_4203, new_AGEMA_signal_4202, new_AGEMA_signal_4201, Midori_rounds_mul_MC1_n8}), .c ({new_AGEMA_signal_4293, new_AGEMA_signal_4292, new_AGEMA_signal_4291, Midori_rounds_SR_Inv_Result[61]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U9 ( .a ({new_AGEMA_signal_4158, new_AGEMA_signal_4157, new_AGEMA_signal_4156, Midori_rounds_mul_input[49]}), .b ({new_AGEMA_signal_4167, new_AGEMA_signal_4166, new_AGEMA_signal_4165, Midori_rounds_mul_input[53]}), .c ({new_AGEMA_signal_4203, new_AGEMA_signal_4202, new_AGEMA_signal_4201, Midori_rounds_mul_MC1_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U6 ( .a ({new_AGEMA_signal_4191, new_AGEMA_signal_4190, new_AGEMA_signal_4189, Midori_rounds_mul_input[63]}), .b ({new_AGEMA_signal_4206, new_AGEMA_signal_4205, new_AGEMA_signal_4204, Midori_rounds_mul_MC1_n2}), .c ({new_AGEMA_signal_4296, new_AGEMA_signal_4295, new_AGEMA_signal_4294, Midori_rounds_SR_Inv_Result[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U5 ( .a ({new_AGEMA_signal_4164, new_AGEMA_signal_4163, new_AGEMA_signal_4162, Midori_rounds_mul_input[51]}), .b ({new_AGEMA_signal_4173, new_AGEMA_signal_4172, new_AGEMA_signal_4171, Midori_rounds_mul_input[55]}), .c ({new_AGEMA_signal_4206, new_AGEMA_signal_4205, new_AGEMA_signal_4204, Midori_rounds_mul_MC1_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U24 ( .a ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, new_AGEMA_signal_4147, Midori_rounds_mul_input[45]}), .b ({new_AGEMA_signal_4221, new_AGEMA_signal_4220, new_AGEMA_signal_4219, Midori_rounds_mul_MC2_n8}), .c ({new_AGEMA_signal_4302, new_AGEMA_signal_4301, new_AGEMA_signal_4300, Midori_rounds_SR_Inv_Result[45]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U22 ( .a ({new_AGEMA_signal_4128, new_AGEMA_signal_4127, new_AGEMA_signal_4126, Midori_rounds_mul_input[35]}), .b ({new_AGEMA_signal_4212, new_AGEMA_signal_4211, new_AGEMA_signal_4210, Midori_rounds_mul_MC2_n6}), .c ({new_AGEMA_signal_4305, new_AGEMA_signal_4304, new_AGEMA_signal_4303, Midori_rounds_SR_Inv_Result[19]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U20 ( .a ({new_AGEMA_signal_4122, new_AGEMA_signal_4121, new_AGEMA_signal_4120, Midori_rounds_mul_input[33]}), .b ({new_AGEMA_signal_4218, new_AGEMA_signal_4217, new_AGEMA_signal_4216, Midori_rounds_mul_MC2_n4}), .c ({new_AGEMA_signal_4311, new_AGEMA_signal_4310, new_AGEMA_signal_4309, Midori_rounds_SR_Inv_Result[17]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U18 ( .a ({new_AGEMA_signal_4137, new_AGEMA_signal_4136, new_AGEMA_signal_4135, Midori_rounds_mul_input[39]}), .b ({new_AGEMA_signal_4212, new_AGEMA_signal_4211, new_AGEMA_signal_4210, Midori_rounds_mul_MC2_n6}), .c ({new_AGEMA_signal_4314, new_AGEMA_signal_4313, new_AGEMA_signal_4312, Midori_rounds_SR_Inv_Result[59]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U17 ( .a ({new_AGEMA_signal_4155, new_AGEMA_signal_4154, new_AGEMA_signal_4153, Midori_rounds_mul_input[47]}), .b ({new_AGEMA_signal_4146, new_AGEMA_signal_4145, new_AGEMA_signal_4144, Midori_rounds_mul_input[43]}), .c ({new_AGEMA_signal_4212, new_AGEMA_signal_4211, new_AGEMA_signal_4210, Midori_rounds_mul_MC2_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U14 ( .a ({new_AGEMA_signal_4131, new_AGEMA_signal_4130, new_AGEMA_signal_4129, Midori_rounds_mul_input[37]}), .b ({new_AGEMA_signal_4218, new_AGEMA_signal_4217, new_AGEMA_signal_4216, Midori_rounds_mul_MC2_n4}), .c ({new_AGEMA_signal_4320, new_AGEMA_signal_4319, new_AGEMA_signal_4318, Midori_rounds_SR_Inv_Result[57]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U13 ( .a ({new_AGEMA_signal_4140, new_AGEMA_signal_4139, new_AGEMA_signal_4138, Midori_rounds_mul_input[41]}), .b ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, new_AGEMA_signal_4147, Midori_rounds_mul_input[45]}), .c ({new_AGEMA_signal_4218, new_AGEMA_signal_4217, new_AGEMA_signal_4216, Midori_rounds_mul_MC2_n4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U12 ( .a ({new_AGEMA_signal_4146, new_AGEMA_signal_4145, new_AGEMA_signal_4144, Midori_rounds_mul_input[43]}), .b ({new_AGEMA_signal_4224, new_AGEMA_signal_4223, new_AGEMA_signal_4222, Midori_rounds_mul_MC2_n2}), .c ({new_AGEMA_signal_4323, new_AGEMA_signal_4322, new_AGEMA_signal_4321, Midori_rounds_SR_Inv_Result[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U10 ( .a ({new_AGEMA_signal_4140, new_AGEMA_signal_4139, new_AGEMA_signal_4138, Midori_rounds_mul_input[41]}), .b ({new_AGEMA_signal_4221, new_AGEMA_signal_4220, new_AGEMA_signal_4219, Midori_rounds_mul_MC2_n8}), .c ({new_AGEMA_signal_4329, new_AGEMA_signal_4328, new_AGEMA_signal_4327, Midori_rounds_SR_Inv_Result[5]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U9 ( .a ({new_AGEMA_signal_4122, new_AGEMA_signal_4121, new_AGEMA_signal_4120, Midori_rounds_mul_input[33]}), .b ({new_AGEMA_signal_4131, new_AGEMA_signal_4130, new_AGEMA_signal_4129, Midori_rounds_mul_input[37]}), .c ({new_AGEMA_signal_4221, new_AGEMA_signal_4220, new_AGEMA_signal_4219, Midori_rounds_mul_MC2_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U6 ( .a ({new_AGEMA_signal_4155, new_AGEMA_signal_4154, new_AGEMA_signal_4153, Midori_rounds_mul_input[47]}), .b ({new_AGEMA_signal_4224, new_AGEMA_signal_4223, new_AGEMA_signal_4222, Midori_rounds_mul_MC2_n2}), .c ({new_AGEMA_signal_4332, new_AGEMA_signal_4331, new_AGEMA_signal_4330, Midori_rounds_SR_Inv_Result[47]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U5 ( .a ({new_AGEMA_signal_4128, new_AGEMA_signal_4127, new_AGEMA_signal_4126, Midori_rounds_mul_input[35]}), .b ({new_AGEMA_signal_4137, new_AGEMA_signal_4136, new_AGEMA_signal_4135, Midori_rounds_mul_input[39]}), .c ({new_AGEMA_signal_4224, new_AGEMA_signal_4223, new_AGEMA_signal_4222, Midori_rounds_mul_MC2_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U24 ( .a ({new_AGEMA_signal_4113, new_AGEMA_signal_4112, new_AGEMA_signal_4111, Midori_rounds_mul_input[29]}), .b ({new_AGEMA_signal_4239, new_AGEMA_signal_4238, new_AGEMA_signal_4237, Midori_rounds_mul_MC3_n8}), .c ({new_AGEMA_signal_4338, new_AGEMA_signal_4337, new_AGEMA_signal_4336, Midori_rounds_SR_Inv_Result[49]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U22 ( .a ({new_AGEMA_signal_4092, new_AGEMA_signal_4091, new_AGEMA_signal_4090, Midori_rounds_mul_input[19]}), .b ({new_AGEMA_signal_4230, new_AGEMA_signal_4229, new_AGEMA_signal_4228, Midori_rounds_mul_MC3_n6}), .c ({new_AGEMA_signal_4341, new_AGEMA_signal_4340, new_AGEMA_signal_4339, Midori_rounds_SR_Inv_Result[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U20 ( .a ({new_AGEMA_signal_4086, new_AGEMA_signal_4085, new_AGEMA_signal_4084, Midori_rounds_mul_input[17]}), .b ({new_AGEMA_signal_4236, new_AGEMA_signal_4235, new_AGEMA_signal_4234, Midori_rounds_mul_MC3_n4}), .c ({new_AGEMA_signal_4347, new_AGEMA_signal_4346, new_AGEMA_signal_4345, Midori_rounds_SR_Inv_Result[13]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U18 ( .a ({new_AGEMA_signal_4101, new_AGEMA_signal_4100, new_AGEMA_signal_4099, Midori_rounds_mul_input[23]}), .b ({new_AGEMA_signal_4230, new_AGEMA_signal_4229, new_AGEMA_signal_4228, Midori_rounds_mul_MC3_n6}), .c ({new_AGEMA_signal_4350, new_AGEMA_signal_4349, new_AGEMA_signal_4348, Midori_rounds_SR_Inv_Result[39]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U17 ( .a ({new_AGEMA_signal_4119, new_AGEMA_signal_4118, new_AGEMA_signal_4117, Midori_rounds_mul_input[31]}), .b ({new_AGEMA_signal_4110, new_AGEMA_signal_4109, new_AGEMA_signal_4108, Midori_rounds_mul_input[27]}), .c ({new_AGEMA_signal_4230, new_AGEMA_signal_4229, new_AGEMA_signal_4228, Midori_rounds_mul_MC3_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U14 ( .a ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, new_AGEMA_signal_4093, Midori_rounds_mul_input[21]}), .b ({new_AGEMA_signal_4236, new_AGEMA_signal_4235, new_AGEMA_signal_4234, Midori_rounds_mul_MC3_n4}), .c ({new_AGEMA_signal_4356, new_AGEMA_signal_4355, new_AGEMA_signal_4354, Midori_rounds_SR_Inv_Result[37]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U13 ( .a ({new_AGEMA_signal_4104, new_AGEMA_signal_4103, new_AGEMA_signal_4102, Midori_rounds_mul_input[25]}), .b ({new_AGEMA_signal_4113, new_AGEMA_signal_4112, new_AGEMA_signal_4111, Midori_rounds_mul_input[29]}), .c ({new_AGEMA_signal_4236, new_AGEMA_signal_4235, new_AGEMA_signal_4234, Midori_rounds_mul_MC3_n4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U12 ( .a ({new_AGEMA_signal_4110, new_AGEMA_signal_4109, new_AGEMA_signal_4108, Midori_rounds_mul_input[27]}), .b ({new_AGEMA_signal_4242, new_AGEMA_signal_4241, new_AGEMA_signal_4240, Midori_rounds_mul_MC3_n2}), .c ({new_AGEMA_signal_4359, new_AGEMA_signal_4358, new_AGEMA_signal_4357, Midori_rounds_SR_Inv_Result[27]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U10 ( .a ({new_AGEMA_signal_4104, new_AGEMA_signal_4103, new_AGEMA_signal_4102, Midori_rounds_mul_input[25]}), .b ({new_AGEMA_signal_4239, new_AGEMA_signal_4238, new_AGEMA_signal_4237, Midori_rounds_mul_MC3_n8}), .c ({new_AGEMA_signal_4365, new_AGEMA_signal_4364, new_AGEMA_signal_4363, Midori_rounds_SR_Inv_Result[25]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U9 ( .a ({new_AGEMA_signal_4086, new_AGEMA_signal_4085, new_AGEMA_signal_4084, Midori_rounds_mul_input[17]}), .b ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, new_AGEMA_signal_4093, Midori_rounds_mul_input[21]}), .c ({new_AGEMA_signal_4239, new_AGEMA_signal_4238, new_AGEMA_signal_4237, Midori_rounds_mul_MC3_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U6 ( .a ({new_AGEMA_signal_4119, new_AGEMA_signal_4118, new_AGEMA_signal_4117, Midori_rounds_mul_input[31]}), .b ({new_AGEMA_signal_4242, new_AGEMA_signal_4241, new_AGEMA_signal_4240, Midori_rounds_mul_MC3_n2}), .c ({new_AGEMA_signal_4368, new_AGEMA_signal_4367, new_AGEMA_signal_4366, Midori_rounds_SR_Inv_Result[51]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U5 ( .a ({new_AGEMA_signal_4092, new_AGEMA_signal_4091, new_AGEMA_signal_4090, Midori_rounds_mul_input[19]}), .b ({new_AGEMA_signal_4101, new_AGEMA_signal_4100, new_AGEMA_signal_4099, Midori_rounds_mul_input[23]}), .c ({new_AGEMA_signal_4242, new_AGEMA_signal_4241, new_AGEMA_signal_4240, Midori_rounds_mul_MC3_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U24 ( .a ({new_AGEMA_signal_4077, new_AGEMA_signal_4076, new_AGEMA_signal_4075, Midori_rounds_mul_input[13]}), .b ({new_AGEMA_signal_4257, new_AGEMA_signal_4256, new_AGEMA_signal_4255, Midori_rounds_mul_MC4_n8}), .c ({new_AGEMA_signal_4374, new_AGEMA_signal_4373, new_AGEMA_signal_4372, Midori_rounds_SR_Inv_Result[9]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U22 ( .a ({new_AGEMA_signal_4056, new_AGEMA_signal_4055, new_AGEMA_signal_4054, Midori_rounds_mul_input[3]}), .b ({new_AGEMA_signal_4248, new_AGEMA_signal_4247, new_AGEMA_signal_4246, Midori_rounds_mul_MC4_n6}), .c ({new_AGEMA_signal_4377, new_AGEMA_signal_4376, new_AGEMA_signal_4375, Midori_rounds_SR_Inv_Result[55]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U20 ( .a ({new_AGEMA_signal_4050, new_AGEMA_signal_4049, new_AGEMA_signal_4048, Midori_rounds_mul_input[1]}), .b ({new_AGEMA_signal_4254, new_AGEMA_signal_4253, new_AGEMA_signal_4252, Midori_rounds_mul_MC4_n4}), .c ({new_AGEMA_signal_4383, new_AGEMA_signal_4382, new_AGEMA_signal_4381, Midori_rounds_SR_Inv_Result[53]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U18 ( .a ({new_AGEMA_signal_4065, new_AGEMA_signal_4064, new_AGEMA_signal_4063, Midori_rounds_mul_input[7]}), .b ({new_AGEMA_signal_4248, new_AGEMA_signal_4247, new_AGEMA_signal_4246, Midori_rounds_mul_MC4_n6}), .c ({new_AGEMA_signal_4386, new_AGEMA_signal_4385, new_AGEMA_signal_4384, Midori_rounds_SR_Inv_Result[31]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U17 ( .a ({new_AGEMA_signal_4083, new_AGEMA_signal_4082, new_AGEMA_signal_4081, Midori_rounds_mul_input[15]}), .b ({new_AGEMA_signal_4074, new_AGEMA_signal_4073, new_AGEMA_signal_4072, Midori_rounds_mul_input[11]}), .c ({new_AGEMA_signal_4248, new_AGEMA_signal_4247, new_AGEMA_signal_4246, Midori_rounds_mul_MC4_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U14 ( .a ({new_AGEMA_signal_4059, new_AGEMA_signal_4058, new_AGEMA_signal_4057, Midori_rounds_mul_input[5]}), .b ({new_AGEMA_signal_4254, new_AGEMA_signal_4253, new_AGEMA_signal_4252, Midori_rounds_mul_MC4_n4}), .c ({new_AGEMA_signal_4392, new_AGEMA_signal_4391, new_AGEMA_signal_4390, Midori_rounds_SR_Inv_Result[29]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U13 ( .a ({new_AGEMA_signal_4068, new_AGEMA_signal_4067, new_AGEMA_signal_4066, Midori_rounds_mul_input[9]}), .b ({new_AGEMA_signal_4077, new_AGEMA_signal_4076, new_AGEMA_signal_4075, Midori_rounds_mul_input[13]}), .c ({new_AGEMA_signal_4254, new_AGEMA_signal_4253, new_AGEMA_signal_4252, Midori_rounds_mul_MC4_n4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U12 ( .a ({new_AGEMA_signal_4074, new_AGEMA_signal_4073, new_AGEMA_signal_4072, Midori_rounds_mul_input[11]}), .b ({new_AGEMA_signal_4260, new_AGEMA_signal_4259, new_AGEMA_signal_4258, Midori_rounds_mul_MC4_n2}), .c ({new_AGEMA_signal_4395, new_AGEMA_signal_4394, new_AGEMA_signal_4393, Midori_rounds_SR_Inv_Result[35]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U10 ( .a ({new_AGEMA_signal_4068, new_AGEMA_signal_4067, new_AGEMA_signal_4066, Midori_rounds_mul_input[9]}), .b ({new_AGEMA_signal_4257, new_AGEMA_signal_4256, new_AGEMA_signal_4255, Midori_rounds_mul_MC4_n8}), .c ({new_AGEMA_signal_4401, new_AGEMA_signal_4400, new_AGEMA_signal_4399, Midori_rounds_SR_Inv_Result[33]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U9 ( .a ({new_AGEMA_signal_4050, new_AGEMA_signal_4049, new_AGEMA_signal_4048, Midori_rounds_mul_input[1]}), .b ({new_AGEMA_signal_4059, new_AGEMA_signal_4058, new_AGEMA_signal_4057, Midori_rounds_mul_input[5]}), .c ({new_AGEMA_signal_4257, new_AGEMA_signal_4256, new_AGEMA_signal_4255, Midori_rounds_mul_MC4_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U6 ( .a ({new_AGEMA_signal_4083, new_AGEMA_signal_4082, new_AGEMA_signal_4081, Midori_rounds_mul_input[15]}), .b ({new_AGEMA_signal_4260, new_AGEMA_signal_4259, new_AGEMA_signal_4258, Midori_rounds_mul_MC4_n2}), .c ({new_AGEMA_signal_4404, new_AGEMA_signal_4403, new_AGEMA_signal_4402, Midori_rounds_SR_Inv_Result[11]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U5 ( .a ({new_AGEMA_signal_4056, new_AGEMA_signal_4055, new_AGEMA_signal_4054, Midori_rounds_mul_input[3]}), .b ({new_AGEMA_signal_4065, new_AGEMA_signal_4064, new_AGEMA_signal_4063, Midori_rounds_mul_input[7]}), .c ({new_AGEMA_signal_4260, new_AGEMA_signal_4259, new_AGEMA_signal_4258, Midori_rounds_mul_MC4_n2}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_1_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4539, new_AGEMA_signal_4538, new_AGEMA_signal_4537, Midori_rounds_mul_ResultXORkey[1]}), .a ({new_AGEMA_signal_4284, new_AGEMA_signal_4283, new_AGEMA_signal_4282, Midori_rounds_SR_Inv_Result[1]}), .c ({new_AGEMA_signal_4608, new_AGEMA_signal_4607, new_AGEMA_signal_4606, Midori_rounds_round_Result[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_3_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4482, new_AGEMA_signal_4481, new_AGEMA_signal_4480, Midori_rounds_mul_ResultXORkey[3]}), .a ({new_AGEMA_signal_4278, new_AGEMA_signal_4277, new_AGEMA_signal_4276, Midori_rounds_SR_Inv_Result[3]}), .c ({new_AGEMA_signal_4614, new_AGEMA_signal_4613, new_AGEMA_signal_4612, Midori_rounds_round_Result[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_5_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4431, new_AGEMA_signal_4430, new_AGEMA_signal_4429, Midori_rounds_mul_ResultXORkey[5]}), .a ({new_AGEMA_signal_4329, new_AGEMA_signal_4328, new_AGEMA_signal_4327, Midori_rounds_SR_Inv_Result[5]}), .c ({new_AGEMA_signal_4617, new_AGEMA_signal_4616, new_AGEMA_signal_4615, Midori_rounds_round_Result[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_7_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4416, new_AGEMA_signal_4415, new_AGEMA_signal_4414, Midori_rounds_mul_ResultXORkey[7]}), .a ({new_AGEMA_signal_4323, new_AGEMA_signal_4322, new_AGEMA_signal_4321, Midori_rounds_SR_Inv_Result[7]}), .c ({new_AGEMA_signal_4623, new_AGEMA_signal_4622, new_AGEMA_signal_4621, Midori_rounds_round_Result[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_9_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4410, new_AGEMA_signal_4409, new_AGEMA_signal_4408, Midori_rounds_mul_ResultXORkey[9]}), .a ({new_AGEMA_signal_4374, new_AGEMA_signal_4373, new_AGEMA_signal_4372, Midori_rounds_SR_Inv_Result[9]}), .c ({new_AGEMA_signal_4626, new_AGEMA_signal_4625, new_AGEMA_signal_4624, Midori_rounds_round_Result[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_11_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4560, new_AGEMA_signal_4559, new_AGEMA_signal_4558, Midori_rounds_mul_ResultXORkey[11]}), .a ({new_AGEMA_signal_4404, new_AGEMA_signal_4403, new_AGEMA_signal_4402, Midori_rounds_SR_Inv_Result[11]}), .c ({new_AGEMA_signal_4632, new_AGEMA_signal_4631, new_AGEMA_signal_4630, Midori_rounds_round_Result[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_13_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, new_AGEMA_signal_4555, Midori_rounds_mul_ResultXORkey[13]}), .a ({new_AGEMA_signal_4347, new_AGEMA_signal_4346, new_AGEMA_signal_4345, Midori_rounds_SR_Inv_Result[13]}), .c ({new_AGEMA_signal_4635, new_AGEMA_signal_4634, new_AGEMA_signal_4633, Midori_rounds_round_Result[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_15_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4551, new_AGEMA_signal_4550, new_AGEMA_signal_4549, Midori_rounds_mul_ResultXORkey[15]}), .a ({new_AGEMA_signal_4341, new_AGEMA_signal_4340, new_AGEMA_signal_4339, Midori_rounds_SR_Inv_Result[15]}), .c ({new_AGEMA_signal_4641, new_AGEMA_signal_4640, new_AGEMA_signal_4639, Midori_rounds_round_Result[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_17_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4548, new_AGEMA_signal_4547, new_AGEMA_signal_4546, Midori_rounds_mul_ResultXORkey[17]}), .a ({new_AGEMA_signal_4311, new_AGEMA_signal_4310, new_AGEMA_signal_4309, Midori_rounds_SR_Inv_Result[17]}), .c ({new_AGEMA_signal_4644, new_AGEMA_signal_4643, new_AGEMA_signal_4642, Midori_rounds_round_Result[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_19_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4542, new_AGEMA_signal_4541, new_AGEMA_signal_4540, Midori_rounds_mul_ResultXORkey[19]}), .a ({new_AGEMA_signal_4305, new_AGEMA_signal_4304, new_AGEMA_signal_4303, Midori_rounds_SR_Inv_Result[19]}), .c ({new_AGEMA_signal_4650, new_AGEMA_signal_4649, new_AGEMA_signal_4648, Midori_rounds_round_Result[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_21_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4533, new_AGEMA_signal_4532, new_AGEMA_signal_4531, Midori_rounds_mul_ResultXORkey[21]}), .a ({new_AGEMA_signal_4266, new_AGEMA_signal_4265, new_AGEMA_signal_4264, Midori_rounds_SR_Inv_Result[21]}), .c ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, new_AGEMA_signal_4651, Midori_rounds_round_Result[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_23_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4527, new_AGEMA_signal_4526, new_AGEMA_signal_4525, Midori_rounds_mul_ResultXORkey[23]}), .a ({new_AGEMA_signal_4296, new_AGEMA_signal_4295, new_AGEMA_signal_4294, Midori_rounds_SR_Inv_Result[23]}), .c ({new_AGEMA_signal_4659, new_AGEMA_signal_4658, new_AGEMA_signal_4657, Midori_rounds_round_Result[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_25_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4524, new_AGEMA_signal_4523, new_AGEMA_signal_4522, Midori_rounds_mul_ResultXORkey[25]}), .a ({new_AGEMA_signal_4365, new_AGEMA_signal_4364, new_AGEMA_signal_4363, Midori_rounds_SR_Inv_Result[25]}), .c ({new_AGEMA_signal_4662, new_AGEMA_signal_4661, new_AGEMA_signal_4660, Midori_rounds_round_Result[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_27_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4518, new_AGEMA_signal_4517, new_AGEMA_signal_4516, Midori_rounds_mul_ResultXORkey[27]}), .a ({new_AGEMA_signal_4359, new_AGEMA_signal_4358, new_AGEMA_signal_4357, Midori_rounds_SR_Inv_Result[27]}), .c ({new_AGEMA_signal_4668, new_AGEMA_signal_4667, new_AGEMA_signal_4666, Midori_rounds_round_Result[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_29_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4515, new_AGEMA_signal_4514, new_AGEMA_signal_4513, Midori_rounds_mul_ResultXORkey[29]}), .a ({new_AGEMA_signal_4392, new_AGEMA_signal_4391, new_AGEMA_signal_4390, Midori_rounds_SR_Inv_Result[29]}), .c ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, new_AGEMA_signal_4669, Midori_rounds_round_Result[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_31_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4506, new_AGEMA_signal_4505, new_AGEMA_signal_4504, Midori_rounds_mul_ResultXORkey[31]}), .a ({new_AGEMA_signal_4386, new_AGEMA_signal_4385, new_AGEMA_signal_4384, Midori_rounds_SR_Inv_Result[31]}), .c ({new_AGEMA_signal_4677, new_AGEMA_signal_4676, new_AGEMA_signal_4675, Midori_rounds_round_Result[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_33_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4503, new_AGEMA_signal_4502, new_AGEMA_signal_4501, Midori_rounds_mul_ResultXORkey[33]}), .a ({new_AGEMA_signal_4401, new_AGEMA_signal_4400, new_AGEMA_signal_4399, Midori_rounds_SR_Inv_Result[33]}), .c ({new_AGEMA_signal_4680, new_AGEMA_signal_4679, new_AGEMA_signal_4678, Midori_rounds_round_Result[33]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_35_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4497, new_AGEMA_signal_4496, new_AGEMA_signal_4495, Midori_rounds_mul_ResultXORkey[35]}), .a ({new_AGEMA_signal_4395, new_AGEMA_signal_4394, new_AGEMA_signal_4393, Midori_rounds_SR_Inv_Result[35]}), .c ({new_AGEMA_signal_4686, new_AGEMA_signal_4685, new_AGEMA_signal_4684, Midori_rounds_round_Result[35]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_37_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4491, new_AGEMA_signal_4490, new_AGEMA_signal_4489, Midori_rounds_mul_ResultXORkey[37]}), .a ({new_AGEMA_signal_4356, new_AGEMA_signal_4355, new_AGEMA_signal_4354, Midori_rounds_SR_Inv_Result[37]}), .c ({new_AGEMA_signal_4689, new_AGEMA_signal_4688, new_AGEMA_signal_4687, Midori_rounds_round_Result[37]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_39_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4485, new_AGEMA_signal_4484, new_AGEMA_signal_4483, Midori_rounds_mul_ResultXORkey[39]}), .a ({new_AGEMA_signal_4350, new_AGEMA_signal_4349, new_AGEMA_signal_4348, Midori_rounds_SR_Inv_Result[39]}), .c ({new_AGEMA_signal_4695, new_AGEMA_signal_4694, new_AGEMA_signal_4693, Midori_rounds_round_Result[39]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_41_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4479, new_AGEMA_signal_4478, new_AGEMA_signal_4477, Midori_rounds_mul_ResultXORkey[41]}), .a ({new_AGEMA_signal_4275, new_AGEMA_signal_4274, new_AGEMA_signal_4273, Midori_rounds_SR_Inv_Result[41]}), .c ({new_AGEMA_signal_4698, new_AGEMA_signal_4697, new_AGEMA_signal_4696, Midori_rounds_round_Result[41]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_43_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4473, new_AGEMA_signal_4472, new_AGEMA_signal_4471, Midori_rounds_mul_ResultXORkey[43]}), .a ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, new_AGEMA_signal_4267, Midori_rounds_SR_Inv_Result[43]}), .c ({new_AGEMA_signal_4704, new_AGEMA_signal_4703, new_AGEMA_signal_4702, Midori_rounds_round_Result[43]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_45_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4467, new_AGEMA_signal_4466, new_AGEMA_signal_4465, Midori_rounds_mul_ResultXORkey[45]}), .a ({new_AGEMA_signal_4302, new_AGEMA_signal_4301, new_AGEMA_signal_4300, Midori_rounds_SR_Inv_Result[45]}), .c ({new_AGEMA_signal_4707, new_AGEMA_signal_4706, new_AGEMA_signal_4705, Midori_rounds_round_Result[45]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_47_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4461, new_AGEMA_signal_4460, new_AGEMA_signal_4459, Midori_rounds_mul_ResultXORkey[47]}), .a ({new_AGEMA_signal_4332, new_AGEMA_signal_4331, new_AGEMA_signal_4330, Midori_rounds_SR_Inv_Result[47]}), .c ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, new_AGEMA_signal_4711, Midori_rounds_round_Result[47]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_49_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4458, new_AGEMA_signal_4457, new_AGEMA_signal_4456, Midori_rounds_mul_ResultXORkey[49]}), .a ({new_AGEMA_signal_4338, new_AGEMA_signal_4337, new_AGEMA_signal_4336, Midori_rounds_SR_Inv_Result[49]}), .c ({new_AGEMA_signal_4716, new_AGEMA_signal_4715, new_AGEMA_signal_4714, Midori_rounds_round_Result[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_51_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4452, new_AGEMA_signal_4451, new_AGEMA_signal_4450, Midori_rounds_mul_ResultXORkey[51]}), .a ({new_AGEMA_signal_4368, new_AGEMA_signal_4367, new_AGEMA_signal_4366, Midori_rounds_SR_Inv_Result[51]}), .c ({new_AGEMA_signal_4722, new_AGEMA_signal_4721, new_AGEMA_signal_4720, Midori_rounds_round_Result[51]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_53_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4449, new_AGEMA_signal_4448, new_AGEMA_signal_4447, Midori_rounds_mul_ResultXORkey[53]}), .a ({new_AGEMA_signal_4383, new_AGEMA_signal_4382, new_AGEMA_signal_4381, Midori_rounds_SR_Inv_Result[53]}), .c ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, new_AGEMA_signal_4723, Midori_rounds_round_Result[53]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_55_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4443, new_AGEMA_signal_4442, new_AGEMA_signal_4441, Midori_rounds_mul_ResultXORkey[55]}), .a ({new_AGEMA_signal_4377, new_AGEMA_signal_4376, new_AGEMA_signal_4375, Midori_rounds_SR_Inv_Result[55]}), .c ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, new_AGEMA_signal_4729, Midori_rounds_round_Result[55]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_57_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4440, new_AGEMA_signal_4439, new_AGEMA_signal_4438, Midori_rounds_mul_ResultXORkey[57]}), .a ({new_AGEMA_signal_4320, new_AGEMA_signal_4319, new_AGEMA_signal_4318, Midori_rounds_SR_Inv_Result[57]}), .c ({new_AGEMA_signal_4734, new_AGEMA_signal_4733, new_AGEMA_signal_4732, Midori_rounds_round_Result[57]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_59_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4434, new_AGEMA_signal_4433, new_AGEMA_signal_4432, Midori_rounds_mul_ResultXORkey[59]}), .a ({new_AGEMA_signal_4314, new_AGEMA_signal_4313, new_AGEMA_signal_4312, Midori_rounds_SR_Inv_Result[59]}), .c ({new_AGEMA_signal_4740, new_AGEMA_signal_4739, new_AGEMA_signal_4738, Midori_rounds_round_Result[59]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_61_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4428, new_AGEMA_signal_4427, new_AGEMA_signal_4426, Midori_rounds_mul_ResultXORkey[61]}), .a ({new_AGEMA_signal_4293, new_AGEMA_signal_4292, new_AGEMA_signal_4291, Midori_rounds_SR_Inv_Result[61]}), .c ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, new_AGEMA_signal_4741, Midori_rounds_round_Result[61]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_63_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4422, new_AGEMA_signal_4421, new_AGEMA_signal_4420, Midori_rounds_mul_ResultXORkey[63]}), .a ({new_AGEMA_signal_4287, new_AGEMA_signal_4286, new_AGEMA_signal_4285, Midori_rounds_SR_Inv_Result[63]}), .c ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, new_AGEMA_signal_4747, Midori_rounds_round_Result[63]}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U127 ( .a ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, new_AGEMA_signal_1471, wk[8]}), .b ({new_AGEMA_signal_3555, new_AGEMA_signal_3554, new_AGEMA_signal_3553, Midori_rounds_SR_Result[8]}), .c ({DataOut_s3[8], DataOut_s2[8], DataOut_s1[8], DataOut_s0[8]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U125 ( .a ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, new_AGEMA_signal_1489, wk[6]}), .b ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, new_AGEMA_signal_3535, Midori_rounds_SR_Result[46]}), .c ({DataOut_s3[6], DataOut_s2[6], DataOut_s1[6], DataOut_s0[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U123 ( .a ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, new_AGEMA_signal_1507, wk[62]}), .b ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, new_AGEMA_signal_3703, Midori_rounds_SR_Result[62]}), .c ({DataOut_s3[62], DataOut_s2[62], DataOut_s1[62], DataOut_s0[62]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U121 ( .a ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, new_AGEMA_signal_1525, wk[60]}), .b ({new_AGEMA_signal_3711, new_AGEMA_signal_3710, new_AGEMA_signal_3709, Midori_rounds_SR_Result[60]}), .c ({DataOut_s3[60], DataOut_s2[60], DataOut_s1[60], DataOut_s0[60]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U118 ( .a ({new_AGEMA_signal_1554, new_AGEMA_signal_1553, new_AGEMA_signal_1552, wk[58]}), .b ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, new_AGEMA_signal_3691, Midori_rounds_SR_Result[34]}), .c ({DataOut_s3[58], DataOut_s2[58], DataOut_s1[58], DataOut_s0[58]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U116 ( .a ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, new_AGEMA_signal_1570, wk[56]}), .b ({new_AGEMA_signal_3699, new_AGEMA_signal_3698, new_AGEMA_signal_3697, Midori_rounds_SR_Result[32]}), .c ({DataOut_s3[56], DataOut_s2[56], DataOut_s1[56], DataOut_s0[56]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U114 ( .a ({new_AGEMA_signal_1590, new_AGEMA_signal_1589, new_AGEMA_signal_1588, wk[54]}), .b ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, new_AGEMA_signal_3679, Midori_rounds_SR_Result[6]}), .c ({DataOut_s3[54], DataOut_s2[54], DataOut_s1[54], DataOut_s0[54]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U112 ( .a ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, new_AGEMA_signal_1606, wk[52]}), .b ({new_AGEMA_signal_3687, new_AGEMA_signal_3686, new_AGEMA_signal_3685, Midori_rounds_SR_Result[4]}), .c ({DataOut_s3[52], DataOut_s2[52], DataOut_s1[52], DataOut_s0[52]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U110 ( .a ({new_AGEMA_signal_1626, new_AGEMA_signal_1625, new_AGEMA_signal_1624, wk[50]}), .b ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, new_AGEMA_signal_3667, Midori_rounds_SR_Result[26]}), .c ({DataOut_s3[50], DataOut_s2[50], DataOut_s1[50], DataOut_s0[50]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U109 ( .a ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, new_AGEMA_signal_1633, wk[4]}), .b ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, new_AGEMA_signal_3541, Midori_rounds_SR_Result[44]}), .c ({DataOut_s3[4], DataOut_s2[4], DataOut_s1[4], DataOut_s0[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U107 ( .a ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, new_AGEMA_signal_1651, wk[48]}), .b ({new_AGEMA_signal_3675, new_AGEMA_signal_3674, new_AGEMA_signal_3673, Midori_rounds_SR_Result[24]}), .c ({DataOut_s3[48], DataOut_s2[48], DataOut_s1[48], DataOut_s0[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U105 ( .a ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, new_AGEMA_signal_1669, wk[46]}), .b ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, new_AGEMA_signal_3655, Midori_rounds_SR_Result[42]}), .c ({DataOut_s3[46], DataOut_s2[46], DataOut_s1[46], DataOut_s0[46]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U103 ( .a ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, new_AGEMA_signal_1687, wk[44]}), .b ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, new_AGEMA_signal_3661, Midori_rounds_SR_Result[40]}), .c ({DataOut_s3[44], DataOut_s2[44], DataOut_s1[44], DataOut_s0[44]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U101 ( .a ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, new_AGEMA_signal_1705, wk[42]}), .b ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, new_AGEMA_signal_3643, Midori_rounds_SR_Result[54]}), .c ({DataOut_s3[42], DataOut_s2[42], DataOut_s1[42], DataOut_s0[42]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U99 ( .a ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, new_AGEMA_signal_1723, wk[40]}), .b ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, new_AGEMA_signal_3649, Midori_rounds_SR_Result[52]}), .c ({DataOut_s3[40], DataOut_s2[40], DataOut_s1[40], DataOut_s0[40]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U96 ( .a ({new_AGEMA_signal_1752, new_AGEMA_signal_1751, new_AGEMA_signal_1750, wk[38]}), .b ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, new_AGEMA_signal_3631, Midori_rounds_SR_Result[18]}), .c ({DataOut_s3[38], DataOut_s2[38], DataOut_s1[38], DataOut_s0[38]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U94 ( .a ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, new_AGEMA_signal_1768, wk[36]}), .b ({new_AGEMA_signal_3639, new_AGEMA_signal_3638, new_AGEMA_signal_3637, Midori_rounds_SR_Result[16]}), .c ({DataOut_s3[36], DataOut_s2[36], DataOut_s1[36], DataOut_s0[36]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U92 ( .a ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, new_AGEMA_signal_1786, wk[34]}), .b ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, new_AGEMA_signal_3619, Midori_rounds_SR_Result[14]}), .c ({DataOut_s3[34], DataOut_s2[34], DataOut_s1[34], DataOut_s0[34]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U90 ( .a ({new_AGEMA_signal_1806, new_AGEMA_signal_1805, new_AGEMA_signal_1804, wk[32]}), .b ({new_AGEMA_signal_3627, new_AGEMA_signal_3626, new_AGEMA_signal_3625, Midori_rounds_SR_Result[12]}), .c ({DataOut_s3[32], DataOut_s2[32], DataOut_s1[32], DataOut_s0[32]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U88 ( .a ({new_AGEMA_signal_1824, new_AGEMA_signal_1823, new_AGEMA_signal_1822, wk[30]}), .b ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, new_AGEMA_signal_3607, Midori_rounds_SR_Result[2]}), .c ({DataOut_s3[30], DataOut_s2[30], DataOut_s1[30], DataOut_s0[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U87 ( .a ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, new_AGEMA_signal_1831, wk[2]}), .b ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, new_AGEMA_signal_3523, Midori_rounds_SR_Result[50]}), .c ({DataOut_s3[2], DataOut_s2[2], DataOut_s1[2], DataOut_s0[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U85 ( .a ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, new_AGEMA_signal_1849, wk[28]}), .b ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, new_AGEMA_signal_3613, Midori_rounds_SR_Result[0]}), .c ({DataOut_s3[28], DataOut_s2[28], DataOut_s1[28], DataOut_s0[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U83 ( .a ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, new_AGEMA_signal_1867, wk[26]}), .b ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, new_AGEMA_signal_3595, Midori_rounds_SR_Result[30]}), .c ({DataOut_s3[26], DataOut_s2[26], DataOut_s1[26], DataOut_s0[26]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U81 ( .a ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, new_AGEMA_signal_1885, wk[24]}), .b ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, new_AGEMA_signal_3601, Midori_rounds_SR_Result[28]}), .c ({DataOut_s3[24], DataOut_s2[24], DataOut_s1[24], DataOut_s0[24]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U79 ( .a ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, new_AGEMA_signal_1903, wk[22]}), .b ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, new_AGEMA_signal_3583, Midori_rounds_SR_Result[58]}), .c ({DataOut_s3[22], DataOut_s2[22], DataOut_s1[22], DataOut_s0[22]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U77 ( .a ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, new_AGEMA_signal_1921, wk[20]}), .b ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, new_AGEMA_signal_3589, Midori_rounds_SR_Result[56]}), .c ({DataOut_s3[20], DataOut_s2[20], DataOut_s1[20], DataOut_s0[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U74 ( .a ({new_AGEMA_signal_1950, new_AGEMA_signal_1949, new_AGEMA_signal_1948, wk[18]}), .b ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, new_AGEMA_signal_3571, Midori_rounds_SR_Result[38]}), .c ({DataOut_s3[18], DataOut_s2[18], DataOut_s1[18], DataOut_s0[18]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U72 ( .a ({new_AGEMA_signal_1968, new_AGEMA_signal_1967, new_AGEMA_signal_1966, wk[16]}), .b ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, new_AGEMA_signal_3577, Midori_rounds_SR_Result[36]}), .c ({DataOut_s3[16], DataOut_s2[16], DataOut_s1[16], DataOut_s0[16]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U70 ( .a ({new_AGEMA_signal_1986, new_AGEMA_signal_1985, new_AGEMA_signal_1984, wk[14]}), .b ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, new_AGEMA_signal_3559, Midori_rounds_SR_Result[22]}), .c ({DataOut_s3[14], DataOut_s2[14], DataOut_s1[14], DataOut_s0[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U68 ( .a ({new_AGEMA_signal_2004, new_AGEMA_signal_2003, new_AGEMA_signal_2002, wk[12]}), .b ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, new_AGEMA_signal_3565, Midori_rounds_SR_Result[20]}), .c ({DataOut_s3[12], DataOut_s2[12], DataOut_s1[12], DataOut_s0[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U66 ( .a ({new_AGEMA_signal_2022, new_AGEMA_signal_2021, new_AGEMA_signal_2020, wk[10]}), .b ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, new_AGEMA_signal_3547, Midori_rounds_SR_Result[10]}), .c ({DataOut_s3[10], DataOut_s2[10], DataOut_s1[10], DataOut_s0[10]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_U65 ( .a ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, new_AGEMA_signal_2029, wk[0]}), .b ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, new_AGEMA_signal_3529, Midori_rounds_SR_Result[48]}), .c ({DataOut_s3[0], DataOut_s2[0], DataOut_s1[0], DataOut_s0[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U143 ( .a ({new_AGEMA_signal_3555, new_AGEMA_signal_3554, new_AGEMA_signal_3553, Midori_rounds_SR_Result[8]}), .b ({new_AGEMA_signal_4413, new_AGEMA_signal_4412, new_AGEMA_signal_4411, Midori_rounds_n16}), .c ({new_AGEMA_signal_4566, new_AGEMA_signal_4565, new_AGEMA_signal_4564, Midori_rounds_sub_ResultXORkey[8]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U141 ( .a ({new_AGEMA_signal_3132, new_AGEMA_signal_3131, new_AGEMA_signal_3130, Midori_rounds_SelectedKey_6_}), .b ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, new_AGEMA_signal_3535, Midori_rounds_SR_Result[46]}), .c ({new_AGEMA_signal_3912, new_AGEMA_signal_3911, new_AGEMA_signal_3910, Midori_rounds_sub_ResultXORkey[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U139 ( .a ({new_AGEMA_signal_3276, new_AGEMA_signal_3275, new_AGEMA_signal_3274, Midori_rounds_SelectedKey_62_}), .b ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, new_AGEMA_signal_3703, Midori_rounds_SR_Result[62]}), .c ({new_AGEMA_signal_3918, new_AGEMA_signal_3917, new_AGEMA_signal_3916, Midori_rounds_sub_ResultXORkey[62]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U137 ( .a ({new_AGEMA_signal_3711, new_AGEMA_signal_3710, new_AGEMA_signal_3709, Midori_rounds_SR_Result[60]}), .b ({new_AGEMA_signal_4578, new_AGEMA_signal_4577, new_AGEMA_signal_4576, Midori_rounds_n15}), .c ({new_AGEMA_signal_4752, new_AGEMA_signal_4751, new_AGEMA_signal_4750, Midori_rounds_sub_ResultXORkey[60]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U134 ( .a ({new_AGEMA_signal_3264, new_AGEMA_signal_3263, new_AGEMA_signal_3262, Midori_rounds_SelectedKey_58_}), .b ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, new_AGEMA_signal_3691, Midori_rounds_SR_Result[34]}), .c ({new_AGEMA_signal_3930, new_AGEMA_signal_3929, new_AGEMA_signal_3928, Midori_rounds_sub_ResultXORkey[58]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U132 ( .a ({new_AGEMA_signal_3699, new_AGEMA_signal_3698, new_AGEMA_signal_3697, Midori_rounds_SR_Result[32]}), .b ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, new_AGEMA_signal_4579, Midori_rounds_n14}), .c ({new_AGEMA_signal_4755, new_AGEMA_signal_4754, new_AGEMA_signal_4753, Midori_rounds_sub_ResultXORkey[56]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U130 ( .a ({new_AGEMA_signal_3252, new_AGEMA_signal_3251, new_AGEMA_signal_3250, Midori_rounds_SelectedKey_54_}), .b ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, new_AGEMA_signal_3679, Midori_rounds_SR_Result[6]}), .c ({new_AGEMA_signal_3939, new_AGEMA_signal_3938, new_AGEMA_signal_3937, Midori_rounds_sub_ResultXORkey[54]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U128 ( .a ({new_AGEMA_signal_3687, new_AGEMA_signal_3686, new_AGEMA_signal_3685, Midori_rounds_SR_Result[4]}), .b ({new_AGEMA_signal_4584, new_AGEMA_signal_4583, new_AGEMA_signal_4582, Midori_rounds_n13}), .c ({new_AGEMA_signal_4758, new_AGEMA_signal_4757, new_AGEMA_signal_4756, Midori_rounds_sub_ResultXORkey[52]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U126 ( .a ({new_AGEMA_signal_3240, new_AGEMA_signal_3239, new_AGEMA_signal_3238, Midori_rounds_SelectedKey_50_}), .b ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, new_AGEMA_signal_3667, Midori_rounds_SR_Result[26]}), .c ({new_AGEMA_signal_3948, new_AGEMA_signal_3947, new_AGEMA_signal_3946, Midori_rounds_sub_ResultXORkey[50]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U125 ( .a ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, new_AGEMA_signal_3541, Midori_rounds_SR_Result[44]}), .b ({new_AGEMA_signal_4587, new_AGEMA_signal_4586, new_AGEMA_signal_4585, Midori_rounds_n12}), .c ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, new_AGEMA_signal_4759, Midori_rounds_sub_ResultXORkey[4]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U123 ( .a ({new_AGEMA_signal_3675, new_AGEMA_signal_3674, new_AGEMA_signal_3673, Midori_rounds_SR_Result[24]}), .b ({new_AGEMA_signal_4944, new_AGEMA_signal_4943, new_AGEMA_signal_4942, Midori_rounds_n11}), .c ({new_AGEMA_signal_4977, new_AGEMA_signal_4976, new_AGEMA_signal_4975, Midori_rounds_sub_ResultXORkey[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U121 ( .a ({new_AGEMA_signal_3228, new_AGEMA_signal_3227, new_AGEMA_signal_3226, Midori_rounds_SelectedKey_46_}), .b ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, new_AGEMA_signal_3655, Midori_rounds_SR_Result[42]}), .c ({new_AGEMA_signal_3957, new_AGEMA_signal_3956, new_AGEMA_signal_3955, Midori_rounds_sub_ResultXORkey[46]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U119 ( .a ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, new_AGEMA_signal_3661, Midori_rounds_SR_Result[40]}), .b ({new_AGEMA_signal_4470, new_AGEMA_signal_4469, new_AGEMA_signal_4468, Midori_rounds_n10}), .c ({new_AGEMA_signal_4569, new_AGEMA_signal_4568, new_AGEMA_signal_4567, Midori_rounds_sub_ResultXORkey[44]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U117 ( .a ({new_AGEMA_signal_3216, new_AGEMA_signal_3215, new_AGEMA_signal_3214, Midori_rounds_SelectedKey_42_}), .b ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, new_AGEMA_signal_3643, Midori_rounds_SR_Result[54]}), .c ({new_AGEMA_signal_3966, new_AGEMA_signal_3965, new_AGEMA_signal_3964, Midori_rounds_sub_ResultXORkey[42]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U115 ( .a ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, new_AGEMA_signal_3649, Midori_rounds_SR_Result[52]}), .b ({new_AGEMA_signal_4590, new_AGEMA_signal_4589, new_AGEMA_signal_4588, Midori_rounds_n9}), .c ({new_AGEMA_signal_4764, new_AGEMA_signal_4763, new_AGEMA_signal_4762, Midori_rounds_sub_ResultXORkey[40]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U112 ( .a ({new_AGEMA_signal_3204, new_AGEMA_signal_3203, new_AGEMA_signal_3202, Midori_rounds_SelectedKey_38_}), .b ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, new_AGEMA_signal_3631, Midori_rounds_SR_Result[18]}), .c ({new_AGEMA_signal_3978, new_AGEMA_signal_3977, new_AGEMA_signal_3976, Midori_rounds_sub_ResultXORkey[38]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U110 ( .a ({new_AGEMA_signal_3639, new_AGEMA_signal_3638, new_AGEMA_signal_3637, Midori_rounds_SR_Result[16]}), .b ({new_AGEMA_signal_4494, new_AGEMA_signal_4493, new_AGEMA_signal_4492, Midori_rounds_n8}), .c ({new_AGEMA_signal_4572, new_AGEMA_signal_4571, new_AGEMA_signal_4570, Midori_rounds_sub_ResultXORkey[36]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U108 ( .a ({new_AGEMA_signal_3192, new_AGEMA_signal_3191, new_AGEMA_signal_3190, Midori_rounds_SelectedKey_34_}), .b ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, new_AGEMA_signal_3619, Midori_rounds_SR_Result[14]}), .c ({new_AGEMA_signal_3987, new_AGEMA_signal_3986, new_AGEMA_signal_3985, Midori_rounds_sub_ResultXORkey[34]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U106 ( .a ({new_AGEMA_signal_3627, new_AGEMA_signal_3626, new_AGEMA_signal_3625, Midori_rounds_SR_Result[12]}), .b ({new_AGEMA_signal_4593, new_AGEMA_signal_4592, new_AGEMA_signal_4591, Midori_rounds_n7}), .c ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, new_AGEMA_signal_4765, Midori_rounds_sub_ResultXORkey[32]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U104 ( .a ({new_AGEMA_signal_3180, new_AGEMA_signal_3179, new_AGEMA_signal_3178, Midori_rounds_SelectedKey_30_}), .b ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, new_AGEMA_signal_3607, Midori_rounds_SR_Result[2]}), .c ({new_AGEMA_signal_3996, new_AGEMA_signal_3995, new_AGEMA_signal_3994, Midori_rounds_sub_ResultXORkey[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U103 ( .a ({new_AGEMA_signal_2040, new_AGEMA_signal_2039, new_AGEMA_signal_2038, Midori_rounds_SelectedKey_2_}), .b ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, new_AGEMA_signal_3523, Midori_rounds_SR_Result[50]}), .c ({new_AGEMA_signal_3999, new_AGEMA_signal_3998, new_AGEMA_signal_3997, Midori_rounds_sub_ResultXORkey[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U101 ( .a ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, new_AGEMA_signal_3613, Midori_rounds_SR_Result[0]}), .b ({new_AGEMA_signal_4782, new_AGEMA_signal_4781, new_AGEMA_signal_4780, Midori_rounds_n6}), .c ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, new_AGEMA_signal_4939, Midori_rounds_sub_ResultXORkey[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U99 ( .a ({new_AGEMA_signal_2070, new_AGEMA_signal_2069, new_AGEMA_signal_2068, Midori_rounds_SelectedKey_26_}), .b ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, new_AGEMA_signal_3595, Midori_rounds_SR_Result[30]}), .c ({new_AGEMA_signal_4008, new_AGEMA_signal_4007, new_AGEMA_signal_4006, Midori_rounds_sub_ResultXORkey[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U97 ( .a ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, new_AGEMA_signal_3601, Midori_rounds_SR_Result[28]}), .b ({new_AGEMA_signal_4596, new_AGEMA_signal_4595, new_AGEMA_signal_4594, Midori_rounds_n5}), .c ({new_AGEMA_signal_4770, new_AGEMA_signal_4769, new_AGEMA_signal_4768, Midori_rounds_sub_ResultXORkey[24]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U95 ( .a ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, new_AGEMA_signal_3157, Midori_rounds_SelectedKey_22_}), .b ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, new_AGEMA_signal_3583, Midori_rounds_SR_Result[58]}), .c ({new_AGEMA_signal_4017, new_AGEMA_signal_4016, new_AGEMA_signal_4015, Midori_rounds_sub_ResultXORkey[22]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U93 ( .a ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, new_AGEMA_signal_3589, Midori_rounds_SR_Result[56]}), .b ({new_AGEMA_signal_4536, new_AGEMA_signal_4535, new_AGEMA_signal_4534, Midori_rounds_n4}), .c ({new_AGEMA_signal_4575, new_AGEMA_signal_4574, new_AGEMA_signal_4573, Midori_rounds_sub_ResultXORkey[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U90 ( .a ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, new_AGEMA_signal_3145, Midori_rounds_SelectedKey_18_}), .b ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, new_AGEMA_signal_3571, Midori_rounds_SR_Result[38]}), .c ({new_AGEMA_signal_4029, new_AGEMA_signal_4028, new_AGEMA_signal_4027, Midori_rounds_sub_ResultXORkey[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U88 ( .a ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, new_AGEMA_signal_3577, Midori_rounds_SR_Result[36]}), .b ({new_AGEMA_signal_4599, new_AGEMA_signal_4598, new_AGEMA_signal_4597, Midori_rounds_n3}), .c ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, new_AGEMA_signal_4771, Midori_rounds_sub_ResultXORkey[16]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U86 ( .a ({new_AGEMA_signal_2064, new_AGEMA_signal_2063, new_AGEMA_signal_2062, Midori_rounds_SelectedKey_14_}), .b ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, new_AGEMA_signal_3559, Midori_rounds_SR_Result[22]}), .c ({new_AGEMA_signal_4038, new_AGEMA_signal_4037, new_AGEMA_signal_4036, Midori_rounds_sub_ResultXORkey[14]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U84 ( .a ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, new_AGEMA_signal_3565, Midori_rounds_SR_Result[20]}), .b ({new_AGEMA_signal_4602, new_AGEMA_signal_4601, new_AGEMA_signal_4600, Midori_rounds_n2}), .c ({new_AGEMA_signal_4776, new_AGEMA_signal_4775, new_AGEMA_signal_4774, Midori_rounds_sub_ResultXORkey[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U82 ( .a ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, new_AGEMA_signal_2053, Midori_rounds_SelectedKey_10_}), .b ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, new_AGEMA_signal_3547, Midori_rounds_SR_Result[10]}), .c ({new_AGEMA_signal_4047, new_AGEMA_signal_4046, new_AGEMA_signal_4045, Midori_rounds_sub_ResultXORkey[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U81 ( .a ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, new_AGEMA_signal_3529, Midori_rounds_SR_Result[48]}), .b ({new_AGEMA_signal_4605, new_AGEMA_signal_4604, new_AGEMA_signal_4603, Midori_rounds_n1}), .c ({new_AGEMA_signal_4779, new_AGEMA_signal_4778, new_AGEMA_signal_4777, Midori_rounds_sub_ResultXORkey[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U79 ( .a ({new_AGEMA_signal_5028, new_AGEMA_signal_5027, new_AGEMA_signal_5026, Midori_rounds_SR_Inv_Result[8]}), .b ({new_AGEMA_signal_4413, new_AGEMA_signal_4412, new_AGEMA_signal_4411, Midori_rounds_n16}), .c ({new_AGEMA_signal_5040, new_AGEMA_signal_5039, new_AGEMA_signal_5038, Midori_rounds_mul_ResultXORkey[8]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U76 ( .a ({new_AGEMA_signal_3132, new_AGEMA_signal_3131, new_AGEMA_signal_3130, Midori_rounds_SelectedKey_6_}), .b ({new_AGEMA_signal_4380, new_AGEMA_signal_4379, new_AGEMA_signal_4378, Midori_rounds_SR_Inv_Result[54]}), .c ({new_AGEMA_signal_4419, new_AGEMA_signal_4418, new_AGEMA_signal_4417, Midori_rounds_mul_ResultXORkey[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U74 ( .a ({new_AGEMA_signal_3276, new_AGEMA_signal_3275, new_AGEMA_signal_3274, Midori_rounds_SelectedKey_62_}), .b ({new_AGEMA_signal_4290, new_AGEMA_signal_4289, new_AGEMA_signal_4288, Midori_rounds_SR_Inv_Result[62]}), .c ({new_AGEMA_signal_4425, new_AGEMA_signal_4424, new_AGEMA_signal_4423, Midori_rounds_mul_ResultXORkey[62]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U72 ( .a ({new_AGEMA_signal_5097, new_AGEMA_signal_5096, new_AGEMA_signal_5095, Midori_rounds_SR_Inv_Result[60]}), .b ({new_AGEMA_signal_4578, new_AGEMA_signal_4577, new_AGEMA_signal_4576, Midori_rounds_n15}), .c ({new_AGEMA_signal_5133, new_AGEMA_signal_5132, new_AGEMA_signal_5131, Midori_rounds_mul_ResultXORkey[60]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U68 ( .a ({new_AGEMA_signal_3264, new_AGEMA_signal_3263, new_AGEMA_signal_3262, Midori_rounds_SelectedKey_58_}), .b ({new_AGEMA_signal_4299, new_AGEMA_signal_4298, new_AGEMA_signal_4297, Midori_rounds_SR_Inv_Result[22]}), .c ({new_AGEMA_signal_4437, new_AGEMA_signal_4436, new_AGEMA_signal_4435, Midori_rounds_mul_ResultXORkey[58]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U66 ( .a ({new_AGEMA_signal_5094, new_AGEMA_signal_5093, new_AGEMA_signal_5092, Midori_rounds_SR_Inv_Result[20]}), .b ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, new_AGEMA_signal_4579, Midori_rounds_n14}), .c ({new_AGEMA_signal_5136, new_AGEMA_signal_5135, new_AGEMA_signal_5134, Midori_rounds_mul_ResultXORkey[56]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U63 ( .a ({new_AGEMA_signal_3252, new_AGEMA_signal_3251, new_AGEMA_signal_3250, Midori_rounds_SelectedKey_54_}), .b ({new_AGEMA_signal_4272, new_AGEMA_signal_4271, new_AGEMA_signal_4270, Midori_rounds_SR_Inv_Result[42]}), .c ({new_AGEMA_signal_4446, new_AGEMA_signal_4445, new_AGEMA_signal_4444, Midori_rounds_mul_ResultXORkey[54]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U61 ( .a ({new_AGEMA_signal_5073, new_AGEMA_signal_5072, new_AGEMA_signal_5071, Midori_rounds_SR_Inv_Result[40]}), .b ({new_AGEMA_signal_4584, new_AGEMA_signal_4583, new_AGEMA_signal_4582, Midori_rounds_n13}), .c ({new_AGEMA_signal_5085, new_AGEMA_signal_5084, new_AGEMA_signal_5083, Midori_rounds_mul_ResultXORkey[52]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U58 ( .a ({new_AGEMA_signal_3240, new_AGEMA_signal_3239, new_AGEMA_signal_3238, Midori_rounds_SelectedKey_50_}), .b ({new_AGEMA_signal_4281, new_AGEMA_signal_4280, new_AGEMA_signal_4279, Midori_rounds_SR_Inv_Result[2]}), .c ({new_AGEMA_signal_4455, new_AGEMA_signal_4454, new_AGEMA_signal_4453, Midori_rounds_mul_ResultXORkey[50]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U57 ( .a ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, new_AGEMA_signal_5029, Midori_rounds_SR_Inv_Result[52]}), .b ({new_AGEMA_signal_4587, new_AGEMA_signal_4586, new_AGEMA_signal_4585, Midori_rounds_n12}), .c ({new_AGEMA_signal_5043, new_AGEMA_signal_5042, new_AGEMA_signal_5041, Midori_rounds_mul_ResultXORkey[4]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U54 ( .a ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, new_AGEMA_signal_5002, Midori_rounds_SR_Inv_Result[0]}), .b ({new_AGEMA_signal_4944, new_AGEMA_signal_4943, new_AGEMA_signal_4942, Midori_rounds_n11}), .c ({new_AGEMA_signal_5046, new_AGEMA_signal_5045, new_AGEMA_signal_5044, Midori_rounds_mul_ResultXORkey[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U51 ( .a ({new_AGEMA_signal_3228, new_AGEMA_signal_3227, new_AGEMA_signal_3226, Midori_rounds_SelectedKey_46_}), .b ({new_AGEMA_signal_4326, new_AGEMA_signal_4325, new_AGEMA_signal_4324, Midori_rounds_SR_Inv_Result[6]}), .c ({new_AGEMA_signal_4464, new_AGEMA_signal_4463, new_AGEMA_signal_4462, Midori_rounds_mul_ResultXORkey[46]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U49 ( .a ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, new_AGEMA_signal_5011, Midori_rounds_SR_Inv_Result[4]}), .b ({new_AGEMA_signal_4470, new_AGEMA_signal_4469, new_AGEMA_signal_4468, Midori_rounds_n10}), .c ({new_AGEMA_signal_5049, new_AGEMA_signal_5048, new_AGEMA_signal_5047, Midori_rounds_mul_ResultXORkey[44]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U46 ( .a ({new_AGEMA_signal_3216, new_AGEMA_signal_3215, new_AGEMA_signal_3214, Midori_rounds_SelectedKey_42_}), .b ({new_AGEMA_signal_4335, new_AGEMA_signal_4334, new_AGEMA_signal_4333, Midori_rounds_SR_Inv_Result[46]}), .c ({new_AGEMA_signal_4476, new_AGEMA_signal_4475, new_AGEMA_signal_4474, Midori_rounds_mul_ResultXORkey[42]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U44 ( .a ({new_AGEMA_signal_5007, new_AGEMA_signal_5006, new_AGEMA_signal_5005, Midori_rounds_SR_Inv_Result[44]}), .b ({new_AGEMA_signal_4590, new_AGEMA_signal_4589, new_AGEMA_signal_4588, Midori_rounds_n9}), .c ({new_AGEMA_signal_5052, new_AGEMA_signal_5051, new_AGEMA_signal_5050, Midori_rounds_mul_ResultXORkey[40]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U40 ( .a ({new_AGEMA_signal_3204, new_AGEMA_signal_3203, new_AGEMA_signal_3202, Midori_rounds_SelectedKey_38_}), .b ({new_AGEMA_signal_4308, new_AGEMA_signal_4307, new_AGEMA_signal_4306, Midori_rounds_SR_Inv_Result[18]}), .c ({new_AGEMA_signal_4488, new_AGEMA_signal_4487, new_AGEMA_signal_4486, Midori_rounds_mul_ResultXORkey[38]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U38 ( .a ({new_AGEMA_signal_5010, new_AGEMA_signal_5009, new_AGEMA_signal_5008, Midori_rounds_SR_Inv_Result[16]}), .b ({new_AGEMA_signal_4494, new_AGEMA_signal_4493, new_AGEMA_signal_4492, Midori_rounds_n8}), .c ({new_AGEMA_signal_5055, new_AGEMA_signal_5054, new_AGEMA_signal_5053, Midori_rounds_mul_ResultXORkey[36]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U35 ( .a ({new_AGEMA_signal_3192, new_AGEMA_signal_3191, new_AGEMA_signal_3190, Midori_rounds_SelectedKey_34_}), .b ({new_AGEMA_signal_4317, new_AGEMA_signal_4316, new_AGEMA_signal_4315, Midori_rounds_SR_Inv_Result[58]}), .c ({new_AGEMA_signal_4500, new_AGEMA_signal_4499, new_AGEMA_signal_4498, Midori_rounds_mul_ResultXORkey[34]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U33 ( .a ({new_AGEMA_signal_5016, new_AGEMA_signal_5015, new_AGEMA_signal_5014, Midori_rounds_SR_Inv_Result[56]}), .b ({new_AGEMA_signal_4593, new_AGEMA_signal_4592, new_AGEMA_signal_4591, Midori_rounds_n7}), .c ({new_AGEMA_signal_5058, new_AGEMA_signal_5057, new_AGEMA_signal_5056, Midori_rounds_mul_ResultXORkey[32]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U30 ( .a ({new_AGEMA_signal_3180, new_AGEMA_signal_3179, new_AGEMA_signal_3178, Midori_rounds_SelectedKey_30_}), .b ({new_AGEMA_signal_4362, new_AGEMA_signal_4361, new_AGEMA_signal_4360, Midori_rounds_SR_Inv_Result[26]}), .c ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, new_AGEMA_signal_4507, Midori_rounds_mul_ResultXORkey[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U29 ( .a ({new_AGEMA_signal_2040, new_AGEMA_signal_2039, new_AGEMA_signal_2038, Midori_rounds_SelectedKey_2_}), .b ({new_AGEMA_signal_4389, new_AGEMA_signal_4388, new_AGEMA_signal_4387, Midori_rounds_SR_Inv_Result[30]}), .c ({new_AGEMA_signal_4512, new_AGEMA_signal_4511, new_AGEMA_signal_4510, Midori_rounds_mul_ResultXORkey[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U27 ( .a ({new_AGEMA_signal_5022, new_AGEMA_signal_5021, new_AGEMA_signal_5020, Midori_rounds_SR_Inv_Result[24]}), .b ({new_AGEMA_signal_4782, new_AGEMA_signal_4781, new_AGEMA_signal_4780, Midori_rounds_n6}), .c ({new_AGEMA_signal_5061, new_AGEMA_signal_5060, new_AGEMA_signal_5059, Midori_rounds_mul_ResultXORkey[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U24 ( .a ({new_AGEMA_signal_2070, new_AGEMA_signal_2069, new_AGEMA_signal_2068, Midori_rounds_SelectedKey_26_}), .b ({new_AGEMA_signal_4371, new_AGEMA_signal_4370, new_AGEMA_signal_4369, Midori_rounds_SR_Inv_Result[50]}), .c ({new_AGEMA_signal_4521, new_AGEMA_signal_4520, new_AGEMA_signal_4519, Midori_rounds_mul_ResultXORkey[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U22 ( .a ({new_AGEMA_signal_5019, new_AGEMA_signal_5018, new_AGEMA_signal_5017, Midori_rounds_SR_Inv_Result[48]}), .b ({new_AGEMA_signal_4596, new_AGEMA_signal_4595, new_AGEMA_signal_4594, Midori_rounds_n5}), .c ({new_AGEMA_signal_5064, new_AGEMA_signal_5063, new_AGEMA_signal_5062, Midori_rounds_mul_ResultXORkey[24]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U19 ( .a ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, new_AGEMA_signal_3157, Midori_rounds_SelectedKey_22_}), .b ({new_AGEMA_signal_4344, new_AGEMA_signal_4343, new_AGEMA_signal_4342, Midori_rounds_SR_Inv_Result[14]}), .c ({new_AGEMA_signal_4530, new_AGEMA_signal_4529, new_AGEMA_signal_4528, Midori_rounds_mul_ResultXORkey[22]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U17 ( .a ({new_AGEMA_signal_5079, new_AGEMA_signal_5078, new_AGEMA_signal_5077, Midori_rounds_SR_Inv_Result[12]}), .b ({new_AGEMA_signal_4536, new_AGEMA_signal_4535, new_AGEMA_signal_4534, Midori_rounds_n4}), .c ({new_AGEMA_signal_5088, new_AGEMA_signal_5087, new_AGEMA_signal_5086, Midori_rounds_mul_ResultXORkey[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U13 ( .a ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, new_AGEMA_signal_3145, Midori_rounds_SelectedKey_18_}), .b ({new_AGEMA_signal_4353, new_AGEMA_signal_4352, new_AGEMA_signal_4351, Midori_rounds_SR_Inv_Result[38]}), .c ({new_AGEMA_signal_4545, new_AGEMA_signal_4544, new_AGEMA_signal_4543, Midori_rounds_mul_ResultXORkey[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U11 ( .a ({new_AGEMA_signal_5082, new_AGEMA_signal_5081, new_AGEMA_signal_5080, Midori_rounds_SR_Inv_Result[36]}), .b ({new_AGEMA_signal_4599, new_AGEMA_signal_4598, new_AGEMA_signal_4597, Midori_rounds_n3}), .c ({new_AGEMA_signal_5091, new_AGEMA_signal_5090, new_AGEMA_signal_5089, Midori_rounds_mul_ResultXORkey[16]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U8 ( .a ({new_AGEMA_signal_2064, new_AGEMA_signal_2063, new_AGEMA_signal_2062, Midori_rounds_SelectedKey_14_}), .b ({new_AGEMA_signal_4398, new_AGEMA_signal_4397, new_AGEMA_signal_4396, Midori_rounds_SR_Inv_Result[34]}), .c ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, Midori_rounds_mul_ResultXORkey[14]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U6 ( .a ({new_AGEMA_signal_5034, new_AGEMA_signal_5033, new_AGEMA_signal_5032, Midori_rounds_SR_Inv_Result[32]}), .b ({new_AGEMA_signal_4602, new_AGEMA_signal_4601, new_AGEMA_signal_4600, Midori_rounds_n2}), .c ({new_AGEMA_signal_5067, new_AGEMA_signal_5066, new_AGEMA_signal_5065, Midori_rounds_mul_ResultXORkey[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U3 ( .a ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, new_AGEMA_signal_2053, Midori_rounds_SelectedKey_10_}), .b ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, new_AGEMA_signal_4405, Midori_rounds_SR_Inv_Result[10]}), .c ({new_AGEMA_signal_4563, new_AGEMA_signal_4562, new_AGEMA_signal_4561, Midori_rounds_mul_ResultXORkey[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_U2 ( .a ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, new_AGEMA_signal_5035, Midori_rounds_SR_Inv_Result[28]}), .b ({new_AGEMA_signal_4605, new_AGEMA_signal_4604, new_AGEMA_signal_4603, Midori_rounds_n1}), .c ({new_AGEMA_signal_5070, new_AGEMA_signal_5069, new_AGEMA_signal_5068, Midori_rounds_mul_ResultXORkey[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_5100, new_AGEMA_signal_5099, new_AGEMA_signal_5098, Midori_rounds_round_Result[0]}), .a ({new_AGEMA_signal_2838, new_AGEMA_signal_2837, new_AGEMA_signal_2836, Midori_add_Result_Start[0]}), .c ({new_AGEMA_signal_5139, new_AGEMA_signal_5138, new_AGEMA_signal_5137, Midori_rounds_roundResult_Reg_SFF_0_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4611, new_AGEMA_signal_4610, new_AGEMA_signal_4609, Midori_rounds_round_Result[2]}), .a ({new_AGEMA_signal_2706, new_AGEMA_signal_2705, new_AGEMA_signal_2704, Midori_add_Result_Start[2]}), .c ({new_AGEMA_signal_4788, new_AGEMA_signal_4787, new_AGEMA_signal_4786, Midori_rounds_roundResult_Reg_SFF_2_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_5103, new_AGEMA_signal_5102, new_AGEMA_signal_5101, Midori_rounds_round_Result[4]}), .a ({new_AGEMA_signal_2574, new_AGEMA_signal_2573, new_AGEMA_signal_2572, Midori_add_Result_Start[4]}), .c ({new_AGEMA_signal_5142, new_AGEMA_signal_5141, new_AGEMA_signal_5140, Midori_rounds_roundResult_Reg_SFF_4_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4620, new_AGEMA_signal_4619, new_AGEMA_signal_4618, Midori_rounds_round_Result[6]}), .a ({new_AGEMA_signal_2478, new_AGEMA_signal_2477, new_AGEMA_signal_2476, Midori_add_Result_Start[6]}), .c ({new_AGEMA_signal_4797, new_AGEMA_signal_4796, new_AGEMA_signal_4795, Midori_rounds_roundResult_Reg_SFF_6_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_5106, new_AGEMA_signal_5105, new_AGEMA_signal_5104, Midori_rounds_round_Result[8]}), .a ({new_AGEMA_signal_2466, new_AGEMA_signal_2465, new_AGEMA_signal_2464, Midori_add_Result_Start[8]}), .c ({new_AGEMA_signal_5145, new_AGEMA_signal_5144, new_AGEMA_signal_5143, Midori_rounds_roundResult_Reg_SFF_8_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4629, new_AGEMA_signal_4628, new_AGEMA_signal_4627, Midori_rounds_round_Result[10]}), .a ({new_AGEMA_signal_2832, new_AGEMA_signal_2831, new_AGEMA_signal_2830, Midori_add_Result_Start[10]}), .c ({new_AGEMA_signal_4806, new_AGEMA_signal_4805, new_AGEMA_signal_4804, Midori_rounds_roundResult_Reg_SFF_10_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_5109, new_AGEMA_signal_5108, new_AGEMA_signal_5107, Midori_rounds_round_Result[12]}), .a ({new_AGEMA_signal_2820, new_AGEMA_signal_2819, new_AGEMA_signal_2818, Midori_add_Result_Start[12]}), .c ({new_AGEMA_signal_5148, new_AGEMA_signal_5147, new_AGEMA_signal_5146, Midori_rounds_roundResult_Reg_SFF_12_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4638, new_AGEMA_signal_4637, new_AGEMA_signal_4636, Midori_rounds_round_Result[14]}), .a ({new_AGEMA_signal_2808, new_AGEMA_signal_2807, new_AGEMA_signal_2806, Midori_add_Result_Start[14]}), .c ({new_AGEMA_signal_4815, new_AGEMA_signal_4814, new_AGEMA_signal_4813, Midori_rounds_roundResult_Reg_SFF_14_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_5172, new_AGEMA_signal_5171, new_AGEMA_signal_5170, Midori_rounds_round_Result[16]}), .a ({new_AGEMA_signal_2796, new_AGEMA_signal_2795, new_AGEMA_signal_2794, Midori_add_Result_Start[16]}), .c ({new_AGEMA_signal_5181, new_AGEMA_signal_5180, new_AGEMA_signal_5179, Midori_rounds_roundResult_Reg_SFF_16_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4647, new_AGEMA_signal_4646, new_AGEMA_signal_4645, Midori_rounds_round_Result[18]}), .a ({new_AGEMA_signal_2784, new_AGEMA_signal_2783, new_AGEMA_signal_2782, Midori_add_Result_Start[18]}), .c ({new_AGEMA_signal_4824, new_AGEMA_signal_4823, new_AGEMA_signal_4822, Midori_rounds_roundResult_Reg_SFF_18_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_5175, new_AGEMA_signal_5174, new_AGEMA_signal_5173, Midori_rounds_round_Result[20]}), .a ({new_AGEMA_signal_2766, new_AGEMA_signal_2765, new_AGEMA_signal_2764, Midori_add_Result_Start[20]}), .c ({new_AGEMA_signal_5184, new_AGEMA_signal_5183, new_AGEMA_signal_5182, Midori_rounds_roundResult_Reg_SFF_20_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4656, new_AGEMA_signal_4655, new_AGEMA_signal_4654, Midori_rounds_round_Result[22]}), .a ({new_AGEMA_signal_2754, new_AGEMA_signal_2753, new_AGEMA_signal_2752, Midori_add_Result_Start[22]}), .c ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, new_AGEMA_signal_4831, Midori_rounds_roundResult_Reg_SFF_22_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_5112, new_AGEMA_signal_5111, new_AGEMA_signal_5110, Midori_rounds_round_Result[24]}), .a ({new_AGEMA_signal_2742, new_AGEMA_signal_2741, new_AGEMA_signal_2740, Midori_add_Result_Start[24]}), .c ({new_AGEMA_signal_5151, new_AGEMA_signal_5150, new_AGEMA_signal_5149, Midori_rounds_roundResult_Reg_SFF_24_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4665, new_AGEMA_signal_4664, new_AGEMA_signal_4663, Midori_rounds_round_Result[26]}), .a ({new_AGEMA_signal_2730, new_AGEMA_signal_2729, new_AGEMA_signal_2728, Midori_add_Result_Start[26]}), .c ({new_AGEMA_signal_4842, new_AGEMA_signal_4841, new_AGEMA_signal_4840, Midori_rounds_roundResult_Reg_SFF_26_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_5115, new_AGEMA_signal_5114, new_AGEMA_signal_5113, Midori_rounds_round_Result[28]}), .a ({new_AGEMA_signal_2718, new_AGEMA_signal_2717, new_AGEMA_signal_2716, Midori_add_Result_Start[28]}), .c ({new_AGEMA_signal_5154, new_AGEMA_signal_5153, new_AGEMA_signal_5152, Midori_rounds_roundResult_Reg_SFF_28_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4674, new_AGEMA_signal_4673, new_AGEMA_signal_4672, Midori_rounds_round_Result[30]}), .a ({new_AGEMA_signal_2700, new_AGEMA_signal_2699, new_AGEMA_signal_2698, Midori_add_Result_Start[30]}), .c ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, new_AGEMA_signal_4849, Midori_rounds_roundResult_Reg_SFF_30_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_5118, new_AGEMA_signal_5117, new_AGEMA_signal_5116, Midori_rounds_round_Result[32]}), .a ({new_AGEMA_signal_2688, new_AGEMA_signal_2687, new_AGEMA_signal_2686, Midori_add_Result_Start[32]}), .c ({new_AGEMA_signal_5157, new_AGEMA_signal_5156, new_AGEMA_signal_5155, Midori_rounds_roundResult_Reg_SFF_32_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4683, new_AGEMA_signal_4682, new_AGEMA_signal_4681, Midori_rounds_round_Result[34]}), .a ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, new_AGEMA_signal_2674, Midori_add_Result_Start[34]}), .c ({new_AGEMA_signal_4860, new_AGEMA_signal_4859, new_AGEMA_signal_4858, Midori_rounds_roundResult_Reg_SFF_34_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_5121, new_AGEMA_signal_5120, new_AGEMA_signal_5119, Midori_rounds_round_Result[36]}), .a ({new_AGEMA_signal_2664, new_AGEMA_signal_2663, new_AGEMA_signal_2662, Midori_add_Result_Start[36]}), .c ({new_AGEMA_signal_5160, new_AGEMA_signal_5159, new_AGEMA_signal_5158, Midori_rounds_roundResult_Reg_SFF_36_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4692, new_AGEMA_signal_4691, new_AGEMA_signal_4690, Midori_rounds_round_Result[38]}), .a ({new_AGEMA_signal_2652, new_AGEMA_signal_2651, new_AGEMA_signal_2650, Midori_add_Result_Start[38]}), .c ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, Midori_rounds_roundResult_Reg_SFF_38_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_5124, new_AGEMA_signal_5123, new_AGEMA_signal_5122, Midori_rounds_round_Result[40]}), .a ({new_AGEMA_signal_2634, new_AGEMA_signal_2633, new_AGEMA_signal_2632, Midori_add_Result_Start[40]}), .c ({new_AGEMA_signal_5163, new_AGEMA_signal_5162, new_AGEMA_signal_5161, Midori_rounds_roundResult_Reg_SFF_40_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4701, new_AGEMA_signal_4700, new_AGEMA_signal_4699, Midori_rounds_round_Result[42]}), .a ({new_AGEMA_signal_2622, new_AGEMA_signal_2621, new_AGEMA_signal_2620, Midori_add_Result_Start[42]}), .c ({new_AGEMA_signal_4878, new_AGEMA_signal_4877, new_AGEMA_signal_4876, Midori_rounds_roundResult_Reg_SFF_42_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_5127, new_AGEMA_signal_5126, new_AGEMA_signal_5125, Midori_rounds_round_Result[44]}), .a ({new_AGEMA_signal_2610, new_AGEMA_signal_2609, new_AGEMA_signal_2608, Midori_add_Result_Start[44]}), .c ({new_AGEMA_signal_5166, new_AGEMA_signal_5165, new_AGEMA_signal_5164, Midori_rounds_roundResult_Reg_SFF_44_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4710, new_AGEMA_signal_4709, new_AGEMA_signal_4708, Midori_rounds_round_Result[46]}), .a ({new_AGEMA_signal_2598, new_AGEMA_signal_2597, new_AGEMA_signal_2596, Midori_add_Result_Start[46]}), .c ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, new_AGEMA_signal_4885, Midori_rounds_roundResult_Reg_SFF_46_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_5130, new_AGEMA_signal_5129, new_AGEMA_signal_5128, Midori_rounds_round_Result[48]}), .a ({new_AGEMA_signal_2586, new_AGEMA_signal_2585, new_AGEMA_signal_2584, Midori_add_Result_Start[48]}), .c ({new_AGEMA_signal_5169, new_AGEMA_signal_5168, new_AGEMA_signal_5167, Midori_rounds_roundResult_Reg_SFF_48_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4719, new_AGEMA_signal_4718, new_AGEMA_signal_4717, Midori_rounds_round_Result[50]}), .a ({new_AGEMA_signal_2568, new_AGEMA_signal_2567, new_AGEMA_signal_2566, Midori_add_Result_Start[50]}), .c ({new_AGEMA_signal_4896, new_AGEMA_signal_4895, new_AGEMA_signal_4894, Midori_rounds_roundResult_Reg_SFF_50_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_5178, new_AGEMA_signal_5177, new_AGEMA_signal_5176, Midori_rounds_round_Result[52]}), .a ({new_AGEMA_signal_2556, new_AGEMA_signal_2555, new_AGEMA_signal_2554, Midori_add_Result_Start[52]}), .c ({new_AGEMA_signal_5187, new_AGEMA_signal_5186, new_AGEMA_signal_5185, Midori_rounds_roundResult_Reg_SFF_52_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4728, new_AGEMA_signal_4727, new_AGEMA_signal_4726, Midori_rounds_round_Result[54]}), .a ({new_AGEMA_signal_2544, new_AGEMA_signal_2543, new_AGEMA_signal_2542, Midori_add_Result_Start[54]}), .c ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, new_AGEMA_signal_4903, Midori_rounds_roundResult_Reg_SFF_54_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_5190, new_AGEMA_signal_5189, new_AGEMA_signal_5188, Midori_rounds_round_Result[56]}), .a ({new_AGEMA_signal_2532, new_AGEMA_signal_2531, new_AGEMA_signal_2530, Midori_add_Result_Start[56]}), .c ({new_AGEMA_signal_5196, new_AGEMA_signal_5195, new_AGEMA_signal_5194, Midori_rounds_roundResult_Reg_SFF_56_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4737, new_AGEMA_signal_4736, new_AGEMA_signal_4735, Midori_rounds_round_Result[58]}), .a ({new_AGEMA_signal_2520, new_AGEMA_signal_2519, new_AGEMA_signal_2518, Midori_add_Result_Start[58]}), .c ({new_AGEMA_signal_4914, new_AGEMA_signal_4913, new_AGEMA_signal_4912, Midori_rounds_roundResult_Reg_SFF_58_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_5193, new_AGEMA_signal_5192, new_AGEMA_signal_5191, Midori_rounds_round_Result[60]}), .a ({new_AGEMA_signal_2502, new_AGEMA_signal_2501, new_AGEMA_signal_2500, Midori_add_Result_Start[60]}), .c ({new_AGEMA_signal_5199, new_AGEMA_signal_5198, new_AGEMA_signal_5197, Midori_rounds_roundResult_Reg_SFF_60_DQ}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_4746, new_AGEMA_signal_4745, new_AGEMA_signal_4744, Midori_rounds_round_Result[62]}), .a ({new_AGEMA_signal_2490, new_AGEMA_signal_2489, new_AGEMA_signal_2488, Midori_add_Result_Start[62]}), .c ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, new_AGEMA_signal_4921, Midori_rounds_roundResult_Reg_SFF_62_DQ}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U17 ( .a ({new_AGEMA_signal_2844, new_AGEMA_signal_2843, new_AGEMA_signal_2842, Midori_rounds_sub_sBox_PRINCE_0_n15}), .b ({new_AGEMA_signal_3288, new_AGEMA_signal_3287, new_AGEMA_signal_3286, Midori_rounds_sub_sBox_PRINCE_0_n12}), .clk (clk), .r ({Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, new_AGEMA_signal_3523, Midori_rounds_SR_Result[50]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U8 ( .a ({new_AGEMA_signal_2856, new_AGEMA_signal_2855, new_AGEMA_signal_2854, Midori_rounds_sub_sBox_PRINCE_0_n13}), .b ({new_AGEMA_signal_3294, new_AGEMA_signal_3293, new_AGEMA_signal_3292, Midori_rounds_sub_sBox_PRINCE_0_n3}), .clk (clk), .r ({Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, new_AGEMA_signal_3529, Midori_rounds_SR_Result[48]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U17 ( .a ({new_AGEMA_signal_2862, new_AGEMA_signal_2861, new_AGEMA_signal_2860, Midori_rounds_sub_sBox_PRINCE_1_n15}), .b ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, new_AGEMA_signal_3301, Midori_rounds_sub_sBox_PRINCE_1_n12}), .clk (clk), .r ({Fresh[1361], Fresh[1360], Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, new_AGEMA_signal_3535, Midori_rounds_SR_Result[46]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U8 ( .a ({new_AGEMA_signal_2874, new_AGEMA_signal_2873, new_AGEMA_signal_2872, Midori_rounds_sub_sBox_PRINCE_1_n13}), .b ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, new_AGEMA_signal_3307, Midori_rounds_sub_sBox_PRINCE_1_n3}), .clk (clk), .r ({Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362]}), .c ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, new_AGEMA_signal_3541, Midori_rounds_SR_Result[44]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U17 ( .a ({new_AGEMA_signal_2880, new_AGEMA_signal_2879, new_AGEMA_signal_2878, Midori_rounds_sub_sBox_PRINCE_2_n15}), .b ({new_AGEMA_signal_3318, new_AGEMA_signal_3317, new_AGEMA_signal_3316, Midori_rounds_sub_sBox_PRINCE_2_n12}), .clk (clk), .r ({Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, new_AGEMA_signal_3547, Midori_rounds_SR_Result[10]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U8 ( .a ({new_AGEMA_signal_2892, new_AGEMA_signal_2891, new_AGEMA_signal_2890, Midori_rounds_sub_sBox_PRINCE_2_n13}), .b ({new_AGEMA_signal_3324, new_AGEMA_signal_3323, new_AGEMA_signal_3322, Midori_rounds_sub_sBox_PRINCE_2_n3}), .clk (clk), .r ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374]}), .c ({new_AGEMA_signal_3555, new_AGEMA_signal_3554, new_AGEMA_signal_3553, Midori_rounds_SR_Result[8]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U17 ( .a ({new_AGEMA_signal_2898, new_AGEMA_signal_2897, new_AGEMA_signal_2896, Midori_rounds_sub_sBox_PRINCE_3_n15}), .b ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, new_AGEMA_signal_3331, Midori_rounds_sub_sBox_PRINCE_3_n12}), .clk (clk), .r ({Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, new_AGEMA_signal_3559, Midori_rounds_SR_Result[22]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U8 ( .a ({new_AGEMA_signal_2910, new_AGEMA_signal_2909, new_AGEMA_signal_2908, Midori_rounds_sub_sBox_PRINCE_3_n13}), .b ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, new_AGEMA_signal_3337, Midori_rounds_sub_sBox_PRINCE_3_n3}), .clk (clk), .r ({Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386]}), .c ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, new_AGEMA_signal_3565, Midori_rounds_SR_Result[20]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U17 ( .a ({new_AGEMA_signal_2916, new_AGEMA_signal_2915, new_AGEMA_signal_2914, Midori_rounds_sub_sBox_PRINCE_4_n15}), .b ({new_AGEMA_signal_3348, new_AGEMA_signal_3347, new_AGEMA_signal_3346, Midori_rounds_sub_sBox_PRINCE_4_n12}), .clk (clk), .r ({Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, new_AGEMA_signal_3571, Midori_rounds_SR_Result[38]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U8 ( .a ({new_AGEMA_signal_2928, new_AGEMA_signal_2927, new_AGEMA_signal_2926, Midori_rounds_sub_sBox_PRINCE_4_n13}), .b ({new_AGEMA_signal_3354, new_AGEMA_signal_3353, new_AGEMA_signal_3352, Midori_rounds_sub_sBox_PRINCE_4_n3}), .clk (clk), .r ({Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400], Fresh[1399], Fresh[1398]}), .c ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, new_AGEMA_signal_3577, Midori_rounds_SR_Result[36]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U17 ( .a ({new_AGEMA_signal_2934, new_AGEMA_signal_2933, new_AGEMA_signal_2932, Midori_rounds_sub_sBox_PRINCE_5_n15}), .b ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, new_AGEMA_signal_3361, Midori_rounds_sub_sBox_PRINCE_5_n12}), .clk (clk), .r ({Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, new_AGEMA_signal_3583, Midori_rounds_SR_Result[58]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U8 ( .a ({new_AGEMA_signal_2946, new_AGEMA_signal_2945, new_AGEMA_signal_2944, Midori_rounds_sub_sBox_PRINCE_5_n13}), .b ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, new_AGEMA_signal_3367, Midori_rounds_sub_sBox_PRINCE_5_n3}), .clk (clk), .r ({Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, new_AGEMA_signal_3589, Midori_rounds_SR_Result[56]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U17 ( .a ({new_AGEMA_signal_2952, new_AGEMA_signal_2951, new_AGEMA_signal_2950, Midori_rounds_sub_sBox_PRINCE_6_n15}), .b ({new_AGEMA_signal_3378, new_AGEMA_signal_3377, new_AGEMA_signal_3376, Midori_rounds_sub_sBox_PRINCE_6_n12}), .clk (clk), .r ({Fresh[1421], Fresh[1420], Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, new_AGEMA_signal_3595, Midori_rounds_SR_Result[30]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U8 ( .a ({new_AGEMA_signal_2964, new_AGEMA_signal_2963, new_AGEMA_signal_2962, Midori_rounds_sub_sBox_PRINCE_6_n13}), .b ({new_AGEMA_signal_3384, new_AGEMA_signal_3383, new_AGEMA_signal_3382, Midori_rounds_sub_sBox_PRINCE_6_n3}), .clk (clk), .r ({Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422]}), .c ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, new_AGEMA_signal_3601, Midori_rounds_SR_Result[28]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U17 ( .a ({new_AGEMA_signal_2970, new_AGEMA_signal_2969, new_AGEMA_signal_2968, Midori_rounds_sub_sBox_PRINCE_7_n15}), .b ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, new_AGEMA_signal_3391, Midori_rounds_sub_sBox_PRINCE_7_n12}), .clk (clk), .r ({Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, new_AGEMA_signal_3607, Midori_rounds_SR_Result[2]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U8 ( .a ({new_AGEMA_signal_2982, new_AGEMA_signal_2981, new_AGEMA_signal_2980, Midori_rounds_sub_sBox_PRINCE_7_n13}), .b ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, new_AGEMA_signal_3397, Midori_rounds_sub_sBox_PRINCE_7_n3}), .clk (clk), .r ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434]}), .c ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, new_AGEMA_signal_3613, Midori_rounds_SR_Result[0]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U17 ( .a ({new_AGEMA_signal_2988, new_AGEMA_signal_2987, new_AGEMA_signal_2986, Midori_rounds_sub_sBox_PRINCE_8_n15}), .b ({new_AGEMA_signal_3408, new_AGEMA_signal_3407, new_AGEMA_signal_3406, Midori_rounds_sub_sBox_PRINCE_8_n12}), .clk (clk), .r ({Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, new_AGEMA_signal_3619, Midori_rounds_SR_Result[14]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U8 ( .a ({new_AGEMA_signal_3000, new_AGEMA_signal_2999, new_AGEMA_signal_2998, Midori_rounds_sub_sBox_PRINCE_8_n13}), .b ({new_AGEMA_signal_3414, new_AGEMA_signal_3413, new_AGEMA_signal_3412, Midori_rounds_sub_sBox_PRINCE_8_n3}), .clk (clk), .r ({Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446]}), .c ({new_AGEMA_signal_3627, new_AGEMA_signal_3626, new_AGEMA_signal_3625, Midori_rounds_SR_Result[12]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U17 ( .a ({new_AGEMA_signal_3006, new_AGEMA_signal_3005, new_AGEMA_signal_3004, Midori_rounds_sub_sBox_PRINCE_9_n15}), .b ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, new_AGEMA_signal_3421, Midori_rounds_sub_sBox_PRINCE_9_n12}), .clk (clk), .r ({Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, new_AGEMA_signal_3631, Midori_rounds_SR_Result[18]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U8 ( .a ({new_AGEMA_signal_3018, new_AGEMA_signal_3017, new_AGEMA_signal_3016, Midori_rounds_sub_sBox_PRINCE_9_n13}), .b ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, new_AGEMA_signal_3427, Midori_rounds_sub_sBox_PRINCE_9_n3}), .clk (clk), .r ({Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460], Fresh[1459], Fresh[1458]}), .c ({new_AGEMA_signal_3639, new_AGEMA_signal_3638, new_AGEMA_signal_3637, Midori_rounds_SR_Result[16]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U17 ( .a ({new_AGEMA_signal_3024, new_AGEMA_signal_3023, new_AGEMA_signal_3022, Midori_rounds_sub_sBox_PRINCE_10_n15}), .b ({new_AGEMA_signal_3438, new_AGEMA_signal_3437, new_AGEMA_signal_3436, Midori_rounds_sub_sBox_PRINCE_10_n12}), .clk (clk), .r ({Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, new_AGEMA_signal_3643, Midori_rounds_SR_Result[54]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U8 ( .a ({new_AGEMA_signal_3036, new_AGEMA_signal_3035, new_AGEMA_signal_3034, Midori_rounds_sub_sBox_PRINCE_10_n13}), .b ({new_AGEMA_signal_3444, new_AGEMA_signal_3443, new_AGEMA_signal_3442, Midori_rounds_sub_sBox_PRINCE_10_n3}), .clk (clk), .r ({Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, new_AGEMA_signal_3649, Midori_rounds_SR_Result[52]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U17 ( .a ({new_AGEMA_signal_3042, new_AGEMA_signal_3041, new_AGEMA_signal_3040, Midori_rounds_sub_sBox_PRINCE_11_n15}), .b ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, new_AGEMA_signal_3451, Midori_rounds_sub_sBox_PRINCE_11_n12}), .clk (clk), .r ({Fresh[1481], Fresh[1480], Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, new_AGEMA_signal_3655, Midori_rounds_SR_Result[42]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U8 ( .a ({new_AGEMA_signal_3054, new_AGEMA_signal_3053, new_AGEMA_signal_3052, Midori_rounds_sub_sBox_PRINCE_11_n13}), .b ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, new_AGEMA_signal_3457, Midori_rounds_sub_sBox_PRINCE_11_n3}), .clk (clk), .r ({Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482]}), .c ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, new_AGEMA_signal_3661, Midori_rounds_SR_Result[40]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U17 ( .a ({new_AGEMA_signal_3060, new_AGEMA_signal_3059, new_AGEMA_signal_3058, Midori_rounds_sub_sBox_PRINCE_12_n15}), .b ({new_AGEMA_signal_3468, new_AGEMA_signal_3467, new_AGEMA_signal_3466, Midori_rounds_sub_sBox_PRINCE_12_n12}), .clk (clk), .r ({Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, new_AGEMA_signal_3667, Midori_rounds_SR_Result[26]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U8 ( .a ({new_AGEMA_signal_3072, new_AGEMA_signal_3071, new_AGEMA_signal_3070, Midori_rounds_sub_sBox_PRINCE_12_n13}), .b ({new_AGEMA_signal_3474, new_AGEMA_signal_3473, new_AGEMA_signal_3472, Midori_rounds_sub_sBox_PRINCE_12_n3}), .clk (clk), .r ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494]}), .c ({new_AGEMA_signal_3675, new_AGEMA_signal_3674, new_AGEMA_signal_3673, Midori_rounds_SR_Result[24]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U17 ( .a ({new_AGEMA_signal_3078, new_AGEMA_signal_3077, new_AGEMA_signal_3076, Midori_rounds_sub_sBox_PRINCE_13_n15}), .b ({new_AGEMA_signal_3483, new_AGEMA_signal_3482, new_AGEMA_signal_3481, Midori_rounds_sub_sBox_PRINCE_13_n12}), .clk (clk), .r ({Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, new_AGEMA_signal_3679, Midori_rounds_SR_Result[6]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U8 ( .a ({new_AGEMA_signal_3090, new_AGEMA_signal_3089, new_AGEMA_signal_3088, Midori_rounds_sub_sBox_PRINCE_13_n13}), .b ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, new_AGEMA_signal_3487, Midori_rounds_sub_sBox_PRINCE_13_n3}), .clk (clk), .r ({Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506]}), .c ({new_AGEMA_signal_3687, new_AGEMA_signal_3686, new_AGEMA_signal_3685, Midori_rounds_SR_Result[4]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U17 ( .a ({new_AGEMA_signal_3096, new_AGEMA_signal_3095, new_AGEMA_signal_3094, Midori_rounds_sub_sBox_PRINCE_14_n15}), .b ({new_AGEMA_signal_3498, new_AGEMA_signal_3497, new_AGEMA_signal_3496, Midori_rounds_sub_sBox_PRINCE_14_n12}), .clk (clk), .r ({Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, new_AGEMA_signal_3691, Midori_rounds_SR_Result[34]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U8 ( .a ({new_AGEMA_signal_3108, new_AGEMA_signal_3107, new_AGEMA_signal_3106, Midori_rounds_sub_sBox_PRINCE_14_n13}), .b ({new_AGEMA_signal_3504, new_AGEMA_signal_3503, new_AGEMA_signal_3502, Midori_rounds_sub_sBox_PRINCE_14_n3}), .clk (clk), .r ({Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520], Fresh[1519], Fresh[1518]}), .c ({new_AGEMA_signal_3699, new_AGEMA_signal_3698, new_AGEMA_signal_3697, Midori_rounds_SR_Result[32]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U17 ( .a ({new_AGEMA_signal_3114, new_AGEMA_signal_3113, new_AGEMA_signal_3112, Midori_rounds_sub_sBox_PRINCE_15_n15}), .b ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, new_AGEMA_signal_3511, Midori_rounds_sub_sBox_PRINCE_15_n12}), .clk (clk), .r ({Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, new_AGEMA_signal_3703, Midori_rounds_SR_Result[62]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U8 ( .a ({new_AGEMA_signal_3126, new_AGEMA_signal_3125, new_AGEMA_signal_3124, Midori_rounds_sub_sBox_PRINCE_15_n13}), .b ({new_AGEMA_signal_3519, new_AGEMA_signal_3518, new_AGEMA_signal_3517, Midori_rounds_sub_sBox_PRINCE_15_n3}), .clk (clk), .r ({Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({new_AGEMA_signal_3711, new_AGEMA_signal_3710, new_AGEMA_signal_3709, Midori_rounds_SR_Result[60]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_0_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, new_AGEMA_signal_3613, Midori_rounds_SR_Result[0]}), .a ({new_AGEMA_signal_4779, new_AGEMA_signal_4778, new_AGEMA_signal_4777, Midori_rounds_sub_ResultXORkey[0]}), .c ({new_AGEMA_signal_4947, new_AGEMA_signal_4946, new_AGEMA_signal_4945, Midori_rounds_mul_input[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_2_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, new_AGEMA_signal_3607, Midori_rounds_SR_Result[2]}), .a ({new_AGEMA_signal_3999, new_AGEMA_signal_3998, new_AGEMA_signal_3997, Midori_rounds_sub_ResultXORkey[2]}), .c ({new_AGEMA_signal_4053, new_AGEMA_signal_4052, new_AGEMA_signal_4051, Midori_rounds_mul_input[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_4_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3687, new_AGEMA_signal_3686, new_AGEMA_signal_3685, Midori_rounds_SR_Result[4]}), .a ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, new_AGEMA_signal_4759, Midori_rounds_sub_ResultXORkey[4]}), .c ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, Midori_rounds_mul_input[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_6_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, new_AGEMA_signal_3679, Midori_rounds_SR_Result[6]}), .a ({new_AGEMA_signal_3912, new_AGEMA_signal_3911, new_AGEMA_signal_3910, Midori_rounds_sub_ResultXORkey[6]}), .c ({new_AGEMA_signal_4062, new_AGEMA_signal_4061, new_AGEMA_signal_4060, Midori_rounds_mul_input[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_8_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3555, new_AGEMA_signal_3554, new_AGEMA_signal_3553, Midori_rounds_SR_Result[8]}), .a ({new_AGEMA_signal_4566, new_AGEMA_signal_4565, new_AGEMA_signal_4564, Midori_rounds_sub_ResultXORkey[8]}), .c ({new_AGEMA_signal_4929, new_AGEMA_signal_4928, new_AGEMA_signal_4927, Midori_rounds_mul_input[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_10_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, new_AGEMA_signal_3547, Midori_rounds_SR_Result[10]}), .a ({new_AGEMA_signal_4047, new_AGEMA_signal_4046, new_AGEMA_signal_4045, Midori_rounds_sub_ResultXORkey[10]}), .c ({new_AGEMA_signal_4071, new_AGEMA_signal_4070, new_AGEMA_signal_4069, Midori_rounds_mul_input[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_12_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3627, new_AGEMA_signal_3626, new_AGEMA_signal_3625, Midori_rounds_SR_Result[12]}), .a ({new_AGEMA_signal_4776, new_AGEMA_signal_4775, new_AGEMA_signal_4774, Midori_rounds_sub_ResultXORkey[12]}), .c ({new_AGEMA_signal_4953, new_AGEMA_signal_4952, new_AGEMA_signal_4951, Midori_rounds_mul_input[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_14_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, new_AGEMA_signal_3619, Midori_rounds_SR_Result[14]}), .a ({new_AGEMA_signal_4038, new_AGEMA_signal_4037, new_AGEMA_signal_4036, Midori_rounds_sub_ResultXORkey[14]}), .c ({new_AGEMA_signal_4080, new_AGEMA_signal_4079, new_AGEMA_signal_4078, Midori_rounds_mul_input[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_16_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3639, new_AGEMA_signal_3638, new_AGEMA_signal_3637, Midori_rounds_SR_Result[16]}), .a ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, new_AGEMA_signal_4771, Midori_rounds_sub_ResultXORkey[16]}), .c ({new_AGEMA_signal_4956, new_AGEMA_signal_4955, new_AGEMA_signal_4954, Midori_rounds_mul_input[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_18_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, new_AGEMA_signal_3631, Midori_rounds_SR_Result[18]}), .a ({new_AGEMA_signal_4029, new_AGEMA_signal_4028, new_AGEMA_signal_4027, Midori_rounds_sub_ResultXORkey[18]}), .c ({new_AGEMA_signal_4089, new_AGEMA_signal_4088, new_AGEMA_signal_4087, Midori_rounds_mul_input[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_20_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, new_AGEMA_signal_3565, Midori_rounds_SR_Result[20]}), .a ({new_AGEMA_signal_4575, new_AGEMA_signal_4574, new_AGEMA_signal_4573, Midori_rounds_sub_ResultXORkey[20]}), .c ({new_AGEMA_signal_4932, new_AGEMA_signal_4931, new_AGEMA_signal_4930, Midori_rounds_mul_input[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_22_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, new_AGEMA_signal_3559, Midori_rounds_SR_Result[22]}), .a ({new_AGEMA_signal_4017, new_AGEMA_signal_4016, new_AGEMA_signal_4015, Midori_rounds_sub_ResultXORkey[22]}), .c ({new_AGEMA_signal_4098, new_AGEMA_signal_4097, new_AGEMA_signal_4096, Midori_rounds_mul_input[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_24_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3675, new_AGEMA_signal_3674, new_AGEMA_signal_3673, Midori_rounds_SR_Result[24]}), .a ({new_AGEMA_signal_4770, new_AGEMA_signal_4769, new_AGEMA_signal_4768, Midori_rounds_sub_ResultXORkey[24]}), .c ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, new_AGEMA_signal_4957, Midori_rounds_mul_input[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_26_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, new_AGEMA_signal_3667, Midori_rounds_SR_Result[26]}), .a ({new_AGEMA_signal_4008, new_AGEMA_signal_4007, new_AGEMA_signal_4006, Midori_rounds_sub_ResultXORkey[26]}), .c ({new_AGEMA_signal_4107, new_AGEMA_signal_4106, new_AGEMA_signal_4105, Midori_rounds_mul_input[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_28_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, new_AGEMA_signal_3601, Midori_rounds_SR_Result[28]}), .a ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, new_AGEMA_signal_4939, Midori_rounds_sub_ResultXORkey[28]}), .c ({new_AGEMA_signal_4980, new_AGEMA_signal_4979, new_AGEMA_signal_4978, Midori_rounds_mul_input[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_30_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, new_AGEMA_signal_3595, Midori_rounds_SR_Result[30]}), .a ({new_AGEMA_signal_3996, new_AGEMA_signal_3995, new_AGEMA_signal_3994, Midori_rounds_sub_ResultXORkey[30]}), .c ({new_AGEMA_signal_4116, new_AGEMA_signal_4115, new_AGEMA_signal_4114, Midori_rounds_mul_input[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_32_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3699, new_AGEMA_signal_3698, new_AGEMA_signal_3697, Midori_rounds_SR_Result[32]}), .a ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, new_AGEMA_signal_4765, Midori_rounds_sub_ResultXORkey[32]}), .c ({new_AGEMA_signal_4962, new_AGEMA_signal_4961, new_AGEMA_signal_4960, Midori_rounds_mul_input[32]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_34_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, new_AGEMA_signal_3691, Midori_rounds_SR_Result[34]}), .a ({new_AGEMA_signal_3987, new_AGEMA_signal_3986, new_AGEMA_signal_3985, Midori_rounds_sub_ResultXORkey[34]}), .c ({new_AGEMA_signal_4125, new_AGEMA_signal_4124, new_AGEMA_signal_4123, Midori_rounds_mul_input[34]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_36_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, new_AGEMA_signal_3577, Midori_rounds_SR_Result[36]}), .a ({new_AGEMA_signal_4572, new_AGEMA_signal_4571, new_AGEMA_signal_4570, Midori_rounds_sub_ResultXORkey[36]}), .c ({new_AGEMA_signal_4935, new_AGEMA_signal_4934, new_AGEMA_signal_4933, Midori_rounds_mul_input[36]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_38_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, new_AGEMA_signal_3571, Midori_rounds_SR_Result[38]}), .a ({new_AGEMA_signal_3978, new_AGEMA_signal_3977, new_AGEMA_signal_3976, Midori_rounds_sub_ResultXORkey[38]}), .c ({new_AGEMA_signal_4134, new_AGEMA_signal_4133, new_AGEMA_signal_4132, Midori_rounds_mul_input[38]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_40_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, new_AGEMA_signal_3661, Midori_rounds_SR_Result[40]}), .a ({new_AGEMA_signal_4764, new_AGEMA_signal_4763, new_AGEMA_signal_4762, Midori_rounds_sub_ResultXORkey[40]}), .c ({new_AGEMA_signal_4965, new_AGEMA_signal_4964, new_AGEMA_signal_4963, Midori_rounds_mul_input[40]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_42_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, new_AGEMA_signal_3655, Midori_rounds_SR_Result[42]}), .a ({new_AGEMA_signal_3966, new_AGEMA_signal_3965, new_AGEMA_signal_3964, Midori_rounds_sub_ResultXORkey[42]}), .c ({new_AGEMA_signal_4143, new_AGEMA_signal_4142, new_AGEMA_signal_4141, Midori_rounds_mul_input[42]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_44_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, new_AGEMA_signal_3541, Midori_rounds_SR_Result[44]}), .a ({new_AGEMA_signal_4569, new_AGEMA_signal_4568, new_AGEMA_signal_4567, Midori_rounds_sub_ResultXORkey[44]}), .c ({new_AGEMA_signal_4938, new_AGEMA_signal_4937, new_AGEMA_signal_4936, Midori_rounds_mul_input[44]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_46_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, new_AGEMA_signal_3535, Midori_rounds_SR_Result[46]}), .a ({new_AGEMA_signal_3957, new_AGEMA_signal_3956, new_AGEMA_signal_3955, Midori_rounds_sub_ResultXORkey[46]}), .c ({new_AGEMA_signal_4152, new_AGEMA_signal_4151, new_AGEMA_signal_4150, Midori_rounds_mul_input[46]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_48_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, new_AGEMA_signal_3529, Midori_rounds_SR_Result[48]}), .a ({new_AGEMA_signal_4977, new_AGEMA_signal_4976, new_AGEMA_signal_4975, Midori_rounds_sub_ResultXORkey[48]}), .c ({new_AGEMA_signal_5001, new_AGEMA_signal_5000, new_AGEMA_signal_4999, Midori_rounds_mul_input[48]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_50_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, new_AGEMA_signal_3523, Midori_rounds_SR_Result[50]}), .a ({new_AGEMA_signal_3948, new_AGEMA_signal_3947, new_AGEMA_signal_3946, Midori_rounds_sub_ResultXORkey[50]}), .c ({new_AGEMA_signal_4161, new_AGEMA_signal_4160, new_AGEMA_signal_4159, Midori_rounds_mul_input[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_52_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, new_AGEMA_signal_3649, Midori_rounds_SR_Result[52]}), .a ({new_AGEMA_signal_4758, new_AGEMA_signal_4757, new_AGEMA_signal_4756, Midori_rounds_sub_ResultXORkey[52]}), .c ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, new_AGEMA_signal_4966, Midori_rounds_mul_input[52]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_54_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, new_AGEMA_signal_3643, Midori_rounds_SR_Result[54]}), .a ({new_AGEMA_signal_3939, new_AGEMA_signal_3938, new_AGEMA_signal_3937, Midori_rounds_sub_ResultXORkey[54]}), .c ({new_AGEMA_signal_4170, new_AGEMA_signal_4169, new_AGEMA_signal_4168, Midori_rounds_mul_input[54]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_56_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, new_AGEMA_signal_3589, Midori_rounds_SR_Result[56]}), .a ({new_AGEMA_signal_4755, new_AGEMA_signal_4754, new_AGEMA_signal_4753, Midori_rounds_sub_ResultXORkey[56]}), .c ({new_AGEMA_signal_4971, new_AGEMA_signal_4970, new_AGEMA_signal_4969, Midori_rounds_mul_input[56]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_58_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, new_AGEMA_signal_3583, Midori_rounds_SR_Result[58]}), .a ({new_AGEMA_signal_3930, new_AGEMA_signal_3929, new_AGEMA_signal_3928, Midori_rounds_sub_ResultXORkey[58]}), .c ({new_AGEMA_signal_4179, new_AGEMA_signal_4178, new_AGEMA_signal_4177, Midori_rounds_mul_input[58]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_60_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3711, new_AGEMA_signal_3710, new_AGEMA_signal_3709, Midori_rounds_SR_Result[60]}), .a ({new_AGEMA_signal_4752, new_AGEMA_signal_4751, new_AGEMA_signal_4750, Midori_rounds_sub_ResultXORkey[60]}), .c ({new_AGEMA_signal_4974, new_AGEMA_signal_4973, new_AGEMA_signal_4972, Midori_rounds_mul_input[60]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_62_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, new_AGEMA_signal_3703, Midori_rounds_SR_Result[62]}), .a ({new_AGEMA_signal_3918, new_AGEMA_signal_3917, new_AGEMA_signal_3916, Midori_rounds_sub_ResultXORkey[62]}), .c ({new_AGEMA_signal_4188, new_AGEMA_signal_4187, new_AGEMA_signal_4186, Midori_rounds_mul_input[62]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U23 ( .a ({new_AGEMA_signal_4974, new_AGEMA_signal_4973, new_AGEMA_signal_4972, Midori_rounds_mul_input[60]}), .b ({new_AGEMA_signal_5076, new_AGEMA_signal_5075, new_AGEMA_signal_5074, Midori_rounds_mul_MC1_n7}), .c ({new_AGEMA_signal_5094, new_AGEMA_signal_5093, new_AGEMA_signal_5092, Midori_rounds_SR_Inv_Result[20]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U21 ( .a ({new_AGEMA_signal_4161, new_AGEMA_signal_4160, new_AGEMA_signal_4159, Midori_rounds_mul_input[50]}), .b ({new_AGEMA_signal_4197, new_AGEMA_signal_4196, new_AGEMA_signal_4195, Midori_rounds_mul_MC1_n5}), .c ({new_AGEMA_signal_4272, new_AGEMA_signal_4271, new_AGEMA_signal_4270, Midori_rounds_SR_Inv_Result[42]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U19 ( .a ({new_AGEMA_signal_5001, new_AGEMA_signal_5000, new_AGEMA_signal_4999, Midori_rounds_mul_input[48]}), .b ({new_AGEMA_signal_4983, new_AGEMA_signal_4982, new_AGEMA_signal_4981, Midori_rounds_mul_MC1_n3}), .c ({new_AGEMA_signal_5073, new_AGEMA_signal_5072, new_AGEMA_signal_5071, Midori_rounds_SR_Inv_Result[40]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U16 ( .a ({new_AGEMA_signal_4170, new_AGEMA_signal_4169, new_AGEMA_signal_4168, Midori_rounds_mul_input[54]}), .b ({new_AGEMA_signal_4197, new_AGEMA_signal_4196, new_AGEMA_signal_4195, Midori_rounds_mul_MC1_n5}), .c ({new_AGEMA_signal_4281, new_AGEMA_signal_4280, new_AGEMA_signal_4279, Midori_rounds_SR_Inv_Result[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U15 ( .a ({new_AGEMA_signal_4188, new_AGEMA_signal_4187, new_AGEMA_signal_4186, Midori_rounds_mul_input[62]}), .b ({new_AGEMA_signal_4179, new_AGEMA_signal_4178, new_AGEMA_signal_4177, Midori_rounds_mul_input[58]}), .c ({new_AGEMA_signal_4197, new_AGEMA_signal_4196, new_AGEMA_signal_4195, Midori_rounds_mul_MC1_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U11 ( .a ({new_AGEMA_signal_4179, new_AGEMA_signal_4178, new_AGEMA_signal_4177, Midori_rounds_mul_input[58]}), .b ({new_AGEMA_signal_4209, new_AGEMA_signal_4208, new_AGEMA_signal_4207, Midori_rounds_mul_MC1_n1}), .c ({new_AGEMA_signal_4290, new_AGEMA_signal_4289, new_AGEMA_signal_4288, Midori_rounds_SR_Inv_Result[62]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U8 ( .a ({new_AGEMA_signal_4971, new_AGEMA_signal_4970, new_AGEMA_signal_4969, Midori_rounds_mul_input[56]}), .b ({new_AGEMA_signal_5076, new_AGEMA_signal_5075, new_AGEMA_signal_5074, Midori_rounds_mul_MC1_n7}), .c ({new_AGEMA_signal_5097, new_AGEMA_signal_5096, new_AGEMA_signal_5095, Midori_rounds_SR_Inv_Result[60]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U7 ( .a ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, new_AGEMA_signal_4966, Midori_rounds_mul_input[52]}), .b ({new_AGEMA_signal_5001, new_AGEMA_signal_5000, new_AGEMA_signal_4999, Midori_rounds_mul_input[48]}), .c ({new_AGEMA_signal_5076, new_AGEMA_signal_5075, new_AGEMA_signal_5074, Midori_rounds_mul_MC1_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U4 ( .a ({new_AGEMA_signal_4188, new_AGEMA_signal_4187, new_AGEMA_signal_4186, Midori_rounds_mul_input[62]}), .b ({new_AGEMA_signal_4209, new_AGEMA_signal_4208, new_AGEMA_signal_4207, Midori_rounds_mul_MC1_n1}), .c ({new_AGEMA_signal_4299, new_AGEMA_signal_4298, new_AGEMA_signal_4297, Midori_rounds_SR_Inv_Result[22]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U3 ( .a ({new_AGEMA_signal_4161, new_AGEMA_signal_4160, new_AGEMA_signal_4159, Midori_rounds_mul_input[50]}), .b ({new_AGEMA_signal_4170, new_AGEMA_signal_4169, new_AGEMA_signal_4168, Midori_rounds_mul_input[54]}), .c ({new_AGEMA_signal_4209, new_AGEMA_signal_4208, new_AGEMA_signal_4207, Midori_rounds_mul_MC1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U2 ( .a ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, new_AGEMA_signal_4966, Midori_rounds_mul_input[52]}), .b ({new_AGEMA_signal_4983, new_AGEMA_signal_4982, new_AGEMA_signal_4981, Midori_rounds_mul_MC1_n3}), .c ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, new_AGEMA_signal_5002, Midori_rounds_SR_Inv_Result[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC1_U1 ( .a ({new_AGEMA_signal_4974, new_AGEMA_signal_4973, new_AGEMA_signal_4972, Midori_rounds_mul_input[60]}), .b ({new_AGEMA_signal_4971, new_AGEMA_signal_4970, new_AGEMA_signal_4969, Midori_rounds_mul_input[56]}), .c ({new_AGEMA_signal_4983, new_AGEMA_signal_4982, new_AGEMA_signal_4981, Midori_rounds_mul_MC1_n3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U23 ( .a ({new_AGEMA_signal_4938, new_AGEMA_signal_4937, new_AGEMA_signal_4936, Midori_rounds_mul_input[44]}), .b ({new_AGEMA_signal_4986, new_AGEMA_signal_4985, new_AGEMA_signal_4984, Midori_rounds_mul_MC2_n7}), .c ({new_AGEMA_signal_5007, new_AGEMA_signal_5006, new_AGEMA_signal_5005, Midori_rounds_SR_Inv_Result[44]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U21 ( .a ({new_AGEMA_signal_4125, new_AGEMA_signal_4124, new_AGEMA_signal_4123, Midori_rounds_mul_input[34]}), .b ({new_AGEMA_signal_4215, new_AGEMA_signal_4214, new_AGEMA_signal_4213, Midori_rounds_mul_MC2_n5}), .c ({new_AGEMA_signal_4308, new_AGEMA_signal_4307, new_AGEMA_signal_4306, Midori_rounds_SR_Inv_Result[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U19 ( .a ({new_AGEMA_signal_4962, new_AGEMA_signal_4961, new_AGEMA_signal_4960, Midori_rounds_mul_input[32]}), .b ({new_AGEMA_signal_4989, new_AGEMA_signal_4988, new_AGEMA_signal_4987, Midori_rounds_mul_MC2_n3}), .c ({new_AGEMA_signal_5010, new_AGEMA_signal_5009, new_AGEMA_signal_5008, Midori_rounds_SR_Inv_Result[16]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U16 ( .a ({new_AGEMA_signal_4134, new_AGEMA_signal_4133, new_AGEMA_signal_4132, Midori_rounds_mul_input[38]}), .b ({new_AGEMA_signal_4215, new_AGEMA_signal_4214, new_AGEMA_signal_4213, Midori_rounds_mul_MC2_n5}), .c ({new_AGEMA_signal_4317, new_AGEMA_signal_4316, new_AGEMA_signal_4315, Midori_rounds_SR_Inv_Result[58]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U15 ( .a ({new_AGEMA_signal_4152, new_AGEMA_signal_4151, new_AGEMA_signal_4150, Midori_rounds_mul_input[46]}), .b ({new_AGEMA_signal_4143, new_AGEMA_signal_4142, new_AGEMA_signal_4141, Midori_rounds_mul_input[42]}), .c ({new_AGEMA_signal_4215, new_AGEMA_signal_4214, new_AGEMA_signal_4213, Midori_rounds_mul_MC2_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U11 ( .a ({new_AGEMA_signal_4143, new_AGEMA_signal_4142, new_AGEMA_signal_4141, Midori_rounds_mul_input[42]}), .b ({new_AGEMA_signal_4227, new_AGEMA_signal_4226, new_AGEMA_signal_4225, Midori_rounds_mul_MC2_n1}), .c ({new_AGEMA_signal_4326, new_AGEMA_signal_4325, new_AGEMA_signal_4324, Midori_rounds_SR_Inv_Result[6]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U8 ( .a ({new_AGEMA_signal_4965, new_AGEMA_signal_4964, new_AGEMA_signal_4963, Midori_rounds_mul_input[40]}), .b ({new_AGEMA_signal_4986, new_AGEMA_signal_4985, new_AGEMA_signal_4984, Midori_rounds_mul_MC2_n7}), .c ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, new_AGEMA_signal_5011, Midori_rounds_SR_Inv_Result[4]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U7 ( .a ({new_AGEMA_signal_4935, new_AGEMA_signal_4934, new_AGEMA_signal_4933, Midori_rounds_mul_input[36]}), .b ({new_AGEMA_signal_4962, new_AGEMA_signal_4961, new_AGEMA_signal_4960, Midori_rounds_mul_input[32]}), .c ({new_AGEMA_signal_4986, new_AGEMA_signal_4985, new_AGEMA_signal_4984, Midori_rounds_mul_MC2_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U4 ( .a ({new_AGEMA_signal_4152, new_AGEMA_signal_4151, new_AGEMA_signal_4150, Midori_rounds_mul_input[46]}), .b ({new_AGEMA_signal_4227, new_AGEMA_signal_4226, new_AGEMA_signal_4225, Midori_rounds_mul_MC2_n1}), .c ({new_AGEMA_signal_4335, new_AGEMA_signal_4334, new_AGEMA_signal_4333, Midori_rounds_SR_Inv_Result[46]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U3 ( .a ({new_AGEMA_signal_4125, new_AGEMA_signal_4124, new_AGEMA_signal_4123, Midori_rounds_mul_input[34]}), .b ({new_AGEMA_signal_4134, new_AGEMA_signal_4133, new_AGEMA_signal_4132, Midori_rounds_mul_input[38]}), .c ({new_AGEMA_signal_4227, new_AGEMA_signal_4226, new_AGEMA_signal_4225, Midori_rounds_mul_MC2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U2 ( .a ({new_AGEMA_signal_4935, new_AGEMA_signal_4934, new_AGEMA_signal_4933, Midori_rounds_mul_input[36]}), .b ({new_AGEMA_signal_4989, new_AGEMA_signal_4988, new_AGEMA_signal_4987, Midori_rounds_mul_MC2_n3}), .c ({new_AGEMA_signal_5016, new_AGEMA_signal_5015, new_AGEMA_signal_5014, Midori_rounds_SR_Inv_Result[56]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC2_U1 ( .a ({new_AGEMA_signal_4938, new_AGEMA_signal_4937, new_AGEMA_signal_4936, Midori_rounds_mul_input[44]}), .b ({new_AGEMA_signal_4965, new_AGEMA_signal_4964, new_AGEMA_signal_4963, Midori_rounds_mul_input[40]}), .c ({new_AGEMA_signal_4989, new_AGEMA_signal_4988, new_AGEMA_signal_4987, Midori_rounds_mul_MC2_n3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U23 ( .a ({new_AGEMA_signal_4980, new_AGEMA_signal_4979, new_AGEMA_signal_4978, Midori_rounds_mul_input[28]}), .b ({new_AGEMA_signal_4992, new_AGEMA_signal_4991, new_AGEMA_signal_4990, Midori_rounds_mul_MC3_n7}), .c ({new_AGEMA_signal_5019, new_AGEMA_signal_5018, new_AGEMA_signal_5017, Midori_rounds_SR_Inv_Result[48]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U21 ( .a ({new_AGEMA_signal_4089, new_AGEMA_signal_4088, new_AGEMA_signal_4087, Midori_rounds_mul_input[18]}), .b ({new_AGEMA_signal_4233, new_AGEMA_signal_4232, new_AGEMA_signal_4231, Midori_rounds_mul_MC3_n5}), .c ({new_AGEMA_signal_4344, new_AGEMA_signal_4343, new_AGEMA_signal_4342, Midori_rounds_SR_Inv_Result[14]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U19 ( .a ({new_AGEMA_signal_4956, new_AGEMA_signal_4955, new_AGEMA_signal_4954, Midori_rounds_mul_input[16]}), .b ({new_AGEMA_signal_5025, new_AGEMA_signal_5024, new_AGEMA_signal_5023, Midori_rounds_mul_MC3_n3}), .c ({new_AGEMA_signal_5079, new_AGEMA_signal_5078, new_AGEMA_signal_5077, Midori_rounds_SR_Inv_Result[12]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U16 ( .a ({new_AGEMA_signal_4098, new_AGEMA_signal_4097, new_AGEMA_signal_4096, Midori_rounds_mul_input[22]}), .b ({new_AGEMA_signal_4233, new_AGEMA_signal_4232, new_AGEMA_signal_4231, Midori_rounds_mul_MC3_n5}), .c ({new_AGEMA_signal_4353, new_AGEMA_signal_4352, new_AGEMA_signal_4351, Midori_rounds_SR_Inv_Result[38]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U15 ( .a ({new_AGEMA_signal_4116, new_AGEMA_signal_4115, new_AGEMA_signal_4114, Midori_rounds_mul_input[30]}), .b ({new_AGEMA_signal_4107, new_AGEMA_signal_4106, new_AGEMA_signal_4105, Midori_rounds_mul_input[26]}), .c ({new_AGEMA_signal_4233, new_AGEMA_signal_4232, new_AGEMA_signal_4231, Midori_rounds_mul_MC3_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U11 ( .a ({new_AGEMA_signal_4107, new_AGEMA_signal_4106, new_AGEMA_signal_4105, Midori_rounds_mul_input[26]}), .b ({new_AGEMA_signal_4245, new_AGEMA_signal_4244, new_AGEMA_signal_4243, Midori_rounds_mul_MC3_n1}), .c ({new_AGEMA_signal_4362, new_AGEMA_signal_4361, new_AGEMA_signal_4360, Midori_rounds_SR_Inv_Result[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U8 ( .a ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, new_AGEMA_signal_4957, Midori_rounds_mul_input[24]}), .b ({new_AGEMA_signal_4992, new_AGEMA_signal_4991, new_AGEMA_signal_4990, Midori_rounds_mul_MC3_n7}), .c ({new_AGEMA_signal_5022, new_AGEMA_signal_5021, new_AGEMA_signal_5020, Midori_rounds_SR_Inv_Result[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U7 ( .a ({new_AGEMA_signal_4932, new_AGEMA_signal_4931, new_AGEMA_signal_4930, Midori_rounds_mul_input[20]}), .b ({new_AGEMA_signal_4956, new_AGEMA_signal_4955, new_AGEMA_signal_4954, Midori_rounds_mul_input[16]}), .c ({new_AGEMA_signal_4992, new_AGEMA_signal_4991, new_AGEMA_signal_4990, Midori_rounds_mul_MC3_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U4 ( .a ({new_AGEMA_signal_4116, new_AGEMA_signal_4115, new_AGEMA_signal_4114, Midori_rounds_mul_input[30]}), .b ({new_AGEMA_signal_4245, new_AGEMA_signal_4244, new_AGEMA_signal_4243, Midori_rounds_mul_MC3_n1}), .c ({new_AGEMA_signal_4371, new_AGEMA_signal_4370, new_AGEMA_signal_4369, Midori_rounds_SR_Inv_Result[50]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U3 ( .a ({new_AGEMA_signal_4089, new_AGEMA_signal_4088, new_AGEMA_signal_4087, Midori_rounds_mul_input[18]}), .b ({new_AGEMA_signal_4098, new_AGEMA_signal_4097, new_AGEMA_signal_4096, Midori_rounds_mul_input[22]}), .c ({new_AGEMA_signal_4245, new_AGEMA_signal_4244, new_AGEMA_signal_4243, Midori_rounds_mul_MC3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U2 ( .a ({new_AGEMA_signal_4932, new_AGEMA_signal_4931, new_AGEMA_signal_4930, Midori_rounds_mul_input[20]}), .b ({new_AGEMA_signal_5025, new_AGEMA_signal_5024, new_AGEMA_signal_5023, Midori_rounds_mul_MC3_n3}), .c ({new_AGEMA_signal_5082, new_AGEMA_signal_5081, new_AGEMA_signal_5080, Midori_rounds_SR_Inv_Result[36]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC3_U1 ( .a ({new_AGEMA_signal_4980, new_AGEMA_signal_4979, new_AGEMA_signal_4978, Midori_rounds_mul_input[28]}), .b ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, new_AGEMA_signal_4957, Midori_rounds_mul_input[24]}), .c ({new_AGEMA_signal_5025, new_AGEMA_signal_5024, new_AGEMA_signal_5023, Midori_rounds_mul_MC3_n3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U23 ( .a ({new_AGEMA_signal_4953, new_AGEMA_signal_4952, new_AGEMA_signal_4951, Midori_rounds_mul_input[12]}), .b ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, new_AGEMA_signal_4993, Midori_rounds_mul_MC4_n7}), .c ({new_AGEMA_signal_5028, new_AGEMA_signal_5027, new_AGEMA_signal_5026, Midori_rounds_SR_Inv_Result[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U21 ( .a ({new_AGEMA_signal_4053, new_AGEMA_signal_4052, new_AGEMA_signal_4051, Midori_rounds_mul_input[2]}), .b ({new_AGEMA_signal_4251, new_AGEMA_signal_4250, new_AGEMA_signal_4249, Midori_rounds_mul_MC4_n5}), .c ({new_AGEMA_signal_4380, new_AGEMA_signal_4379, new_AGEMA_signal_4378, Midori_rounds_SR_Inv_Result[54]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U19 ( .a ({new_AGEMA_signal_4947, new_AGEMA_signal_4946, new_AGEMA_signal_4945, Midori_rounds_mul_input[0]}), .b ({new_AGEMA_signal_4998, new_AGEMA_signal_4997, new_AGEMA_signal_4996, Midori_rounds_mul_MC4_n3}), .c ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, new_AGEMA_signal_5029, Midori_rounds_SR_Inv_Result[52]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U16 ( .a ({new_AGEMA_signal_4062, new_AGEMA_signal_4061, new_AGEMA_signal_4060, Midori_rounds_mul_input[6]}), .b ({new_AGEMA_signal_4251, new_AGEMA_signal_4250, new_AGEMA_signal_4249, Midori_rounds_mul_MC4_n5}), .c ({new_AGEMA_signal_4389, new_AGEMA_signal_4388, new_AGEMA_signal_4387, Midori_rounds_SR_Inv_Result[30]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U15 ( .a ({new_AGEMA_signal_4080, new_AGEMA_signal_4079, new_AGEMA_signal_4078, Midori_rounds_mul_input[14]}), .b ({new_AGEMA_signal_4071, new_AGEMA_signal_4070, new_AGEMA_signal_4069, Midori_rounds_mul_input[10]}), .c ({new_AGEMA_signal_4251, new_AGEMA_signal_4250, new_AGEMA_signal_4249, Midori_rounds_mul_MC4_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U11 ( .a ({new_AGEMA_signal_4071, new_AGEMA_signal_4070, new_AGEMA_signal_4069, Midori_rounds_mul_input[10]}), .b ({new_AGEMA_signal_4263, new_AGEMA_signal_4262, new_AGEMA_signal_4261, Midori_rounds_mul_MC4_n1}), .c ({new_AGEMA_signal_4398, new_AGEMA_signal_4397, new_AGEMA_signal_4396, Midori_rounds_SR_Inv_Result[34]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U8 ( .a ({new_AGEMA_signal_4929, new_AGEMA_signal_4928, new_AGEMA_signal_4927, Midori_rounds_mul_input[8]}), .b ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, new_AGEMA_signal_4993, Midori_rounds_mul_MC4_n7}), .c ({new_AGEMA_signal_5034, new_AGEMA_signal_5033, new_AGEMA_signal_5032, Midori_rounds_SR_Inv_Result[32]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U7 ( .a ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, Midori_rounds_mul_input[4]}), .b ({new_AGEMA_signal_4947, new_AGEMA_signal_4946, new_AGEMA_signal_4945, Midori_rounds_mul_input[0]}), .c ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, new_AGEMA_signal_4993, Midori_rounds_mul_MC4_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U4 ( .a ({new_AGEMA_signal_4080, new_AGEMA_signal_4079, new_AGEMA_signal_4078, Midori_rounds_mul_input[14]}), .b ({new_AGEMA_signal_4263, new_AGEMA_signal_4262, new_AGEMA_signal_4261, Midori_rounds_mul_MC4_n1}), .c ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, new_AGEMA_signal_4405, Midori_rounds_SR_Inv_Result[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U3 ( .a ({new_AGEMA_signal_4053, new_AGEMA_signal_4052, new_AGEMA_signal_4051, Midori_rounds_mul_input[2]}), .b ({new_AGEMA_signal_4062, new_AGEMA_signal_4061, new_AGEMA_signal_4060, Midori_rounds_mul_input[6]}), .c ({new_AGEMA_signal_4263, new_AGEMA_signal_4262, new_AGEMA_signal_4261, Midori_rounds_mul_MC4_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U2 ( .a ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, Midori_rounds_mul_input[4]}), .b ({new_AGEMA_signal_4998, new_AGEMA_signal_4997, new_AGEMA_signal_4996, Midori_rounds_mul_MC4_n3}), .c ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, new_AGEMA_signal_5035, Midori_rounds_SR_Inv_Result[28]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) Midori_rounds_mul_MC4_U1 ( .a ({new_AGEMA_signal_4953, new_AGEMA_signal_4952, new_AGEMA_signal_4951, Midori_rounds_mul_input[12]}), .b ({new_AGEMA_signal_4929, new_AGEMA_signal_4928, new_AGEMA_signal_4927, Midori_rounds_mul_input[8]}), .c ({new_AGEMA_signal_4998, new_AGEMA_signal_4997, new_AGEMA_signal_4996, Midori_rounds_mul_MC4_n3}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_0_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_5070, new_AGEMA_signal_5069, new_AGEMA_signal_5068, Midori_rounds_mul_ResultXORkey[0]}), .a ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, new_AGEMA_signal_5002, Midori_rounds_SR_Inv_Result[0]}), .c ({new_AGEMA_signal_5100, new_AGEMA_signal_5099, new_AGEMA_signal_5098, Midori_rounds_round_Result[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_2_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4512, new_AGEMA_signal_4511, new_AGEMA_signal_4510, Midori_rounds_mul_ResultXORkey[2]}), .a ({new_AGEMA_signal_4281, new_AGEMA_signal_4280, new_AGEMA_signal_4279, Midori_rounds_SR_Inv_Result[2]}), .c ({new_AGEMA_signal_4611, new_AGEMA_signal_4610, new_AGEMA_signal_4609, Midori_rounds_round_Result[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_4_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_5043, new_AGEMA_signal_5042, new_AGEMA_signal_5041, Midori_rounds_mul_ResultXORkey[4]}), .a ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, new_AGEMA_signal_5011, Midori_rounds_SR_Inv_Result[4]}), .c ({new_AGEMA_signal_5103, new_AGEMA_signal_5102, new_AGEMA_signal_5101, Midori_rounds_round_Result[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_6_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4419, new_AGEMA_signal_4418, new_AGEMA_signal_4417, Midori_rounds_mul_ResultXORkey[6]}), .a ({new_AGEMA_signal_4326, new_AGEMA_signal_4325, new_AGEMA_signal_4324, Midori_rounds_SR_Inv_Result[6]}), .c ({new_AGEMA_signal_4620, new_AGEMA_signal_4619, new_AGEMA_signal_4618, Midori_rounds_round_Result[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_8_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_5040, new_AGEMA_signal_5039, new_AGEMA_signal_5038, Midori_rounds_mul_ResultXORkey[8]}), .a ({new_AGEMA_signal_5028, new_AGEMA_signal_5027, new_AGEMA_signal_5026, Midori_rounds_SR_Inv_Result[8]}), .c ({new_AGEMA_signal_5106, new_AGEMA_signal_5105, new_AGEMA_signal_5104, Midori_rounds_round_Result[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_10_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4563, new_AGEMA_signal_4562, new_AGEMA_signal_4561, Midori_rounds_mul_ResultXORkey[10]}), .a ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, new_AGEMA_signal_4405, Midori_rounds_SR_Inv_Result[10]}), .c ({new_AGEMA_signal_4629, new_AGEMA_signal_4628, new_AGEMA_signal_4627, Midori_rounds_round_Result[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_12_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_5067, new_AGEMA_signal_5066, new_AGEMA_signal_5065, Midori_rounds_mul_ResultXORkey[12]}), .a ({new_AGEMA_signal_5079, new_AGEMA_signal_5078, new_AGEMA_signal_5077, Midori_rounds_SR_Inv_Result[12]}), .c ({new_AGEMA_signal_5109, new_AGEMA_signal_5108, new_AGEMA_signal_5107, Midori_rounds_round_Result[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_14_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, Midori_rounds_mul_ResultXORkey[14]}), .a ({new_AGEMA_signal_4344, new_AGEMA_signal_4343, new_AGEMA_signal_4342, Midori_rounds_SR_Inv_Result[14]}), .c ({new_AGEMA_signal_4638, new_AGEMA_signal_4637, new_AGEMA_signal_4636, Midori_rounds_round_Result[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_16_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_5091, new_AGEMA_signal_5090, new_AGEMA_signal_5089, Midori_rounds_mul_ResultXORkey[16]}), .a ({new_AGEMA_signal_5010, new_AGEMA_signal_5009, new_AGEMA_signal_5008, Midori_rounds_SR_Inv_Result[16]}), .c ({new_AGEMA_signal_5172, new_AGEMA_signal_5171, new_AGEMA_signal_5170, Midori_rounds_round_Result[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_18_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4545, new_AGEMA_signal_4544, new_AGEMA_signal_4543, Midori_rounds_mul_ResultXORkey[18]}), .a ({new_AGEMA_signal_4308, new_AGEMA_signal_4307, new_AGEMA_signal_4306, Midori_rounds_SR_Inv_Result[18]}), .c ({new_AGEMA_signal_4647, new_AGEMA_signal_4646, new_AGEMA_signal_4645, Midori_rounds_round_Result[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_20_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_5088, new_AGEMA_signal_5087, new_AGEMA_signal_5086, Midori_rounds_mul_ResultXORkey[20]}), .a ({new_AGEMA_signal_5094, new_AGEMA_signal_5093, new_AGEMA_signal_5092, Midori_rounds_SR_Inv_Result[20]}), .c ({new_AGEMA_signal_5175, new_AGEMA_signal_5174, new_AGEMA_signal_5173, Midori_rounds_round_Result[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_22_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4530, new_AGEMA_signal_4529, new_AGEMA_signal_4528, Midori_rounds_mul_ResultXORkey[22]}), .a ({new_AGEMA_signal_4299, new_AGEMA_signal_4298, new_AGEMA_signal_4297, Midori_rounds_SR_Inv_Result[22]}), .c ({new_AGEMA_signal_4656, new_AGEMA_signal_4655, new_AGEMA_signal_4654, Midori_rounds_round_Result[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_24_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_5064, new_AGEMA_signal_5063, new_AGEMA_signal_5062, Midori_rounds_mul_ResultXORkey[24]}), .a ({new_AGEMA_signal_5022, new_AGEMA_signal_5021, new_AGEMA_signal_5020, Midori_rounds_SR_Inv_Result[24]}), .c ({new_AGEMA_signal_5112, new_AGEMA_signal_5111, new_AGEMA_signal_5110, Midori_rounds_round_Result[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_26_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4521, new_AGEMA_signal_4520, new_AGEMA_signal_4519, Midori_rounds_mul_ResultXORkey[26]}), .a ({new_AGEMA_signal_4362, new_AGEMA_signal_4361, new_AGEMA_signal_4360, Midori_rounds_SR_Inv_Result[26]}), .c ({new_AGEMA_signal_4665, new_AGEMA_signal_4664, new_AGEMA_signal_4663, Midori_rounds_round_Result[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_28_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_5061, new_AGEMA_signal_5060, new_AGEMA_signal_5059, Midori_rounds_mul_ResultXORkey[28]}), .a ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, new_AGEMA_signal_5035, Midori_rounds_SR_Inv_Result[28]}), .c ({new_AGEMA_signal_5115, new_AGEMA_signal_5114, new_AGEMA_signal_5113, Midori_rounds_round_Result[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_30_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, new_AGEMA_signal_4507, Midori_rounds_mul_ResultXORkey[30]}), .a ({new_AGEMA_signal_4389, new_AGEMA_signal_4388, new_AGEMA_signal_4387, Midori_rounds_SR_Inv_Result[30]}), .c ({new_AGEMA_signal_4674, new_AGEMA_signal_4673, new_AGEMA_signal_4672, Midori_rounds_round_Result[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_32_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_5058, new_AGEMA_signal_5057, new_AGEMA_signal_5056, Midori_rounds_mul_ResultXORkey[32]}), .a ({new_AGEMA_signal_5034, new_AGEMA_signal_5033, new_AGEMA_signal_5032, Midori_rounds_SR_Inv_Result[32]}), .c ({new_AGEMA_signal_5118, new_AGEMA_signal_5117, new_AGEMA_signal_5116, Midori_rounds_round_Result[32]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_34_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4500, new_AGEMA_signal_4499, new_AGEMA_signal_4498, Midori_rounds_mul_ResultXORkey[34]}), .a ({new_AGEMA_signal_4398, new_AGEMA_signal_4397, new_AGEMA_signal_4396, Midori_rounds_SR_Inv_Result[34]}), .c ({new_AGEMA_signal_4683, new_AGEMA_signal_4682, new_AGEMA_signal_4681, Midori_rounds_round_Result[34]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_36_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_5055, new_AGEMA_signal_5054, new_AGEMA_signal_5053, Midori_rounds_mul_ResultXORkey[36]}), .a ({new_AGEMA_signal_5082, new_AGEMA_signal_5081, new_AGEMA_signal_5080, Midori_rounds_SR_Inv_Result[36]}), .c ({new_AGEMA_signal_5121, new_AGEMA_signal_5120, new_AGEMA_signal_5119, Midori_rounds_round_Result[36]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_38_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4488, new_AGEMA_signal_4487, new_AGEMA_signal_4486, Midori_rounds_mul_ResultXORkey[38]}), .a ({new_AGEMA_signal_4353, new_AGEMA_signal_4352, new_AGEMA_signal_4351, Midori_rounds_SR_Inv_Result[38]}), .c ({new_AGEMA_signal_4692, new_AGEMA_signal_4691, new_AGEMA_signal_4690, Midori_rounds_round_Result[38]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_40_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_5052, new_AGEMA_signal_5051, new_AGEMA_signal_5050, Midori_rounds_mul_ResultXORkey[40]}), .a ({new_AGEMA_signal_5073, new_AGEMA_signal_5072, new_AGEMA_signal_5071, Midori_rounds_SR_Inv_Result[40]}), .c ({new_AGEMA_signal_5124, new_AGEMA_signal_5123, new_AGEMA_signal_5122, Midori_rounds_round_Result[40]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_42_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4476, new_AGEMA_signal_4475, new_AGEMA_signal_4474, Midori_rounds_mul_ResultXORkey[42]}), .a ({new_AGEMA_signal_4272, new_AGEMA_signal_4271, new_AGEMA_signal_4270, Midori_rounds_SR_Inv_Result[42]}), .c ({new_AGEMA_signal_4701, new_AGEMA_signal_4700, new_AGEMA_signal_4699, Midori_rounds_round_Result[42]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_44_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_5049, new_AGEMA_signal_5048, new_AGEMA_signal_5047, Midori_rounds_mul_ResultXORkey[44]}), .a ({new_AGEMA_signal_5007, new_AGEMA_signal_5006, new_AGEMA_signal_5005, Midori_rounds_SR_Inv_Result[44]}), .c ({new_AGEMA_signal_5127, new_AGEMA_signal_5126, new_AGEMA_signal_5125, Midori_rounds_round_Result[44]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_46_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4464, new_AGEMA_signal_4463, new_AGEMA_signal_4462, Midori_rounds_mul_ResultXORkey[46]}), .a ({new_AGEMA_signal_4335, new_AGEMA_signal_4334, new_AGEMA_signal_4333, Midori_rounds_SR_Inv_Result[46]}), .c ({new_AGEMA_signal_4710, new_AGEMA_signal_4709, new_AGEMA_signal_4708, Midori_rounds_round_Result[46]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_48_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_5046, new_AGEMA_signal_5045, new_AGEMA_signal_5044, Midori_rounds_mul_ResultXORkey[48]}), .a ({new_AGEMA_signal_5019, new_AGEMA_signal_5018, new_AGEMA_signal_5017, Midori_rounds_SR_Inv_Result[48]}), .c ({new_AGEMA_signal_5130, new_AGEMA_signal_5129, new_AGEMA_signal_5128, Midori_rounds_round_Result[48]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_50_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4455, new_AGEMA_signal_4454, new_AGEMA_signal_4453, Midori_rounds_mul_ResultXORkey[50]}), .a ({new_AGEMA_signal_4371, new_AGEMA_signal_4370, new_AGEMA_signal_4369, Midori_rounds_SR_Inv_Result[50]}), .c ({new_AGEMA_signal_4719, new_AGEMA_signal_4718, new_AGEMA_signal_4717, Midori_rounds_round_Result[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_52_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_5085, new_AGEMA_signal_5084, new_AGEMA_signal_5083, Midori_rounds_mul_ResultXORkey[52]}), .a ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, new_AGEMA_signal_5029, Midori_rounds_SR_Inv_Result[52]}), .c ({new_AGEMA_signal_5178, new_AGEMA_signal_5177, new_AGEMA_signal_5176, Midori_rounds_round_Result[52]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_54_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4446, new_AGEMA_signal_4445, new_AGEMA_signal_4444, Midori_rounds_mul_ResultXORkey[54]}), .a ({new_AGEMA_signal_4380, new_AGEMA_signal_4379, new_AGEMA_signal_4378, Midori_rounds_SR_Inv_Result[54]}), .c ({new_AGEMA_signal_4728, new_AGEMA_signal_4727, new_AGEMA_signal_4726, Midori_rounds_round_Result[54]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_56_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_5136, new_AGEMA_signal_5135, new_AGEMA_signal_5134, Midori_rounds_mul_ResultXORkey[56]}), .a ({new_AGEMA_signal_5016, new_AGEMA_signal_5015, new_AGEMA_signal_5014, Midori_rounds_SR_Inv_Result[56]}), .c ({new_AGEMA_signal_5190, new_AGEMA_signal_5189, new_AGEMA_signal_5188, Midori_rounds_round_Result[56]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_58_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4437, new_AGEMA_signal_4436, new_AGEMA_signal_4435, Midori_rounds_mul_ResultXORkey[58]}), .a ({new_AGEMA_signal_4317, new_AGEMA_signal_4316, new_AGEMA_signal_4315, Midori_rounds_SR_Inv_Result[58]}), .c ({new_AGEMA_signal_4737, new_AGEMA_signal_4736, new_AGEMA_signal_4735, Midori_rounds_round_Result[58]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_60_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_5133, new_AGEMA_signal_5132, new_AGEMA_signal_5131, Midori_rounds_mul_ResultXORkey[60]}), .a ({new_AGEMA_signal_5097, new_AGEMA_signal_5096, new_AGEMA_signal_5095, Midori_rounds_SR_Inv_Result[60]}), .c ({new_AGEMA_signal_5193, new_AGEMA_signal_5192, new_AGEMA_signal_5191, Midori_rounds_round_Result[60]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_62_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_4425, new_AGEMA_signal_4424, new_AGEMA_signal_4423, Midori_rounds_mul_ResultXORkey[62]}), .a ({new_AGEMA_signal_4290, new_AGEMA_signal_4289, new_AGEMA_signal_4288, Midori_rounds_SR_Inv_Result[62]}), .c ({new_AGEMA_signal_4746, new_AGEMA_signal_4745, new_AGEMA_signal_4744, Midori_rounds_round_Result[62]}) ) ;

    /* register cells */
    DFF_X1 controller_roundCounter_count_reg_0__FF_FF ( .CK (clk_gated), .D (controller_roundCounter_N7), .Q (round_Signal[0]), .QN () ) ;
    DFF_X1 controller_roundCounter_count_reg_1__FF_FF ( .CK (clk_gated), .D (controller_roundCounter_N8), .Q (round_Signal[1]), .QN () ) ;
    DFF_X1 controller_roundCounter_count_reg_2__FF_FF ( .CK (clk_gated), .D (controller_roundCounter_n2), .Q (round_Signal[2]), .QN () ) ;
    DFF_X1 controller_roundCounter_count_reg_3__FF_FF ( .CK (clk_gated), .D (controller_roundCounter_N10), .Q (round_Signal[3]), .QN () ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5139, new_AGEMA_signal_5138, new_AGEMA_signal_5137, Midori_rounds_roundResult_Reg_SFF_0_DQ}), .Q ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, new_AGEMA_signal_2071, Midori_rounds_roundReg_out[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4785, new_AGEMA_signal_4784, new_AGEMA_signal_4783, Midori_rounds_roundResult_Reg_SFF_1_DQ}), .Q ({new_AGEMA_signal_3282, new_AGEMA_signal_3281, new_AGEMA_signal_3280, Midori_rounds_roundReg_out[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4788, new_AGEMA_signal_4787, new_AGEMA_signal_4786, Midori_rounds_roundResult_Reg_SFF_2_DQ}), .Q ({new_AGEMA_signal_2082, new_AGEMA_signal_2081, new_AGEMA_signal_2080, Midori_rounds_roundReg_out[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4791, new_AGEMA_signal_4790, new_AGEMA_signal_4789, Midori_rounds_roundResult_Reg_SFF_3_DQ}), .Q ({new_AGEMA_signal_2076, new_AGEMA_signal_2075, new_AGEMA_signal_2074, Midori_rounds_roundReg_out[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5142, new_AGEMA_signal_5141, new_AGEMA_signal_5140, Midori_rounds_roundResult_Reg_SFF_4_DQ}), .Q ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, new_AGEMA_signal_2095, Midori_rounds_roundReg_out[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4794, new_AGEMA_signal_4793, new_AGEMA_signal_4792, Midori_rounds_roundResult_Reg_SFF_5_DQ}), .Q ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, new_AGEMA_signal_3295, Midori_rounds_roundReg_out[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4797, new_AGEMA_signal_4796, new_AGEMA_signal_4795, Midori_rounds_roundResult_Reg_SFF_6_DQ}), .Q ({new_AGEMA_signal_2106, new_AGEMA_signal_2105, new_AGEMA_signal_2104, Midori_rounds_roundReg_out[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4800, new_AGEMA_signal_4799, new_AGEMA_signal_4798, Midori_rounds_roundResult_Reg_SFF_7_DQ}), .Q ({new_AGEMA_signal_2100, new_AGEMA_signal_2099, new_AGEMA_signal_2098, Midori_rounds_roundReg_out[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_8_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5145, new_AGEMA_signal_5144, new_AGEMA_signal_5143, Midori_rounds_roundResult_Reg_SFF_8_DQ}), .Q ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, new_AGEMA_signal_2119, Midori_rounds_roundReg_out[8]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_9_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4803, new_AGEMA_signal_4802, new_AGEMA_signal_4801, Midori_rounds_roundResult_Reg_SFF_9_DQ}), .Q ({new_AGEMA_signal_3312, new_AGEMA_signal_3311, new_AGEMA_signal_3310, Midori_rounds_roundReg_out[9]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_10_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4806, new_AGEMA_signal_4805, new_AGEMA_signal_4804, Midori_rounds_roundResult_Reg_SFF_10_DQ}), .Q ({new_AGEMA_signal_2130, new_AGEMA_signal_2129, new_AGEMA_signal_2128, Midori_rounds_roundReg_out[10]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_11_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4809, new_AGEMA_signal_4808, new_AGEMA_signal_4807, Midori_rounds_roundResult_Reg_SFF_11_DQ}), .Q ({new_AGEMA_signal_2124, new_AGEMA_signal_2123, new_AGEMA_signal_2122, Midori_rounds_roundReg_out[11]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_12_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5148, new_AGEMA_signal_5147, new_AGEMA_signal_5146, Midori_rounds_roundResult_Reg_SFF_12_DQ}), .Q ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, new_AGEMA_signal_2143, Midori_rounds_roundReg_out[12]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_13_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4812, new_AGEMA_signal_4811, new_AGEMA_signal_4810, Midori_rounds_roundResult_Reg_SFF_13_DQ}), .Q ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, new_AGEMA_signal_3325, Midori_rounds_roundReg_out[13]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_14_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4815, new_AGEMA_signal_4814, new_AGEMA_signal_4813, Midori_rounds_roundResult_Reg_SFF_14_DQ}), .Q ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, new_AGEMA_signal_2152, Midori_rounds_roundReg_out[14]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_15_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4818, new_AGEMA_signal_4817, new_AGEMA_signal_4816, Midori_rounds_roundResult_Reg_SFF_15_DQ}), .Q ({new_AGEMA_signal_2148, new_AGEMA_signal_2147, new_AGEMA_signal_2146, Midori_rounds_roundReg_out[15]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_16_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5181, new_AGEMA_signal_5180, new_AGEMA_signal_5179, Midori_rounds_roundResult_Reg_SFF_16_DQ}), .Q ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, new_AGEMA_signal_2167, Midori_rounds_roundReg_out[16]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_17_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4821, new_AGEMA_signal_4820, new_AGEMA_signal_4819, Midori_rounds_roundResult_Reg_SFF_17_DQ}), .Q ({new_AGEMA_signal_3342, new_AGEMA_signal_3341, new_AGEMA_signal_3340, Midori_rounds_roundReg_out[17]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_18_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4824, new_AGEMA_signal_4823, new_AGEMA_signal_4822, Midori_rounds_roundResult_Reg_SFF_18_DQ}), .Q ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, new_AGEMA_signal_2176, Midori_rounds_roundReg_out[18]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_19_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4827, new_AGEMA_signal_4826, new_AGEMA_signal_4825, Midori_rounds_roundResult_Reg_SFF_19_DQ}), .Q ({new_AGEMA_signal_2172, new_AGEMA_signal_2171, new_AGEMA_signal_2170, Midori_rounds_roundReg_out[19]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_20_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5184, new_AGEMA_signal_5183, new_AGEMA_signal_5182, Midori_rounds_roundResult_Reg_SFF_20_DQ}), .Q ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, new_AGEMA_signal_2191, Midori_rounds_roundReg_out[20]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_21_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4830, new_AGEMA_signal_4829, new_AGEMA_signal_4828, Midori_rounds_roundResult_Reg_SFF_21_DQ}), .Q ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, new_AGEMA_signal_3355, Midori_rounds_roundReg_out[21]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_22_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, new_AGEMA_signal_4831, Midori_rounds_roundResult_Reg_SFF_22_DQ}), .Q ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, new_AGEMA_signal_2200, Midori_rounds_roundReg_out[22]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_23_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4836, new_AGEMA_signal_4835, new_AGEMA_signal_4834, Midori_rounds_roundResult_Reg_SFF_23_DQ}), .Q ({new_AGEMA_signal_2196, new_AGEMA_signal_2195, new_AGEMA_signal_2194, Midori_rounds_roundReg_out[23]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_24_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5151, new_AGEMA_signal_5150, new_AGEMA_signal_5149, Midori_rounds_roundResult_Reg_SFF_24_DQ}), .Q ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, new_AGEMA_signal_2215, Midori_rounds_roundReg_out[24]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_25_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4839, new_AGEMA_signal_4838, new_AGEMA_signal_4837, Midori_rounds_roundResult_Reg_SFF_25_DQ}), .Q ({new_AGEMA_signal_3372, new_AGEMA_signal_3371, new_AGEMA_signal_3370, Midori_rounds_roundReg_out[25]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_26_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4842, new_AGEMA_signal_4841, new_AGEMA_signal_4840, Midori_rounds_roundResult_Reg_SFF_26_DQ}), .Q ({new_AGEMA_signal_2226, new_AGEMA_signal_2225, new_AGEMA_signal_2224, Midori_rounds_roundReg_out[26]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_27_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4845, new_AGEMA_signal_4844, new_AGEMA_signal_4843, Midori_rounds_roundResult_Reg_SFF_27_DQ}), .Q ({new_AGEMA_signal_2220, new_AGEMA_signal_2219, new_AGEMA_signal_2218, Midori_rounds_roundReg_out[27]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_28_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5154, new_AGEMA_signal_5153, new_AGEMA_signal_5152, Midori_rounds_roundResult_Reg_SFF_28_DQ}), .Q ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, new_AGEMA_signal_2239, Midori_rounds_roundReg_out[28]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_29_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4848, new_AGEMA_signal_4847, new_AGEMA_signal_4846, Midori_rounds_roundResult_Reg_SFF_29_DQ}), .Q ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, new_AGEMA_signal_3385, Midori_rounds_roundReg_out[29]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_30_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, new_AGEMA_signal_4849, Midori_rounds_roundResult_Reg_SFF_30_DQ}), .Q ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, new_AGEMA_signal_2248, Midori_rounds_roundReg_out[30]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_31_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4854, new_AGEMA_signal_4853, new_AGEMA_signal_4852, Midori_rounds_roundResult_Reg_SFF_31_DQ}), .Q ({new_AGEMA_signal_2244, new_AGEMA_signal_2243, new_AGEMA_signal_2242, Midori_rounds_roundReg_out[31]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_32_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5157, new_AGEMA_signal_5156, new_AGEMA_signal_5155, Midori_rounds_roundResult_Reg_SFF_32_DQ}), .Q ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, new_AGEMA_signal_2263, Midori_rounds_roundReg_out[32]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_33_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4857, new_AGEMA_signal_4856, new_AGEMA_signal_4855, Midori_rounds_roundResult_Reg_SFF_33_DQ}), .Q ({new_AGEMA_signal_3402, new_AGEMA_signal_3401, new_AGEMA_signal_3400, Midori_rounds_roundReg_out[33]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_34_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4860, new_AGEMA_signal_4859, new_AGEMA_signal_4858, Midori_rounds_roundResult_Reg_SFF_34_DQ}), .Q ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, new_AGEMA_signal_2272, Midori_rounds_roundReg_out[34]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_35_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4863, new_AGEMA_signal_4862, new_AGEMA_signal_4861, Midori_rounds_roundResult_Reg_SFF_35_DQ}), .Q ({new_AGEMA_signal_2268, new_AGEMA_signal_2267, new_AGEMA_signal_2266, Midori_rounds_roundReg_out[35]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_36_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5160, new_AGEMA_signal_5159, new_AGEMA_signal_5158, Midori_rounds_roundResult_Reg_SFF_36_DQ}), .Q ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, new_AGEMA_signal_2287, Midori_rounds_roundReg_out[36]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_37_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4866, new_AGEMA_signal_4865, new_AGEMA_signal_4864, Midori_rounds_roundResult_Reg_SFF_37_DQ}), .Q ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, new_AGEMA_signal_3415, Midori_rounds_roundReg_out[37]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_38_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, Midori_rounds_roundResult_Reg_SFF_38_DQ}), .Q ({new_AGEMA_signal_2298, new_AGEMA_signal_2297, new_AGEMA_signal_2296, Midori_rounds_roundReg_out[38]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_39_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4872, new_AGEMA_signal_4871, new_AGEMA_signal_4870, Midori_rounds_roundResult_Reg_SFF_39_DQ}), .Q ({new_AGEMA_signal_2292, new_AGEMA_signal_2291, new_AGEMA_signal_2290, Midori_rounds_roundReg_out[39]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_40_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5163, new_AGEMA_signal_5162, new_AGEMA_signal_5161, Midori_rounds_roundResult_Reg_SFF_40_DQ}), .Q ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, new_AGEMA_signal_2311, Midori_rounds_roundReg_out[40]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_41_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4875, new_AGEMA_signal_4874, new_AGEMA_signal_4873, Midori_rounds_roundResult_Reg_SFF_41_DQ}), .Q ({new_AGEMA_signal_3432, new_AGEMA_signal_3431, new_AGEMA_signal_3430, Midori_rounds_roundReg_out[41]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_42_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4878, new_AGEMA_signal_4877, new_AGEMA_signal_4876, Midori_rounds_roundResult_Reg_SFF_42_DQ}), .Q ({new_AGEMA_signal_2322, new_AGEMA_signal_2321, new_AGEMA_signal_2320, Midori_rounds_roundReg_out[42]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_43_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4881, new_AGEMA_signal_4880, new_AGEMA_signal_4879, Midori_rounds_roundResult_Reg_SFF_43_DQ}), .Q ({new_AGEMA_signal_2316, new_AGEMA_signal_2315, new_AGEMA_signal_2314, Midori_rounds_roundReg_out[43]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_44_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5166, new_AGEMA_signal_5165, new_AGEMA_signal_5164, Midori_rounds_roundResult_Reg_SFF_44_DQ}), .Q ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, new_AGEMA_signal_2335, Midori_rounds_roundReg_out[44]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_45_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4884, new_AGEMA_signal_4883, new_AGEMA_signal_4882, Midori_rounds_roundResult_Reg_SFF_45_DQ}), .Q ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, new_AGEMA_signal_3445, Midori_rounds_roundReg_out[45]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_46_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, new_AGEMA_signal_4885, Midori_rounds_roundResult_Reg_SFF_46_DQ}), .Q ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, new_AGEMA_signal_2344, Midori_rounds_roundReg_out[46]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_47_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4890, new_AGEMA_signal_4889, new_AGEMA_signal_4888, Midori_rounds_roundResult_Reg_SFF_47_DQ}), .Q ({new_AGEMA_signal_2340, new_AGEMA_signal_2339, new_AGEMA_signal_2338, Midori_rounds_roundReg_out[47]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_48_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5169, new_AGEMA_signal_5168, new_AGEMA_signal_5167, Midori_rounds_roundResult_Reg_SFF_48_DQ}), .Q ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, new_AGEMA_signal_2359, Midori_rounds_roundReg_out[48]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_49_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4893, new_AGEMA_signal_4892, new_AGEMA_signal_4891, Midori_rounds_roundResult_Reg_SFF_49_DQ}), .Q ({new_AGEMA_signal_3462, new_AGEMA_signal_3461, new_AGEMA_signal_3460, Midori_rounds_roundReg_out[49]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_50_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4896, new_AGEMA_signal_4895, new_AGEMA_signal_4894, Midori_rounds_roundResult_Reg_SFF_50_DQ}), .Q ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, new_AGEMA_signal_2368, Midori_rounds_roundReg_out[50]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_51_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4899, new_AGEMA_signal_4898, new_AGEMA_signal_4897, Midori_rounds_roundResult_Reg_SFF_51_DQ}), .Q ({new_AGEMA_signal_2364, new_AGEMA_signal_2363, new_AGEMA_signal_2362, Midori_rounds_roundReg_out[51]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_52_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5187, new_AGEMA_signal_5186, new_AGEMA_signal_5185, Midori_rounds_roundResult_Reg_SFF_52_DQ}), .Q ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, new_AGEMA_signal_2383, Midori_rounds_roundReg_out[52]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_53_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4902, new_AGEMA_signal_4901, new_AGEMA_signal_4900, Midori_rounds_roundResult_Reg_SFF_53_DQ}), .Q ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, new_AGEMA_signal_3475, Midori_rounds_roundReg_out[53]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_54_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, new_AGEMA_signal_4903, Midori_rounds_roundResult_Reg_SFF_54_DQ}), .Q ({new_AGEMA_signal_2394, new_AGEMA_signal_2393, new_AGEMA_signal_2392, Midori_rounds_roundReg_out[54]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_55_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4908, new_AGEMA_signal_4907, new_AGEMA_signal_4906, Midori_rounds_roundResult_Reg_SFF_55_DQ}), .Q ({new_AGEMA_signal_2388, new_AGEMA_signal_2387, new_AGEMA_signal_2386, Midori_rounds_roundReg_out[55]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_56_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5196, new_AGEMA_signal_5195, new_AGEMA_signal_5194, Midori_rounds_roundResult_Reg_SFF_56_DQ}), .Q ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, new_AGEMA_signal_2407, Midori_rounds_roundReg_out[56]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_57_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4911, new_AGEMA_signal_4910, new_AGEMA_signal_4909, Midori_rounds_roundResult_Reg_SFF_57_DQ}), .Q ({new_AGEMA_signal_3492, new_AGEMA_signal_3491, new_AGEMA_signal_3490, Midori_rounds_roundReg_out[57]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_58_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4914, new_AGEMA_signal_4913, new_AGEMA_signal_4912, Midori_rounds_roundResult_Reg_SFF_58_DQ}), .Q ({new_AGEMA_signal_2418, new_AGEMA_signal_2417, new_AGEMA_signal_2416, Midori_rounds_roundReg_out[58]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_59_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4917, new_AGEMA_signal_4916, new_AGEMA_signal_4915, Midori_rounds_roundResult_Reg_SFF_59_DQ}), .Q ({new_AGEMA_signal_2412, new_AGEMA_signal_2411, new_AGEMA_signal_2410, Midori_rounds_roundReg_out[59]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_60_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_5199, new_AGEMA_signal_5198, new_AGEMA_signal_5197, Midori_rounds_roundResult_Reg_SFF_60_DQ}), .Q ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, new_AGEMA_signal_2431, Midori_rounds_roundReg_out[60]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_61_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4920, new_AGEMA_signal_4919, new_AGEMA_signal_4918, Midori_rounds_roundResult_Reg_SFF_61_DQ}), .Q ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, new_AGEMA_signal_3505, Midori_rounds_roundReg_out[61]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_62_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, new_AGEMA_signal_4921, Midori_rounds_roundResult_Reg_SFF_62_DQ}), .Q ({new_AGEMA_signal_2442, new_AGEMA_signal_2441, new_AGEMA_signal_2440, Midori_rounds_roundReg_out[62]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_63_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4926, new_AGEMA_signal_4925, new_AGEMA_signal_4924, Midori_rounds_roundResult_Reg_SFF_63_DQ}), .Q ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, new_AGEMA_signal_2434, Midori_rounds_roundReg_out[63]}) ) ;
endmodule
