////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module CRAFT in file /AGEMA/Designs/CRAFT_round-based/AGEMA/CRAFT.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module CRAFT_HPC2_ClockGating_d2 (plaintext_s0, key_s0, clk, rst, key_s1, key_s2, plaintext_s1, plaintext_s2, Fresh, ciphertext_s0, done, ciphertext_s1, ciphertext_s2, Synch);
    input [63:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input rst ;
    input [127:0] key_s1 ;
    input [127:0] key_s2 ;
    input [63:0] plaintext_s1 ;
    input [63:0] plaintext_s2 ;
    input [767:0] Fresh ;
    output [63:0] ciphertext_s0 ;
    output done ;
    output [63:0] ciphertext_s1 ;
    output [63:0] ciphertext_s2 ;
    output Synch ;
    wire RoundConstant_4_ ;
    wire RoundConstant_0 ;
    wire done_internal ;
    wire MCInst_XOR_r0_Inst_0_n2 ;
    wire MCInst_XOR_r0_Inst_0_n1 ;
    wire MCInst_XOR_r1_Inst_0_n1 ;
    wire MCInst_XOR_r0_Inst_1_n2 ;
    wire MCInst_XOR_r0_Inst_1_n1 ;
    wire MCInst_XOR_r1_Inst_1_n1 ;
    wire MCInst_XOR_r0_Inst_2_n2 ;
    wire MCInst_XOR_r0_Inst_2_n1 ;
    wire MCInst_XOR_r1_Inst_2_n1 ;
    wire MCInst_XOR_r0_Inst_3_n2 ;
    wire MCInst_XOR_r0_Inst_3_n1 ;
    wire MCInst_XOR_r1_Inst_3_n1 ;
    wire MCInst_XOR_r0_Inst_4_n2 ;
    wire MCInst_XOR_r0_Inst_4_n1 ;
    wire MCInst_XOR_r1_Inst_4_n1 ;
    wire MCInst_XOR_r0_Inst_5_n2 ;
    wire MCInst_XOR_r0_Inst_5_n1 ;
    wire MCInst_XOR_r1_Inst_5_n1 ;
    wire MCInst_XOR_r0_Inst_6_n2 ;
    wire MCInst_XOR_r0_Inst_6_n1 ;
    wire MCInst_XOR_r1_Inst_6_n1 ;
    wire MCInst_XOR_r0_Inst_7_n2 ;
    wire MCInst_XOR_r0_Inst_7_n1 ;
    wire MCInst_XOR_r1_Inst_7_n1 ;
    wire MCInst_XOR_r0_Inst_8_n2 ;
    wire MCInst_XOR_r0_Inst_8_n1 ;
    wire MCInst_XOR_r1_Inst_8_n1 ;
    wire MCInst_XOR_r0_Inst_9_n2 ;
    wire MCInst_XOR_r0_Inst_9_n1 ;
    wire MCInst_XOR_r1_Inst_9_n1 ;
    wire MCInst_XOR_r0_Inst_10_n2 ;
    wire MCInst_XOR_r0_Inst_10_n1 ;
    wire MCInst_XOR_r1_Inst_10_n1 ;
    wire MCInst_XOR_r0_Inst_11_n2 ;
    wire MCInst_XOR_r0_Inst_11_n1 ;
    wire MCInst_XOR_r1_Inst_11_n1 ;
    wire MCInst_XOR_r0_Inst_12_n2 ;
    wire MCInst_XOR_r0_Inst_12_n1 ;
    wire MCInst_XOR_r1_Inst_12_n1 ;
    wire MCInst_XOR_r0_Inst_13_n2 ;
    wire MCInst_XOR_r0_Inst_13_n1 ;
    wire MCInst_XOR_r1_Inst_13_n1 ;
    wire MCInst_XOR_r0_Inst_14_n2 ;
    wire MCInst_XOR_r0_Inst_14_n1 ;
    wire MCInst_XOR_r1_Inst_14_n1 ;
    wire MCInst_XOR_r0_Inst_15_n2 ;
    wire MCInst_XOR_r0_Inst_15_n1 ;
    wire MCInst_XOR_r1_Inst_15_n1 ;
    wire AddKeyXOR1_XORInst_0_0_n1 ;
    wire AddKeyXOR1_XORInst_0_1_n1 ;
    wire AddKeyXOR1_XORInst_0_2_n1 ;
    wire AddKeyXOR1_XORInst_0_3_n1 ;
    wire AddKeyXOR1_XORInst_1_0_n1 ;
    wire AddKeyXOR1_XORInst_1_1_n1 ;
    wire AddKeyXOR1_XORInst_1_2_n1 ;
    wire AddKeyXOR1_XORInst_1_3_n1 ;
    wire AddKeyXOR1_XORInst_2_0_n1 ;
    wire AddKeyXOR1_XORInst_2_1_n1 ;
    wire AddKeyXOR1_XORInst_2_2_n1 ;
    wire AddKeyXOR1_XORInst_2_3_n1 ;
    wire AddKeyXOR1_XORInst_3_0_n1 ;
    wire AddKeyXOR1_XORInst_3_1_n1 ;
    wire AddKeyXOR1_XORInst_3_2_n1 ;
    wire AddKeyXOR1_XORInst_3_3_n1 ;
    wire AddKeyConstXOR_XORInst_0_0_n2 ;
    wire AddKeyConstXOR_XORInst_0_0_n1 ;
    wire AddKeyConstXOR_XORInst_0_1_n2 ;
    wire AddKeyConstXOR_XORInst_0_1_n1 ;
    wire AddKeyConstXOR_XORInst_0_2_n2 ;
    wire AddKeyConstXOR_XORInst_0_2_n1 ;
    wire AddKeyConstXOR_XORInst_0_3_n2 ;
    wire AddKeyConstXOR_XORInst_0_3_n1 ;
    wire AddKeyConstXOR_XORInst_1_0_n2 ;
    wire AddKeyConstXOR_XORInst_1_0_n1 ;
    wire AddKeyConstXOR_XORInst_1_1_n2 ;
    wire AddKeyConstXOR_XORInst_1_1_n1 ;
    wire AddKeyConstXOR_XORInst_1_2_n2 ;
    wire AddKeyConstXOR_XORInst_1_2_n1 ;
    wire AddKeyConstXOR_XORInst_1_3_n2 ;
    wire AddKeyConstXOR_XORInst_1_3_n1 ;
    wire AddKeyXOR2_XORInst_0_0_n1 ;
    wire AddKeyXOR2_XORInst_0_1_n1 ;
    wire AddKeyXOR2_XORInst_0_2_n1 ;
    wire AddKeyXOR2_XORInst_0_3_n1 ;
    wire AddKeyXOR2_XORInst_1_0_n1 ;
    wire AddKeyXOR2_XORInst_1_1_n1 ;
    wire AddKeyXOR2_XORInst_1_2_n1 ;
    wire AddKeyXOR2_XORInst_1_3_n1 ;
    wire AddKeyXOR2_XORInst_2_0_n1 ;
    wire AddKeyXOR2_XORInst_2_1_n1 ;
    wire AddKeyXOR2_XORInst_2_2_n1 ;
    wire AddKeyXOR2_XORInst_2_3_n1 ;
    wire AddKeyXOR2_XORInst_3_0_n1 ;
    wire AddKeyXOR2_XORInst_3_1_n1 ;
    wire AddKeyXOR2_XORInst_3_2_n1 ;
    wire AddKeyXOR2_XORInst_3_3_n1 ;
    wire AddKeyXOR2_XORInst_4_0_n1 ;
    wire AddKeyXOR2_XORInst_4_1_n1 ;
    wire AddKeyXOR2_XORInst_4_2_n1 ;
    wire AddKeyXOR2_XORInst_4_3_n1 ;
    wire AddKeyXOR2_XORInst_5_0_n1 ;
    wire AddKeyXOR2_XORInst_5_1_n1 ;
    wire AddKeyXOR2_XORInst_5_2_n1 ;
    wire AddKeyXOR2_XORInst_5_3_n1 ;
    wire AddKeyXOR2_XORInst_6_0_n1 ;
    wire AddKeyXOR2_XORInst_6_1_n1 ;
    wire AddKeyXOR2_XORInst_6_2_n1 ;
    wire AddKeyXOR2_XORInst_6_3_n1 ;
    wire AddKeyXOR2_XORInst_7_0_n1 ;
    wire AddKeyXOR2_XORInst_7_1_n1 ;
    wire AddKeyXOR2_XORInst_7_2_n1 ;
    wire AddKeyXOR2_XORInst_7_3_n1 ;
    wire AddKeyXOR2_XORInst_8_0_n1 ;
    wire AddKeyXOR2_XORInst_8_1_n1 ;
    wire AddKeyXOR2_XORInst_8_2_n1 ;
    wire AddKeyXOR2_XORInst_8_3_n1 ;
    wire AddKeyXOR2_XORInst_9_0_n1 ;
    wire AddKeyXOR2_XORInst_9_1_n1 ;
    wire AddKeyXOR2_XORInst_9_2_n1 ;
    wire AddKeyXOR2_XORInst_9_3_n1 ;
    wire SubCellInst_SboxInst_0_n15 ;
    wire SubCellInst_SboxInst_0_n14 ;
    wire SubCellInst_SboxInst_0_n13 ;
    wire SubCellInst_SboxInst_0_n12 ;
    wire SubCellInst_SboxInst_0_n11 ;
    wire SubCellInst_SboxInst_0_n10 ;
    wire SubCellInst_SboxInst_0_n9 ;
    wire SubCellInst_SboxInst_0_n8 ;
    wire SubCellInst_SboxInst_0_n7 ;
    wire SubCellInst_SboxInst_0_n6 ;
    wire SubCellInst_SboxInst_0_n5 ;
    wire SubCellInst_SboxInst_0_n4 ;
    wire SubCellInst_SboxInst_0_n3 ;
    wire SubCellInst_SboxInst_0_n2 ;
    wire SubCellInst_SboxInst_0_n1 ;
    wire SubCellInst_SboxInst_1_n15 ;
    wire SubCellInst_SboxInst_1_n14 ;
    wire SubCellInst_SboxInst_1_n13 ;
    wire SubCellInst_SboxInst_1_n12 ;
    wire SubCellInst_SboxInst_1_n11 ;
    wire SubCellInst_SboxInst_1_n10 ;
    wire SubCellInst_SboxInst_1_n9 ;
    wire SubCellInst_SboxInst_1_n8 ;
    wire SubCellInst_SboxInst_1_n7 ;
    wire SubCellInst_SboxInst_1_n6 ;
    wire SubCellInst_SboxInst_1_n5 ;
    wire SubCellInst_SboxInst_1_n4 ;
    wire SubCellInst_SboxInst_1_n3 ;
    wire SubCellInst_SboxInst_1_n2 ;
    wire SubCellInst_SboxInst_1_n1 ;
    wire SubCellInst_SboxInst_2_n15 ;
    wire SubCellInst_SboxInst_2_n14 ;
    wire SubCellInst_SboxInst_2_n13 ;
    wire SubCellInst_SboxInst_2_n12 ;
    wire SubCellInst_SboxInst_2_n11 ;
    wire SubCellInst_SboxInst_2_n10 ;
    wire SubCellInst_SboxInst_2_n9 ;
    wire SubCellInst_SboxInst_2_n8 ;
    wire SubCellInst_SboxInst_2_n7 ;
    wire SubCellInst_SboxInst_2_n6 ;
    wire SubCellInst_SboxInst_2_n5 ;
    wire SubCellInst_SboxInst_2_n4 ;
    wire SubCellInst_SboxInst_2_n3 ;
    wire SubCellInst_SboxInst_2_n2 ;
    wire SubCellInst_SboxInst_2_n1 ;
    wire SubCellInst_SboxInst_3_n15 ;
    wire SubCellInst_SboxInst_3_n14 ;
    wire SubCellInst_SboxInst_3_n13 ;
    wire SubCellInst_SboxInst_3_n12 ;
    wire SubCellInst_SboxInst_3_n11 ;
    wire SubCellInst_SboxInst_3_n10 ;
    wire SubCellInst_SboxInst_3_n9 ;
    wire SubCellInst_SboxInst_3_n8 ;
    wire SubCellInst_SboxInst_3_n7 ;
    wire SubCellInst_SboxInst_3_n6 ;
    wire SubCellInst_SboxInst_3_n5 ;
    wire SubCellInst_SboxInst_3_n4 ;
    wire SubCellInst_SboxInst_3_n3 ;
    wire SubCellInst_SboxInst_3_n2 ;
    wire SubCellInst_SboxInst_3_n1 ;
    wire SubCellInst_SboxInst_4_n15 ;
    wire SubCellInst_SboxInst_4_n14 ;
    wire SubCellInst_SboxInst_4_n13 ;
    wire SubCellInst_SboxInst_4_n12 ;
    wire SubCellInst_SboxInst_4_n11 ;
    wire SubCellInst_SboxInst_4_n10 ;
    wire SubCellInst_SboxInst_4_n9 ;
    wire SubCellInst_SboxInst_4_n8 ;
    wire SubCellInst_SboxInst_4_n7 ;
    wire SubCellInst_SboxInst_4_n6 ;
    wire SubCellInst_SboxInst_4_n5 ;
    wire SubCellInst_SboxInst_4_n4 ;
    wire SubCellInst_SboxInst_4_n3 ;
    wire SubCellInst_SboxInst_4_n2 ;
    wire SubCellInst_SboxInst_4_n1 ;
    wire SubCellInst_SboxInst_5_n15 ;
    wire SubCellInst_SboxInst_5_n14 ;
    wire SubCellInst_SboxInst_5_n13 ;
    wire SubCellInst_SboxInst_5_n12 ;
    wire SubCellInst_SboxInst_5_n11 ;
    wire SubCellInst_SboxInst_5_n10 ;
    wire SubCellInst_SboxInst_5_n9 ;
    wire SubCellInst_SboxInst_5_n8 ;
    wire SubCellInst_SboxInst_5_n7 ;
    wire SubCellInst_SboxInst_5_n6 ;
    wire SubCellInst_SboxInst_5_n5 ;
    wire SubCellInst_SboxInst_5_n4 ;
    wire SubCellInst_SboxInst_5_n3 ;
    wire SubCellInst_SboxInst_5_n2 ;
    wire SubCellInst_SboxInst_5_n1 ;
    wire SubCellInst_SboxInst_6_n15 ;
    wire SubCellInst_SboxInst_6_n14 ;
    wire SubCellInst_SboxInst_6_n13 ;
    wire SubCellInst_SboxInst_6_n12 ;
    wire SubCellInst_SboxInst_6_n11 ;
    wire SubCellInst_SboxInst_6_n10 ;
    wire SubCellInst_SboxInst_6_n9 ;
    wire SubCellInst_SboxInst_6_n8 ;
    wire SubCellInst_SboxInst_6_n7 ;
    wire SubCellInst_SboxInst_6_n6 ;
    wire SubCellInst_SboxInst_6_n5 ;
    wire SubCellInst_SboxInst_6_n4 ;
    wire SubCellInst_SboxInst_6_n3 ;
    wire SubCellInst_SboxInst_6_n2 ;
    wire SubCellInst_SboxInst_6_n1 ;
    wire SubCellInst_SboxInst_7_n15 ;
    wire SubCellInst_SboxInst_7_n14 ;
    wire SubCellInst_SboxInst_7_n13 ;
    wire SubCellInst_SboxInst_7_n12 ;
    wire SubCellInst_SboxInst_7_n11 ;
    wire SubCellInst_SboxInst_7_n10 ;
    wire SubCellInst_SboxInst_7_n9 ;
    wire SubCellInst_SboxInst_7_n8 ;
    wire SubCellInst_SboxInst_7_n7 ;
    wire SubCellInst_SboxInst_7_n6 ;
    wire SubCellInst_SboxInst_7_n5 ;
    wire SubCellInst_SboxInst_7_n4 ;
    wire SubCellInst_SboxInst_7_n3 ;
    wire SubCellInst_SboxInst_7_n2 ;
    wire SubCellInst_SboxInst_7_n1 ;
    wire SubCellInst_SboxInst_8_n15 ;
    wire SubCellInst_SboxInst_8_n14 ;
    wire SubCellInst_SboxInst_8_n13 ;
    wire SubCellInst_SboxInst_8_n12 ;
    wire SubCellInst_SboxInst_8_n11 ;
    wire SubCellInst_SboxInst_8_n10 ;
    wire SubCellInst_SboxInst_8_n9 ;
    wire SubCellInst_SboxInst_8_n8 ;
    wire SubCellInst_SboxInst_8_n7 ;
    wire SubCellInst_SboxInst_8_n6 ;
    wire SubCellInst_SboxInst_8_n5 ;
    wire SubCellInst_SboxInst_8_n4 ;
    wire SubCellInst_SboxInst_8_n3 ;
    wire SubCellInst_SboxInst_8_n2 ;
    wire SubCellInst_SboxInst_8_n1 ;
    wire SubCellInst_SboxInst_9_n15 ;
    wire SubCellInst_SboxInst_9_n14 ;
    wire SubCellInst_SboxInst_9_n13 ;
    wire SubCellInst_SboxInst_9_n12 ;
    wire SubCellInst_SboxInst_9_n11 ;
    wire SubCellInst_SboxInst_9_n10 ;
    wire SubCellInst_SboxInst_9_n9 ;
    wire SubCellInst_SboxInst_9_n8 ;
    wire SubCellInst_SboxInst_9_n7 ;
    wire SubCellInst_SboxInst_9_n6 ;
    wire SubCellInst_SboxInst_9_n5 ;
    wire SubCellInst_SboxInst_9_n4 ;
    wire SubCellInst_SboxInst_9_n3 ;
    wire SubCellInst_SboxInst_9_n2 ;
    wire SubCellInst_SboxInst_9_n1 ;
    wire SubCellInst_SboxInst_10_n15 ;
    wire SubCellInst_SboxInst_10_n14 ;
    wire SubCellInst_SboxInst_10_n13 ;
    wire SubCellInst_SboxInst_10_n12 ;
    wire SubCellInst_SboxInst_10_n11 ;
    wire SubCellInst_SboxInst_10_n10 ;
    wire SubCellInst_SboxInst_10_n9 ;
    wire SubCellInst_SboxInst_10_n8 ;
    wire SubCellInst_SboxInst_10_n7 ;
    wire SubCellInst_SboxInst_10_n6 ;
    wire SubCellInst_SboxInst_10_n5 ;
    wire SubCellInst_SboxInst_10_n4 ;
    wire SubCellInst_SboxInst_10_n3 ;
    wire SubCellInst_SboxInst_10_n2 ;
    wire SubCellInst_SboxInst_10_n1 ;
    wire SubCellInst_SboxInst_11_n15 ;
    wire SubCellInst_SboxInst_11_n14 ;
    wire SubCellInst_SboxInst_11_n13 ;
    wire SubCellInst_SboxInst_11_n12 ;
    wire SubCellInst_SboxInst_11_n11 ;
    wire SubCellInst_SboxInst_11_n10 ;
    wire SubCellInst_SboxInst_11_n9 ;
    wire SubCellInst_SboxInst_11_n8 ;
    wire SubCellInst_SboxInst_11_n7 ;
    wire SubCellInst_SboxInst_11_n6 ;
    wire SubCellInst_SboxInst_11_n5 ;
    wire SubCellInst_SboxInst_11_n4 ;
    wire SubCellInst_SboxInst_11_n3 ;
    wire SubCellInst_SboxInst_11_n2 ;
    wire SubCellInst_SboxInst_11_n1 ;
    wire SubCellInst_SboxInst_12_n15 ;
    wire SubCellInst_SboxInst_12_n14 ;
    wire SubCellInst_SboxInst_12_n13 ;
    wire SubCellInst_SboxInst_12_n12 ;
    wire SubCellInst_SboxInst_12_n11 ;
    wire SubCellInst_SboxInst_12_n10 ;
    wire SubCellInst_SboxInst_12_n9 ;
    wire SubCellInst_SboxInst_12_n8 ;
    wire SubCellInst_SboxInst_12_n7 ;
    wire SubCellInst_SboxInst_12_n6 ;
    wire SubCellInst_SboxInst_12_n5 ;
    wire SubCellInst_SboxInst_12_n4 ;
    wire SubCellInst_SboxInst_12_n3 ;
    wire SubCellInst_SboxInst_12_n2 ;
    wire SubCellInst_SboxInst_12_n1 ;
    wire SubCellInst_SboxInst_13_n15 ;
    wire SubCellInst_SboxInst_13_n14 ;
    wire SubCellInst_SboxInst_13_n13 ;
    wire SubCellInst_SboxInst_13_n12 ;
    wire SubCellInst_SboxInst_13_n11 ;
    wire SubCellInst_SboxInst_13_n10 ;
    wire SubCellInst_SboxInst_13_n9 ;
    wire SubCellInst_SboxInst_13_n8 ;
    wire SubCellInst_SboxInst_13_n7 ;
    wire SubCellInst_SboxInst_13_n6 ;
    wire SubCellInst_SboxInst_13_n5 ;
    wire SubCellInst_SboxInst_13_n4 ;
    wire SubCellInst_SboxInst_13_n3 ;
    wire SubCellInst_SboxInst_13_n2 ;
    wire SubCellInst_SboxInst_13_n1 ;
    wire SubCellInst_SboxInst_14_n15 ;
    wire SubCellInst_SboxInst_14_n14 ;
    wire SubCellInst_SboxInst_14_n13 ;
    wire SubCellInst_SboxInst_14_n12 ;
    wire SubCellInst_SboxInst_14_n11 ;
    wire SubCellInst_SboxInst_14_n10 ;
    wire SubCellInst_SboxInst_14_n9 ;
    wire SubCellInst_SboxInst_14_n8 ;
    wire SubCellInst_SboxInst_14_n7 ;
    wire SubCellInst_SboxInst_14_n6 ;
    wire SubCellInst_SboxInst_14_n5 ;
    wire SubCellInst_SboxInst_14_n4 ;
    wire SubCellInst_SboxInst_14_n3 ;
    wire SubCellInst_SboxInst_14_n2 ;
    wire SubCellInst_SboxInst_14_n1 ;
    wire SubCellInst_SboxInst_15_n15 ;
    wire SubCellInst_SboxInst_15_n14 ;
    wire SubCellInst_SboxInst_15_n13 ;
    wire SubCellInst_SboxInst_15_n12 ;
    wire SubCellInst_SboxInst_15_n11 ;
    wire SubCellInst_SboxInst_15_n10 ;
    wire SubCellInst_SboxInst_15_n9 ;
    wire SubCellInst_SboxInst_15_n8 ;
    wire SubCellInst_SboxInst_15_n7 ;
    wire SubCellInst_SboxInst_15_n6 ;
    wire SubCellInst_SboxInst_15_n5 ;
    wire SubCellInst_SboxInst_15_n4 ;
    wire SubCellInst_SboxInst_15_n3 ;
    wire SubCellInst_SboxInst_15_n2 ;
    wire SubCellInst_SboxInst_15_n1 ;
    wire KeyMUX_n9 ;
    wire KeyMUX_n8 ;
    wire KeyMUX_n7 ;
    wire FSMSignalsInst_n5 ;
    wire FSMSignalsInst_n4 ;
    wire FSMSignalsInst_n3 ;
    wire FSMSignalsInst_n2 ;
    wire FSMSignalsInst_n1 ;
    wire selectsUpdateInst_n3 ;
    wire [63:0] Feedback ;
    wire [63:32] MCInput ;
    wire [63:0] MCOutput ;
    wire [63:0] SelectedKey ;
    wire [63:0] AddRoundKeyOutput ;
    wire [1:0] selects ;
    wire [6:0] FSMReg ;
    wire [6:0] FSMUpdate ;
    wire [1:0] selectsReg ;
    wire [1:0] selectsNext ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire clk_gated ;

    /* cells in depth 0 */
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2030, new_AGEMA_signal_2029, SelectedKey[40]}), .b ({1'b0, 1'b0, RoundConstant_0}), .c ({new_AGEMA_signal_2396, new_AGEMA_signal_2395, AddKeyConstXOR_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2036, new_AGEMA_signal_2035, SelectedKey[41]}), .b ({1'b0, 1'b0, FSMUpdate[0]}), .c ({new_AGEMA_signal_2398, new_AGEMA_signal_2397, AddKeyConstXOR_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2042, new_AGEMA_signal_2041, SelectedKey[42]}), .b ({1'b0, 1'b0, FSMUpdate[1]}), .c ({new_AGEMA_signal_2400, new_AGEMA_signal_2399, AddKeyConstXOR_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2048, new_AGEMA_signal_2047, SelectedKey[43]}), .b ({1'b0, 1'b0, 1'b0}), .c ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, AddKeyConstXOR_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, SelectedKey[44]}), .b ({1'b0, 1'b0, RoundConstant_4_}), .c ({new_AGEMA_signal_2404, new_AGEMA_signal_2403, AddKeyConstXOR_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2060, new_AGEMA_signal_2059, SelectedKey[45]}), .b ({1'b0, 1'b0, FSMUpdate[3]}), .c ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, AddKeyConstXOR_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2066, new_AGEMA_signal_2065, SelectedKey[46]}), .b ({1'b0, 1'b0, FSMUpdate[4]}), .c ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, AddKeyConstXOR_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, SelectedKey[47]}), .b ({1'b0, 1'b0, FSMUpdate[5]}), .c ({new_AGEMA_signal_2410, new_AGEMA_signal_2409, AddKeyConstXOR_XORInst_1_3_n1}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U4 ( .a ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_1030, new_AGEMA_signal_1029, SubCellInst_SboxInst_0_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U2 ( .a ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_1032, new_AGEMA_signal_1031, SubCellInst_SboxInst_0_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U1 ( .a ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, SubCellInst_SboxInst_0_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U4 ( .a ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, SubCellInst_SboxInst_1_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U2 ( .a ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .b ({new_AGEMA_signal_1048, new_AGEMA_signal_1047, SubCellInst_SboxInst_1_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U1 ( .a ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .b ({new_AGEMA_signal_1050, new_AGEMA_signal_1049, SubCellInst_SboxInst_1_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U4 ( .a ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .b ({new_AGEMA_signal_1062, new_AGEMA_signal_1061, SubCellInst_SboxInst_2_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U2 ( .a ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, SubCellInst_SboxInst_2_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U1 ( .a ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({new_AGEMA_signal_1066, new_AGEMA_signal_1065, SubCellInst_SboxInst_2_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U4 ( .a ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_1078, new_AGEMA_signal_1077, SubCellInst_SboxInst_3_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U2 ( .a ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_1080, new_AGEMA_signal_1079, SubCellInst_SboxInst_3_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U1 ( .a ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .b ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, SubCellInst_SboxInst_3_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U4 ( .a ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, SubCellInst_SboxInst_4_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U2 ( .a ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .b ({new_AGEMA_signal_1096, new_AGEMA_signal_1095, SubCellInst_SboxInst_4_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U1 ( .a ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .b ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, SubCellInst_SboxInst_4_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U4 ( .a ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .b ({new_AGEMA_signal_1110, new_AGEMA_signal_1109, SubCellInst_SboxInst_5_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U2 ( .a ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, SubCellInst_SboxInst_5_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U1 ( .a ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, SubCellInst_SboxInst_5_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U4 ( .a ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_1126, new_AGEMA_signal_1125, SubCellInst_SboxInst_6_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U2 ( .a ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .b ({new_AGEMA_signal_1128, new_AGEMA_signal_1127, SubCellInst_SboxInst_6_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U1 ( .a ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .b ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, SubCellInst_SboxInst_6_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U4 ( .a ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .b ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, SubCellInst_SboxInst_7_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U2 ( .a ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, SubCellInst_SboxInst_7_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U1 ( .a ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({new_AGEMA_signal_1146, new_AGEMA_signal_1145, SubCellInst_SboxInst_7_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U4 ( .a ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, SubCellInst_SboxInst_8_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U2 ( .a ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .b ({new_AGEMA_signal_1160, new_AGEMA_signal_1159, SubCellInst_SboxInst_8_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U1 ( .a ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .b ({new_AGEMA_signal_1162, new_AGEMA_signal_1161, SubCellInst_SboxInst_8_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U4 ( .a ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_1174, new_AGEMA_signal_1173, SubCellInst_SboxInst_9_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U2 ( .a ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_1176, new_AGEMA_signal_1175, SubCellInst_SboxInst_9_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U1 ( .a ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, SubCellInst_SboxInst_9_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U4 ( .a ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, SubCellInst_SboxInst_10_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U2 ( .a ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_1192, new_AGEMA_signal_1191, SubCellInst_SboxInst_10_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U1 ( .a ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .b ({new_AGEMA_signal_1194, new_AGEMA_signal_1193, SubCellInst_SboxInst_10_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U4 ( .a ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .b ({new_AGEMA_signal_1206, new_AGEMA_signal_1205, SubCellInst_SboxInst_11_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U2 ( .a ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, SubCellInst_SboxInst_11_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U1 ( .a ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({new_AGEMA_signal_1210, new_AGEMA_signal_1209, SubCellInst_SboxInst_11_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U4 ( .a ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .b ({new_AGEMA_signal_1222, new_AGEMA_signal_1221, SubCellInst_SboxInst_12_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U2 ( .a ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({new_AGEMA_signal_1224, new_AGEMA_signal_1223, SubCellInst_SboxInst_12_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U1 ( .a ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({new_AGEMA_signal_1226, new_AGEMA_signal_1225, SubCellInst_SboxInst_12_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U4 ( .a ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, SubCellInst_SboxInst_13_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U2 ( .a ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .b ({new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_13_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U1 ( .a ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .b ({new_AGEMA_signal_1242, new_AGEMA_signal_1241, SubCellInst_SboxInst_13_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U4 ( .a ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .b ({new_AGEMA_signal_1254, new_AGEMA_signal_1253, SubCellInst_SboxInst_14_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U2 ( .a ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, SubCellInst_SboxInst_14_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U1 ( .a ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_14_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U4 ( .a ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_1270, new_AGEMA_signal_1269, SubCellInst_SboxInst_15_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U2 ( .a ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .b ({new_AGEMA_signal_1272, new_AGEMA_signal_1271, SubCellInst_SboxInst_15_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U1 ( .a ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .b ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, SubCellInst_SboxInst_15_n9}) ) ;
    INV_X1 KeyMUX_U3 ( .A (selects[0]), .ZN (KeyMUX_n9) ) ;
    INV_X1 KeyMUX_U2 ( .A (KeyMUX_n9), .ZN (KeyMUX_n8) ) ;
    INV_X1 KeyMUX_U1 ( .A (KeyMUX_n9), .ZN (KeyMUX_n7) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_0_U1 ( .s (selects[0]), .b ({key_s2[64], key_s1[64], key_s0[64]}), .a ({key_s2[0], key_s1[0], key_s0[0]}), .c ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, SelectedKey[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_1_U1 ( .s (KeyMUX_n8), .b ({key_s2[65], key_s1[65], key_s0[65]}), .a ({key_s2[1], key_s1[1], key_s0[1]}), .c ({new_AGEMA_signal_1856, new_AGEMA_signal_1855, SelectedKey[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_2_U1 ( .s (selects[0]), .b ({key_s2[66], key_s1[66], key_s0[66]}), .a ({key_s2[2], key_s1[2], key_s0[2]}), .c ({new_AGEMA_signal_1478, new_AGEMA_signal_1477, SelectedKey[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_3_U1 ( .s (KeyMUX_n8), .b ({key_s2[67], key_s1[67], key_s0[67]}), .a ({key_s2[3], key_s1[3], key_s0[3]}), .c ({new_AGEMA_signal_1862, new_AGEMA_signal_1861, SelectedKey[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_4_U1 ( .s (KeyMUX_n8), .b ({key_s2[68], key_s1[68], key_s0[68]}), .a ({key_s2[4], key_s1[4], key_s0[4]}), .c ({new_AGEMA_signal_1868, new_AGEMA_signal_1867, SelectedKey[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_5_U1 ( .s (KeyMUX_n8), .b ({key_s2[69], key_s1[69], key_s0[69]}), .a ({key_s2[5], key_s1[5], key_s0[5]}), .c ({new_AGEMA_signal_1874, new_AGEMA_signal_1873, SelectedKey[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_6_U1 ( .s (KeyMUX_n8), .b ({key_s2[70], key_s1[70], key_s0[70]}), .a ({key_s2[6], key_s1[6], key_s0[6]}), .c ({new_AGEMA_signal_1880, new_AGEMA_signal_1879, SelectedKey[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_7_U1 ( .s (KeyMUX_n8), .b ({key_s2[71], key_s1[71], key_s0[71]}), .a ({key_s2[7], key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_1886, new_AGEMA_signal_1885, SelectedKey[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_8_U1 ( .s (KeyMUX_n8), .b ({key_s2[72], key_s1[72], key_s0[72]}), .a ({key_s2[8], key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_1892, new_AGEMA_signal_1891, SelectedKey[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_9_U1 ( .s (KeyMUX_n8), .b ({key_s2[73], key_s1[73], key_s0[73]}), .a ({key_s2[9], key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_1898, new_AGEMA_signal_1897, SelectedKey[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_10_U1 ( .s (KeyMUX_n8), .b ({key_s2[74], key_s1[74], key_s0[74]}), .a ({key_s2[10], key_s1[10], key_s0[10]}), .c ({new_AGEMA_signal_1904, new_AGEMA_signal_1903, SelectedKey[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_11_U1 ( .s (KeyMUX_n8), .b ({key_s2[75], key_s1[75], key_s0[75]}), .a ({key_s2[11], key_s1[11], key_s0[11]}), .c ({new_AGEMA_signal_1910, new_AGEMA_signal_1909, SelectedKey[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_12_U1 ( .s (KeyMUX_n8), .b ({key_s2[76], key_s1[76], key_s0[76]}), .a ({key_s2[12], key_s1[12], key_s0[12]}), .c ({new_AGEMA_signal_1916, new_AGEMA_signal_1915, SelectedKey[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_13_U1 ( .s (KeyMUX_n8), .b ({key_s2[77], key_s1[77], key_s0[77]}), .a ({key_s2[13], key_s1[13], key_s0[13]}), .c ({new_AGEMA_signal_1922, new_AGEMA_signal_1921, SelectedKey[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_14_U1 ( .s (KeyMUX_n8), .b ({key_s2[78], key_s1[78], key_s0[78]}), .a ({key_s2[14], key_s1[14], key_s0[14]}), .c ({new_AGEMA_signal_1928, new_AGEMA_signal_1927, SelectedKey[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_15_U1 ( .s (KeyMUX_n8), .b ({key_s2[79], key_s1[79], key_s0[79]}), .a ({key_s2[15], key_s1[15], key_s0[15]}), .c ({new_AGEMA_signal_1934, new_AGEMA_signal_1933, SelectedKey[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_16_U1 ( .s (KeyMUX_n8), .b ({key_s2[80], key_s1[80], key_s0[80]}), .a ({key_s2[16], key_s1[16], key_s0[16]}), .c ({new_AGEMA_signal_1940, new_AGEMA_signal_1939, SelectedKey[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_17_U1 ( .s (KeyMUX_n8), .b ({key_s2[81], key_s1[81], key_s0[81]}), .a ({key_s2[17], key_s1[17], key_s0[17]}), .c ({new_AGEMA_signal_1946, new_AGEMA_signal_1945, SelectedKey[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_18_U1 ( .s (KeyMUX_n8), .b ({key_s2[82], key_s1[82], key_s0[82]}), .a ({key_s2[18], key_s1[18], key_s0[18]}), .c ({new_AGEMA_signal_1952, new_AGEMA_signal_1951, SelectedKey[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_19_U1 ( .s (KeyMUX_n8), .b ({key_s2[83], key_s1[83], key_s0[83]}), .a ({key_s2[19], key_s1[19], key_s0[19]}), .c ({new_AGEMA_signal_1958, new_AGEMA_signal_1957, SelectedKey[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_20_U1 ( .s (KeyMUX_n8), .b ({key_s2[84], key_s1[84], key_s0[84]}), .a ({key_s2[20], key_s1[20], key_s0[20]}), .c ({new_AGEMA_signal_1964, new_AGEMA_signal_1963, SelectedKey[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_21_U1 ( .s (KeyMUX_n8), .b ({key_s2[85], key_s1[85], key_s0[85]}), .a ({key_s2[21], key_s1[21], key_s0[21]}), .c ({new_AGEMA_signal_1970, new_AGEMA_signal_1969, SelectedKey[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_22_U1 ( .s (selects[0]), .b ({key_s2[86], key_s1[86], key_s0[86]}), .a ({key_s2[22], key_s1[22], key_s0[22]}), .c ({new_AGEMA_signal_1484, new_AGEMA_signal_1483, SelectedKey[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_23_U1 ( .s (selects[0]), .b ({key_s2[87], key_s1[87], key_s0[87]}), .a ({key_s2[23], key_s1[23], key_s0[23]}), .c ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, SelectedKey[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_24_U1 ( .s (selects[0]), .b ({key_s2[88], key_s1[88], key_s0[88]}), .a ({key_s2[24], key_s1[24], key_s0[24]}), .c ({new_AGEMA_signal_1496, new_AGEMA_signal_1495, SelectedKey[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_25_U1 ( .s (selects[0]), .b ({key_s2[89], key_s1[89], key_s0[89]}), .a ({key_s2[25], key_s1[25], key_s0[25]}), .c ({new_AGEMA_signal_1502, new_AGEMA_signal_1501, SelectedKey[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_26_U1 ( .s (selects[0]), .b ({key_s2[90], key_s1[90], key_s0[90]}), .a ({key_s2[26], key_s1[26], key_s0[26]}), .c ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, SelectedKey[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_27_U1 ( .s (selects[0]), .b ({key_s2[91], key_s1[91], key_s0[91]}), .a ({key_s2[27], key_s1[27], key_s0[27]}), .c ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, SelectedKey[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_28_U1 ( .s (KeyMUX_n7), .b ({key_s2[92], key_s1[92], key_s0[92]}), .a ({key_s2[28], key_s1[28], key_s0[28]}), .c ({new_AGEMA_signal_1976, new_AGEMA_signal_1975, SelectedKey[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_29_U1 ( .s (KeyMUX_n7), .b ({key_s2[93], key_s1[93], key_s0[93]}), .a ({key_s2[29], key_s1[29], key_s0[29]}), .c ({new_AGEMA_signal_1982, new_AGEMA_signal_1981, SelectedKey[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_30_U1 ( .s (KeyMUX_n7), .b ({key_s2[94], key_s1[94], key_s0[94]}), .a ({key_s2[30], key_s1[30], key_s0[30]}), .c ({new_AGEMA_signal_1988, new_AGEMA_signal_1987, SelectedKey[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_31_U1 ( .s (KeyMUX_n7), .b ({key_s2[95], key_s1[95], key_s0[95]}), .a ({key_s2[31], key_s1[31], key_s0[31]}), .c ({new_AGEMA_signal_1994, new_AGEMA_signal_1993, SelectedKey[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_32_U1 ( .s (KeyMUX_n7), .b ({key_s2[96], key_s1[96], key_s0[96]}), .a ({key_s2[32], key_s1[32], key_s0[32]}), .c ({new_AGEMA_signal_2000, new_AGEMA_signal_1999, SelectedKey[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_33_U1 ( .s (selects[0]), .b ({key_s2[97], key_s1[97], key_s0[97]}), .a ({key_s2[33], key_s1[33], key_s0[33]}), .c ({new_AGEMA_signal_1520, new_AGEMA_signal_1519, SelectedKey[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_34_U1 ( .s (KeyMUX_n7), .b ({key_s2[98], key_s1[98], key_s0[98]}), .a ({key_s2[34], key_s1[34], key_s0[34]}), .c ({new_AGEMA_signal_2006, new_AGEMA_signal_2005, SelectedKey[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_35_U1 ( .s (KeyMUX_n7), .b ({key_s2[99], key_s1[99], key_s0[99]}), .a ({key_s2[35], key_s1[35], key_s0[35]}), .c ({new_AGEMA_signal_2012, new_AGEMA_signal_2011, SelectedKey[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_36_U1 ( .s (selects[0]), .b ({key_s2[100], key_s1[100], key_s0[100]}), .a ({key_s2[36], key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, SelectedKey[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_37_U1 ( .s (KeyMUX_n7), .b ({key_s2[101], key_s1[101], key_s0[101]}), .a ({key_s2[37], key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_2018, new_AGEMA_signal_2017, SelectedKey[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_38_U1 ( .s (KeyMUX_n7), .b ({key_s2[102], key_s1[102], key_s0[102]}), .a ({key_s2[38], key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_2024, new_AGEMA_signal_2023, SelectedKey[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_39_U1 ( .s (selects[0]), .b ({key_s2[103], key_s1[103], key_s0[103]}), .a ({key_s2[39], key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_1532, new_AGEMA_signal_1531, SelectedKey[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_40_U1 ( .s (KeyMUX_n7), .b ({key_s2[104], key_s1[104], key_s0[104]}), .a ({key_s2[40], key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_2030, new_AGEMA_signal_2029, SelectedKey[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_41_U1 ( .s (KeyMUX_n7), .b ({key_s2[105], key_s1[105], key_s0[105]}), .a ({key_s2[41], key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_2036, new_AGEMA_signal_2035, SelectedKey[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_42_U1 ( .s (KeyMUX_n7), .b ({key_s2[106], key_s1[106], key_s0[106]}), .a ({key_s2[42], key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_2042, new_AGEMA_signal_2041, SelectedKey[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_43_U1 ( .s (KeyMUX_n7), .b ({key_s2[107], key_s1[107], key_s0[107]}), .a ({key_s2[43], key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_2048, new_AGEMA_signal_2047, SelectedKey[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_44_U1 ( .s (KeyMUX_n7), .b ({key_s2[108], key_s1[108], key_s0[108]}), .a ({key_s2[44], key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, SelectedKey[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_45_U1 ( .s (KeyMUX_n7), .b ({key_s2[109], key_s1[109], key_s0[109]}), .a ({key_s2[45], key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_2060, new_AGEMA_signal_2059, SelectedKey[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_46_U1 ( .s (KeyMUX_n7), .b ({key_s2[110], key_s1[110], key_s0[110]}), .a ({key_s2[46], key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_2066, new_AGEMA_signal_2065, SelectedKey[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_47_U1 ( .s (KeyMUX_n7), .b ({key_s2[111], key_s1[111], key_s0[111]}), .a ({key_s2[47], key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, SelectedKey[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_48_U1 ( .s (KeyMUX_n7), .b ({key_s2[112], key_s1[112], key_s0[112]}), .a ({key_s2[48], key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, SelectedKey[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_49_U1 ( .s (KeyMUX_n7), .b ({key_s2[113], key_s1[113], key_s0[113]}), .a ({key_s2[49], key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_2084, new_AGEMA_signal_2083, SelectedKey[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_50_U1 ( .s (KeyMUX_n7), .b ({key_s2[114], key_s1[114], key_s0[114]}), .a ({key_s2[50], key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, SelectedKey[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_51_U1 ( .s (KeyMUX_n7), .b ({key_s2[115], key_s1[115], key_s0[115]}), .a ({key_s2[51], key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_2096, new_AGEMA_signal_2095, SelectedKey[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_52_U1 ( .s (KeyMUX_n7), .b ({key_s2[116], key_s1[116], key_s0[116]}), .a ({key_s2[52], key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_2102, new_AGEMA_signal_2101, SelectedKey[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_53_U1 ( .s (selects[0]), .b ({key_s2[117], key_s1[117], key_s0[117]}), .a ({key_s2[53], key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_1538, new_AGEMA_signal_1537, SelectedKey[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_54_U1 ( .s (selects[0]), .b ({key_s2[118], key_s1[118], key_s0[118]}), .a ({key_s2[54], key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, SelectedKey[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_55_U1 ( .s (KeyMUX_n7), .b ({key_s2[119], key_s1[119], key_s0[119]}), .a ({key_s2[55], key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_2108, new_AGEMA_signal_2107, SelectedKey[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_56_U1 ( .s (selects[0]), .b ({key_s2[120], key_s1[120], key_s0[120]}), .a ({key_s2[56], key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, SelectedKey[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_57_U1 ( .s (KeyMUX_n7), .b ({key_s2[121], key_s1[121], key_s0[121]}), .a ({key_s2[57], key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, SelectedKey[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_58_U1 ( .s (KeyMUX_n7), .b ({key_s2[122], key_s1[122], key_s0[122]}), .a ({key_s2[58], key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_2120, new_AGEMA_signal_2119, SelectedKey[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_59_U1 ( .s (selects[0]), .b ({key_s2[123], key_s1[123], key_s0[123]}), .a ({key_s2[59], key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, SelectedKey[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_60_U1 ( .s (KeyMUX_n7), .b ({key_s2[124], key_s1[124], key_s0[124]}), .a ({key_s2[60], key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, SelectedKey[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_61_U1 ( .s (KeyMUX_n7), .b ({key_s2[125], key_s1[125], key_s0[125]}), .a ({key_s2[61], key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_2132, new_AGEMA_signal_2131, SelectedKey[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_62_U1 ( .s (selects[0]), .b ({key_s2[126], key_s1[126], key_s0[126]}), .a ({key_s2[62], key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, SelectedKey[62]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyMUX_MUXInst_63_U1 ( .s (KeyMUX_n7), .b ({key_s2[127], key_s1[127], key_s0[127]}), .a ({key_s2[63], key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_2138, new_AGEMA_signal_2137, SelectedKey[63]}) ) ;
    MUX2_X1 FSMMUX_MUXInst_0_U1 ( .S (rst), .A (FSMReg[0]), .B (1'b1), .Z (RoundConstant_0) ) ;
    MUX2_X1 FSMMUX_MUXInst_1_U1 ( .S (rst), .A (FSMReg[1]), .B (1'b0), .Z (FSMUpdate[0]) ) ;
    MUX2_X1 FSMMUX_MUXInst_2_U1 ( .S (rst), .A (FSMReg[2]), .B (1'b0), .Z (FSMUpdate[1]) ) ;
    MUX2_X1 FSMMUX_MUXInst_3_U1 ( .S (rst), .A (FSMReg[3]), .B (1'b1), .Z (RoundConstant_4_) ) ;
    MUX2_X1 FSMMUX_MUXInst_4_U1 ( .S (rst), .A (FSMReg[4]), .B (1'b0), .Z (FSMUpdate[3]) ) ;
    MUX2_X1 FSMMUX_MUXInst_5_U1 ( .S (rst), .A (FSMReg[5]), .B (1'b0), .Z (FSMUpdate[4]) ) ;
    MUX2_X1 FSMMUX_MUXInst_6_U1 ( .S (rst), .A (FSMReg[6]), .B (1'b0), .Z (FSMUpdate[5]) ) ;
    XOR2_X1 FSMUpdateInst_U2 ( .A (RoundConstant_4_), .B (FSMUpdate[3]), .Z (FSMUpdate[6]) ) ;
    XOR2_X1 FSMUpdateInst_U1 ( .A (FSMUpdate[0]), .B (RoundConstant_0), .Z (FSMUpdate[2]) ) ;
    AND2_X1 FSMSignalsInst_U6 ( .A1 (FSMUpdate[5]), .A2 (FSMSignalsInst_n5), .ZN (done_internal) ) ;
    NOR2_X1 FSMSignalsInst_U5 ( .A1 (FSMSignalsInst_n4), .A2 (FSMSignalsInst_n3), .ZN (FSMSignalsInst_n5) ) ;
    NAND2_X1 FSMSignalsInst_U4 ( .A1 (FSMSignalsInst_n2), .A2 (FSMSignalsInst_n1), .ZN (FSMSignalsInst_n3) ) ;
    NOR2_X1 FSMSignalsInst_U3 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdate[4]), .ZN (FSMSignalsInst_n1) ) ;
    NOR2_X1 FSMSignalsInst_U2 ( .A1 (FSMUpdate[0]), .A2 (RoundConstant_4_), .ZN (FSMSignalsInst_n2) ) ;
    NAND2_X1 FSMSignalsInst_U1 ( .A1 (RoundConstant_0), .A2 (FSMUpdate[1]), .ZN (FSMSignalsInst_n4) ) ;
    MUX2_X1 selectsMUX_MUXInst_0_U1 ( .S (rst), .A (selectsReg[0]), .B (1'b0), .Z (selects[0]) ) ;
    MUX2_X1 selectsMUX_MUXInst_1_U1 ( .S (rst), .A (selectsReg[1]), .B (1'b0), .Z (selects[1]) ) ;
    XNOR2_X1 selectsUpdateInst_U3 ( .A (selectsUpdateInst_n3), .B (selects[1]), .ZN (selectsNext[1]) ) ;
    XNOR2_X1 selectsUpdateInst_U2 ( .A (selects[0]), .B (1'b0), .ZN (selectsUpdateInst_n3) ) ;
    INV_X1 selectsUpdateInst_U1 ( .A (selects[0]), .ZN (selectsNext[0]) ) ;
    ClockGatingController #(9) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U14 ( .a ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_1024, new_AGEMA_signal_1023, SubCellInst_SboxInst_0_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U13 ( .a ({new_AGEMA_signal_1032, new_AGEMA_signal_1031, SubCellInst_SboxInst_0_n8}), .b ({new_AGEMA_signal_1030, new_AGEMA_signal_1029, SubCellInst_SboxInst_0_n7}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, SubCellInst_SboxInst_0_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U10 ( .a ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, SubCellInst_SboxInst_0_n9}), .clk (clk), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, SubCellInst_SboxInst_0_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U9 ( .a ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_1032, new_AGEMA_signal_1031, SubCellInst_SboxInst_0_n8}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({new_AGEMA_signal_1282, new_AGEMA_signal_1281, SubCellInst_SboxInst_0_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U5 ( .a ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, SubCellInst_SboxInst_0_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U3 ( .a ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, SubCellInst_SboxInst_0_n9}), .b ({new_AGEMA_signal_1032, new_AGEMA_signal_1031, SubCellInst_SboxInst_0_n8}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, SubCellInst_SboxInst_0_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U14 ( .a ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .b ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .clk (clk), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_1040, new_AGEMA_signal_1039, SubCellInst_SboxInst_1_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U13 ( .a ({new_AGEMA_signal_1048, new_AGEMA_signal_1047, SubCellInst_SboxInst_1_n8}), .b ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, SubCellInst_SboxInst_1_n7}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({new_AGEMA_signal_1290, new_AGEMA_signal_1289, SubCellInst_SboxInst_1_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U10 ( .a ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .b ({new_AGEMA_signal_1050, new_AGEMA_signal_1049, SubCellInst_SboxInst_1_n9}), .clk (clk), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, SubCellInst_SboxInst_1_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U9 ( .a ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .b ({new_AGEMA_signal_1048, new_AGEMA_signal_1047, SubCellInst_SboxInst_1_n8}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({new_AGEMA_signal_1294, new_AGEMA_signal_1293, SubCellInst_SboxInst_1_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U5 ( .a ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .b ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .clk (clk), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_1044, new_AGEMA_signal_1043, SubCellInst_SboxInst_1_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U3 ( .a ({new_AGEMA_signal_1050, new_AGEMA_signal_1049, SubCellInst_SboxInst_1_n9}), .b ({new_AGEMA_signal_1048, new_AGEMA_signal_1047, SubCellInst_SboxInst_1_n8}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({new_AGEMA_signal_1298, new_AGEMA_signal_1297, SubCellInst_SboxInst_1_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U14 ( .a ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_1056, new_AGEMA_signal_1055, SubCellInst_SboxInst_2_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U13 ( .a ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, SubCellInst_SboxInst_2_n8}), .b ({new_AGEMA_signal_1062, new_AGEMA_signal_1061, SubCellInst_SboxInst_2_n7}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({new_AGEMA_signal_1302, new_AGEMA_signal_1301, SubCellInst_SboxInst_2_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U10 ( .a ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({new_AGEMA_signal_1066, new_AGEMA_signal_1065, SubCellInst_SboxInst_2_n9}), .clk (clk), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, SubCellInst_SboxInst_2_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U9 ( .a ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, SubCellInst_SboxInst_2_n8}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({new_AGEMA_signal_1306, new_AGEMA_signal_1305, SubCellInst_SboxInst_2_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U5 ( .a ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_1060, new_AGEMA_signal_1059, SubCellInst_SboxInst_2_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U3 ( .a ({new_AGEMA_signal_1066, new_AGEMA_signal_1065, SubCellInst_SboxInst_2_n9}), .b ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, SubCellInst_SboxInst_2_n8}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({new_AGEMA_signal_1310, new_AGEMA_signal_1309, SubCellInst_SboxInst_2_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U14 ( .a ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .clk (clk), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_1072, new_AGEMA_signal_1071, SubCellInst_SboxInst_3_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U13 ( .a ({new_AGEMA_signal_1080, new_AGEMA_signal_1079, SubCellInst_SboxInst_3_n8}), .b ({new_AGEMA_signal_1078, new_AGEMA_signal_1077, SubCellInst_SboxInst_3_n7}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({new_AGEMA_signal_1314, new_AGEMA_signal_1313, SubCellInst_SboxInst_3_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U10 ( .a ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, SubCellInst_SboxInst_3_n9}), .clk (clk), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, SubCellInst_SboxInst_3_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U9 ( .a ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .b ({new_AGEMA_signal_1080, new_AGEMA_signal_1079, SubCellInst_SboxInst_3_n8}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({new_AGEMA_signal_1318, new_AGEMA_signal_1317, SubCellInst_SboxInst_3_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U5 ( .a ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .clk (clk), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, SubCellInst_SboxInst_3_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U3 ( .a ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, SubCellInst_SboxInst_3_n9}), .b ({new_AGEMA_signal_1080, new_AGEMA_signal_1079, SubCellInst_SboxInst_3_n8}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, SubCellInst_SboxInst_3_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U14 ( .a ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .b ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .clk (clk), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, SubCellInst_SboxInst_4_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U13 ( .a ({new_AGEMA_signal_1096, new_AGEMA_signal_1095, SubCellInst_SboxInst_4_n8}), .b ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, SubCellInst_SboxInst_4_n7}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({new_AGEMA_signal_1326, new_AGEMA_signal_1325, SubCellInst_SboxInst_4_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U10 ( .a ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .b ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, SubCellInst_SboxInst_4_n9}), .clk (clk), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, SubCellInst_SboxInst_4_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U9 ( .a ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .b ({new_AGEMA_signal_1096, new_AGEMA_signal_1095, SubCellInst_SboxInst_4_n8}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({new_AGEMA_signal_1330, new_AGEMA_signal_1329, SubCellInst_SboxInst_4_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U5 ( .a ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .b ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .clk (clk), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_1092, new_AGEMA_signal_1091, SubCellInst_SboxInst_4_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U3 ( .a ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, SubCellInst_SboxInst_4_n9}), .b ({new_AGEMA_signal_1096, new_AGEMA_signal_1095, SubCellInst_SboxInst_4_n8}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({new_AGEMA_signal_1334, new_AGEMA_signal_1333, SubCellInst_SboxInst_4_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U14 ( .a ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_1104, new_AGEMA_signal_1103, SubCellInst_SboxInst_5_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U13 ( .a ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, SubCellInst_SboxInst_5_n8}), .b ({new_AGEMA_signal_1110, new_AGEMA_signal_1109, SubCellInst_SboxInst_5_n7}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({new_AGEMA_signal_1338, new_AGEMA_signal_1337, SubCellInst_SboxInst_5_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U10 ( .a ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, SubCellInst_SboxInst_5_n9}), .clk (clk), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, SubCellInst_SboxInst_5_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U9 ( .a ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, SubCellInst_SboxInst_5_n8}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({new_AGEMA_signal_1342, new_AGEMA_signal_1341, SubCellInst_SboxInst_5_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U5 ( .a ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r ({Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_1108, new_AGEMA_signal_1107, SubCellInst_SboxInst_5_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U3 ( .a ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, SubCellInst_SboxInst_5_n9}), .b ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, SubCellInst_SboxInst_5_n8}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105]}), .c ({new_AGEMA_signal_1346, new_AGEMA_signal_1345, SubCellInst_SboxInst_5_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U14 ( .a ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .b ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .clk (clk), .r ({Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_1120, new_AGEMA_signal_1119, SubCellInst_SboxInst_6_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U13 ( .a ({new_AGEMA_signal_1128, new_AGEMA_signal_1127, SubCellInst_SboxInst_6_n8}), .b ({new_AGEMA_signal_1126, new_AGEMA_signal_1125, SubCellInst_SboxInst_6_n7}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111]}), .c ({new_AGEMA_signal_1350, new_AGEMA_signal_1349, SubCellInst_SboxInst_6_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U10 ( .a ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .b ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, SubCellInst_SboxInst_6_n9}), .clk (clk), .r ({Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_1352, new_AGEMA_signal_1351, SubCellInst_SboxInst_6_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U9 ( .a ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .b ({new_AGEMA_signal_1128, new_AGEMA_signal_1127, SubCellInst_SboxInst_6_n8}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117]}), .c ({new_AGEMA_signal_1354, new_AGEMA_signal_1353, SubCellInst_SboxInst_6_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U5 ( .a ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .b ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .clk (clk), .r ({Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, SubCellInst_SboxInst_6_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U3 ( .a ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, SubCellInst_SboxInst_6_n9}), .b ({new_AGEMA_signal_1128, new_AGEMA_signal_1127, SubCellInst_SboxInst_6_n8}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123]}), .c ({new_AGEMA_signal_1358, new_AGEMA_signal_1357, SubCellInst_SboxInst_6_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U14 ( .a ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r ({Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, SubCellInst_SboxInst_7_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U13 ( .a ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, SubCellInst_SboxInst_7_n8}), .b ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, SubCellInst_SboxInst_7_n7}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129]}), .c ({new_AGEMA_signal_1362, new_AGEMA_signal_1361, SubCellInst_SboxInst_7_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U10 ( .a ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({new_AGEMA_signal_1146, new_AGEMA_signal_1145, SubCellInst_SboxInst_7_n9}), .clk (clk), .r ({Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_1364, new_AGEMA_signal_1363, SubCellInst_SboxInst_7_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U9 ( .a ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, SubCellInst_SboxInst_7_n8}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135]}), .c ({new_AGEMA_signal_1366, new_AGEMA_signal_1365, SubCellInst_SboxInst_7_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U5 ( .a ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r ({Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_1140, new_AGEMA_signal_1139, SubCellInst_SboxInst_7_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U3 ( .a ({new_AGEMA_signal_1146, new_AGEMA_signal_1145, SubCellInst_SboxInst_7_n9}), .b ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, SubCellInst_SboxInst_7_n8}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141]}), .c ({new_AGEMA_signal_1370, new_AGEMA_signal_1369, SubCellInst_SboxInst_7_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U14 ( .a ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .b ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .clk (clk), .r ({Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_1152, new_AGEMA_signal_1151, SubCellInst_SboxInst_8_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U13 ( .a ({new_AGEMA_signal_1160, new_AGEMA_signal_1159, SubCellInst_SboxInst_8_n8}), .b ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, SubCellInst_SboxInst_8_n7}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147]}), .c ({new_AGEMA_signal_1374, new_AGEMA_signal_1373, SubCellInst_SboxInst_8_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U10 ( .a ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .b ({new_AGEMA_signal_1162, new_AGEMA_signal_1161, SubCellInst_SboxInst_8_n9}), .clk (clk), .r ({Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_1376, new_AGEMA_signal_1375, SubCellInst_SboxInst_8_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U9 ( .a ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .b ({new_AGEMA_signal_1160, new_AGEMA_signal_1159, SubCellInst_SboxInst_8_n8}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153]}), .c ({new_AGEMA_signal_1378, new_AGEMA_signal_1377, SubCellInst_SboxInst_8_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U5 ( .a ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .b ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .clk (clk), .r ({Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_1156, new_AGEMA_signal_1155, SubCellInst_SboxInst_8_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U3 ( .a ({new_AGEMA_signal_1162, new_AGEMA_signal_1161, SubCellInst_SboxInst_8_n9}), .b ({new_AGEMA_signal_1160, new_AGEMA_signal_1159, SubCellInst_SboxInst_8_n8}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159]}), .c ({new_AGEMA_signal_1382, new_AGEMA_signal_1381, SubCellInst_SboxInst_8_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U14 ( .a ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r ({Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_1168, new_AGEMA_signal_1167, SubCellInst_SboxInst_9_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U13 ( .a ({new_AGEMA_signal_1176, new_AGEMA_signal_1175, SubCellInst_SboxInst_9_n8}), .b ({new_AGEMA_signal_1174, new_AGEMA_signal_1173, SubCellInst_SboxInst_9_n7}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165]}), .c ({new_AGEMA_signal_1386, new_AGEMA_signal_1385, SubCellInst_SboxInst_9_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U10 ( .a ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, SubCellInst_SboxInst_9_n9}), .clk (clk), .r ({Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_1388, new_AGEMA_signal_1387, SubCellInst_SboxInst_9_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U9 ( .a ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_1176, new_AGEMA_signal_1175, SubCellInst_SboxInst_9_n8}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171]}), .c ({new_AGEMA_signal_1390, new_AGEMA_signal_1389, SubCellInst_SboxInst_9_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U5 ( .a ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r ({Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_1172, new_AGEMA_signal_1171, SubCellInst_SboxInst_9_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U3 ( .a ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, SubCellInst_SboxInst_9_n9}), .b ({new_AGEMA_signal_1176, new_AGEMA_signal_1175, SubCellInst_SboxInst_9_n8}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177]}), .c ({new_AGEMA_signal_1394, new_AGEMA_signal_1393, SubCellInst_SboxInst_9_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U14 ( .a ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .clk (clk), .r ({Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_1184, new_AGEMA_signal_1183, SubCellInst_SboxInst_10_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U13 ( .a ({new_AGEMA_signal_1192, new_AGEMA_signal_1191, SubCellInst_SboxInst_10_n8}), .b ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, SubCellInst_SboxInst_10_n7}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183]}), .c ({new_AGEMA_signal_1398, new_AGEMA_signal_1397, SubCellInst_SboxInst_10_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U10 ( .a ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_1194, new_AGEMA_signal_1193, SubCellInst_SboxInst_10_n9}), .clk (clk), .r ({Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_1400, new_AGEMA_signal_1399, SubCellInst_SboxInst_10_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U9 ( .a ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .b ({new_AGEMA_signal_1192, new_AGEMA_signal_1191, SubCellInst_SboxInst_10_n8}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189]}), .c ({new_AGEMA_signal_1402, new_AGEMA_signal_1401, SubCellInst_SboxInst_10_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U5 ( .a ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .clk (clk), .r ({Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_1188, new_AGEMA_signal_1187, SubCellInst_SboxInst_10_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U3 ( .a ({new_AGEMA_signal_1194, new_AGEMA_signal_1193, SubCellInst_SboxInst_10_n9}), .b ({new_AGEMA_signal_1192, new_AGEMA_signal_1191, SubCellInst_SboxInst_10_n8}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195]}), .c ({new_AGEMA_signal_1406, new_AGEMA_signal_1405, SubCellInst_SboxInst_10_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U14 ( .a ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r ({Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_1200, new_AGEMA_signal_1199, SubCellInst_SboxInst_11_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U13 ( .a ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, SubCellInst_SboxInst_11_n8}), .b ({new_AGEMA_signal_1206, new_AGEMA_signal_1205, SubCellInst_SboxInst_11_n7}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201]}), .c ({new_AGEMA_signal_1410, new_AGEMA_signal_1409, SubCellInst_SboxInst_11_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U10 ( .a ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({new_AGEMA_signal_1210, new_AGEMA_signal_1209, SubCellInst_SboxInst_11_n9}), .clk (clk), .r ({Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_1412, new_AGEMA_signal_1411, SubCellInst_SboxInst_11_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U9 ( .a ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, SubCellInst_SboxInst_11_n8}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207]}), .c ({new_AGEMA_signal_1414, new_AGEMA_signal_1413, SubCellInst_SboxInst_11_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U5 ( .a ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r ({Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_1204, new_AGEMA_signal_1203, SubCellInst_SboxInst_11_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U3 ( .a ({new_AGEMA_signal_1210, new_AGEMA_signal_1209, SubCellInst_SboxInst_11_n9}), .b ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, SubCellInst_SboxInst_11_n8}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213]}), .c ({new_AGEMA_signal_1418, new_AGEMA_signal_1417, SubCellInst_SboxInst_11_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U14 ( .a ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r ({Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_1216, new_AGEMA_signal_1215, SubCellInst_SboxInst_12_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U13 ( .a ({new_AGEMA_signal_1224, new_AGEMA_signal_1223, SubCellInst_SboxInst_12_n8}), .b ({new_AGEMA_signal_1222, new_AGEMA_signal_1221, SubCellInst_SboxInst_12_n7}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219]}), .c ({new_AGEMA_signal_1422, new_AGEMA_signal_1421, SubCellInst_SboxInst_12_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U10 ( .a ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({new_AGEMA_signal_1226, new_AGEMA_signal_1225, SubCellInst_SboxInst_12_n9}), .clk (clk), .r ({Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_1424, new_AGEMA_signal_1423, SubCellInst_SboxInst_12_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U9 ( .a ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({new_AGEMA_signal_1224, new_AGEMA_signal_1223, SubCellInst_SboxInst_12_n8}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225]}), .c ({new_AGEMA_signal_1426, new_AGEMA_signal_1425, SubCellInst_SboxInst_12_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U5 ( .a ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r ({Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, SubCellInst_SboxInst_12_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U3 ( .a ({new_AGEMA_signal_1226, new_AGEMA_signal_1225, SubCellInst_SboxInst_12_n9}), .b ({new_AGEMA_signal_1224, new_AGEMA_signal_1223, SubCellInst_SboxInst_12_n8}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231]}), .c ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, SubCellInst_SboxInst_12_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U14 ( .a ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .b ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .clk (clk), .r ({Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, SubCellInst_SboxInst_13_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U13 ( .a ({new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_13_n8}), .b ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, SubCellInst_SboxInst_13_n7}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237]}), .c ({new_AGEMA_signal_1434, new_AGEMA_signal_1433, SubCellInst_SboxInst_13_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U10 ( .a ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .b ({new_AGEMA_signal_1242, new_AGEMA_signal_1241, SubCellInst_SboxInst_13_n9}), .clk (clk), .r ({Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_1436, new_AGEMA_signal_1435, SubCellInst_SboxInst_13_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U9 ( .a ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .b ({new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_13_n8}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243]}), .c ({new_AGEMA_signal_1438, new_AGEMA_signal_1437, SubCellInst_SboxInst_13_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U5 ( .a ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .b ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .clk (clk), .r ({Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_1236, new_AGEMA_signal_1235, SubCellInst_SboxInst_13_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U3 ( .a ({new_AGEMA_signal_1242, new_AGEMA_signal_1241, SubCellInst_SboxInst_13_n9}), .b ({new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_13_n8}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249]}), .c ({new_AGEMA_signal_1442, new_AGEMA_signal_1441, SubCellInst_SboxInst_13_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U14 ( .a ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r ({Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_1248, new_AGEMA_signal_1247, SubCellInst_SboxInst_14_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U13 ( .a ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, SubCellInst_SboxInst_14_n8}), .b ({new_AGEMA_signal_1254, new_AGEMA_signal_1253, SubCellInst_SboxInst_14_n7}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255]}), .c ({new_AGEMA_signal_1446, new_AGEMA_signal_1445, SubCellInst_SboxInst_14_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U10 ( .a ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_14_n9}), .clk (clk), .r ({Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_1448, new_AGEMA_signal_1447, SubCellInst_SboxInst_14_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U9 ( .a ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, SubCellInst_SboxInst_14_n8}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261]}), .c ({new_AGEMA_signal_1450, new_AGEMA_signal_1449, SubCellInst_SboxInst_14_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U5 ( .a ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r ({Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_1252, new_AGEMA_signal_1251, SubCellInst_SboxInst_14_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U3 ( .a ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_14_n9}), .b ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, SubCellInst_SboxInst_14_n8}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267]}), .c ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, SubCellInst_SboxInst_14_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U14 ( .a ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .b ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .clk (clk), .r ({Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_1264, new_AGEMA_signal_1263, SubCellInst_SboxInst_15_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U13 ( .a ({new_AGEMA_signal_1272, new_AGEMA_signal_1271, SubCellInst_SboxInst_15_n8}), .b ({new_AGEMA_signal_1270, new_AGEMA_signal_1269, SubCellInst_SboxInst_15_n7}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273]}), .c ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, SubCellInst_SboxInst_15_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U10 ( .a ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .b ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, SubCellInst_SboxInst_15_n9}), .clk (clk), .r ({Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_1460, new_AGEMA_signal_1459, SubCellInst_SboxInst_15_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U9 ( .a ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .b ({new_AGEMA_signal_1272, new_AGEMA_signal_1271, SubCellInst_SboxInst_15_n8}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279]}), .c ({new_AGEMA_signal_1462, new_AGEMA_signal_1461, SubCellInst_SboxInst_15_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U5 ( .a ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .b ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .clk (clk), .r ({Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, SubCellInst_SboxInst_15_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U3 ( .a ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, SubCellInst_SboxInst_15_n9}), .b ({new_AGEMA_signal_1272, new_AGEMA_signal_1271, SubCellInst_SboxInst_15_n8}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285]}), .c ({new_AGEMA_signal_1466, new_AGEMA_signal_1465, SubCellInst_SboxInst_15_n13}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    or_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U18 ( .a ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, SubCellInst_SboxInst_0_n13}), .b ({ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r ({Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_1566, new_AGEMA_signal_1565, SubCellInst_SboxInst_0_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U15 ( .a ({new_AGEMA_signal_1024, new_AGEMA_signal_1023, SubCellInst_SboxInst_0_n10}), .b ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, SubCellInst_SboxInst_0_n9}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291]}), .c ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_0_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U11 ( .a ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, SubCellInst_SboxInst_0_n4}), .clk (clk), .r ({Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_1570, new_AGEMA_signal_1569, SubCellInst_SboxInst_0_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U6 ( .a ({new_AGEMA_signal_1030, new_AGEMA_signal_1029, SubCellInst_SboxInst_0_n7}), .b ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, SubCellInst_SboxInst_0_n1}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297]}), .c ({new_AGEMA_signal_1284, new_AGEMA_signal_1283, SubCellInst_SboxInst_0_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U18 ( .a ({new_AGEMA_signal_1298, new_AGEMA_signal_1297, SubCellInst_SboxInst_1_n13}), .b ({ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .clk (clk), .r ({Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_1576, new_AGEMA_signal_1575, SubCellInst_SboxInst_1_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U15 ( .a ({new_AGEMA_signal_1040, new_AGEMA_signal_1039, SubCellInst_SboxInst_1_n10}), .b ({new_AGEMA_signal_1050, new_AGEMA_signal_1049, SubCellInst_SboxInst_1_n9}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303]}), .c ({new_AGEMA_signal_1288, new_AGEMA_signal_1287, SubCellInst_SboxInst_1_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U11 ( .a ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, SubCellInst_SboxInst_1_n4}), .clk (clk), .r ({Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_1580, new_AGEMA_signal_1579, SubCellInst_SboxInst_1_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U6 ( .a ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, SubCellInst_SboxInst_1_n7}), .b ({new_AGEMA_signal_1044, new_AGEMA_signal_1043, SubCellInst_SboxInst_1_n1}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309]}), .c ({new_AGEMA_signal_1296, new_AGEMA_signal_1295, SubCellInst_SboxInst_1_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U18 ( .a ({new_AGEMA_signal_1310, new_AGEMA_signal_1309, SubCellInst_SboxInst_2_n13}), .b ({ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r ({Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, SubCellInst_SboxInst_2_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U15 ( .a ({new_AGEMA_signal_1056, new_AGEMA_signal_1055, SubCellInst_SboxInst_2_n10}), .b ({new_AGEMA_signal_1066, new_AGEMA_signal_1065, SubCellInst_SboxInst_2_n9}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315]}), .c ({new_AGEMA_signal_1300, new_AGEMA_signal_1299, SubCellInst_SboxInst_2_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U11 ( .a ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .b ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, SubCellInst_SboxInst_2_n4}), .clk (clk), .r ({Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_1590, new_AGEMA_signal_1589, SubCellInst_SboxInst_2_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U6 ( .a ({new_AGEMA_signal_1062, new_AGEMA_signal_1061, SubCellInst_SboxInst_2_n7}), .b ({new_AGEMA_signal_1060, new_AGEMA_signal_1059, SubCellInst_SboxInst_2_n1}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321]}), .c ({new_AGEMA_signal_1308, new_AGEMA_signal_1307, SubCellInst_SboxInst_2_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U18 ( .a ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, SubCellInst_SboxInst_3_n13}), .b ({ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .clk (clk), .r ({Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_1596, new_AGEMA_signal_1595, SubCellInst_SboxInst_3_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U15 ( .a ({new_AGEMA_signal_1072, new_AGEMA_signal_1071, SubCellInst_SboxInst_3_n10}), .b ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, SubCellInst_SboxInst_3_n9}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327]}), .c ({new_AGEMA_signal_1312, new_AGEMA_signal_1311, SubCellInst_SboxInst_3_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U11 ( .a ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, SubCellInst_SboxInst_3_n4}), .clk (clk), .r ({Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_1600, new_AGEMA_signal_1599, SubCellInst_SboxInst_3_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U6 ( .a ({new_AGEMA_signal_1078, new_AGEMA_signal_1077, SubCellInst_SboxInst_3_n7}), .b ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, SubCellInst_SboxInst_3_n1}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333]}), .c ({new_AGEMA_signal_1320, new_AGEMA_signal_1319, SubCellInst_SboxInst_3_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U18 ( .a ({new_AGEMA_signal_1334, new_AGEMA_signal_1333, SubCellInst_SboxInst_4_n13}), .b ({ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .clk (clk), .r ({Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_1606, new_AGEMA_signal_1605, SubCellInst_SboxInst_4_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U15 ( .a ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, SubCellInst_SboxInst_4_n10}), .b ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, SubCellInst_SboxInst_4_n9}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339]}), .c ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, SubCellInst_SboxInst_4_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U11 ( .a ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, SubCellInst_SboxInst_4_n4}), .clk (clk), .r ({Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_1610, new_AGEMA_signal_1609, SubCellInst_SboxInst_4_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U6 ( .a ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, SubCellInst_SboxInst_4_n7}), .b ({new_AGEMA_signal_1092, new_AGEMA_signal_1091, SubCellInst_SboxInst_4_n1}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345]}), .c ({new_AGEMA_signal_1332, new_AGEMA_signal_1331, SubCellInst_SboxInst_4_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U18 ( .a ({new_AGEMA_signal_1346, new_AGEMA_signal_1345, SubCellInst_SboxInst_5_n13}), .b ({ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r ({Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_1616, new_AGEMA_signal_1615, SubCellInst_SboxInst_5_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U15 ( .a ({new_AGEMA_signal_1104, new_AGEMA_signal_1103, SubCellInst_SboxInst_5_n10}), .b ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, SubCellInst_SboxInst_5_n9}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351]}), .c ({new_AGEMA_signal_1336, new_AGEMA_signal_1335, SubCellInst_SboxInst_5_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U11 ( .a ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .b ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, SubCellInst_SboxInst_5_n4}), .clk (clk), .r ({Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_1620, new_AGEMA_signal_1619, SubCellInst_SboxInst_5_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U6 ( .a ({new_AGEMA_signal_1110, new_AGEMA_signal_1109, SubCellInst_SboxInst_5_n7}), .b ({new_AGEMA_signal_1108, new_AGEMA_signal_1107, SubCellInst_SboxInst_5_n1}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357]}), .c ({new_AGEMA_signal_1344, new_AGEMA_signal_1343, SubCellInst_SboxInst_5_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U18 ( .a ({new_AGEMA_signal_1358, new_AGEMA_signal_1357, SubCellInst_SboxInst_6_n13}), .b ({ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .clk (clk), .r ({Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_1626, new_AGEMA_signal_1625, SubCellInst_SboxInst_6_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U15 ( .a ({new_AGEMA_signal_1120, new_AGEMA_signal_1119, SubCellInst_SboxInst_6_n10}), .b ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, SubCellInst_SboxInst_6_n9}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363]}), .c ({new_AGEMA_signal_1348, new_AGEMA_signal_1347, SubCellInst_SboxInst_6_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U11 ( .a ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_1352, new_AGEMA_signal_1351, SubCellInst_SboxInst_6_n4}), .clk (clk), .r ({Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_1630, new_AGEMA_signal_1629, SubCellInst_SboxInst_6_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U6 ( .a ({new_AGEMA_signal_1126, new_AGEMA_signal_1125, SubCellInst_SboxInst_6_n7}), .b ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, SubCellInst_SboxInst_6_n1}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369]}), .c ({new_AGEMA_signal_1356, new_AGEMA_signal_1355, SubCellInst_SboxInst_6_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U18 ( .a ({new_AGEMA_signal_1370, new_AGEMA_signal_1369, SubCellInst_SboxInst_7_n13}), .b ({ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r ({Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_1636, new_AGEMA_signal_1635, SubCellInst_SboxInst_7_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U15 ( .a ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, SubCellInst_SboxInst_7_n10}), .b ({new_AGEMA_signal_1146, new_AGEMA_signal_1145, SubCellInst_SboxInst_7_n9}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375]}), .c ({new_AGEMA_signal_1360, new_AGEMA_signal_1359, SubCellInst_SboxInst_7_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U11 ( .a ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .b ({new_AGEMA_signal_1364, new_AGEMA_signal_1363, SubCellInst_SboxInst_7_n4}), .clk (clk), .r ({Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_1640, new_AGEMA_signal_1639, SubCellInst_SboxInst_7_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U6 ( .a ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, SubCellInst_SboxInst_7_n7}), .b ({new_AGEMA_signal_1140, new_AGEMA_signal_1139, SubCellInst_SboxInst_7_n1}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381]}), .c ({new_AGEMA_signal_1368, new_AGEMA_signal_1367, SubCellInst_SboxInst_7_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U18 ( .a ({new_AGEMA_signal_1382, new_AGEMA_signal_1381, SubCellInst_SboxInst_8_n13}), .b ({ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .clk (clk), .r ({Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_1646, new_AGEMA_signal_1645, SubCellInst_SboxInst_8_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U15 ( .a ({new_AGEMA_signal_1152, new_AGEMA_signal_1151, SubCellInst_SboxInst_8_n10}), .b ({new_AGEMA_signal_1162, new_AGEMA_signal_1161, SubCellInst_SboxInst_8_n9}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387]}), .c ({new_AGEMA_signal_1372, new_AGEMA_signal_1371, SubCellInst_SboxInst_8_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U11 ( .a ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_1376, new_AGEMA_signal_1375, SubCellInst_SboxInst_8_n4}), .clk (clk), .r ({Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_1650, new_AGEMA_signal_1649, SubCellInst_SboxInst_8_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U6 ( .a ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, SubCellInst_SboxInst_8_n7}), .b ({new_AGEMA_signal_1156, new_AGEMA_signal_1155, SubCellInst_SboxInst_8_n1}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393]}), .c ({new_AGEMA_signal_1380, new_AGEMA_signal_1379, SubCellInst_SboxInst_8_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U18 ( .a ({new_AGEMA_signal_1394, new_AGEMA_signal_1393, SubCellInst_SboxInst_9_n13}), .b ({ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r ({Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_1656, new_AGEMA_signal_1655, SubCellInst_SboxInst_9_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U15 ( .a ({new_AGEMA_signal_1168, new_AGEMA_signal_1167, SubCellInst_SboxInst_9_n10}), .b ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, SubCellInst_SboxInst_9_n9}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399]}), .c ({new_AGEMA_signal_1384, new_AGEMA_signal_1383, SubCellInst_SboxInst_9_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U11 ( .a ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_1388, new_AGEMA_signal_1387, SubCellInst_SboxInst_9_n4}), .clk (clk), .r ({Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_1660, new_AGEMA_signal_1659, SubCellInst_SboxInst_9_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U6 ( .a ({new_AGEMA_signal_1174, new_AGEMA_signal_1173, SubCellInst_SboxInst_9_n7}), .b ({new_AGEMA_signal_1172, new_AGEMA_signal_1171, SubCellInst_SboxInst_9_n1}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405]}), .c ({new_AGEMA_signal_1392, new_AGEMA_signal_1391, SubCellInst_SboxInst_9_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U18 ( .a ({new_AGEMA_signal_1406, new_AGEMA_signal_1405, SubCellInst_SboxInst_10_n13}), .b ({ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .clk (clk), .r ({Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_1666, new_AGEMA_signal_1665, SubCellInst_SboxInst_10_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U15 ( .a ({new_AGEMA_signal_1184, new_AGEMA_signal_1183, SubCellInst_SboxInst_10_n10}), .b ({new_AGEMA_signal_1194, new_AGEMA_signal_1193, SubCellInst_SboxInst_10_n9}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411]}), .c ({new_AGEMA_signal_1396, new_AGEMA_signal_1395, SubCellInst_SboxInst_10_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U11 ( .a ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_1400, new_AGEMA_signal_1399, SubCellInst_SboxInst_10_n4}), .clk (clk), .r ({Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_1670, new_AGEMA_signal_1669, SubCellInst_SboxInst_10_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U6 ( .a ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, SubCellInst_SboxInst_10_n7}), .b ({new_AGEMA_signal_1188, new_AGEMA_signal_1187, SubCellInst_SboxInst_10_n1}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417]}), .c ({new_AGEMA_signal_1404, new_AGEMA_signal_1403, SubCellInst_SboxInst_10_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U18 ( .a ({new_AGEMA_signal_1418, new_AGEMA_signal_1417, SubCellInst_SboxInst_11_n13}), .b ({ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r ({Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, SubCellInst_SboxInst_11_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U15 ( .a ({new_AGEMA_signal_1200, new_AGEMA_signal_1199, SubCellInst_SboxInst_11_n10}), .b ({new_AGEMA_signal_1210, new_AGEMA_signal_1209, SubCellInst_SboxInst_11_n9}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423]}), .c ({new_AGEMA_signal_1408, new_AGEMA_signal_1407, SubCellInst_SboxInst_11_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U11 ( .a ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .b ({new_AGEMA_signal_1412, new_AGEMA_signal_1411, SubCellInst_SboxInst_11_n4}), .clk (clk), .r ({Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_1680, new_AGEMA_signal_1679, SubCellInst_SboxInst_11_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U6 ( .a ({new_AGEMA_signal_1206, new_AGEMA_signal_1205, SubCellInst_SboxInst_11_n7}), .b ({new_AGEMA_signal_1204, new_AGEMA_signal_1203, SubCellInst_SboxInst_11_n1}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429]}), .c ({new_AGEMA_signal_1416, new_AGEMA_signal_1415, SubCellInst_SboxInst_11_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U18 ( .a ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, SubCellInst_SboxInst_12_n13}), .b ({ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r ({Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_1686, new_AGEMA_signal_1685, SubCellInst_SboxInst_12_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U15 ( .a ({new_AGEMA_signal_1216, new_AGEMA_signal_1215, SubCellInst_SboxInst_12_n10}), .b ({new_AGEMA_signal_1226, new_AGEMA_signal_1225, SubCellInst_SboxInst_12_n9}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435]}), .c ({new_AGEMA_signal_1420, new_AGEMA_signal_1419, SubCellInst_SboxInst_12_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U11 ( .a ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .b ({new_AGEMA_signal_1424, new_AGEMA_signal_1423, SubCellInst_SboxInst_12_n4}), .clk (clk), .r ({Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_1690, new_AGEMA_signal_1689, SubCellInst_SboxInst_12_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U6 ( .a ({new_AGEMA_signal_1222, new_AGEMA_signal_1221, SubCellInst_SboxInst_12_n7}), .b ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, SubCellInst_SboxInst_12_n1}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441]}), .c ({new_AGEMA_signal_1428, new_AGEMA_signal_1427, SubCellInst_SboxInst_12_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U18 ( .a ({new_AGEMA_signal_1442, new_AGEMA_signal_1441, SubCellInst_SboxInst_13_n13}), .b ({ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .clk (clk), .r ({Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_1696, new_AGEMA_signal_1695, SubCellInst_SboxInst_13_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U15 ( .a ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, SubCellInst_SboxInst_13_n10}), .b ({new_AGEMA_signal_1242, new_AGEMA_signal_1241, SubCellInst_SboxInst_13_n9}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447]}), .c ({new_AGEMA_signal_1432, new_AGEMA_signal_1431, SubCellInst_SboxInst_13_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U11 ( .a ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_1436, new_AGEMA_signal_1435, SubCellInst_SboxInst_13_n4}), .clk (clk), .r ({Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_1700, new_AGEMA_signal_1699, SubCellInst_SboxInst_13_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U6 ( .a ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, SubCellInst_SboxInst_13_n7}), .b ({new_AGEMA_signal_1236, new_AGEMA_signal_1235, SubCellInst_SboxInst_13_n1}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453]}), .c ({new_AGEMA_signal_1440, new_AGEMA_signal_1439, SubCellInst_SboxInst_13_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U18 ( .a ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, SubCellInst_SboxInst_14_n13}), .b ({ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r ({Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, SubCellInst_SboxInst_14_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U15 ( .a ({new_AGEMA_signal_1248, new_AGEMA_signal_1247, SubCellInst_SboxInst_14_n10}), .b ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_14_n9}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459]}), .c ({new_AGEMA_signal_1444, new_AGEMA_signal_1443, SubCellInst_SboxInst_14_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U11 ( .a ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .b ({new_AGEMA_signal_1448, new_AGEMA_signal_1447, SubCellInst_SboxInst_14_n4}), .clk (clk), .r ({Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_1710, new_AGEMA_signal_1709, SubCellInst_SboxInst_14_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U6 ( .a ({new_AGEMA_signal_1254, new_AGEMA_signal_1253, SubCellInst_SboxInst_14_n7}), .b ({new_AGEMA_signal_1252, new_AGEMA_signal_1251, SubCellInst_SboxInst_14_n1}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465]}), .c ({new_AGEMA_signal_1452, new_AGEMA_signal_1451, SubCellInst_SboxInst_14_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U18 ( .a ({new_AGEMA_signal_1466, new_AGEMA_signal_1465, SubCellInst_SboxInst_15_n13}), .b ({ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .clk (clk), .r ({Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_1716, new_AGEMA_signal_1715, SubCellInst_SboxInst_15_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U15 ( .a ({new_AGEMA_signal_1264, new_AGEMA_signal_1263, SubCellInst_SboxInst_15_n10}), .b ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, SubCellInst_SboxInst_15_n9}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471]}), .c ({new_AGEMA_signal_1456, new_AGEMA_signal_1455, SubCellInst_SboxInst_15_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U11 ( .a ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_1460, new_AGEMA_signal_1459, SubCellInst_SboxInst_15_n4}), .clk (clk), .r ({Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_1720, new_AGEMA_signal_1719, SubCellInst_SboxInst_15_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U6 ( .a ({new_AGEMA_signal_1270, new_AGEMA_signal_1269, SubCellInst_SboxInst_15_n7}), .b ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, SubCellInst_SboxInst_15_n1}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477]}), .c ({new_AGEMA_signal_1464, new_AGEMA_signal_1463, SubCellInst_SboxInst_15_n2}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_1_U1 ( .s (rst), .b ({new_AGEMA_signal_1728, new_AGEMA_signal_1727, Feedback[1]}), .a ({plaintext_s2[1], plaintext_s1[1], plaintext_s0[1]}), .c ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, MCOutput[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_3_U1 ( .s (rst), .b ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, Feedback[3]}), .a ({plaintext_s2[3], plaintext_s1[3], plaintext_s0[3]}), .c ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, MCOutput[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_5_U1 ( .s (rst), .b ({new_AGEMA_signal_1736, new_AGEMA_signal_1735, Feedback[5]}), .a ({plaintext_s2[5], plaintext_s1[5], plaintext_s0[5]}), .c ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, MCOutput[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_7_U1 ( .s (rst), .b ({new_AGEMA_signal_1732, new_AGEMA_signal_1731, Feedback[7]}), .a ({plaintext_s2[7], plaintext_s1[7], plaintext_s0[7]}), .c ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, MCOutput[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_9_U1 ( .s (rst), .b ({new_AGEMA_signal_1744, new_AGEMA_signal_1743, Feedback[9]}), .a ({plaintext_s2[9], plaintext_s1[9], plaintext_s0[9]}), .c ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, MCOutput[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_11_U1 ( .s (rst), .b ({new_AGEMA_signal_1740, new_AGEMA_signal_1739, Feedback[11]}), .a ({plaintext_s2[11], plaintext_s1[11], plaintext_s0[11]}), .c ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, MCOutput[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_13_U1 ( .s (rst), .b ({new_AGEMA_signal_1752, new_AGEMA_signal_1751, Feedback[13]}), .a ({plaintext_s2[13], plaintext_s1[13], plaintext_s0[13]}), .c ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, MCOutput[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_15_U1 ( .s (rst), .b ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, Feedback[15]}), .a ({plaintext_s2[15], plaintext_s1[15], plaintext_s0[15]}), .c ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, MCOutput[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_17_U1 ( .s (rst), .b ({new_AGEMA_signal_1760, new_AGEMA_signal_1759, Feedback[17]}), .a ({plaintext_s2[17], plaintext_s1[17], plaintext_s0[17]}), .c ({new_AGEMA_signal_2210, new_AGEMA_signal_2209, MCOutput[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_19_U1 ( .s (rst), .b ({new_AGEMA_signal_1756, new_AGEMA_signal_1755, Feedback[19]}), .a ({plaintext_s2[19], plaintext_s1[19], plaintext_s0[19]}), .c ({new_AGEMA_signal_2218, new_AGEMA_signal_2217, MCOutput[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_21_U1 ( .s (rst), .b ({new_AGEMA_signal_1768, new_AGEMA_signal_1767, Feedback[21]}), .a ({plaintext_s2[21], plaintext_s1[21], plaintext_s0[21]}), .c ({new_AGEMA_signal_2226, new_AGEMA_signal_2225, MCOutput[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_23_U1 ( .s (rst), .b ({new_AGEMA_signal_1764, new_AGEMA_signal_1763, Feedback[23]}), .a ({plaintext_s2[23], plaintext_s1[23], plaintext_s0[23]}), .c ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, MCOutput[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_25_U1 ( .s (rst), .b ({new_AGEMA_signal_1776, new_AGEMA_signal_1775, Feedback[25]}), .a ({plaintext_s2[25], plaintext_s1[25], plaintext_s0[25]}), .c ({new_AGEMA_signal_2242, new_AGEMA_signal_2241, MCOutput[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_27_U1 ( .s (rst), .b ({new_AGEMA_signal_1772, new_AGEMA_signal_1771, Feedback[27]}), .a ({plaintext_s2[27], plaintext_s1[27], plaintext_s0[27]}), .c ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, MCOutput[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_29_U1 ( .s (rst), .b ({new_AGEMA_signal_1784, new_AGEMA_signal_1783, Feedback[29]}), .a ({plaintext_s2[29], plaintext_s1[29], plaintext_s0[29]}), .c ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, MCOutput[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_31_U1 ( .s (rst), .b ({new_AGEMA_signal_1780, new_AGEMA_signal_1779, Feedback[31]}), .a ({plaintext_s2[31], plaintext_s1[31], plaintext_s0[31]}), .c ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, MCOutput[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_33_U1 ( .s (rst), .b ({new_AGEMA_signal_1792, new_AGEMA_signal_1791, Feedback[33]}), .a ({plaintext_s2[33], plaintext_s1[33], plaintext_s0[33]}), .c ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, MCInput[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_35_U1 ( .s (rst), .b ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, Feedback[35]}), .a ({plaintext_s2[35], plaintext_s1[35], plaintext_s0[35]}), .c ({new_AGEMA_signal_2282, new_AGEMA_signal_2281, MCInput[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_37_U1 ( .s (rst), .b ({new_AGEMA_signal_1800, new_AGEMA_signal_1799, Feedback[37]}), .a ({plaintext_s2[37], plaintext_s1[37], plaintext_s0[37]}), .c ({new_AGEMA_signal_2290, new_AGEMA_signal_2289, MCInput[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_39_U1 ( .s (rst), .b ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, Feedback[39]}), .a ({plaintext_s2[39], plaintext_s1[39], plaintext_s0[39]}), .c ({new_AGEMA_signal_2298, new_AGEMA_signal_2297, MCInput[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_41_U1 ( .s (rst), .b ({new_AGEMA_signal_1808, new_AGEMA_signal_1807, Feedback[41]}), .a ({plaintext_s2[41], plaintext_s1[41], plaintext_s0[41]}), .c ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, MCInput[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_43_U1 ( .s (rst), .b ({new_AGEMA_signal_1804, new_AGEMA_signal_1803, Feedback[43]}), .a ({plaintext_s2[43], plaintext_s1[43], plaintext_s0[43]}), .c ({new_AGEMA_signal_2314, new_AGEMA_signal_2313, MCInput[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_45_U1 ( .s (rst), .b ({new_AGEMA_signal_1816, new_AGEMA_signal_1815, Feedback[45]}), .a ({plaintext_s2[45], plaintext_s1[45], plaintext_s0[45]}), .c ({new_AGEMA_signal_2322, new_AGEMA_signal_2321, MCInput[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_47_U1 ( .s (rst), .b ({new_AGEMA_signal_1812, new_AGEMA_signal_1811, Feedback[47]}), .a ({plaintext_s2[47], plaintext_s1[47], plaintext_s0[47]}), .c ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, MCInput[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_49_U1 ( .s (rst), .b ({new_AGEMA_signal_1824, new_AGEMA_signal_1823, Feedback[49]}), .a ({plaintext_s2[49], plaintext_s1[49], plaintext_s0[49]}), .c ({new_AGEMA_signal_2338, new_AGEMA_signal_2337, MCInput[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_51_U1 ( .s (rst), .b ({new_AGEMA_signal_1820, new_AGEMA_signal_1819, Feedback[51]}), .a ({plaintext_s2[51], plaintext_s1[51], plaintext_s0[51]}), .c ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, MCInput[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_53_U1 ( .s (rst), .b ({new_AGEMA_signal_1832, new_AGEMA_signal_1831, Feedback[53]}), .a ({plaintext_s2[53], plaintext_s1[53], plaintext_s0[53]}), .c ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, MCInput[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_55_U1 ( .s (rst), .b ({new_AGEMA_signal_1828, new_AGEMA_signal_1827, Feedback[55]}), .a ({plaintext_s2[55], plaintext_s1[55], plaintext_s0[55]}), .c ({new_AGEMA_signal_2362, new_AGEMA_signal_2361, MCInput[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_57_U1 ( .s (rst), .b ({new_AGEMA_signal_1840, new_AGEMA_signal_1839, Feedback[57]}), .a ({plaintext_s2[57], plaintext_s1[57], plaintext_s0[57]}), .c ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, MCInput[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_59_U1 ( .s (rst), .b ({new_AGEMA_signal_1836, new_AGEMA_signal_1835, Feedback[59]}), .a ({plaintext_s2[59], plaintext_s1[59], plaintext_s0[59]}), .c ({new_AGEMA_signal_2378, new_AGEMA_signal_2377, MCInput[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_61_U1 ( .s (rst), .b ({new_AGEMA_signal_1848, new_AGEMA_signal_1847, Feedback[61]}), .a ({plaintext_s2[61], plaintext_s1[61], plaintext_s0[61]}), .c ({new_AGEMA_signal_2386, new_AGEMA_signal_2385, MCInput[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_63_U1 ( .s (rst), .b ({new_AGEMA_signal_1844, new_AGEMA_signal_1843, Feedback[63]}), .a ({plaintext_s2[63], plaintext_s1[63], plaintext_s0[63]}), .c ({new_AGEMA_signal_2394, new_AGEMA_signal_2393, MCInput[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_1_U3 ( .a ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, MCInst_XOR_r0_Inst_1_n2}), .b ({new_AGEMA_signal_2418, new_AGEMA_signal_2417, MCInst_XOR_r0_Inst_1_n1}), .c ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, MCOutput[49]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_1_U2 ( .a ({new_AGEMA_signal_2210, new_AGEMA_signal_2209, MCOutput[17]}), .b ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, MCOutput[1]}), .c ({new_AGEMA_signal_2418, new_AGEMA_signal_2417, MCInst_XOR_r0_Inst_1_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2338, new_AGEMA_signal_2337, MCInput[49]}), .c ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, MCInst_XOR_r0_Inst_1_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_1_U2 ( .a ({new_AGEMA_signal_2422, new_AGEMA_signal_2421, MCInst_XOR_r1_Inst_1_n1}), .b ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, MCOutput[1]}), .c ({new_AGEMA_signal_2578, new_AGEMA_signal_2577, MCOutput[33]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, MCInput[33]}), .c ({new_AGEMA_signal_2422, new_AGEMA_signal_2421, MCInst_XOR_r1_Inst_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_3_U3 ( .a ({new_AGEMA_signal_2432, new_AGEMA_signal_2431, MCInst_XOR_r0_Inst_3_n2}), .b ({new_AGEMA_signal_2430, new_AGEMA_signal_2429, MCInst_XOR_r0_Inst_3_n1}), .c ({new_AGEMA_signal_2584, new_AGEMA_signal_2583, MCOutput[51]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_3_U2 ( .a ({new_AGEMA_signal_2218, new_AGEMA_signal_2217, MCOutput[19]}), .b ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, MCOutput[3]}), .c ({new_AGEMA_signal_2430, new_AGEMA_signal_2429, MCInst_XOR_r0_Inst_3_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, MCInput[51]}), .c ({new_AGEMA_signal_2432, new_AGEMA_signal_2431, MCInst_XOR_r0_Inst_3_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_3_U2 ( .a ({new_AGEMA_signal_2434, new_AGEMA_signal_2433, MCInst_XOR_r1_Inst_3_n1}), .b ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, MCOutput[3]}), .c ({new_AGEMA_signal_2586, new_AGEMA_signal_2585, MCOutput[35]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2282, new_AGEMA_signal_2281, MCInput[35]}), .c ({new_AGEMA_signal_2434, new_AGEMA_signal_2433, MCInst_XOR_r1_Inst_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_5_U3 ( .a ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, MCInst_XOR_r0_Inst_5_n2}), .b ({new_AGEMA_signal_2442, new_AGEMA_signal_2441, MCInst_XOR_r0_Inst_5_n1}), .c ({new_AGEMA_signal_2592, new_AGEMA_signal_2591, MCOutput[53]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_5_U2 ( .a ({new_AGEMA_signal_2226, new_AGEMA_signal_2225, MCOutput[21]}), .b ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, MCOutput[5]}), .c ({new_AGEMA_signal_2442, new_AGEMA_signal_2441, MCInst_XOR_r0_Inst_5_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_5_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, MCInput[53]}), .c ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, MCInst_XOR_r0_Inst_5_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_5_U2 ( .a ({new_AGEMA_signal_2446, new_AGEMA_signal_2445, MCInst_XOR_r1_Inst_5_n1}), .b ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, MCOutput[5]}), .c ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, MCOutput[37]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_5_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2290, new_AGEMA_signal_2289, MCInput[37]}), .c ({new_AGEMA_signal_2446, new_AGEMA_signal_2445, MCInst_XOR_r1_Inst_5_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_7_U3 ( .a ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, MCInst_XOR_r0_Inst_7_n2}), .b ({new_AGEMA_signal_2454, new_AGEMA_signal_2453, MCInst_XOR_r0_Inst_7_n1}), .c ({new_AGEMA_signal_2600, new_AGEMA_signal_2599, MCOutput[55]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_7_U2 ( .a ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, MCOutput[23]}), .b ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, MCOutput[7]}), .c ({new_AGEMA_signal_2454, new_AGEMA_signal_2453, MCInst_XOR_r0_Inst_7_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_7_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2362, new_AGEMA_signal_2361, MCInput[55]}), .c ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, MCInst_XOR_r0_Inst_7_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_7_U2 ( .a ({new_AGEMA_signal_2458, new_AGEMA_signal_2457, MCInst_XOR_r1_Inst_7_n1}), .b ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, MCOutput[7]}), .c ({new_AGEMA_signal_2602, new_AGEMA_signal_2601, MCOutput[39]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_7_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2298, new_AGEMA_signal_2297, MCInput[39]}), .c ({new_AGEMA_signal_2458, new_AGEMA_signal_2457, MCInst_XOR_r1_Inst_7_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_9_U3 ( .a ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, MCInst_XOR_r0_Inst_9_n2}), .b ({new_AGEMA_signal_2466, new_AGEMA_signal_2465, MCInst_XOR_r0_Inst_9_n1}), .c ({new_AGEMA_signal_2608, new_AGEMA_signal_2607, MCOutput[57]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_9_U2 ( .a ({new_AGEMA_signal_2242, new_AGEMA_signal_2241, MCOutput[25]}), .b ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, MCOutput[9]}), .c ({new_AGEMA_signal_2466, new_AGEMA_signal_2465, MCInst_XOR_r0_Inst_9_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_9_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, MCInput[57]}), .c ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, MCInst_XOR_r0_Inst_9_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_9_U2 ( .a ({new_AGEMA_signal_2470, new_AGEMA_signal_2469, MCInst_XOR_r1_Inst_9_n1}), .b ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, MCOutput[9]}), .c ({new_AGEMA_signal_2610, new_AGEMA_signal_2609, MCOutput[41]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_9_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, MCInput[41]}), .c ({new_AGEMA_signal_2470, new_AGEMA_signal_2469, MCInst_XOR_r1_Inst_9_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_11_U3 ( .a ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, MCInst_XOR_r0_Inst_11_n2}), .b ({new_AGEMA_signal_2478, new_AGEMA_signal_2477, MCInst_XOR_r0_Inst_11_n1}), .c ({new_AGEMA_signal_2616, new_AGEMA_signal_2615, MCOutput[59]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_11_U2 ( .a ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, MCOutput[27]}), .b ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, MCOutput[11]}), .c ({new_AGEMA_signal_2478, new_AGEMA_signal_2477, MCInst_XOR_r0_Inst_11_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_11_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2378, new_AGEMA_signal_2377, MCInput[59]}), .c ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, MCInst_XOR_r0_Inst_11_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_11_U2 ( .a ({new_AGEMA_signal_2482, new_AGEMA_signal_2481, MCInst_XOR_r1_Inst_11_n1}), .b ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, MCOutput[11]}), .c ({new_AGEMA_signal_2618, new_AGEMA_signal_2617, MCOutput[43]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_11_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2314, new_AGEMA_signal_2313, MCInput[43]}), .c ({new_AGEMA_signal_2482, new_AGEMA_signal_2481, MCInst_XOR_r1_Inst_11_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_13_U3 ( .a ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, MCInst_XOR_r0_Inst_13_n2}), .b ({new_AGEMA_signal_2490, new_AGEMA_signal_2489, MCInst_XOR_r0_Inst_13_n1}), .c ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, MCOutput[61]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_13_U2 ( .a ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, MCOutput[29]}), .b ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, MCOutput[13]}), .c ({new_AGEMA_signal_2490, new_AGEMA_signal_2489, MCInst_XOR_r0_Inst_13_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_13_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2386, new_AGEMA_signal_2385, MCInput[61]}), .c ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, MCInst_XOR_r0_Inst_13_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_13_U2 ( .a ({new_AGEMA_signal_2494, new_AGEMA_signal_2493, MCInst_XOR_r1_Inst_13_n1}), .b ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, MCOutput[13]}), .c ({new_AGEMA_signal_2626, new_AGEMA_signal_2625, MCOutput[45]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_13_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2322, new_AGEMA_signal_2321, MCInput[45]}), .c ({new_AGEMA_signal_2494, new_AGEMA_signal_2493, MCInst_XOR_r1_Inst_13_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_15_U3 ( .a ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, MCInst_XOR_r0_Inst_15_n2}), .b ({new_AGEMA_signal_2502, new_AGEMA_signal_2501, MCInst_XOR_r0_Inst_15_n1}), .c ({new_AGEMA_signal_2632, new_AGEMA_signal_2631, MCOutput[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_15_U2 ( .a ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, MCOutput[31]}), .b ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, MCOutput[15]}), .c ({new_AGEMA_signal_2502, new_AGEMA_signal_2501, MCInst_XOR_r0_Inst_15_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_15_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2394, new_AGEMA_signal_2393, MCInput[63]}), .c ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, MCInst_XOR_r0_Inst_15_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_15_U2 ( .a ({new_AGEMA_signal_2506, new_AGEMA_signal_2505, MCInst_XOR_r1_Inst_15_n1}), .b ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, MCOutput[15]}), .c ({new_AGEMA_signal_2634, new_AGEMA_signal_2633, MCOutput[47]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_15_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, MCInput[47]}), .c ({new_AGEMA_signal_2506, new_AGEMA_signal_2505, MCInst_XOR_r1_Inst_15_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2702, new_AGEMA_signal_2701, AddKeyXOR1_XORInst_0_1_n1}), .b ({new_AGEMA_signal_2084, new_AGEMA_signal_2083, SelectedKey[49]}), .c ({new_AGEMA_signal_2766, new_AGEMA_signal_2765, AddRoundKeyOutput[49]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, MCOutput[49]}), .c ({new_AGEMA_signal_2702, new_AGEMA_signal_2701, AddKeyXOR1_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2706, new_AGEMA_signal_2705, AddKeyXOR1_XORInst_0_3_n1}), .b ({new_AGEMA_signal_2096, new_AGEMA_signal_2095, SelectedKey[51]}), .c ({new_AGEMA_signal_2770, new_AGEMA_signal_2769, AddRoundKeyOutput[51]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2584, new_AGEMA_signal_2583, MCOutput[51]}), .c ({new_AGEMA_signal_2706, new_AGEMA_signal_2705, AddKeyXOR1_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, AddKeyXOR1_XORInst_1_1_n1}), .b ({new_AGEMA_signal_1538, new_AGEMA_signal_1537, SelectedKey[53]}), .c ({new_AGEMA_signal_2774, new_AGEMA_signal_2773, AddRoundKeyOutput[53]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2592, new_AGEMA_signal_2591, MCOutput[53]}), .c ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, AddKeyXOR1_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, AddKeyXOR1_XORInst_1_3_n1}), .b ({new_AGEMA_signal_2108, new_AGEMA_signal_2107, SelectedKey[55]}), .c ({new_AGEMA_signal_2778, new_AGEMA_signal_2777, AddRoundKeyOutput[55]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2600, new_AGEMA_signal_2599, MCOutput[55]}), .c ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, AddKeyXOR1_XORInst_1_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_2718, new_AGEMA_signal_2717, AddKeyXOR1_XORInst_2_1_n1}), .b ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, SelectedKey[57]}), .c ({new_AGEMA_signal_2782, new_AGEMA_signal_2781, AddRoundKeyOutput[57]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2608, new_AGEMA_signal_2607, MCOutput[57]}), .c ({new_AGEMA_signal_2718, new_AGEMA_signal_2717, AddKeyXOR1_XORInst_2_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_2722, new_AGEMA_signal_2721, AddKeyXOR1_XORInst_2_3_n1}), .b ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, SelectedKey[59]}), .c ({new_AGEMA_signal_2786, new_AGEMA_signal_2785, AddRoundKeyOutput[59]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2616, new_AGEMA_signal_2615, MCOutput[59]}), .c ({new_AGEMA_signal_2722, new_AGEMA_signal_2721, AddKeyXOR1_XORInst_2_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, AddKeyXOR1_XORInst_3_1_n1}), .b ({new_AGEMA_signal_2132, new_AGEMA_signal_2131, SelectedKey[61]}), .c ({new_AGEMA_signal_2790, new_AGEMA_signal_2789, AddRoundKeyOutput[61]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, MCOutput[61]}), .c ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, AddKeyXOR1_XORInst_3_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_2730, new_AGEMA_signal_2729, AddKeyXOR1_XORInst_3_3_n1}), .b ({new_AGEMA_signal_2138, new_AGEMA_signal_2137, SelectedKey[63]}), .c ({new_AGEMA_signal_2794, new_AGEMA_signal_2793, AddRoundKeyOutput[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2632, new_AGEMA_signal_2631, MCOutput[63]}), .c ({new_AGEMA_signal_2730, new_AGEMA_signal_2729, AddKeyXOR1_XORInst_3_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_0_1_U3 ( .a ({new_AGEMA_signal_2734, new_AGEMA_signal_2733, AddKeyConstXOR_XORInst_0_1_n2}), .b ({new_AGEMA_signal_2398, new_AGEMA_signal_2397, AddKeyConstXOR_XORInst_0_1_n1}), .c ({new_AGEMA_signal_2798, new_AGEMA_signal_2797, AddRoundKeyOutput[41]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2610, new_AGEMA_signal_2609, MCOutput[41]}), .c ({new_AGEMA_signal_2734, new_AGEMA_signal_2733, AddKeyConstXOR_XORInst_0_1_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_0_3_U3 ( .a ({new_AGEMA_signal_2738, new_AGEMA_signal_2737, AddKeyConstXOR_XORInst_0_3_n2}), .b ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, AddKeyConstXOR_XORInst_0_3_n1}), .c ({new_AGEMA_signal_2802, new_AGEMA_signal_2801, AddRoundKeyOutput[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2618, new_AGEMA_signal_2617, MCOutput[43]}), .c ({new_AGEMA_signal_2738, new_AGEMA_signal_2737, AddKeyConstXOR_XORInst_0_3_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_1_1_U3 ( .a ({new_AGEMA_signal_2742, new_AGEMA_signal_2741, AddKeyConstXOR_XORInst_1_1_n2}), .b ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, AddKeyConstXOR_XORInst_1_1_n1}), .c ({new_AGEMA_signal_2806, new_AGEMA_signal_2805, AddRoundKeyOutput[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2626, new_AGEMA_signal_2625, MCOutput[45]}), .c ({new_AGEMA_signal_2742, new_AGEMA_signal_2741, AddKeyConstXOR_XORInst_1_1_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_1_3_U3 ( .a ({new_AGEMA_signal_2746, new_AGEMA_signal_2745, AddKeyConstXOR_XORInst_1_3_n2}), .b ({new_AGEMA_signal_2410, new_AGEMA_signal_2409, AddKeyConstXOR_XORInst_1_3_n1}), .c ({new_AGEMA_signal_2810, new_AGEMA_signal_2809, AddRoundKeyOutput[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2634, new_AGEMA_signal_2633, MCOutput[47]}), .c ({new_AGEMA_signal_2746, new_AGEMA_signal_2745, AddKeyConstXOR_XORInst_1_3_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, AddKeyXOR2_XORInst_0_1_n1}), .b ({new_AGEMA_signal_1856, new_AGEMA_signal_1855, SelectedKey[1]}), .c ({new_AGEMA_signal_2638, new_AGEMA_signal_2637, AddRoundKeyOutput[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, MCOutput[1]}), .c ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, AddKeyXOR2_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2514, new_AGEMA_signal_2513, AddKeyXOR2_XORInst_0_3_n1}), .b ({new_AGEMA_signal_1862, new_AGEMA_signal_1861, SelectedKey[3]}), .c ({new_AGEMA_signal_2642, new_AGEMA_signal_2641, AddRoundKeyOutput[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, MCOutput[3]}), .c ({new_AGEMA_signal_2514, new_AGEMA_signal_2513, AddKeyXOR2_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2518, new_AGEMA_signal_2517, AddKeyXOR2_XORInst_1_1_n1}), .b ({new_AGEMA_signal_1874, new_AGEMA_signal_1873, SelectedKey[5]}), .c ({new_AGEMA_signal_2646, new_AGEMA_signal_2645, AddRoundKeyOutput[5]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, MCOutput[5]}), .c ({new_AGEMA_signal_2518, new_AGEMA_signal_2517, AddKeyXOR2_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, AddKeyXOR2_XORInst_1_3_n1}), .b ({new_AGEMA_signal_1886, new_AGEMA_signal_1885, SelectedKey[7]}), .c ({new_AGEMA_signal_2650, new_AGEMA_signal_2649, AddRoundKeyOutput[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, MCOutput[7]}), .c ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, AddKeyXOR2_XORInst_1_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_2526, new_AGEMA_signal_2525, AddKeyXOR2_XORInst_2_1_n1}), .b ({new_AGEMA_signal_1898, new_AGEMA_signal_1897, SelectedKey[9]}), .c ({new_AGEMA_signal_2654, new_AGEMA_signal_2653, AddRoundKeyOutput[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, MCOutput[9]}), .c ({new_AGEMA_signal_2526, new_AGEMA_signal_2525, AddKeyXOR2_XORInst_2_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_2530, new_AGEMA_signal_2529, AddKeyXOR2_XORInst_2_3_n1}), .b ({new_AGEMA_signal_1910, new_AGEMA_signal_1909, SelectedKey[11]}), .c ({new_AGEMA_signal_2658, new_AGEMA_signal_2657, AddRoundKeyOutput[11]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, MCOutput[11]}), .c ({new_AGEMA_signal_2530, new_AGEMA_signal_2529, AddKeyXOR2_XORInst_2_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, AddKeyXOR2_XORInst_3_1_n1}), .b ({new_AGEMA_signal_1922, new_AGEMA_signal_1921, SelectedKey[13]}), .c ({new_AGEMA_signal_2662, new_AGEMA_signal_2661, AddRoundKeyOutput[13]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, MCOutput[13]}), .c ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, AddKeyXOR2_XORInst_3_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_2538, new_AGEMA_signal_2537, AddKeyXOR2_XORInst_3_3_n1}), .b ({new_AGEMA_signal_1934, new_AGEMA_signal_1933, SelectedKey[15]}), .c ({new_AGEMA_signal_2666, new_AGEMA_signal_2665, AddRoundKeyOutput[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, MCOutput[15]}), .c ({new_AGEMA_signal_2538, new_AGEMA_signal_2537, AddKeyXOR2_XORInst_3_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_4_1_U2 ( .a ({new_AGEMA_signal_2542, new_AGEMA_signal_2541, AddKeyXOR2_XORInst_4_1_n1}), .b ({new_AGEMA_signal_1946, new_AGEMA_signal_1945, SelectedKey[17]}), .c ({new_AGEMA_signal_2670, new_AGEMA_signal_2669, AddRoundKeyOutput[17]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_4_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2210, new_AGEMA_signal_2209, MCOutput[17]}), .c ({new_AGEMA_signal_2542, new_AGEMA_signal_2541, AddKeyXOR2_XORInst_4_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_4_3_U2 ( .a ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, AddKeyXOR2_XORInst_4_3_n1}), .b ({new_AGEMA_signal_1958, new_AGEMA_signal_1957, SelectedKey[19]}), .c ({new_AGEMA_signal_2674, new_AGEMA_signal_2673, AddRoundKeyOutput[19]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_4_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2218, new_AGEMA_signal_2217, MCOutput[19]}), .c ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, AddKeyXOR2_XORInst_4_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_5_1_U2 ( .a ({new_AGEMA_signal_2550, new_AGEMA_signal_2549, AddKeyXOR2_XORInst_5_1_n1}), .b ({new_AGEMA_signal_1970, new_AGEMA_signal_1969, SelectedKey[21]}), .c ({new_AGEMA_signal_2678, new_AGEMA_signal_2677, AddRoundKeyOutput[21]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_5_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2226, new_AGEMA_signal_2225, MCOutput[21]}), .c ({new_AGEMA_signal_2550, new_AGEMA_signal_2549, AddKeyXOR2_XORInst_5_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_5_3_U2 ( .a ({new_AGEMA_signal_2554, new_AGEMA_signal_2553, AddKeyXOR2_XORInst_5_3_n1}), .b ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, SelectedKey[23]}), .c ({new_AGEMA_signal_2682, new_AGEMA_signal_2681, AddRoundKeyOutput[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_5_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, MCOutput[23]}), .c ({new_AGEMA_signal_2554, new_AGEMA_signal_2553, AddKeyXOR2_XORInst_5_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_6_1_U2 ( .a ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, AddKeyXOR2_XORInst_6_1_n1}), .b ({new_AGEMA_signal_1502, new_AGEMA_signal_1501, SelectedKey[25]}), .c ({new_AGEMA_signal_2686, new_AGEMA_signal_2685, AddRoundKeyOutput[25]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_6_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2242, new_AGEMA_signal_2241, MCOutput[25]}), .c ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, AddKeyXOR2_XORInst_6_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_6_3_U2 ( .a ({new_AGEMA_signal_2562, new_AGEMA_signal_2561, AddKeyXOR2_XORInst_6_3_n1}), .b ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, SelectedKey[27]}), .c ({new_AGEMA_signal_2690, new_AGEMA_signal_2689, AddRoundKeyOutput[27]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_6_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, MCOutput[27]}), .c ({new_AGEMA_signal_2562, new_AGEMA_signal_2561, AddKeyXOR2_XORInst_6_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_7_1_U2 ( .a ({new_AGEMA_signal_2566, new_AGEMA_signal_2565, AddKeyXOR2_XORInst_7_1_n1}), .b ({new_AGEMA_signal_1982, new_AGEMA_signal_1981, SelectedKey[29]}), .c ({new_AGEMA_signal_2694, new_AGEMA_signal_2693, AddRoundKeyOutput[29]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_7_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, MCOutput[29]}), .c ({new_AGEMA_signal_2566, new_AGEMA_signal_2565, AddKeyXOR2_XORInst_7_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_7_3_U2 ( .a ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, AddKeyXOR2_XORInst_7_3_n1}), .b ({new_AGEMA_signal_1994, new_AGEMA_signal_1993, SelectedKey[31]}), .c ({new_AGEMA_signal_2698, new_AGEMA_signal_2697, AddRoundKeyOutput[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_7_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, MCOutput[31]}), .c ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, AddKeyXOR2_XORInst_7_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_8_1_U2 ( .a ({new_AGEMA_signal_2750, new_AGEMA_signal_2749, AddKeyXOR2_XORInst_8_1_n1}), .b ({new_AGEMA_signal_1520, new_AGEMA_signal_1519, SelectedKey[33]}), .c ({new_AGEMA_signal_2814, new_AGEMA_signal_2813, AddRoundKeyOutput[33]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_8_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2578, new_AGEMA_signal_2577, MCOutput[33]}), .c ({new_AGEMA_signal_2750, new_AGEMA_signal_2749, AddKeyXOR2_XORInst_8_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_8_3_U2 ( .a ({new_AGEMA_signal_2754, new_AGEMA_signal_2753, AddKeyXOR2_XORInst_8_3_n1}), .b ({new_AGEMA_signal_2012, new_AGEMA_signal_2011, SelectedKey[35]}), .c ({new_AGEMA_signal_2818, new_AGEMA_signal_2817, AddRoundKeyOutput[35]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_8_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2586, new_AGEMA_signal_2585, MCOutput[35]}), .c ({new_AGEMA_signal_2754, new_AGEMA_signal_2753, AddKeyXOR2_XORInst_8_3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_9_1_U2 ( .a ({new_AGEMA_signal_2758, new_AGEMA_signal_2757, AddKeyXOR2_XORInst_9_1_n1}), .b ({new_AGEMA_signal_2018, new_AGEMA_signal_2017, SelectedKey[37]}), .c ({new_AGEMA_signal_2822, new_AGEMA_signal_2821, AddRoundKeyOutput[37]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_9_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, MCOutput[37]}), .c ({new_AGEMA_signal_2758, new_AGEMA_signal_2757, AddKeyXOR2_XORInst_9_1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_9_3_U2 ( .a ({new_AGEMA_signal_2762, new_AGEMA_signal_2761, AddKeyXOR2_XORInst_9_3_n1}), .b ({new_AGEMA_signal_1532, new_AGEMA_signal_1531, SelectedKey[39]}), .c ({new_AGEMA_signal_2826, new_AGEMA_signal_2825, AddRoundKeyOutput[39]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_9_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2602, new_AGEMA_signal_2601, MCOutput[39]}), .c ({new_AGEMA_signal_2762, new_AGEMA_signal_2761, AddKeyXOR2_XORInst_9_3_n1}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U19 ( .a ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, SubCellInst_SboxInst_0_n15}), .b ({new_AGEMA_signal_1566, new_AGEMA_signal_1565, SubCellInst_SboxInst_0_n14}), .clk (clk), .r ({Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, Feedback[3]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U16 ( .a ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_0_n11}), .b ({ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483]}), .c ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, SubCellInst_SboxInst_0_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U12 ( .a ({new_AGEMA_signal_1282, new_AGEMA_signal_1281, SubCellInst_SboxInst_0_n6}), .b ({new_AGEMA_signal_1570, new_AGEMA_signal_1569, SubCellInst_SboxInst_0_n5}), .clk (clk), .r ({Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_1728, new_AGEMA_signal_1727, Feedback[1]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U7 ( .a ({ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .b ({new_AGEMA_signal_1284, new_AGEMA_signal_1283, SubCellInst_SboxInst_0_n2}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489]}), .c ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, SubCellInst_SboxInst_0_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U19 ( .a ({new_AGEMA_signal_1290, new_AGEMA_signal_1289, SubCellInst_SboxInst_1_n15}), .b ({new_AGEMA_signal_1576, new_AGEMA_signal_1575, SubCellInst_SboxInst_1_n14}), .clk (clk), .r ({Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_1732, new_AGEMA_signal_1731, Feedback[7]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U16 ( .a ({new_AGEMA_signal_1288, new_AGEMA_signal_1287, SubCellInst_SboxInst_1_n11}), .b ({ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495]}), .c ({new_AGEMA_signal_1578, new_AGEMA_signal_1577, SubCellInst_SboxInst_1_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U12 ( .a ({new_AGEMA_signal_1294, new_AGEMA_signal_1293, SubCellInst_SboxInst_1_n6}), .b ({new_AGEMA_signal_1580, new_AGEMA_signal_1579, SubCellInst_SboxInst_1_n5}), .clk (clk), .r ({Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_1736, new_AGEMA_signal_1735, Feedback[5]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U7 ( .a ({ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .b ({new_AGEMA_signal_1296, new_AGEMA_signal_1295, SubCellInst_SboxInst_1_n2}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501]}), .c ({new_AGEMA_signal_1582, new_AGEMA_signal_1581, SubCellInst_SboxInst_1_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U19 ( .a ({new_AGEMA_signal_1302, new_AGEMA_signal_1301, SubCellInst_SboxInst_2_n15}), .b ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, SubCellInst_SboxInst_2_n14}), .clk (clk), .r ({Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_1740, new_AGEMA_signal_1739, Feedback[11]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U16 ( .a ({new_AGEMA_signal_1300, new_AGEMA_signal_1299, SubCellInst_SboxInst_2_n11}), .b ({ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507]}), .c ({new_AGEMA_signal_1588, new_AGEMA_signal_1587, SubCellInst_SboxInst_2_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U12 ( .a ({new_AGEMA_signal_1306, new_AGEMA_signal_1305, SubCellInst_SboxInst_2_n6}), .b ({new_AGEMA_signal_1590, new_AGEMA_signal_1589, SubCellInst_SboxInst_2_n5}), .clk (clk), .r ({Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_1744, new_AGEMA_signal_1743, Feedback[9]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U7 ( .a ({ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .b ({new_AGEMA_signal_1308, new_AGEMA_signal_1307, SubCellInst_SboxInst_2_n2}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513]}), .c ({new_AGEMA_signal_1592, new_AGEMA_signal_1591, SubCellInst_SboxInst_2_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U19 ( .a ({new_AGEMA_signal_1314, new_AGEMA_signal_1313, SubCellInst_SboxInst_3_n15}), .b ({new_AGEMA_signal_1596, new_AGEMA_signal_1595, SubCellInst_SboxInst_3_n14}), .clk (clk), .r ({Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, Feedback[15]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U16 ( .a ({new_AGEMA_signal_1312, new_AGEMA_signal_1311, SubCellInst_SboxInst_3_n11}), .b ({ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519]}), .c ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, SubCellInst_SboxInst_3_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U12 ( .a ({new_AGEMA_signal_1318, new_AGEMA_signal_1317, SubCellInst_SboxInst_3_n6}), .b ({new_AGEMA_signal_1600, new_AGEMA_signal_1599, SubCellInst_SboxInst_3_n5}), .clk (clk), .r ({Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_1752, new_AGEMA_signal_1751, Feedback[13]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U7 ( .a ({ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .b ({new_AGEMA_signal_1320, new_AGEMA_signal_1319, SubCellInst_SboxInst_3_n2}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525]}), .c ({new_AGEMA_signal_1602, new_AGEMA_signal_1601, SubCellInst_SboxInst_3_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U19 ( .a ({new_AGEMA_signal_1326, new_AGEMA_signal_1325, SubCellInst_SboxInst_4_n15}), .b ({new_AGEMA_signal_1606, new_AGEMA_signal_1605, SubCellInst_SboxInst_4_n14}), .clk (clk), .r ({Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_1756, new_AGEMA_signal_1755, Feedback[19]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U16 ( .a ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, SubCellInst_SboxInst_4_n11}), .b ({ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531]}), .c ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, SubCellInst_SboxInst_4_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U12 ( .a ({new_AGEMA_signal_1330, new_AGEMA_signal_1329, SubCellInst_SboxInst_4_n6}), .b ({new_AGEMA_signal_1610, new_AGEMA_signal_1609, SubCellInst_SboxInst_4_n5}), .clk (clk), .r ({Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_1760, new_AGEMA_signal_1759, Feedback[17]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U7 ( .a ({ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .b ({new_AGEMA_signal_1332, new_AGEMA_signal_1331, SubCellInst_SboxInst_4_n2}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537]}), .c ({new_AGEMA_signal_1612, new_AGEMA_signal_1611, SubCellInst_SboxInst_4_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U19 ( .a ({new_AGEMA_signal_1338, new_AGEMA_signal_1337, SubCellInst_SboxInst_5_n15}), .b ({new_AGEMA_signal_1616, new_AGEMA_signal_1615, SubCellInst_SboxInst_5_n14}), .clk (clk), .r ({Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_1764, new_AGEMA_signal_1763, Feedback[23]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U16 ( .a ({new_AGEMA_signal_1336, new_AGEMA_signal_1335, SubCellInst_SboxInst_5_n11}), .b ({ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543]}), .c ({new_AGEMA_signal_1618, new_AGEMA_signal_1617, SubCellInst_SboxInst_5_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U12 ( .a ({new_AGEMA_signal_1342, new_AGEMA_signal_1341, SubCellInst_SboxInst_5_n6}), .b ({new_AGEMA_signal_1620, new_AGEMA_signal_1619, SubCellInst_SboxInst_5_n5}), .clk (clk), .r ({Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_1768, new_AGEMA_signal_1767, Feedback[21]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U7 ( .a ({ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .b ({new_AGEMA_signal_1344, new_AGEMA_signal_1343, SubCellInst_SboxInst_5_n2}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549]}), .c ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, SubCellInst_SboxInst_5_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U19 ( .a ({new_AGEMA_signal_1350, new_AGEMA_signal_1349, SubCellInst_SboxInst_6_n15}), .b ({new_AGEMA_signal_1626, new_AGEMA_signal_1625, SubCellInst_SboxInst_6_n14}), .clk (clk), .r ({Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_1772, new_AGEMA_signal_1771, Feedback[27]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U16 ( .a ({new_AGEMA_signal_1348, new_AGEMA_signal_1347, SubCellInst_SboxInst_6_n11}), .b ({ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555]}), .c ({new_AGEMA_signal_1628, new_AGEMA_signal_1627, SubCellInst_SboxInst_6_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U12 ( .a ({new_AGEMA_signal_1354, new_AGEMA_signal_1353, SubCellInst_SboxInst_6_n6}), .b ({new_AGEMA_signal_1630, new_AGEMA_signal_1629, SubCellInst_SboxInst_6_n5}), .clk (clk), .r ({Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_1776, new_AGEMA_signal_1775, Feedback[25]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U7 ( .a ({ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .b ({new_AGEMA_signal_1356, new_AGEMA_signal_1355, SubCellInst_SboxInst_6_n2}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561]}), .c ({new_AGEMA_signal_1632, new_AGEMA_signal_1631, SubCellInst_SboxInst_6_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U19 ( .a ({new_AGEMA_signal_1362, new_AGEMA_signal_1361, SubCellInst_SboxInst_7_n15}), .b ({new_AGEMA_signal_1636, new_AGEMA_signal_1635, SubCellInst_SboxInst_7_n14}), .clk (clk), .r ({Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_1780, new_AGEMA_signal_1779, Feedback[31]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U16 ( .a ({new_AGEMA_signal_1360, new_AGEMA_signal_1359, SubCellInst_SboxInst_7_n11}), .b ({ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567]}), .c ({new_AGEMA_signal_1638, new_AGEMA_signal_1637, SubCellInst_SboxInst_7_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U12 ( .a ({new_AGEMA_signal_1366, new_AGEMA_signal_1365, SubCellInst_SboxInst_7_n6}), .b ({new_AGEMA_signal_1640, new_AGEMA_signal_1639, SubCellInst_SboxInst_7_n5}), .clk (clk), .r ({Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_1784, new_AGEMA_signal_1783, Feedback[29]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U7 ( .a ({ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .b ({new_AGEMA_signal_1368, new_AGEMA_signal_1367, SubCellInst_SboxInst_7_n2}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573]}), .c ({new_AGEMA_signal_1642, new_AGEMA_signal_1641, SubCellInst_SboxInst_7_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U19 ( .a ({new_AGEMA_signal_1374, new_AGEMA_signal_1373, SubCellInst_SboxInst_8_n15}), .b ({new_AGEMA_signal_1646, new_AGEMA_signal_1645, SubCellInst_SboxInst_8_n14}), .clk (clk), .r ({Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, Feedback[35]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U16 ( .a ({new_AGEMA_signal_1372, new_AGEMA_signal_1371, SubCellInst_SboxInst_8_n11}), .b ({ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579]}), .c ({new_AGEMA_signal_1648, new_AGEMA_signal_1647, SubCellInst_SboxInst_8_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U12 ( .a ({new_AGEMA_signal_1378, new_AGEMA_signal_1377, SubCellInst_SboxInst_8_n6}), .b ({new_AGEMA_signal_1650, new_AGEMA_signal_1649, SubCellInst_SboxInst_8_n5}), .clk (clk), .r ({Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_1792, new_AGEMA_signal_1791, Feedback[33]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U7 ( .a ({ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .b ({new_AGEMA_signal_1380, new_AGEMA_signal_1379, SubCellInst_SboxInst_8_n2}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585]}), .c ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, SubCellInst_SboxInst_8_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U19 ( .a ({new_AGEMA_signal_1386, new_AGEMA_signal_1385, SubCellInst_SboxInst_9_n15}), .b ({new_AGEMA_signal_1656, new_AGEMA_signal_1655, SubCellInst_SboxInst_9_n14}), .clk (clk), .r ({Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, Feedback[39]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U16 ( .a ({new_AGEMA_signal_1384, new_AGEMA_signal_1383, SubCellInst_SboxInst_9_n11}), .b ({ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591]}), .c ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, SubCellInst_SboxInst_9_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U12 ( .a ({new_AGEMA_signal_1390, new_AGEMA_signal_1389, SubCellInst_SboxInst_9_n6}), .b ({new_AGEMA_signal_1660, new_AGEMA_signal_1659, SubCellInst_SboxInst_9_n5}), .clk (clk), .r ({Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_1800, new_AGEMA_signal_1799, Feedback[37]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U7 ( .a ({ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .b ({new_AGEMA_signal_1392, new_AGEMA_signal_1391, SubCellInst_SboxInst_9_n2}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597]}), .c ({new_AGEMA_signal_1662, new_AGEMA_signal_1661, SubCellInst_SboxInst_9_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U19 ( .a ({new_AGEMA_signal_1398, new_AGEMA_signal_1397, SubCellInst_SboxInst_10_n15}), .b ({new_AGEMA_signal_1666, new_AGEMA_signal_1665, SubCellInst_SboxInst_10_n14}), .clk (clk), .r ({Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_1804, new_AGEMA_signal_1803, Feedback[43]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U16 ( .a ({new_AGEMA_signal_1396, new_AGEMA_signal_1395, SubCellInst_SboxInst_10_n11}), .b ({ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603]}), .c ({new_AGEMA_signal_1668, new_AGEMA_signal_1667, SubCellInst_SboxInst_10_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U12 ( .a ({new_AGEMA_signal_1402, new_AGEMA_signal_1401, SubCellInst_SboxInst_10_n6}), .b ({new_AGEMA_signal_1670, new_AGEMA_signal_1669, SubCellInst_SboxInst_10_n5}), .clk (clk), .r ({Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_1808, new_AGEMA_signal_1807, Feedback[41]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U7 ( .a ({ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .b ({new_AGEMA_signal_1404, new_AGEMA_signal_1403, SubCellInst_SboxInst_10_n2}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609]}), .c ({new_AGEMA_signal_1672, new_AGEMA_signal_1671, SubCellInst_SboxInst_10_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U19 ( .a ({new_AGEMA_signal_1410, new_AGEMA_signal_1409, SubCellInst_SboxInst_11_n15}), .b ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, SubCellInst_SboxInst_11_n14}), .clk (clk), .r ({Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_1812, new_AGEMA_signal_1811, Feedback[47]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U16 ( .a ({new_AGEMA_signal_1408, new_AGEMA_signal_1407, SubCellInst_SboxInst_11_n11}), .b ({ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615]}), .c ({new_AGEMA_signal_1678, new_AGEMA_signal_1677, SubCellInst_SboxInst_11_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U12 ( .a ({new_AGEMA_signal_1414, new_AGEMA_signal_1413, SubCellInst_SboxInst_11_n6}), .b ({new_AGEMA_signal_1680, new_AGEMA_signal_1679, SubCellInst_SboxInst_11_n5}), .clk (clk), .r ({Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_1816, new_AGEMA_signal_1815, Feedback[45]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U7 ( .a ({ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .b ({new_AGEMA_signal_1416, new_AGEMA_signal_1415, SubCellInst_SboxInst_11_n2}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621]}), .c ({new_AGEMA_signal_1682, new_AGEMA_signal_1681, SubCellInst_SboxInst_11_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U19 ( .a ({new_AGEMA_signal_1422, new_AGEMA_signal_1421, SubCellInst_SboxInst_12_n15}), .b ({new_AGEMA_signal_1686, new_AGEMA_signal_1685, SubCellInst_SboxInst_12_n14}), .clk (clk), .r ({Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_1820, new_AGEMA_signal_1819, Feedback[51]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U16 ( .a ({new_AGEMA_signal_1420, new_AGEMA_signal_1419, SubCellInst_SboxInst_12_n11}), .b ({ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627]}), .c ({new_AGEMA_signal_1688, new_AGEMA_signal_1687, SubCellInst_SboxInst_12_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U12 ( .a ({new_AGEMA_signal_1426, new_AGEMA_signal_1425, SubCellInst_SboxInst_12_n6}), .b ({new_AGEMA_signal_1690, new_AGEMA_signal_1689, SubCellInst_SboxInst_12_n5}), .clk (clk), .r ({Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_1824, new_AGEMA_signal_1823, Feedback[49]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U7 ( .a ({ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .b ({new_AGEMA_signal_1428, new_AGEMA_signal_1427, SubCellInst_SboxInst_12_n2}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633]}), .c ({new_AGEMA_signal_1692, new_AGEMA_signal_1691, SubCellInst_SboxInst_12_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U19 ( .a ({new_AGEMA_signal_1434, new_AGEMA_signal_1433, SubCellInst_SboxInst_13_n15}), .b ({new_AGEMA_signal_1696, new_AGEMA_signal_1695, SubCellInst_SboxInst_13_n14}), .clk (clk), .r ({Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_1828, new_AGEMA_signal_1827, Feedback[55]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U16 ( .a ({new_AGEMA_signal_1432, new_AGEMA_signal_1431, SubCellInst_SboxInst_13_n11}), .b ({ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639]}), .c ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, SubCellInst_SboxInst_13_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U12 ( .a ({new_AGEMA_signal_1438, new_AGEMA_signal_1437, SubCellInst_SboxInst_13_n6}), .b ({new_AGEMA_signal_1700, new_AGEMA_signal_1699, SubCellInst_SboxInst_13_n5}), .clk (clk), .r ({Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_1832, new_AGEMA_signal_1831, Feedback[53]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U7 ( .a ({ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .b ({new_AGEMA_signal_1440, new_AGEMA_signal_1439, SubCellInst_SboxInst_13_n2}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645]}), .c ({new_AGEMA_signal_1702, new_AGEMA_signal_1701, SubCellInst_SboxInst_13_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U19 ( .a ({new_AGEMA_signal_1446, new_AGEMA_signal_1445, SubCellInst_SboxInst_14_n15}), .b ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, SubCellInst_SboxInst_14_n14}), .clk (clk), .r ({Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_1836, new_AGEMA_signal_1835, Feedback[59]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U16 ( .a ({new_AGEMA_signal_1444, new_AGEMA_signal_1443, SubCellInst_SboxInst_14_n11}), .b ({ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651]}), .c ({new_AGEMA_signal_1708, new_AGEMA_signal_1707, SubCellInst_SboxInst_14_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U12 ( .a ({new_AGEMA_signal_1450, new_AGEMA_signal_1449, SubCellInst_SboxInst_14_n6}), .b ({new_AGEMA_signal_1710, new_AGEMA_signal_1709, SubCellInst_SboxInst_14_n5}), .clk (clk), .r ({Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_1840, new_AGEMA_signal_1839, Feedback[57]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U7 ( .a ({ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .b ({new_AGEMA_signal_1452, new_AGEMA_signal_1451, SubCellInst_SboxInst_14_n2}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657]}), .c ({new_AGEMA_signal_1712, new_AGEMA_signal_1711, SubCellInst_SboxInst_14_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U19 ( .a ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, SubCellInst_SboxInst_15_n15}), .b ({new_AGEMA_signal_1716, new_AGEMA_signal_1715, SubCellInst_SboxInst_15_n14}), .clk (clk), .r ({Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_1844, new_AGEMA_signal_1843, Feedback[63]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U16 ( .a ({new_AGEMA_signal_1456, new_AGEMA_signal_1455, SubCellInst_SboxInst_15_n11}), .b ({ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663]}), .c ({new_AGEMA_signal_1718, new_AGEMA_signal_1717, SubCellInst_SboxInst_15_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U12 ( .a ({new_AGEMA_signal_1462, new_AGEMA_signal_1461, SubCellInst_SboxInst_15_n6}), .b ({new_AGEMA_signal_1720, new_AGEMA_signal_1719, SubCellInst_SboxInst_15_n5}), .clk (clk), .r ({Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_1848, new_AGEMA_signal_1847, Feedback[61]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U7 ( .a ({ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .b ({new_AGEMA_signal_1464, new_AGEMA_signal_1463, SubCellInst_SboxInst_15_n2}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669]}), .c ({new_AGEMA_signal_1722, new_AGEMA_signal_1721, SubCellInst_SboxInst_15_n3}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_0_U1 ( .s (rst), .b ({new_AGEMA_signal_1730, new_AGEMA_signal_1729, Feedback[0]}), .a ({plaintext_s2[0], plaintext_s1[0], plaintext_s0[0]}), .c ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, MCOutput[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_2_U1 ( .s (rst), .b ({new_AGEMA_signal_1726, new_AGEMA_signal_1725, Feedback[2]}), .a ({plaintext_s2[2], plaintext_s1[2], plaintext_s0[2]}), .c ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, MCOutput[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_4_U1 ( .s (rst), .b ({new_AGEMA_signal_1738, new_AGEMA_signal_1737, Feedback[4]}), .a ({plaintext_s2[4], plaintext_s1[4], plaintext_s0[4]}), .c ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, MCOutput[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_6_U1 ( .s (rst), .b ({new_AGEMA_signal_1734, new_AGEMA_signal_1733, Feedback[6]}), .a ({plaintext_s2[6], plaintext_s1[6], plaintext_s0[6]}), .c ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, MCOutput[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_8_U1 ( .s (rst), .b ({new_AGEMA_signal_1746, new_AGEMA_signal_1745, Feedback[8]}), .a ({plaintext_s2[8], plaintext_s1[8], plaintext_s0[8]}), .c ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, MCOutput[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_10_U1 ( .s (rst), .b ({new_AGEMA_signal_1742, new_AGEMA_signal_1741, Feedback[10]}), .a ({plaintext_s2[10], plaintext_s1[10], plaintext_s0[10]}), .c ({new_AGEMA_signal_2182, new_AGEMA_signal_2181, MCOutput[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_12_U1 ( .s (rst), .b ({new_AGEMA_signal_1754, new_AGEMA_signal_1753, Feedback[12]}), .a ({plaintext_s2[12], plaintext_s1[12], plaintext_s0[12]}), .c ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, MCOutput[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_14_U1 ( .s (rst), .b ({new_AGEMA_signal_1750, new_AGEMA_signal_1749, Feedback[14]}), .a ({plaintext_s2[14], plaintext_s1[14], plaintext_s0[14]}), .c ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, MCOutput[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_16_U1 ( .s (rst), .b ({new_AGEMA_signal_1762, new_AGEMA_signal_1761, Feedback[16]}), .a ({plaintext_s2[16], plaintext_s1[16], plaintext_s0[16]}), .c ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, MCOutput[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_18_U1 ( .s (rst), .b ({new_AGEMA_signal_1758, new_AGEMA_signal_1757, Feedback[18]}), .a ({plaintext_s2[18], plaintext_s1[18], plaintext_s0[18]}), .c ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, MCOutput[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_20_U1 ( .s (rst), .b ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, Feedback[20]}), .a ({plaintext_s2[20], plaintext_s1[20], plaintext_s0[20]}), .c ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, MCOutput[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_22_U1 ( .s (rst), .b ({new_AGEMA_signal_1766, new_AGEMA_signal_1765, Feedback[22]}), .a ({plaintext_s2[22], plaintext_s1[22], plaintext_s0[22]}), .c ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, MCOutput[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_24_U1 ( .s (rst), .b ({new_AGEMA_signal_1778, new_AGEMA_signal_1777, Feedback[24]}), .a ({plaintext_s2[24], plaintext_s1[24], plaintext_s0[24]}), .c ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, MCOutput[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_26_U1 ( .s (rst), .b ({new_AGEMA_signal_1774, new_AGEMA_signal_1773, Feedback[26]}), .a ({plaintext_s2[26], plaintext_s1[26], plaintext_s0[26]}), .c ({new_AGEMA_signal_2246, new_AGEMA_signal_2245, MCOutput[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_28_U1 ( .s (rst), .b ({new_AGEMA_signal_1786, new_AGEMA_signal_1785, Feedback[28]}), .a ({plaintext_s2[28], plaintext_s1[28], plaintext_s0[28]}), .c ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, MCOutput[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_30_U1 ( .s (rst), .b ({new_AGEMA_signal_1782, new_AGEMA_signal_1781, Feedback[30]}), .a ({plaintext_s2[30], plaintext_s1[30], plaintext_s0[30]}), .c ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, MCOutput[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_32_U1 ( .s (rst), .b ({new_AGEMA_signal_1794, new_AGEMA_signal_1793, Feedback[32]}), .a ({plaintext_s2[32], plaintext_s1[32], plaintext_s0[32]}), .c ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, MCInput[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_34_U1 ( .s (rst), .b ({new_AGEMA_signal_1790, new_AGEMA_signal_1789, Feedback[34]}), .a ({plaintext_s2[34], plaintext_s1[34], plaintext_s0[34]}), .c ({new_AGEMA_signal_2278, new_AGEMA_signal_2277, MCInput[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_36_U1 ( .s (rst), .b ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, Feedback[36]}), .a ({plaintext_s2[36], plaintext_s1[36], plaintext_s0[36]}), .c ({new_AGEMA_signal_2286, new_AGEMA_signal_2285, MCInput[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_38_U1 ( .s (rst), .b ({new_AGEMA_signal_1798, new_AGEMA_signal_1797, Feedback[38]}), .a ({plaintext_s2[38], plaintext_s1[38], plaintext_s0[38]}), .c ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, MCInput[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_40_U1 ( .s (rst), .b ({new_AGEMA_signal_1810, new_AGEMA_signal_1809, Feedback[40]}), .a ({plaintext_s2[40], plaintext_s1[40], plaintext_s0[40]}), .c ({new_AGEMA_signal_2302, new_AGEMA_signal_2301, MCInput[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_42_U1 ( .s (rst), .b ({new_AGEMA_signal_1806, new_AGEMA_signal_1805, Feedback[42]}), .a ({plaintext_s2[42], plaintext_s1[42], plaintext_s0[42]}), .c ({new_AGEMA_signal_2310, new_AGEMA_signal_2309, MCInput[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_44_U1 ( .s (rst), .b ({new_AGEMA_signal_1818, new_AGEMA_signal_1817, Feedback[44]}), .a ({plaintext_s2[44], plaintext_s1[44], plaintext_s0[44]}), .c ({new_AGEMA_signal_2318, new_AGEMA_signal_2317, MCInput[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_46_U1 ( .s (rst), .b ({new_AGEMA_signal_1814, new_AGEMA_signal_1813, Feedback[46]}), .a ({plaintext_s2[46], plaintext_s1[46], plaintext_s0[46]}), .c ({new_AGEMA_signal_2326, new_AGEMA_signal_2325, MCInput[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_48_U1 ( .s (rst), .b ({new_AGEMA_signal_1826, new_AGEMA_signal_1825, Feedback[48]}), .a ({plaintext_s2[48], plaintext_s1[48], plaintext_s0[48]}), .c ({new_AGEMA_signal_2334, new_AGEMA_signal_2333, MCInput[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_50_U1 ( .s (rst), .b ({new_AGEMA_signal_1822, new_AGEMA_signal_1821, Feedback[50]}), .a ({plaintext_s2[50], plaintext_s1[50], plaintext_s0[50]}), .c ({new_AGEMA_signal_2342, new_AGEMA_signal_2341, MCInput[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_52_U1 ( .s (rst), .b ({new_AGEMA_signal_1834, new_AGEMA_signal_1833, Feedback[52]}), .a ({plaintext_s2[52], plaintext_s1[52], plaintext_s0[52]}), .c ({new_AGEMA_signal_2350, new_AGEMA_signal_2349, MCInput[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_54_U1 ( .s (rst), .b ({new_AGEMA_signal_1830, new_AGEMA_signal_1829, Feedback[54]}), .a ({plaintext_s2[54], plaintext_s1[54], plaintext_s0[54]}), .c ({new_AGEMA_signal_2358, new_AGEMA_signal_2357, MCInput[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_56_U1 ( .s (rst), .b ({new_AGEMA_signal_1842, new_AGEMA_signal_1841, Feedback[56]}), .a ({plaintext_s2[56], plaintext_s1[56], plaintext_s0[56]}), .c ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, MCInput[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_58_U1 ( .s (rst), .b ({new_AGEMA_signal_1838, new_AGEMA_signal_1837, Feedback[58]}), .a ({plaintext_s2[58], plaintext_s1[58], plaintext_s0[58]}), .c ({new_AGEMA_signal_2374, new_AGEMA_signal_2373, MCInput[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_60_U1 ( .s (rst), .b ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, Feedback[60]}), .a ({plaintext_s2[60], plaintext_s1[60], plaintext_s0[60]}), .c ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, MCInput[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) InputMUX_MUXInst_62_U1 ( .s (rst), .b ({new_AGEMA_signal_1846, new_AGEMA_signal_1845, Feedback[62]}), .a ({plaintext_s2[62], plaintext_s1[62], plaintext_s0[62]}), .c ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, MCInput[62]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_0_U3 ( .a ({new_AGEMA_signal_2414, new_AGEMA_signal_2413, MCInst_XOR_r0_Inst_0_n2}), .b ({new_AGEMA_signal_2412, new_AGEMA_signal_2411, MCInst_XOR_r0_Inst_0_n1}), .c ({new_AGEMA_signal_2572, new_AGEMA_signal_2571, MCOutput[48]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_0_U2 ( .a ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, MCOutput[16]}), .b ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, MCOutput[0]}), .c ({new_AGEMA_signal_2412, new_AGEMA_signal_2411, MCInst_XOR_r0_Inst_0_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2334, new_AGEMA_signal_2333, MCInput[48]}), .c ({new_AGEMA_signal_2414, new_AGEMA_signal_2413, MCInst_XOR_r0_Inst_0_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_0_U2 ( .a ({new_AGEMA_signal_2416, new_AGEMA_signal_2415, MCInst_XOR_r1_Inst_0_n1}), .b ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, MCOutput[0]}), .c ({new_AGEMA_signal_2574, new_AGEMA_signal_2573, MCOutput[32]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, MCInput[32]}), .c ({new_AGEMA_signal_2416, new_AGEMA_signal_2415, MCInst_XOR_r1_Inst_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_2_U3 ( .a ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, MCInst_XOR_r0_Inst_2_n2}), .b ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, MCInst_XOR_r0_Inst_2_n1}), .c ({new_AGEMA_signal_2580, new_AGEMA_signal_2579, MCOutput[50]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_2_U2 ( .a ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, MCOutput[18]}), .b ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, MCOutput[2]}), .c ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, MCInst_XOR_r0_Inst_2_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2342, new_AGEMA_signal_2341, MCInput[50]}), .c ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, MCInst_XOR_r0_Inst_2_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_2_U2 ( .a ({new_AGEMA_signal_2428, new_AGEMA_signal_2427, MCInst_XOR_r1_Inst_2_n1}), .b ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, MCOutput[2]}), .c ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, MCOutput[34]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2278, new_AGEMA_signal_2277, MCInput[34]}), .c ({new_AGEMA_signal_2428, new_AGEMA_signal_2427, MCInst_XOR_r1_Inst_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_4_U3 ( .a ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, MCInst_XOR_r0_Inst_4_n2}), .b ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, MCInst_XOR_r0_Inst_4_n1}), .c ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, MCOutput[52]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_4_U2 ( .a ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, MCOutput[20]}), .b ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, MCOutput[4]}), .c ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, MCInst_XOR_r0_Inst_4_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_4_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2350, new_AGEMA_signal_2349, MCInput[52]}), .c ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, MCInst_XOR_r0_Inst_4_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_4_U2 ( .a ({new_AGEMA_signal_2440, new_AGEMA_signal_2439, MCInst_XOR_r1_Inst_4_n1}), .b ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, MCOutput[4]}), .c ({new_AGEMA_signal_2590, new_AGEMA_signal_2589, MCOutput[36]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_4_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2286, new_AGEMA_signal_2285, MCInput[36]}), .c ({new_AGEMA_signal_2440, new_AGEMA_signal_2439, MCInst_XOR_r1_Inst_4_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_6_U3 ( .a ({new_AGEMA_signal_2450, new_AGEMA_signal_2449, MCInst_XOR_r0_Inst_6_n2}), .b ({new_AGEMA_signal_2448, new_AGEMA_signal_2447, MCInst_XOR_r0_Inst_6_n1}), .c ({new_AGEMA_signal_2596, new_AGEMA_signal_2595, MCOutput[54]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_6_U2 ( .a ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, MCOutput[22]}), .b ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, MCOutput[6]}), .c ({new_AGEMA_signal_2448, new_AGEMA_signal_2447, MCInst_XOR_r0_Inst_6_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_6_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2358, new_AGEMA_signal_2357, MCInput[54]}), .c ({new_AGEMA_signal_2450, new_AGEMA_signal_2449, MCInst_XOR_r0_Inst_6_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_6_U2 ( .a ({new_AGEMA_signal_2452, new_AGEMA_signal_2451, MCInst_XOR_r1_Inst_6_n1}), .b ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, MCOutput[6]}), .c ({new_AGEMA_signal_2598, new_AGEMA_signal_2597, MCOutput[38]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_6_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, MCInput[38]}), .c ({new_AGEMA_signal_2452, new_AGEMA_signal_2451, MCInst_XOR_r1_Inst_6_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_8_U3 ( .a ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, MCInst_XOR_r0_Inst_8_n2}), .b ({new_AGEMA_signal_2460, new_AGEMA_signal_2459, MCInst_XOR_r0_Inst_8_n1}), .c ({new_AGEMA_signal_2604, new_AGEMA_signal_2603, MCOutput[56]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_8_U2 ( .a ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, MCOutput[24]}), .b ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, MCOutput[8]}), .c ({new_AGEMA_signal_2460, new_AGEMA_signal_2459, MCInst_XOR_r0_Inst_8_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_8_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, MCInput[56]}), .c ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, MCInst_XOR_r0_Inst_8_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_8_U2 ( .a ({new_AGEMA_signal_2464, new_AGEMA_signal_2463, MCInst_XOR_r1_Inst_8_n1}), .b ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, MCOutput[8]}), .c ({new_AGEMA_signal_2606, new_AGEMA_signal_2605, MCOutput[40]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_8_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2302, new_AGEMA_signal_2301, MCInput[40]}), .c ({new_AGEMA_signal_2464, new_AGEMA_signal_2463, MCInst_XOR_r1_Inst_8_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_10_U3 ( .a ({new_AGEMA_signal_2474, new_AGEMA_signal_2473, MCInst_XOR_r0_Inst_10_n2}), .b ({new_AGEMA_signal_2472, new_AGEMA_signal_2471, MCInst_XOR_r0_Inst_10_n1}), .c ({new_AGEMA_signal_2612, new_AGEMA_signal_2611, MCOutput[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_10_U2 ( .a ({new_AGEMA_signal_2246, new_AGEMA_signal_2245, MCOutput[26]}), .b ({new_AGEMA_signal_2182, new_AGEMA_signal_2181, MCOutput[10]}), .c ({new_AGEMA_signal_2472, new_AGEMA_signal_2471, MCInst_XOR_r0_Inst_10_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_10_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2374, new_AGEMA_signal_2373, MCInput[58]}), .c ({new_AGEMA_signal_2474, new_AGEMA_signal_2473, MCInst_XOR_r0_Inst_10_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_10_U2 ( .a ({new_AGEMA_signal_2476, new_AGEMA_signal_2475, MCInst_XOR_r1_Inst_10_n1}), .b ({new_AGEMA_signal_2182, new_AGEMA_signal_2181, MCOutput[10]}), .c ({new_AGEMA_signal_2614, new_AGEMA_signal_2613, MCOutput[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_10_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2310, new_AGEMA_signal_2309, MCInput[42]}), .c ({new_AGEMA_signal_2476, new_AGEMA_signal_2475, MCInst_XOR_r1_Inst_10_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_12_U3 ( .a ({new_AGEMA_signal_2486, new_AGEMA_signal_2485, MCInst_XOR_r0_Inst_12_n2}), .b ({new_AGEMA_signal_2484, new_AGEMA_signal_2483, MCInst_XOR_r0_Inst_12_n1}), .c ({new_AGEMA_signal_2620, new_AGEMA_signal_2619, MCOutput[60]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_12_U2 ( .a ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, MCOutput[28]}), .b ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, MCOutput[12]}), .c ({new_AGEMA_signal_2484, new_AGEMA_signal_2483, MCInst_XOR_r0_Inst_12_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_12_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, MCInput[60]}), .c ({new_AGEMA_signal_2486, new_AGEMA_signal_2485, MCInst_XOR_r0_Inst_12_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_12_U2 ( .a ({new_AGEMA_signal_2488, new_AGEMA_signal_2487, MCInst_XOR_r1_Inst_12_n1}), .b ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, MCOutput[12]}), .c ({new_AGEMA_signal_2622, new_AGEMA_signal_2621, MCOutput[44]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_12_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2318, new_AGEMA_signal_2317, MCInput[44]}), .c ({new_AGEMA_signal_2488, new_AGEMA_signal_2487, MCInst_XOR_r1_Inst_12_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_14_U3 ( .a ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, MCInst_XOR_r0_Inst_14_n2}), .b ({new_AGEMA_signal_2496, new_AGEMA_signal_2495, MCInst_XOR_r0_Inst_14_n1}), .c ({new_AGEMA_signal_2628, new_AGEMA_signal_2627, MCOutput[62]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_14_U2 ( .a ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, MCOutput[30]}), .b ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, MCOutput[14]}), .c ({new_AGEMA_signal_2496, new_AGEMA_signal_2495, MCInst_XOR_r0_Inst_14_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r0_Inst_14_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, MCInput[62]}), .c ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, MCInst_XOR_r0_Inst_14_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_14_U2 ( .a ({new_AGEMA_signal_2500, new_AGEMA_signal_2499, MCInst_XOR_r1_Inst_14_n1}), .b ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, MCOutput[14]}), .c ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, MCOutput[46]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MCInst_XOR_r1_Inst_14_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2326, new_AGEMA_signal_2325, MCInput[46]}), .c ({new_AGEMA_signal_2500, new_AGEMA_signal_2499, MCInst_XOR_r1_Inst_14_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2700, new_AGEMA_signal_2699, AddKeyXOR1_XORInst_0_0_n1}), .b ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, SelectedKey[48]}), .c ({new_AGEMA_signal_2764, new_AGEMA_signal_2763, AddRoundKeyOutput[48]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2572, new_AGEMA_signal_2571, MCOutput[48]}), .c ({new_AGEMA_signal_2700, new_AGEMA_signal_2699, AddKeyXOR1_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, AddKeyXOR1_XORInst_0_2_n1}), .b ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, SelectedKey[50]}), .c ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, AddRoundKeyOutput[50]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2580, new_AGEMA_signal_2579, MCOutput[50]}), .c ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, AddKeyXOR1_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2708, new_AGEMA_signal_2707, AddKeyXOR1_XORInst_1_0_n1}), .b ({new_AGEMA_signal_2102, new_AGEMA_signal_2101, SelectedKey[52]}), .c ({new_AGEMA_signal_2772, new_AGEMA_signal_2771, AddRoundKeyOutput[52]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, MCOutput[52]}), .c ({new_AGEMA_signal_2708, new_AGEMA_signal_2707, AddKeyXOR1_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2712, new_AGEMA_signal_2711, AddKeyXOR1_XORInst_1_2_n1}), .b ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, SelectedKey[54]}), .c ({new_AGEMA_signal_2776, new_AGEMA_signal_2775, AddRoundKeyOutput[54]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2596, new_AGEMA_signal_2595, MCOutput[54]}), .c ({new_AGEMA_signal_2712, new_AGEMA_signal_2711, AddKeyXOR1_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_2716, new_AGEMA_signal_2715, AddKeyXOR1_XORInst_2_0_n1}), .b ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, SelectedKey[56]}), .c ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, AddRoundKeyOutput[56]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2604, new_AGEMA_signal_2603, MCOutput[56]}), .c ({new_AGEMA_signal_2716, new_AGEMA_signal_2715, AddKeyXOR1_XORInst_2_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_2720, new_AGEMA_signal_2719, AddKeyXOR1_XORInst_2_2_n1}), .b ({new_AGEMA_signal_2120, new_AGEMA_signal_2119, SelectedKey[58]}), .c ({new_AGEMA_signal_2784, new_AGEMA_signal_2783, AddRoundKeyOutput[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2612, new_AGEMA_signal_2611, MCOutput[58]}), .c ({new_AGEMA_signal_2720, new_AGEMA_signal_2719, AddKeyXOR1_XORInst_2_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_2724, new_AGEMA_signal_2723, AddKeyXOR1_XORInst_3_0_n1}), .b ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, SelectedKey[60]}), .c ({new_AGEMA_signal_2788, new_AGEMA_signal_2787, AddRoundKeyOutput[60]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2620, new_AGEMA_signal_2619, MCOutput[60]}), .c ({new_AGEMA_signal_2724, new_AGEMA_signal_2723, AddKeyXOR1_XORInst_3_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_2728, new_AGEMA_signal_2727, AddKeyXOR1_XORInst_3_2_n1}), .b ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, SelectedKey[62]}), .c ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, AddRoundKeyOutput[62]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR1_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2628, new_AGEMA_signal_2627, MCOutput[62]}), .c ({new_AGEMA_signal_2728, new_AGEMA_signal_2727, AddKeyXOR1_XORInst_3_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_0_0_U3 ( .a ({new_AGEMA_signal_2732, new_AGEMA_signal_2731, AddKeyConstXOR_XORInst_0_0_n2}), .b ({new_AGEMA_signal_2396, new_AGEMA_signal_2395, AddKeyConstXOR_XORInst_0_0_n1}), .c ({new_AGEMA_signal_2796, new_AGEMA_signal_2795, AddRoundKeyOutput[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2606, new_AGEMA_signal_2605, MCOutput[40]}), .c ({new_AGEMA_signal_2732, new_AGEMA_signal_2731, AddKeyConstXOR_XORInst_0_0_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_0_2_U3 ( .a ({new_AGEMA_signal_2736, new_AGEMA_signal_2735, AddKeyConstXOR_XORInst_0_2_n2}), .b ({new_AGEMA_signal_2400, new_AGEMA_signal_2399, AddKeyConstXOR_XORInst_0_2_n1}), .c ({new_AGEMA_signal_2800, new_AGEMA_signal_2799, AddRoundKeyOutput[42]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2614, new_AGEMA_signal_2613, MCOutput[42]}), .c ({new_AGEMA_signal_2736, new_AGEMA_signal_2735, AddKeyConstXOR_XORInst_0_2_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_1_0_U3 ( .a ({new_AGEMA_signal_2740, new_AGEMA_signal_2739, AddKeyConstXOR_XORInst_1_0_n2}), .b ({new_AGEMA_signal_2404, new_AGEMA_signal_2403, AddKeyConstXOR_XORInst_1_0_n1}), .c ({new_AGEMA_signal_2804, new_AGEMA_signal_2803, AddRoundKeyOutput[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2622, new_AGEMA_signal_2621, MCOutput[44]}), .c ({new_AGEMA_signal_2740, new_AGEMA_signal_2739, AddKeyConstXOR_XORInst_1_0_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_1_2_U3 ( .a ({new_AGEMA_signal_2744, new_AGEMA_signal_2743, AddKeyConstXOR_XORInst_1_2_n2}), .b ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, AddKeyConstXOR_XORInst_1_2_n1}), .c ({new_AGEMA_signal_2808, new_AGEMA_signal_2807, AddRoundKeyOutput[46]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyConstXOR_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, MCOutput[46]}), .c ({new_AGEMA_signal_2744, new_AGEMA_signal_2743, AddKeyConstXOR_XORInst_1_2_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2508, new_AGEMA_signal_2507, AddKeyXOR2_XORInst_0_0_n1}), .b ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, SelectedKey[0]}), .c ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, AddRoundKeyOutput[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, MCOutput[0]}), .c ({new_AGEMA_signal_2508, new_AGEMA_signal_2507, AddKeyXOR2_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2512, new_AGEMA_signal_2511, AddKeyXOR2_XORInst_0_2_n1}), .b ({new_AGEMA_signal_1478, new_AGEMA_signal_1477, SelectedKey[2]}), .c ({new_AGEMA_signal_2640, new_AGEMA_signal_2639, AddRoundKeyOutput[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, MCOutput[2]}), .c ({new_AGEMA_signal_2512, new_AGEMA_signal_2511, AddKeyXOR2_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, AddKeyXOR2_XORInst_1_0_n1}), .b ({new_AGEMA_signal_1868, new_AGEMA_signal_1867, SelectedKey[4]}), .c ({new_AGEMA_signal_2644, new_AGEMA_signal_2643, AddRoundKeyOutput[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, MCOutput[4]}), .c ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, AddKeyXOR2_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2520, new_AGEMA_signal_2519, AddKeyXOR2_XORInst_1_2_n1}), .b ({new_AGEMA_signal_1880, new_AGEMA_signal_1879, SelectedKey[6]}), .c ({new_AGEMA_signal_2648, new_AGEMA_signal_2647, AddRoundKeyOutput[6]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, MCOutput[6]}), .c ({new_AGEMA_signal_2520, new_AGEMA_signal_2519, AddKeyXOR2_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_2524, new_AGEMA_signal_2523, AddKeyXOR2_XORInst_2_0_n1}), .b ({new_AGEMA_signal_1892, new_AGEMA_signal_1891, SelectedKey[8]}), .c ({new_AGEMA_signal_2652, new_AGEMA_signal_2651, AddRoundKeyOutput[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, MCOutput[8]}), .c ({new_AGEMA_signal_2524, new_AGEMA_signal_2523, AddKeyXOR2_XORInst_2_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_2528, new_AGEMA_signal_2527, AddKeyXOR2_XORInst_2_2_n1}), .b ({new_AGEMA_signal_1904, new_AGEMA_signal_1903, SelectedKey[10]}), .c ({new_AGEMA_signal_2656, new_AGEMA_signal_2655, AddRoundKeyOutput[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2182, new_AGEMA_signal_2181, MCOutput[10]}), .c ({new_AGEMA_signal_2528, new_AGEMA_signal_2527, AddKeyXOR2_XORInst_2_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_2532, new_AGEMA_signal_2531, AddKeyXOR2_XORInst_3_0_n1}), .b ({new_AGEMA_signal_1916, new_AGEMA_signal_1915, SelectedKey[12]}), .c ({new_AGEMA_signal_2660, new_AGEMA_signal_2659, AddRoundKeyOutput[12]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, MCOutput[12]}), .c ({new_AGEMA_signal_2532, new_AGEMA_signal_2531, AddKeyXOR2_XORInst_3_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_2536, new_AGEMA_signal_2535, AddKeyXOR2_XORInst_3_2_n1}), .b ({new_AGEMA_signal_1928, new_AGEMA_signal_1927, SelectedKey[14]}), .c ({new_AGEMA_signal_2664, new_AGEMA_signal_2663, AddRoundKeyOutput[14]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, MCOutput[14]}), .c ({new_AGEMA_signal_2536, new_AGEMA_signal_2535, AddKeyXOR2_XORInst_3_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_4_0_U2 ( .a ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, AddKeyXOR2_XORInst_4_0_n1}), .b ({new_AGEMA_signal_1940, new_AGEMA_signal_1939, SelectedKey[16]}), .c ({new_AGEMA_signal_2668, new_AGEMA_signal_2667, AddRoundKeyOutput[16]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_4_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, MCOutput[16]}), .c ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, AddKeyXOR2_XORInst_4_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_4_2_U2 ( .a ({new_AGEMA_signal_2544, new_AGEMA_signal_2543, AddKeyXOR2_XORInst_4_2_n1}), .b ({new_AGEMA_signal_1952, new_AGEMA_signal_1951, SelectedKey[18]}), .c ({new_AGEMA_signal_2672, new_AGEMA_signal_2671, AddRoundKeyOutput[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_4_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, MCOutput[18]}), .c ({new_AGEMA_signal_2544, new_AGEMA_signal_2543, AddKeyXOR2_XORInst_4_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_5_0_U2 ( .a ({new_AGEMA_signal_2548, new_AGEMA_signal_2547, AddKeyXOR2_XORInst_5_0_n1}), .b ({new_AGEMA_signal_1964, new_AGEMA_signal_1963, SelectedKey[20]}), .c ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, AddRoundKeyOutput[20]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_5_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, MCOutput[20]}), .c ({new_AGEMA_signal_2548, new_AGEMA_signal_2547, AddKeyXOR2_XORInst_5_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_5_2_U2 ( .a ({new_AGEMA_signal_2552, new_AGEMA_signal_2551, AddKeyXOR2_XORInst_5_2_n1}), .b ({new_AGEMA_signal_1484, new_AGEMA_signal_1483, SelectedKey[22]}), .c ({new_AGEMA_signal_2680, new_AGEMA_signal_2679, AddRoundKeyOutput[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_5_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, MCOutput[22]}), .c ({new_AGEMA_signal_2552, new_AGEMA_signal_2551, AddKeyXOR2_XORInst_5_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_6_0_U2 ( .a ({new_AGEMA_signal_2556, new_AGEMA_signal_2555, AddKeyXOR2_XORInst_6_0_n1}), .b ({new_AGEMA_signal_1496, new_AGEMA_signal_1495, SelectedKey[24]}), .c ({new_AGEMA_signal_2684, new_AGEMA_signal_2683, AddRoundKeyOutput[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_6_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, MCOutput[24]}), .c ({new_AGEMA_signal_2556, new_AGEMA_signal_2555, AddKeyXOR2_XORInst_6_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_6_2_U2 ( .a ({new_AGEMA_signal_2560, new_AGEMA_signal_2559, AddKeyXOR2_XORInst_6_2_n1}), .b ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, SelectedKey[26]}), .c ({new_AGEMA_signal_2688, new_AGEMA_signal_2687, AddRoundKeyOutput[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_6_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2246, new_AGEMA_signal_2245, MCOutput[26]}), .c ({new_AGEMA_signal_2560, new_AGEMA_signal_2559, AddKeyXOR2_XORInst_6_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_7_0_U2 ( .a ({new_AGEMA_signal_2564, new_AGEMA_signal_2563, AddKeyXOR2_XORInst_7_0_n1}), .b ({new_AGEMA_signal_1976, new_AGEMA_signal_1975, SelectedKey[28]}), .c ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, AddRoundKeyOutput[28]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_7_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, MCOutput[28]}), .c ({new_AGEMA_signal_2564, new_AGEMA_signal_2563, AddKeyXOR2_XORInst_7_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_7_2_U2 ( .a ({new_AGEMA_signal_2568, new_AGEMA_signal_2567, AddKeyXOR2_XORInst_7_2_n1}), .b ({new_AGEMA_signal_1988, new_AGEMA_signal_1987, SelectedKey[30]}), .c ({new_AGEMA_signal_2696, new_AGEMA_signal_2695, AddRoundKeyOutput[30]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_7_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, MCOutput[30]}), .c ({new_AGEMA_signal_2568, new_AGEMA_signal_2567, AddKeyXOR2_XORInst_7_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_8_0_U2 ( .a ({new_AGEMA_signal_2748, new_AGEMA_signal_2747, AddKeyXOR2_XORInst_8_0_n1}), .b ({new_AGEMA_signal_2000, new_AGEMA_signal_1999, SelectedKey[32]}), .c ({new_AGEMA_signal_2812, new_AGEMA_signal_2811, AddRoundKeyOutput[32]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_8_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2574, new_AGEMA_signal_2573, MCOutput[32]}), .c ({new_AGEMA_signal_2748, new_AGEMA_signal_2747, AddKeyXOR2_XORInst_8_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_8_2_U2 ( .a ({new_AGEMA_signal_2752, new_AGEMA_signal_2751, AddKeyXOR2_XORInst_8_2_n1}), .b ({new_AGEMA_signal_2006, new_AGEMA_signal_2005, SelectedKey[34]}), .c ({new_AGEMA_signal_2816, new_AGEMA_signal_2815, AddRoundKeyOutput[34]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_8_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, MCOutput[34]}), .c ({new_AGEMA_signal_2752, new_AGEMA_signal_2751, AddKeyXOR2_XORInst_8_2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_9_0_U2 ( .a ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, AddKeyXOR2_XORInst_9_0_n1}), .b ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, SelectedKey[36]}), .c ({new_AGEMA_signal_2820, new_AGEMA_signal_2819, AddRoundKeyOutput[36]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_9_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2590, new_AGEMA_signal_2589, MCOutput[36]}), .c ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, AddKeyXOR2_XORInst_9_0_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_9_2_U2 ( .a ({new_AGEMA_signal_2760, new_AGEMA_signal_2759, AddKeyXOR2_XORInst_9_2_n1}), .b ({new_AGEMA_signal_2024, new_AGEMA_signal_2023, SelectedKey[38]}), .c ({new_AGEMA_signal_2824, new_AGEMA_signal_2823, AddRoundKeyOutput[38]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) AddKeyXOR2_XORInst_9_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2598, new_AGEMA_signal_2597, MCOutput[38]}), .c ({new_AGEMA_signal_2760, new_AGEMA_signal_2759, AddKeyXOR2_XORInst_9_2_n1}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U17 ( .a ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, SubCellInst_SboxInst_0_n15}), .b ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, SubCellInst_SboxInst_0_n12}), .clk (clk), .r ({Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_1726, new_AGEMA_signal_1725, Feedback[2]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U8 ( .a ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, SubCellInst_SboxInst_0_n13}), .b ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, SubCellInst_SboxInst_0_n3}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675]}), .c ({new_AGEMA_signal_1730, new_AGEMA_signal_1729, Feedback[0]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U17 ( .a ({new_AGEMA_signal_1290, new_AGEMA_signal_1289, SubCellInst_SboxInst_1_n15}), .b ({new_AGEMA_signal_1578, new_AGEMA_signal_1577, SubCellInst_SboxInst_1_n12}), .clk (clk), .r ({Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_1734, new_AGEMA_signal_1733, Feedback[6]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U8 ( .a ({new_AGEMA_signal_1298, new_AGEMA_signal_1297, SubCellInst_SboxInst_1_n13}), .b ({new_AGEMA_signal_1582, new_AGEMA_signal_1581, SubCellInst_SboxInst_1_n3}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681]}), .c ({new_AGEMA_signal_1738, new_AGEMA_signal_1737, Feedback[4]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U17 ( .a ({new_AGEMA_signal_1302, new_AGEMA_signal_1301, SubCellInst_SboxInst_2_n15}), .b ({new_AGEMA_signal_1588, new_AGEMA_signal_1587, SubCellInst_SboxInst_2_n12}), .clk (clk), .r ({Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_1742, new_AGEMA_signal_1741, Feedback[10]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U8 ( .a ({new_AGEMA_signal_1310, new_AGEMA_signal_1309, SubCellInst_SboxInst_2_n13}), .b ({new_AGEMA_signal_1592, new_AGEMA_signal_1591, SubCellInst_SboxInst_2_n3}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687]}), .c ({new_AGEMA_signal_1746, new_AGEMA_signal_1745, Feedback[8]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U17 ( .a ({new_AGEMA_signal_1314, new_AGEMA_signal_1313, SubCellInst_SboxInst_3_n15}), .b ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, SubCellInst_SboxInst_3_n12}), .clk (clk), .r ({Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_1750, new_AGEMA_signal_1749, Feedback[14]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U8 ( .a ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, SubCellInst_SboxInst_3_n13}), .b ({new_AGEMA_signal_1602, new_AGEMA_signal_1601, SubCellInst_SboxInst_3_n3}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693]}), .c ({new_AGEMA_signal_1754, new_AGEMA_signal_1753, Feedback[12]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U17 ( .a ({new_AGEMA_signal_1326, new_AGEMA_signal_1325, SubCellInst_SboxInst_4_n15}), .b ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, SubCellInst_SboxInst_4_n12}), .clk (clk), .r ({Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_1758, new_AGEMA_signal_1757, Feedback[18]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U8 ( .a ({new_AGEMA_signal_1334, new_AGEMA_signal_1333, SubCellInst_SboxInst_4_n13}), .b ({new_AGEMA_signal_1612, new_AGEMA_signal_1611, SubCellInst_SboxInst_4_n3}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699]}), .c ({new_AGEMA_signal_1762, new_AGEMA_signal_1761, Feedback[16]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U17 ( .a ({new_AGEMA_signal_1338, new_AGEMA_signal_1337, SubCellInst_SboxInst_5_n15}), .b ({new_AGEMA_signal_1618, new_AGEMA_signal_1617, SubCellInst_SboxInst_5_n12}), .clk (clk), .r ({Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_1766, new_AGEMA_signal_1765, Feedback[22]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U8 ( .a ({new_AGEMA_signal_1346, new_AGEMA_signal_1345, SubCellInst_SboxInst_5_n13}), .b ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, SubCellInst_SboxInst_5_n3}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705]}), .c ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, Feedback[20]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U17 ( .a ({new_AGEMA_signal_1350, new_AGEMA_signal_1349, SubCellInst_SboxInst_6_n15}), .b ({new_AGEMA_signal_1628, new_AGEMA_signal_1627, SubCellInst_SboxInst_6_n12}), .clk (clk), .r ({Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_1774, new_AGEMA_signal_1773, Feedback[26]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U8 ( .a ({new_AGEMA_signal_1358, new_AGEMA_signal_1357, SubCellInst_SboxInst_6_n13}), .b ({new_AGEMA_signal_1632, new_AGEMA_signal_1631, SubCellInst_SboxInst_6_n3}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711]}), .c ({new_AGEMA_signal_1778, new_AGEMA_signal_1777, Feedback[24]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U17 ( .a ({new_AGEMA_signal_1362, new_AGEMA_signal_1361, SubCellInst_SboxInst_7_n15}), .b ({new_AGEMA_signal_1638, new_AGEMA_signal_1637, SubCellInst_SboxInst_7_n12}), .clk (clk), .r ({Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_1782, new_AGEMA_signal_1781, Feedback[30]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U8 ( .a ({new_AGEMA_signal_1370, new_AGEMA_signal_1369, SubCellInst_SboxInst_7_n13}), .b ({new_AGEMA_signal_1642, new_AGEMA_signal_1641, SubCellInst_SboxInst_7_n3}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717]}), .c ({new_AGEMA_signal_1786, new_AGEMA_signal_1785, Feedback[28]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U17 ( .a ({new_AGEMA_signal_1374, new_AGEMA_signal_1373, SubCellInst_SboxInst_8_n15}), .b ({new_AGEMA_signal_1648, new_AGEMA_signal_1647, SubCellInst_SboxInst_8_n12}), .clk (clk), .r ({Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_1790, new_AGEMA_signal_1789, Feedback[34]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U8 ( .a ({new_AGEMA_signal_1382, new_AGEMA_signal_1381, SubCellInst_SboxInst_8_n13}), .b ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, SubCellInst_SboxInst_8_n3}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723]}), .c ({new_AGEMA_signal_1794, new_AGEMA_signal_1793, Feedback[32]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U17 ( .a ({new_AGEMA_signal_1386, new_AGEMA_signal_1385, SubCellInst_SboxInst_9_n15}), .b ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, SubCellInst_SboxInst_9_n12}), .clk (clk), .r ({Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_1798, new_AGEMA_signal_1797, Feedback[38]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U8 ( .a ({new_AGEMA_signal_1394, new_AGEMA_signal_1393, SubCellInst_SboxInst_9_n13}), .b ({new_AGEMA_signal_1662, new_AGEMA_signal_1661, SubCellInst_SboxInst_9_n3}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729]}), .c ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, Feedback[36]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U17 ( .a ({new_AGEMA_signal_1398, new_AGEMA_signal_1397, SubCellInst_SboxInst_10_n15}), .b ({new_AGEMA_signal_1668, new_AGEMA_signal_1667, SubCellInst_SboxInst_10_n12}), .clk (clk), .r ({Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_1806, new_AGEMA_signal_1805, Feedback[42]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U8 ( .a ({new_AGEMA_signal_1406, new_AGEMA_signal_1405, SubCellInst_SboxInst_10_n13}), .b ({new_AGEMA_signal_1672, new_AGEMA_signal_1671, SubCellInst_SboxInst_10_n3}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735]}), .c ({new_AGEMA_signal_1810, new_AGEMA_signal_1809, Feedback[40]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U17 ( .a ({new_AGEMA_signal_1410, new_AGEMA_signal_1409, SubCellInst_SboxInst_11_n15}), .b ({new_AGEMA_signal_1678, new_AGEMA_signal_1677, SubCellInst_SboxInst_11_n12}), .clk (clk), .r ({Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_1814, new_AGEMA_signal_1813, Feedback[46]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U8 ( .a ({new_AGEMA_signal_1418, new_AGEMA_signal_1417, SubCellInst_SboxInst_11_n13}), .b ({new_AGEMA_signal_1682, new_AGEMA_signal_1681, SubCellInst_SboxInst_11_n3}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741]}), .c ({new_AGEMA_signal_1818, new_AGEMA_signal_1817, Feedback[44]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U17 ( .a ({new_AGEMA_signal_1422, new_AGEMA_signal_1421, SubCellInst_SboxInst_12_n15}), .b ({new_AGEMA_signal_1688, new_AGEMA_signal_1687, SubCellInst_SboxInst_12_n12}), .clk (clk), .r ({Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_1822, new_AGEMA_signal_1821, Feedback[50]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U8 ( .a ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, SubCellInst_SboxInst_12_n13}), .b ({new_AGEMA_signal_1692, new_AGEMA_signal_1691, SubCellInst_SboxInst_12_n3}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747]}), .c ({new_AGEMA_signal_1826, new_AGEMA_signal_1825, Feedback[48]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U17 ( .a ({new_AGEMA_signal_1434, new_AGEMA_signal_1433, SubCellInst_SboxInst_13_n15}), .b ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, SubCellInst_SboxInst_13_n12}), .clk (clk), .r ({Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_1830, new_AGEMA_signal_1829, Feedback[54]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U8 ( .a ({new_AGEMA_signal_1442, new_AGEMA_signal_1441, SubCellInst_SboxInst_13_n13}), .b ({new_AGEMA_signal_1702, new_AGEMA_signal_1701, SubCellInst_SboxInst_13_n3}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753]}), .c ({new_AGEMA_signal_1834, new_AGEMA_signal_1833, Feedback[52]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U17 ( .a ({new_AGEMA_signal_1446, new_AGEMA_signal_1445, SubCellInst_SboxInst_14_n15}), .b ({new_AGEMA_signal_1708, new_AGEMA_signal_1707, SubCellInst_SboxInst_14_n12}), .clk (clk), .r ({Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_1838, new_AGEMA_signal_1837, Feedback[58]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U8 ( .a ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, SubCellInst_SboxInst_14_n13}), .b ({new_AGEMA_signal_1712, new_AGEMA_signal_1711, SubCellInst_SboxInst_14_n3}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759]}), .c ({new_AGEMA_signal_1842, new_AGEMA_signal_1841, Feedback[56]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U17 ( .a ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, SubCellInst_SboxInst_15_n15}), .b ({new_AGEMA_signal_1718, new_AGEMA_signal_1717, SubCellInst_SboxInst_15_n12}), .clk (clk), .r ({Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_1846, new_AGEMA_signal_1845, Feedback[62]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U8 ( .a ({new_AGEMA_signal_1466, new_AGEMA_signal_1465, SubCellInst_SboxInst_15_n13}), .b ({new_AGEMA_signal_1722, new_AGEMA_signal_1721, SubCellInst_SboxInst_15_n3}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765]}), .c ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, Feedback[60]}) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_63__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2794, new_AGEMA_signal_2793, AddRoundKeyOutput[63]}), .Q ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_62__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, AddRoundKeyOutput[62]}), .Q ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_61__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2790, new_AGEMA_signal_2789, AddRoundKeyOutput[61]}), .Q ({ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_60__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2788, new_AGEMA_signal_2787, AddRoundKeyOutput[60]}), .Q ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_59__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2786, new_AGEMA_signal_2785, AddRoundKeyOutput[59]}), .Q ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_58__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2784, new_AGEMA_signal_2783, AddRoundKeyOutput[58]}), .Q ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_57__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2782, new_AGEMA_signal_2781, AddRoundKeyOutput[57]}), .Q ({ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_56__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, AddRoundKeyOutput[56]}), .Q ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_55__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2778, new_AGEMA_signal_2777, AddRoundKeyOutput[55]}), .Q ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_54__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2776, new_AGEMA_signal_2775, AddRoundKeyOutput[54]}), .Q ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_53__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2774, new_AGEMA_signal_2773, AddRoundKeyOutput[53]}), .Q ({ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_52__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2772, new_AGEMA_signal_2771, AddRoundKeyOutput[52]}), .Q ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_51__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2770, new_AGEMA_signal_2769, AddRoundKeyOutput[51]}), .Q ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_50__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, AddRoundKeyOutput[50]}), .Q ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_49__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2766, new_AGEMA_signal_2765, AddRoundKeyOutput[49]}), .Q ({ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_48__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2764, new_AGEMA_signal_2763, AddRoundKeyOutput[48]}), .Q ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_47__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2810, new_AGEMA_signal_2809, AddRoundKeyOutput[47]}), .Q ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_46__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2808, new_AGEMA_signal_2807, AddRoundKeyOutput[46]}), .Q ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_45__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2806, new_AGEMA_signal_2805, AddRoundKeyOutput[45]}), .Q ({ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_44__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2804, new_AGEMA_signal_2803, AddRoundKeyOutput[44]}), .Q ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_43__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2802, new_AGEMA_signal_2801, AddRoundKeyOutput[43]}), .Q ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_42__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2800, new_AGEMA_signal_2799, AddRoundKeyOutput[42]}), .Q ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_41__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2798, new_AGEMA_signal_2797, AddRoundKeyOutput[41]}), .Q ({ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_40__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2796, new_AGEMA_signal_2795, AddRoundKeyOutput[40]}), .Q ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_39__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2826, new_AGEMA_signal_2825, AddRoundKeyOutput[39]}), .Q ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_38__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2824, new_AGEMA_signal_2823, AddRoundKeyOutput[38]}), .Q ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_37__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2822, new_AGEMA_signal_2821, AddRoundKeyOutput[37]}), .Q ({ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_36__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2820, new_AGEMA_signal_2819, AddRoundKeyOutput[36]}), .Q ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_35__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2818, new_AGEMA_signal_2817, AddRoundKeyOutput[35]}), .Q ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_34__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2816, new_AGEMA_signal_2815, AddRoundKeyOutput[34]}), .Q ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_33__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2814, new_AGEMA_signal_2813, AddRoundKeyOutput[33]}), .Q ({ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_32__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2812, new_AGEMA_signal_2811, AddRoundKeyOutput[32]}), .Q ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_31__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2698, new_AGEMA_signal_2697, AddRoundKeyOutput[31]}), .Q ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_30__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2696, new_AGEMA_signal_2695, AddRoundKeyOutput[30]}), .Q ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_29__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2694, new_AGEMA_signal_2693, AddRoundKeyOutput[29]}), .Q ({ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_28__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, AddRoundKeyOutput[28]}), .Q ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_27__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2690, new_AGEMA_signal_2689, AddRoundKeyOutput[27]}), .Q ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_26__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2688, new_AGEMA_signal_2687, AddRoundKeyOutput[26]}), .Q ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_25__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2686, new_AGEMA_signal_2685, AddRoundKeyOutput[25]}), .Q ({ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_24__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2684, new_AGEMA_signal_2683, AddRoundKeyOutput[24]}), .Q ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_23__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2682, new_AGEMA_signal_2681, AddRoundKeyOutput[23]}), .Q ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_22__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2680, new_AGEMA_signal_2679, AddRoundKeyOutput[22]}), .Q ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_21__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2678, new_AGEMA_signal_2677, AddRoundKeyOutput[21]}), .Q ({ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_20__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, AddRoundKeyOutput[20]}), .Q ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_19__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2674, new_AGEMA_signal_2673, AddRoundKeyOutput[19]}), .Q ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_18__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2672, new_AGEMA_signal_2671, AddRoundKeyOutput[18]}), .Q ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_17__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2670, new_AGEMA_signal_2669, AddRoundKeyOutput[17]}), .Q ({ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_16__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2668, new_AGEMA_signal_2667, AddRoundKeyOutput[16]}), .Q ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_15__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2666, new_AGEMA_signal_2665, AddRoundKeyOutput[15]}), .Q ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_14__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2664, new_AGEMA_signal_2663, AddRoundKeyOutput[14]}), .Q ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_13__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2662, new_AGEMA_signal_2661, AddRoundKeyOutput[13]}), .Q ({ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_12__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2660, new_AGEMA_signal_2659, AddRoundKeyOutput[12]}), .Q ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_11__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2658, new_AGEMA_signal_2657, AddRoundKeyOutput[11]}), .Q ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_10__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2656, new_AGEMA_signal_2655, AddRoundKeyOutput[10]}), .Q ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_9__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2654, new_AGEMA_signal_2653, AddRoundKeyOutput[9]}), .Q ({ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_8__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2652, new_AGEMA_signal_2651, AddRoundKeyOutput[8]}), .Q ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_7__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2650, new_AGEMA_signal_2649, AddRoundKeyOutput[7]}), .Q ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_6__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2648, new_AGEMA_signal_2647, AddRoundKeyOutput[6]}), .Q ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_5__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2646, new_AGEMA_signal_2645, AddRoundKeyOutput[5]}), .Q ({ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_4__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2644, new_AGEMA_signal_2643, AddRoundKeyOutput[4]}), .Q ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2642, new_AGEMA_signal_2641, AddRoundKeyOutput[3]}), .Q ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2640, new_AGEMA_signal_2639, AddRoundKeyOutput[2]}), .Q ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2638, new_AGEMA_signal_2637, AddRoundKeyOutput[1]}), .Q ({ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, AddRoundKeyOutput[0]}), .Q ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_6__FF_FF ( .CK (clk_gated), .D (FSMUpdate[6]), .Q (FSMReg[6]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_5__FF_FF ( .CK (clk_gated), .D (FSMUpdate[5]), .Q (FSMReg[5]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_4__FF_FF ( .CK (clk_gated), .D (FSMUpdate[4]), .Q (FSMReg[4]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_3__FF_FF ( .CK (clk_gated), .D (FSMUpdate[3]), .Q (FSMReg[3]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_2__FF_FF ( .CK (clk_gated), .D (FSMUpdate[2]), .Q (FSMReg[2]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_1__FF_FF ( .CK (clk_gated), .D (FSMUpdate[1]), .Q (FSMReg[1]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_0__FF_FF ( .CK (clk_gated), .D (FSMUpdate[0]), .Q (FSMReg[0]), .QN () ) ;
    DFF_X1 selectsRegInst_s_current_state_reg_1__FF_FF ( .CK (clk_gated), .D (selectsNext[1]), .Q (selectsReg[1]), .QN () ) ;
    DFF_X1 selectsRegInst_s_current_state_reg_0__FF_FF ( .CK (clk_gated), .D (selectsNext[0]), .Q (selectsReg[0]), .QN () ) ;
    DFF_X1 done_reg_FF_FF ( .CK (clk_gated), .D (done_internal), .Q (done), .QN () ) ;
endmodule
